//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 1 0 0 1 0 1 1 0 0 1 0 0 0 0 0 1 1 1 0 1 0 1 1 1 1 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:44 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  AOI22_X1  g0006(.A1(G77), .A2(G244), .B1(G87), .B2(G250), .ZN(new_n207));
  INV_X1    g0007(.A(G116), .ZN(new_n208));
  INV_X1    g0008(.A(G270), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n207), .B1(new_n208), .B2(new_n209), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n211));
  INV_X1    g0011(.A(G226), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  OAI221_X1 g0013(.A(new_n211), .B1(new_n201), .B2(new_n212), .C1(new_n203), .C2(new_n213), .ZN(new_n214));
  AOI211_X1 g0014(.A(new_n210), .B(new_n214), .C1(G97), .C2(G257), .ZN(new_n215));
  INV_X1    g0015(.A(G1), .ZN(new_n216));
  INV_X1    g0016(.A(G20), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n215), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(KEYINPUT1), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT64), .ZN(new_n222));
  INV_X1    g0022(.A(G13), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n218), .A2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n217), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n202), .A2(new_n203), .ZN(new_n230));
  NAND2_X1  g0030(.A1(new_n230), .A2(G50), .ZN(new_n231));
  INV_X1    g0031(.A(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n220), .A2(KEYINPUT1), .B1(new_n229), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g0033(.A1(new_n222), .A2(new_n227), .A3(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G50), .B(G58), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT65), .ZN(new_n245));
  XOR2_X1   g0045(.A(G68), .B(G77), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(KEYINPUT73), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n252), .A2(KEYINPUT14), .ZN(new_n253));
  NAND2_X1  g0053(.A1(G33), .A2(G41), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G1), .A3(G13), .ZN(new_n255));
  OAI21_X1  g0055(.A(new_n216), .B1(G41), .B2(G45), .ZN(new_n256));
  AND2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(G238), .ZN(new_n258));
  INV_X1    g0058(.A(G274), .ZN(new_n259));
  OR2_X1    g0059(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  INV_X1    g0061(.A(G97), .ZN(new_n262));
  NOR2_X1   g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT66), .A2(G1698), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G232), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  OAI22_X1  g0068(.A1(new_n266), .A2(new_n212), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT3), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(new_n261), .ZN(new_n271));
  NAND2_X1  g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n263), .B1(new_n269), .B2(new_n273), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n258), .B(new_n260), .C1(new_n274), .C2(new_n255), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT13), .ZN(new_n276));
  INV_X1    g0076(.A(new_n255), .ZN(new_n277));
  XNOR2_X1  g0077(.A(KEYINPUT66), .B(G1698), .ZN(new_n278));
  AOI22_X1  g0078(.A1(new_n278), .A2(G226), .B1(G232), .B2(G1698), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NOR2_X1   g0082(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n283), .B2(new_n263), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT13), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n284), .A2(new_n285), .A3(new_n258), .A4(new_n260), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n276), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G179), .ZN(new_n289));
  NOR2_X1   g0089(.A1(new_n252), .A2(KEYINPUT14), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n291), .B1(new_n287), .B2(G169), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  AOI211_X1 g0093(.A(new_n293), .B(new_n290), .C1(new_n276), .C2(new_n286), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n253), .B(new_n289), .C1(new_n292), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  AND2_X1   g0096(.A1(new_n296), .A2(new_n228), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NOR2_X1   g0098(.A1(G20), .A2(G33), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n217), .A2(G33), .ZN(new_n301));
  INV_X1    g0101(.A(G77), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n300), .A2(new_n201), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n217), .A2(G68), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n298), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  XNOR2_X1  g0105(.A(new_n305), .B(KEYINPUT11), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n216), .A2(G13), .A3(G20), .ZN(new_n307));
  OAI21_X1  g0107(.A(KEYINPUT72), .B1(new_n307), .B2(G68), .ZN(new_n308));
  XOR2_X1   g0108(.A(new_n308), .B(KEYINPUT12), .Z(new_n309));
  OAI21_X1  g0109(.A(new_n297), .B1(G1), .B2(new_n217), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n306), .B(new_n309), .C1(new_n203), .C2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n295), .A2(new_n311), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n307), .A2(G77), .ZN(new_n313));
  XNOR2_X1  g0113(.A(KEYINPUT8), .B(G58), .ZN(new_n314));
  INV_X1    g0114(.A(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(KEYINPUT15), .B(G87), .Z(new_n316));
  INV_X1    g0116(.A(new_n301), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n315), .A2(new_n299), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g0118(.A(new_n318), .B1(new_n217), .B2(new_n302), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n313), .B1(new_n319), .B2(new_n298), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(new_n302), .B2(new_n310), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI221_X1 g0122(.A(new_n273), .B1(new_n213), .B2(new_n268), .C1(new_n266), .C2(new_n267), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n323), .B1(G107), .B2(new_n273), .ZN(new_n324));
  XNOR2_X1  g0124(.A(new_n324), .B(KEYINPUT68), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n277), .ZN(new_n326));
  INV_X1    g0126(.A(new_n260), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n257), .B2(G244), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n326), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G190), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n322), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  XNOR2_X1  g0131(.A(KEYINPUT69), .B(G200), .ZN(new_n332));
  INV_X1    g0132(.A(new_n332), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n333), .B1(new_n326), .B2(new_n328), .ZN(new_n334));
  OR2_X1    g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(G223), .ZN(new_n336));
  INV_X1    g0136(.A(G222), .ZN(new_n337));
  OAI221_X1 g0137(.A(new_n273), .B1(new_n336), .B2(new_n268), .C1(new_n266), .C2(new_n337), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n338), .B(new_n277), .C1(G77), .C2(new_n273), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n257), .A2(G226), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n339), .A2(new_n260), .A3(new_n340), .ZN(new_n341));
  OR2_X1    g0141(.A1(new_n341), .A2(G179), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n315), .A2(new_n317), .B1(G20), .B2(new_n204), .ZN(new_n343));
  INV_X1    g0143(.A(G150), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n343), .B1(new_n344), .B2(new_n300), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(new_n298), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n310), .A2(G50), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n307), .A2(new_n201), .ZN(new_n348));
  AND3_X1   g0148(.A1(new_n347), .A2(KEYINPUT67), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT67), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n346), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n341), .A2(new_n293), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n342), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G179), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n326), .A2(new_n354), .A3(new_n328), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n355), .A2(new_n321), .ZN(new_n356));
  AOI21_X1  g0156(.A(G169), .B1(new_n326), .B2(new_n328), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AND4_X1   g0158(.A1(new_n312), .A2(new_n335), .A3(new_n353), .A4(new_n358), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n271), .A2(new_n217), .A3(new_n272), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT7), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND4_X1  g0162(.A1(new_n271), .A2(KEYINPUT7), .A3(new_n217), .A4(new_n272), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n203), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g0164(.A(G159), .ZN(new_n365));
  NOR2_X1   g0165(.A1(new_n300), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g0166(.A1(G58), .A2(G68), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n367), .A2(KEYINPUT74), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT74), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n369), .A2(G58), .A3(G68), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n370), .A3(new_n230), .ZN(new_n371));
  AND2_X1   g0171(.A1(new_n371), .A2(G20), .ZN(new_n372));
  NOR3_X1   g0172(.A1(new_n364), .A2(new_n366), .A3(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  OAI21_X1  g0174(.A(KEYINPUT16), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(KEYINPUT7), .B1(new_n282), .B2(new_n217), .ZN(new_n376));
  INV_X1    g0176(.A(new_n363), .ZN(new_n377));
  OAI21_X1  g0177(.A(G68), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(new_n372), .ZN(new_n379));
  INV_X1    g0179(.A(new_n366), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT16), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n381), .A2(KEYINPUT75), .A3(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n375), .A2(new_n298), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n257), .A2(G232), .ZN(new_n385));
  INV_X1    g0185(.A(G87), .ZN(new_n386));
  NOR2_X1   g0186(.A1(new_n261), .A2(new_n386), .ZN(new_n387));
  OAI22_X1  g0187(.A1(new_n266), .A2(new_n336), .B1(new_n212), .B2(new_n268), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n273), .ZN(new_n389));
  OAI211_X1 g0189(.A(new_n260), .B(new_n385), .C1(new_n389), .C2(new_n255), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n390), .A2(G200), .ZN(new_n391));
  MUX2_X1   g0191(.A(new_n307), .B(new_n310), .S(new_n315), .Z(new_n392));
  AND3_X1   g0192(.A1(new_n384), .A2(new_n391), .A3(new_n392), .ZN(new_n393));
  OR2_X1    g0193(.A1(new_n390), .A2(new_n330), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n393), .A2(KEYINPUT78), .A3(KEYINPUT17), .A4(new_n394), .ZN(new_n395));
  INV_X1    g0195(.A(KEYINPUT17), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n384), .A2(new_n394), .A3(new_n391), .A4(new_n392), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT78), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n396), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n395), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n384), .A2(new_n392), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n390), .A2(new_n293), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n278), .A2(G223), .B1(G226), .B2(G1698), .ZN(new_n403));
  NOR2_X1   g0203(.A1(new_n403), .A2(new_n282), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n277), .B1(new_n404), .B2(new_n387), .ZN(new_n405));
  NAND4_X1  g0205(.A1(new_n405), .A2(new_n354), .A3(new_n260), .A4(new_n385), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n402), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  AOI21_X1  g0210(.A(KEYINPUT77), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n407), .B1(new_n384), .B2(new_n392), .ZN(new_n412));
  INV_X1    g0212(.A(KEYINPUT77), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT18), .ZN(new_n414));
  NOR2_X1   g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT76), .ZN(new_n416));
  AND3_X1   g0216(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT18), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n416), .B1(new_n412), .B2(KEYINPUT18), .ZN(new_n418));
  NOR2_X1   g0218(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n400), .B1(new_n415), .B2(new_n419), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT9), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n351), .A2(new_n421), .ZN(new_n422));
  OR2_X1    g0222(.A1(new_n341), .A2(new_n330), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n341), .A2(new_n332), .B1(KEYINPUT70), .B2(KEYINPUT10), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n346), .B(KEYINPUT9), .C1(new_n349), .C2(new_n350), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n422), .A2(new_n423), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  NOR2_X1   g0226(.A1(KEYINPUT70), .A2(KEYINPUT10), .ZN(new_n427));
  OR2_X1    g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n427), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT71), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n288), .A2(new_n432), .A3(G190), .ZN(new_n433));
  OAI21_X1  g0233(.A(KEYINPUT71), .B1(new_n287), .B2(new_n330), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n311), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n287), .A2(G200), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  NAND4_X1  g0237(.A1(new_n359), .A2(new_n420), .A3(new_n431), .A4(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  NOR2_X1   g0240(.A1(KEYINPUT5), .A2(G41), .ZN(new_n441));
  AND2_X1   g0241(.A1(KEYINPUT5), .A2(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(G274), .C1(new_n441), .C2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  OAI21_X1  g0244(.A(new_n440), .B1(new_n442), .B2(new_n441), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n445), .A2(new_n255), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n444), .B1(new_n446), .B2(G270), .ZN(new_n447));
  NAND2_X1  g0247(.A1(G264), .A2(G1698), .ZN(new_n448));
  INV_X1    g0248(.A(G257), .ZN(new_n449));
  OAI211_X1 g0249(.A(new_n273), .B(new_n448), .C1(new_n266), .C2(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G303), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n255), .B1(new_n282), .B2(new_n451), .ZN(new_n452));
  AND3_X1   g0252(.A1(new_n450), .A2(new_n452), .A3(KEYINPUT84), .ZN(new_n453));
  AOI21_X1  g0253(.A(KEYINPUT84), .B1(new_n450), .B2(new_n452), .ZN(new_n454));
  OAI211_X1 g0254(.A(G179), .B(new_n447), .C1(new_n453), .C2(new_n454), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n216), .A2(G33), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n307), .A2(new_n456), .A3(new_n228), .A4(new_n296), .ZN(new_n457));
  OR2_X1    g0257(.A1(new_n457), .A2(new_n208), .ZN(new_n458));
  INV_X1    g0258(.A(new_n307), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n208), .ZN(new_n460));
  AOI22_X1  g0260(.A1(new_n296), .A2(new_n228), .B1(G20), .B2(new_n208), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n462), .B(new_n217), .C1(G33), .C2(new_n262), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n461), .A2(KEYINPUT20), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT20), .B1(new_n461), .B2(new_n463), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n458), .B(new_n460), .C1(new_n464), .C2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT85), .B1(new_n455), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n445), .A2(new_n255), .ZN(new_n469));
  OAI21_X1  g0269(.A(new_n443), .B1(new_n469), .B2(new_n209), .ZN(new_n470));
  INV_X1    g0270(.A(KEYINPUT84), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n448), .B1(new_n280), .B2(new_n281), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(G257), .B2(new_n278), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n277), .B1(new_n273), .B2(G303), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n450), .A2(new_n452), .A3(KEYINPUT84), .ZN(new_n476));
  AOI21_X1  g0276(.A(new_n470), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT85), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n477), .A2(new_n478), .A3(G179), .A4(new_n466), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n466), .A2(G169), .ZN(new_n480));
  OAI21_X1  g0280(.A(KEYINPUT21), .B1(new_n477), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n447), .B1(new_n453), .B2(new_n454), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n482), .A2(new_n483), .A3(G169), .A4(new_n466), .ZN(new_n484));
  AOI22_X1  g0284(.A1(new_n468), .A2(new_n479), .B1(new_n481), .B2(new_n484), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n477), .A2(G190), .ZN(new_n486));
  INV_X1    g0286(.A(G200), .ZN(new_n487));
  OAI211_X1 g0287(.A(new_n486), .B(new_n467), .C1(new_n487), .C2(new_n477), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT6), .ZN(new_n490));
  AND2_X1   g0290(.A1(G97), .A2(G107), .ZN(new_n491));
  NOR2_X1   g0291(.A1(G97), .A2(G107), .ZN(new_n492));
  OAI21_X1  g0292(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(KEYINPUT6), .A2(G97), .ZN(new_n494));
  OAI21_X1  g0294(.A(KEYINPUT79), .B1(new_n494), .B2(G107), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT79), .ZN(new_n496));
  INV_X1    g0296(.A(G107), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(new_n497), .A3(KEYINPUT6), .A4(G97), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n493), .A2(new_n495), .A3(new_n498), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n499), .A2(G20), .B1(G77), .B2(new_n299), .ZN(new_n500));
  OAI21_X1  g0300(.A(G107), .B1(new_n376), .B2(new_n377), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n502), .A2(new_n298), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT80), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n297), .A2(new_n504), .A3(new_n307), .A4(new_n456), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G97), .ZN(new_n508));
  NOR2_X1   g0308(.A1(new_n459), .A2(G97), .ZN(new_n509));
  INV_X1    g0309(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT81), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n262), .B1(new_n505), .B2(new_n506), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT81), .ZN(new_n513));
  NOR3_X1   g0313(.A1(new_n512), .A2(new_n513), .A3(new_n509), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n503), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g0315(.A(KEYINPUT4), .ZN(new_n516));
  OAI21_X1  g0316(.A(G244), .B1(new_n280), .B2(new_n281), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n516), .B1(new_n517), .B2(new_n266), .ZN(new_n518));
  INV_X1    g0318(.A(G244), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n519), .B1(new_n271), .B2(new_n272), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(KEYINPUT4), .A3(new_n278), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n273), .A2(G250), .A3(G1698), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n518), .A2(new_n521), .A3(new_n462), .A4(new_n522), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n277), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n446), .A2(G257), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n524), .A2(new_n443), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n293), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n515), .B(new_n527), .C1(G179), .C2(new_n526), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n526), .A2(G200), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n297), .B1(new_n500), .B2(new_n501), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n508), .A2(KEYINPUT81), .A3(new_n510), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n513), .B1(new_n512), .B2(new_n509), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  AOI22_X1  g0333(.A1(new_n523), .A2(new_n277), .B1(G257), .B2(new_n446), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(G190), .A3(new_n443), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n529), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n528), .A2(new_n536), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT24), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n217), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT22), .ZN(new_n540));
  INV_X1    g0340(.A(KEYINPUT22), .ZN(new_n541));
  NAND4_X1  g0341(.A1(new_n273), .A2(new_n541), .A3(new_n217), .A4(G87), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n317), .A2(G116), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n497), .A2(G20), .ZN(new_n545));
  XNOR2_X1  g0345(.A(new_n545), .B(KEYINPUT23), .ZN(new_n546));
  INV_X1    g0346(.A(new_n546), .ZN(new_n547));
  AND4_X1   g0347(.A1(new_n538), .A2(new_n543), .A3(new_n544), .A4(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n540), .B2(new_n542), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n538), .B1(new_n549), .B2(new_n544), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n298), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n507), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT25), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n307), .A2(G107), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n552), .A2(G107), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n554), .A2(new_n553), .ZN(new_n557));
  OAI21_X1  g0357(.A(G250), .B1(new_n264), .B2(new_n265), .ZN(new_n558));
  NAND2_X1  g0358(.A1(G257), .A2(G1698), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n282), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(G294), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n261), .A2(new_n561), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n277), .B1(new_n560), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n446), .A2(G264), .ZN(new_n564));
  NAND3_X1  g0364(.A1(new_n563), .A2(new_n443), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n565), .A2(KEYINPUT86), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT86), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n563), .A2(new_n564), .A3(new_n567), .A4(new_n443), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n293), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n565), .A2(new_n354), .ZN(new_n570));
  OAI22_X1  g0370(.A1(new_n556), .A2(new_n557), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n572), .A2(KEYINPUT24), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n549), .A2(new_n538), .A3(new_n544), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n297), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n555), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n575), .A2(new_n576), .A3(new_n557), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n566), .A2(new_n330), .A3(new_n568), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n565), .A2(new_n487), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n386), .A2(new_n262), .A3(new_n497), .ZN(new_n582));
  OAI211_X1 g0382(.A(KEYINPUT19), .B(new_n582), .C1(new_n263), .C2(G20), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n217), .B(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT19), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n585), .B1(new_n301), .B2(new_n262), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n583), .A2(new_n584), .A3(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(new_n316), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n587), .A2(new_n298), .B1(new_n459), .B2(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  AOI21_X1  g0390(.A(new_n590), .B1(G87), .B2(new_n552), .ZN(new_n591));
  INV_X1    g0391(.A(new_n440), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n592), .A2(G250), .A3(new_n255), .ZN(new_n593));
  OAI21_X1  g0393(.A(new_n593), .B1(new_n259), .B2(new_n592), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n520), .A2(G1698), .B1(G33), .B2(G116), .ZN(new_n595));
  OAI21_X1  g0395(.A(G238), .B1(new_n264), .B2(new_n265), .ZN(new_n596));
  OAI21_X1  g0396(.A(KEYINPUT82), .B1(new_n596), .B2(new_n282), .ZN(new_n597));
  INV_X1    g0397(.A(KEYINPUT82), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n273), .A2(new_n278), .A3(new_n598), .A4(G238), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n595), .A2(new_n597), .A3(new_n599), .ZN(new_n600));
  AOI211_X1 g0400(.A(new_n330), .B(new_n594), .C1(new_n600), .C2(new_n277), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n600), .A2(new_n277), .ZN(new_n602));
  INV_X1    g0402(.A(new_n594), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n601), .B1(new_n332), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n594), .B1(new_n600), .B2(new_n277), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n606), .A2(G169), .ZN(new_n607));
  AOI211_X1 g0407(.A(G179), .B(new_n594), .C1(new_n600), .C2(new_n277), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n505), .A2(new_n506), .A3(new_n316), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n589), .A2(KEYINPUT83), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT83), .B1(new_n589), .B2(new_n610), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n591), .A2(new_n605), .B1(new_n609), .B2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n537), .A2(new_n571), .A3(new_n581), .A4(new_n614), .ZN(new_n615));
  NOR3_X1   g0415(.A1(new_n438), .A2(new_n489), .A3(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n431), .A2(KEYINPUT90), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT90), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n430), .A2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n617), .A2(new_n619), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n356), .A2(new_n357), .ZN(new_n621));
  AOI22_X1  g0421(.A1(new_n437), .A2(new_n621), .B1(new_n311), .B2(new_n295), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n409), .A2(new_n410), .ZN(new_n623));
  NOR2_X1   g0423(.A1(new_n412), .A2(KEYINPUT18), .ZN(new_n624));
  OAI22_X1  g0424(.A1(new_n622), .A2(new_n400), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  AND2_X1   g0426(.A1(new_n626), .A2(new_n353), .ZN(new_n627));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n604), .A2(new_n628), .A3(new_n332), .ZN(new_n629));
  OAI21_X1  g0429(.A(KEYINPUT88), .B1(new_n606), .B2(new_n333), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n629), .A2(new_n591), .A3(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT89), .ZN(new_n632));
  INV_X1    g0432(.A(new_n601), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT89), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n629), .A2(new_n591), .A3(new_n630), .A4(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n633), .A3(new_n635), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n569), .A2(new_n570), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(new_n577), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n468), .A2(new_n479), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n481), .A2(new_n484), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n581), .B(new_n536), .C1(new_n640), .C2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n638), .B1(new_n528), .B2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n614), .ZN(new_n646));
  OAI21_X1  g0446(.A(KEYINPUT26), .B1(new_n646), .B2(new_n528), .ZN(new_n647));
  INV_X1    g0447(.A(new_n607), .ZN(new_n648));
  OR2_X1    g0448(.A1(new_n648), .A2(KEYINPUT87), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n589), .A2(new_n610), .ZN(new_n650));
  INV_X1    g0450(.A(new_n608), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n648), .A2(KEYINPUT87), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n649), .A2(new_n650), .A3(new_n651), .A4(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n645), .A2(new_n654), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n627), .B1(new_n438), .B2(new_n655), .ZN(G369));
  NOR2_X1   g0456(.A1(new_n223), .A2(G20), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(new_n216), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n658), .A2(KEYINPUT27), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(G213), .A3(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G343), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g0463(.A(new_n663), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n664), .A2(new_n467), .ZN(new_n665));
  MUX2_X1   g0465(.A(new_n489), .B(new_n485), .S(new_n665), .Z(new_n666));
  INV_X1    g0466(.A(G330), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  AND2_X1   g0468(.A1(new_n571), .A2(new_n581), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n669), .B1(new_n577), .B2(new_n664), .ZN(new_n670));
  OAI21_X1  g0470(.A(new_n670), .B1(new_n571), .B2(new_n664), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n640), .A2(new_n664), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n485), .A2(new_n663), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n673), .A3(new_n675), .ZN(G399));
  NOR2_X1   g0476(.A1(new_n224), .A2(G41), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(G1), .ZN(new_n679));
  OR2_X1    g0479(.A1(new_n582), .A2(G116), .ZN(new_n680));
  OAI22_X1  g0480(.A1(new_n679), .A2(new_n680), .B1(new_n231), .B2(new_n678), .ZN(new_n681));
  XOR2_X1   g0481(.A(KEYINPUT91), .B(KEYINPUT28), .Z(new_n682));
  XNOR2_X1  g0482(.A(new_n681), .B(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(new_n528), .ZN(new_n684));
  AND3_X1   g0484(.A1(new_n529), .A2(new_n533), .A3(new_n535), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n685), .B1(new_n571), .B2(new_n485), .ZN(new_n686));
  AOI21_X1  g0486(.A(new_n684), .B1(new_n686), .B2(new_n581), .ZN(new_n687));
  OAI211_X1 g0487(.A(new_n647), .B(new_n653), .C1(new_n687), .C2(new_n638), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  AND3_X1   g0489(.A1(new_n688), .A2(new_n689), .A3(new_n664), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n614), .A2(new_n684), .A3(new_n637), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n653), .B1(new_n636), .B2(new_n637), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI221_X4 g0493(.A(new_n685), .B1(new_n577), .B2(new_n580), .C1(new_n571), .C2(new_n485), .ZN(new_n694));
  AOI21_X1  g0494(.A(KEYINPUT26), .B1(new_n694), .B2(new_n636), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n691), .B(new_n693), .C1(new_n695), .C2(new_n684), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(new_n664), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n690), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT92), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n455), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n475), .A2(new_n476), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n702), .A2(KEYINPUT92), .A3(G179), .A4(new_n447), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n565), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n705), .A2(new_n534), .A3(new_n606), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n699), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n705), .A2(new_n534), .A3(new_n606), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n708), .A2(KEYINPUT30), .A3(new_n701), .A4(new_n703), .ZN(new_n709));
  NOR3_X1   g0509(.A1(new_n705), .A2(new_n477), .A3(G179), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n710), .A2(new_n604), .A3(new_n526), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n707), .A2(new_n709), .A3(new_n711), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n712), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT93), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI21_X1  g0515(.A(KEYINPUT31), .B1(new_n712), .B2(new_n663), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  AOI211_X1 g0517(.A(new_n714), .B(KEYINPUT31), .C1(new_n712), .C2(new_n663), .ZN(new_n718));
  OAI21_X1  g0518(.A(KEYINPUT94), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n614), .A2(new_n571), .A3(new_n581), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  INV_X1    g0521(.A(new_n489), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n721), .A2(new_n722), .A3(new_n537), .A4(new_n664), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(KEYINPUT95), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n528), .A2(new_n536), .ZN(new_n725));
  NOR3_X1   g0525(.A1(new_n720), .A2(new_n489), .A3(new_n725), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT95), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n726), .A2(new_n727), .A3(new_n664), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n712), .A2(new_n663), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n732), .A2(new_n714), .A3(new_n713), .ZN(new_n733));
  INV_X1    g0533(.A(new_n718), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT94), .ZN(new_n735));
  NAND3_X1  g0535(.A1(new_n733), .A2(new_n734), .A3(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n719), .A2(new_n729), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n698), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(KEYINPUT96), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n698), .A2(new_n738), .A3(KEYINPUT96), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n683), .B1(new_n743), .B2(G1), .ZN(G364));
  AOI21_X1  g0544(.A(new_n679), .B1(G45), .B2(new_n657), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n666), .A2(new_n667), .ZN(new_n747));
  XOR2_X1   g0547(.A(new_n747), .B(KEYINPUT97), .Z(new_n748));
  OAI21_X1  g0548(.A(new_n746), .B1(new_n748), .B2(new_n668), .ZN(new_n749));
  NOR2_X1   g0549(.A1(G13), .A2(G33), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n751), .A2(G20), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT98), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n666), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n217), .A2(G190), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n354), .A2(G200), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(G311), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(G179), .A2(G200), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n756), .A2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G329), .ZN(new_n763));
  XOR2_X1   g0563(.A(KEYINPUT33), .B(G317), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n354), .A2(new_n487), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(new_n756), .ZN(new_n766));
  OAI221_X1 g0566(.A(new_n282), .B1(new_n762), .B2(new_n763), .C1(new_n764), .C2(new_n766), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n217), .B1(new_n761), .B2(G190), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  AOI211_X1 g0569(.A(new_n760), .B(new_n767), .C1(G294), .C2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n217), .A2(new_n330), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(new_n757), .ZN(new_n772));
  INV_X1    g0572(.A(KEYINPUT99), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n772), .A2(new_n773), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n332), .A2(new_n354), .A3(new_n756), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  AOI22_X1  g0580(.A1(new_n778), .A2(G322), .B1(new_n780), .B2(G283), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n332), .A2(new_n354), .A3(new_n771), .ZN(new_n782));
  INV_X1    g0582(.A(new_n782), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(G303), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n771), .A2(new_n765), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n785), .A2(KEYINPUT100), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(G326), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n770), .A2(new_n781), .A3(new_n784), .A4(new_n790), .ZN(new_n791));
  OAI22_X1  g0591(.A1(new_n788), .A2(new_n201), .B1(new_n386), .B2(new_n782), .ZN(new_n792));
  AOI21_X1  g0592(.A(new_n792), .B1(G107), .B2(new_n780), .ZN(new_n793));
  INV_X1    g0593(.A(new_n762), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(G159), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT32), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n768), .A2(new_n262), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n273), .B1(new_n766), .B2(new_n203), .ZN(new_n799));
  AOI21_X1  g0599(.A(new_n799), .B1(new_n778), .B2(G58), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n793), .A2(new_n798), .A3(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n758), .A2(new_n302), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n791), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n228), .B1(G20), .B2(new_n293), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n754), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n224), .A2(new_n273), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n232), .A2(new_n439), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(new_n247), .C2(new_n439), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n225), .A2(G355), .A3(new_n273), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n808), .B(new_n809), .C1(G116), .C2(new_n225), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n803), .A2(new_n804), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  AND2_X1   g0611(.A1(new_n755), .A2(new_n811), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n749), .B1(new_n746), .B2(new_n812), .ZN(new_n813));
  XOR2_X1   g0613(.A(new_n813), .B(KEYINPUT101), .Z(G396));
  NAND2_X1  g0614(.A1(new_n321), .A2(new_n663), .ZN(new_n815));
  OAI21_X1  g0615(.A(new_n815), .B1(new_n331), .B2(new_n334), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n358), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g0617(.A1(new_n356), .A2(new_n357), .A3(new_n663), .ZN(new_n818));
  INV_X1    g0618(.A(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n817), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n655), .B2(new_n663), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n818), .B1(new_n358), .B2(new_n816), .ZN(new_n822));
  OAI211_X1 g0622(.A(new_n664), .B(new_n822), .C1(new_n645), .C2(new_n654), .ZN(new_n823));
  AND2_X1   g0623(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g0624(.A(new_n738), .B(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n746), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n779), .A2(new_n203), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n273), .B1(new_n202), .B2(new_n768), .C1(new_n782), .C2(new_n201), .ZN(new_n828));
  INV_X1    g0628(.A(new_n758), .ZN(new_n829));
  AOI22_X1  g0629(.A1(new_n789), .A2(G137), .B1(G159), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n778), .A2(G143), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n830), .B(new_n831), .C1(new_n344), .C2(new_n766), .ZN(new_n832));
  INV_X1    g0632(.A(KEYINPUT34), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n827), .B(new_n828), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(G132), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n833), .B2(new_n832), .C1(new_n835), .C2(new_n762), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n777), .A2(new_n561), .ZN(new_n837));
  INV_X1    g0637(.A(G283), .ZN(new_n838));
  OAI221_X1 g0638(.A(new_n282), .B1(new_n758), .B2(new_n208), .C1(new_n838), .C2(new_n766), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n797), .B(new_n839), .C1(G311), .C2(new_n794), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n779), .A2(new_n386), .ZN(new_n841));
  AOI21_X1  g0641(.A(new_n841), .B1(new_n789), .B2(G303), .ZN(new_n842));
  OAI211_X1 g0642(.A(new_n840), .B(new_n842), .C1(new_n497), .C2(new_n782), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n836), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n804), .A2(new_n750), .ZN(new_n845));
  AOI22_X1  g0645(.A1(new_n844), .A2(new_n804), .B1(new_n302), .B2(new_n845), .ZN(new_n846));
  OAI211_X1 g0646(.A(new_n846), .B(new_n745), .C1(new_n751), .C2(new_n822), .ZN(new_n847));
  AND2_X1   g0647(.A1(new_n826), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(G384));
  INV_X1    g0649(.A(KEYINPUT40), .ZN(new_n850));
  INV_X1    g0650(.A(KEYINPUT38), .ZN(new_n851));
  INV_X1    g0651(.A(new_n661), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n401), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT76), .B1(new_n409), .B2(new_n410), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n409), .A2(KEYINPUT77), .A3(new_n410), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n412), .A2(new_n416), .A3(KEYINPUT18), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n413), .B1(new_n412), .B2(KEYINPUT18), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n854), .A2(new_n855), .A3(new_n856), .A4(new_n857), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n395), .A2(new_n399), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n853), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n409), .A2(new_n853), .A3(new_n397), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT37), .ZN(new_n862));
  XNOR2_X1  g0662(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n851), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  XNOR2_X1  g0664(.A(new_n861), .B(KEYINPUT37), .ZN(new_n865));
  OAI211_X1 g0665(.A(KEYINPUT38), .B(new_n865), .C1(new_n420), .C2(new_n853), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n311), .A2(new_n663), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n435), .B2(new_n436), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT103), .ZN(new_n870));
  AND3_X1   g0670(.A1(new_n295), .A2(new_n870), .A3(new_n311), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n870), .B1(new_n295), .B2(new_n311), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n295), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n437), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(new_n868), .ZN(new_n876));
  AOI21_X1  g0676(.A(new_n820), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n727), .B1(new_n726), .B2(new_n664), .ZN(new_n878));
  NOR4_X1   g0678(.A1(new_n615), .A2(KEYINPUT95), .A3(new_n489), .A4(new_n663), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n713), .A2(KEYINPUT104), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(new_n732), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n730), .A2(KEYINPUT104), .A3(new_n731), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n877), .B1(new_n880), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n850), .B1(new_n867), .B2(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n623), .A2(new_n624), .ZN(new_n887));
  OAI211_X1 g0687(.A(new_n401), .B(new_n852), .C1(new_n887), .C2(new_n400), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n888), .A2(new_n865), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(new_n851), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n890), .A2(new_n866), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n882), .B(new_n883), .C1(new_n878), .C2(new_n879), .ZN(new_n892));
  NAND4_X1  g0692(.A1(new_n891), .A2(KEYINPUT40), .A3(new_n892), .A4(new_n877), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n886), .A2(new_n893), .ZN(new_n894));
  XNOR2_X1  g0694(.A(new_n894), .B(KEYINPUT105), .ZN(new_n895));
  INV_X1    g0695(.A(new_n438), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n895), .B(new_n897), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(G330), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n823), .A2(new_n819), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n873), .A2(new_n876), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  OR2_X1    g0702(.A1(new_n867), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n887), .A2(new_n661), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT39), .ZN(new_n905));
  NOR3_X1   g0705(.A1(new_n860), .A2(new_n851), .A3(new_n863), .ZN(new_n906));
  AOI21_X1  g0706(.A(KEYINPUT38), .B1(new_n888), .B2(new_n865), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n312), .A2(KEYINPUT103), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n295), .A2(new_n870), .A3(new_n311), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(new_n663), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT39), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n908), .A2(new_n912), .A3(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n903), .A2(new_n904), .A3(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n626), .A2(new_n353), .ZN(new_n916));
  INV_X1    g0716(.A(new_n690), .ZN(new_n917));
  INV_X1    g0717(.A(new_n636), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n637), .B1(new_n644), .B2(new_n918), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n692), .B1(new_n919), .B2(new_n528), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n663), .B1(new_n920), .B2(new_n691), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n917), .B1(new_n689), .B2(new_n921), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n916), .B1(new_n922), .B2(new_n896), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n915), .B(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n899), .B(new_n924), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n925), .B1(new_n216), .B2(new_n657), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n208), .B1(new_n499), .B2(KEYINPUT35), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n927), .B(new_n229), .C1(KEYINPUT35), .C2(new_n499), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n928), .B(KEYINPUT36), .ZN(new_n929));
  NAND4_X1  g0729(.A1(new_n232), .A2(G77), .A3(new_n370), .A4(new_n368), .ZN(new_n930));
  XNOR2_X1  g0730(.A(new_n930), .B(KEYINPUT102), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(G50), .B2(new_n203), .ZN(new_n932));
  NAND3_X1  g0732(.A1(new_n932), .A2(G1), .A3(new_n223), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n926), .A2(new_n929), .A3(new_n933), .ZN(G367));
  OR2_X1    g0734(.A1(new_n591), .A2(new_n664), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n636), .A2(new_n935), .ZN(new_n936));
  MUX2_X1   g0736(.A(new_n935), .B(new_n936), .S(new_n653), .Z(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT106), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n537), .B1(new_n533), .B2(new_n664), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n528), .B1(new_n939), .B2(new_n571), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(new_n664), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n675), .A2(new_n939), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT42), .ZN(new_n943));
  AOI22_X1  g0743(.A1(new_n938), .A2(KEYINPUT43), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n684), .A2(new_n663), .ZN(new_n945));
  AND2_X1   g0745(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n672), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g0747(.A(new_n944), .B(new_n947), .Z(new_n948));
  NOR2_X1   g0748(.A1(new_n938), .A2(KEYINPUT43), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n948), .B(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(KEYINPUT107), .B(KEYINPUT41), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n677), .B(new_n951), .Z(new_n952));
  INV_X1    g0752(.A(KEYINPUT109), .ZN(new_n953));
  OAI221_X1 g0753(.A(new_n675), .B1(new_n671), .B2(new_n674), .C1(new_n668), .C2(new_n953), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n668), .A2(new_n953), .ZN(new_n955));
  XOR2_X1   g0755(.A(new_n954), .B(new_n955), .Z(new_n956));
  NAND2_X1  g0756(.A1(new_n743), .A2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT110), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n743), .A2(KEYINPUT110), .A3(new_n956), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n675), .A2(new_n673), .ZN(new_n961));
  INV_X1    g0761(.A(KEYINPUT108), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n946), .B(new_n961), .C1(new_n962), .C2(KEYINPUT44), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n962), .A2(KEYINPUT44), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n946), .A2(new_n961), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(new_n672), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n959), .A2(new_n960), .A3(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n952), .B1(new_n970), .B2(new_n743), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n216), .B1(new_n657), .B2(G45), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n950), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  INV_X1    g0774(.A(new_n806), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n805), .B1(new_n225), .B2(new_n588), .C1(new_n242), .C2(new_n975), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n789), .A2(G311), .B1(G97), .B2(new_n780), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n977), .B1(new_n451), .B2(new_n777), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n768), .A2(new_n497), .ZN(new_n979));
  OAI221_X1 g0779(.A(new_n282), .B1(new_n758), .B2(new_n838), .C1(new_n561), .C2(new_n766), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n782), .A2(new_n208), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n980), .C1(KEYINPUT46), .C2(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(KEYINPUT46), .B2(new_n981), .ZN(new_n983));
  AOI211_X1 g0783(.A(new_n978), .B(new_n983), .C1(G317), .C2(new_n794), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n768), .A2(new_n203), .ZN(new_n985));
  OAI221_X1 g0785(.A(new_n273), .B1(new_n758), .B2(new_n201), .C1(new_n365), .C2(new_n766), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G137), .C2(new_n794), .ZN(new_n987));
  AOI22_X1  g0787(.A1(G150), .A2(new_n778), .B1(new_n789), .B2(G143), .ZN(new_n988));
  OAI211_X1 g0788(.A(new_n987), .B(new_n988), .C1(new_n202), .C2(new_n782), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n779), .A2(new_n302), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n984), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g0792(.A(KEYINPUT111), .B(KEYINPUT47), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n992), .B(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n746), .B1(new_n994), .B2(new_n804), .ZN(new_n995));
  OAI211_X1 g0795(.A(new_n976), .B(new_n995), .C1(new_n938), .C2(new_n753), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n974), .A2(new_n996), .ZN(G387));
  NAND2_X1  g0797(.A1(new_n959), .A2(new_n960), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n998), .B(new_n677), .C1(new_n743), .C2(new_n956), .ZN(new_n999));
  INV_X1    g0799(.A(G322), .ZN(new_n1000));
  OAI22_X1  g0800(.A1(new_n788), .A2(new_n1000), .B1(new_n759), .B2(new_n766), .ZN(new_n1001));
  XOR2_X1   g0801(.A(new_n1001), .B(KEYINPUT113), .Z(new_n1002));
  INV_X1    g0802(.A(G317), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1002), .B1(new_n451), .B2(new_n758), .C1(new_n1003), .C2(new_n777), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(new_n1004), .B(KEYINPUT48), .ZN(new_n1005));
  OAI221_X1 g0805(.A(new_n1005), .B1(new_n838), .B2(new_n768), .C1(new_n561), .C2(new_n782), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT49), .ZN(new_n1007));
  OR2_X1    g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n794), .A2(G326), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1010));
  AOI21_X1  g0810(.A(new_n273), .B1(new_n780), .B2(G116), .ZN(new_n1011));
  NAND4_X1  g0811(.A1(new_n1008), .A2(new_n1009), .A3(new_n1010), .A4(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n777), .A2(new_n201), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n588), .A2(new_n768), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n273), .B1(new_n762), .B2(new_n344), .C1(new_n203), .C2(new_n758), .ZN(new_n1015));
  INV_X1    g0815(.A(new_n766), .ZN(new_n1016));
  AOI211_X1 g0816(.A(new_n1014), .B(new_n1015), .C1(new_n315), .C2(new_n1016), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n782), .A2(new_n302), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(G97), .B2(new_n780), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1017), .B(new_n1019), .C1(new_n365), .C2(new_n788), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1012), .B1(new_n1013), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT114), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n804), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n745), .B1(new_n671), .B2(new_n753), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n680), .A2(new_n225), .A3(new_n273), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(G107), .B2(new_n225), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n1026), .B(KEYINPUT112), .Z(new_n1027));
  NAND2_X1  g0827(.A1(new_n315), .A2(new_n201), .ZN(new_n1028));
  OR2_X1    g0828(.A1(new_n1028), .A2(KEYINPUT50), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n680), .B1(new_n1028), .B2(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(G68), .A2(G77), .ZN(new_n1031));
  NAND4_X1  g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n439), .A4(new_n1031), .ZN(new_n1032));
  OAI211_X1 g0832(.A(new_n806), .B(new_n1032), .C1(new_n239), .C2(new_n439), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1024), .B1(new_n805), .B2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n1023), .A2(new_n1035), .B1(new_n973), .B2(new_n956), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n999), .A2(new_n1036), .ZN(G393));
  NAND2_X1  g0837(.A1(new_n969), .A2(new_n973), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n946), .A2(new_n754), .ZN(new_n1039));
  OR2_X1    g0839(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n805), .B1(new_n262), .B2(new_n225), .C1(new_n250), .C2(new_n975), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1039), .A2(KEYINPUT115), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n203), .A2(new_n782), .B1(new_n779), .B2(new_n386), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n282), .B1(new_n794), .B2(G143), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n302), .B2(new_n768), .C1(new_n314), .C2(new_n758), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n365), .A2(new_n777), .B1(new_n788), .B2(new_n344), .ZN(new_n1046));
  INV_X1    g0846(.A(KEYINPUT51), .ZN(new_n1047));
  AOI211_X1 g0847(.A(new_n1043), .B(new_n1045), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1048), .B1(new_n1047), .B2(new_n1046), .C1(new_n201), .C2(new_n766), .ZN(new_n1049));
  OAI22_X1  g0849(.A1(new_n759), .A2(new_n777), .B1(new_n788), .B2(new_n1003), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1050), .B(KEYINPUT52), .ZN(new_n1051));
  OAI221_X1 g0851(.A(new_n282), .B1(new_n758), .B2(new_n561), .C1(new_n451), .C2(new_n766), .ZN(new_n1052));
  OAI22_X1  g0852(.A1(new_n497), .A2(new_n779), .B1(new_n782), .B2(new_n838), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n1052), .B(new_n1053), .C1(G116), .C2(new_n769), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1051), .B(new_n1054), .C1(new_n1000), .C2(new_n762), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1049), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n746), .B1(new_n1056), .B2(new_n804), .ZN(new_n1057));
  NAND4_X1  g0857(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1038), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n969), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n678), .B1(new_n998), .B2(new_n1060), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1059), .B1(new_n1061), .B2(new_n970), .ZN(new_n1062));
  INV_X1    g0862(.A(new_n1062), .ZN(G390));
  NAND3_X1  g0863(.A1(new_n896), .A2(new_n892), .A3(G330), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n627), .B(new_n1064), .C1(new_n698), .C2(new_n438), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n820), .A2(new_n667), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n901), .B1(new_n737), .B2(new_n1066), .ZN(new_n1067));
  AND3_X1   g0867(.A1(new_n892), .A2(new_n901), .A3(new_n1066), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n900), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n737), .A2(new_n901), .A3(new_n1066), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n818), .B1(new_n921), .B2(new_n817), .ZN(new_n1071));
  AND2_X1   g0871(.A1(new_n892), .A2(new_n1066), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1070), .B(new_n1071), .C1(new_n901), .C2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1065), .B1(new_n1069), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1068), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n912), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n906), .B2(new_n907), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n817), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n819), .B1(new_n697), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n1080), .B2(new_n901), .ZN(new_n1081));
  AOI22_X1  g0881(.A1(new_n908), .A2(new_n913), .B1(new_n902), .B2(new_n1077), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1076), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  AOI22_X1  g0883(.A1(new_n911), .A2(new_n869), .B1(new_n868), .B2(new_n875), .ZN(new_n1084));
  OAI211_X1 g0884(.A(new_n1077), .B(new_n891), .C1(new_n1071), .C2(new_n1084), .ZN(new_n1085));
  AND3_X1   g0885(.A1(new_n864), .A2(new_n866), .A3(KEYINPUT39), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT39), .B1(new_n890), .B2(new_n866), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1084), .B1(new_n819), .B2(new_n823), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n1086), .A2(new_n1087), .B1(new_n1088), .B2(new_n912), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1070), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1085), .A2(new_n1089), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1075), .A2(new_n1083), .A3(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1093));
  AND3_X1   g0893(.A1(new_n1093), .A2(KEYINPUT116), .A3(new_n1074), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT116), .B1(new_n1093), .B2(new_n1074), .ZN(new_n1095));
  OAI211_X1 g0895(.A(new_n677), .B(new_n1092), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n750), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n827), .B1(G87), .B2(new_n783), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n1098), .B1(new_n208), .B2(new_n777), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n768), .A2(new_n302), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n758), .A2(new_n262), .ZN(new_n1101));
  OAI221_X1 g0901(.A(new_n282), .B1(new_n762), .B2(new_n561), .C1(new_n497), .C2(new_n766), .ZN(new_n1102));
  NOR4_X1   g0902(.A1(new_n1099), .A2(new_n1100), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OAI21_X1  g0903(.A(new_n1103), .B1(new_n838), .B2(new_n788), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n282), .B1(new_n1016), .B2(G137), .ZN(new_n1105));
  XNOR2_X1  g0905(.A(KEYINPUT54), .B(G143), .ZN(new_n1106));
  OAI221_X1 g0906(.A(new_n1105), .B1(new_n365), .B2(new_n768), .C1(new_n758), .C2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g0907(.A(new_n1107), .B1(G125), .B2(new_n794), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n778), .A2(G132), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n782), .A2(new_n344), .ZN(new_n1110));
  XNOR2_X1  g0910(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(new_n1110), .B(new_n1111), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n789), .A2(G128), .B1(G50), .B2(new_n780), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n1108), .A2(new_n1109), .A3(new_n1112), .A4(new_n1113), .ZN(new_n1114));
  AND2_X1   g0914(.A1(new_n1104), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n1116), .A2(new_n804), .B1(new_n314), .B2(new_n845), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1097), .A2(new_n745), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n1093), .B2(new_n973), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1096), .A2(new_n1119), .ZN(G378));
  AND2_X1   g0920(.A1(new_n677), .A2(KEYINPUT57), .ZN(new_n1121));
  NAND3_X1  g0921(.A1(new_n886), .A2(G330), .A3(new_n893), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n617), .A2(new_n353), .A3(new_n619), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(KEYINPUT55), .ZN(new_n1124));
  INV_X1    g0924(.A(KEYINPUT55), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n617), .A2(new_n1125), .A3(new_n353), .A4(new_n619), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n351), .A2(new_n852), .ZN(new_n1127));
  XOR2_X1   g0927(.A(new_n1127), .B(KEYINPUT56), .Z(new_n1128));
  AND3_X1   g0928(.A1(new_n1124), .A2(new_n1126), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1128), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1122), .A2(new_n1132), .ZN(new_n1133));
  NAND4_X1  g0933(.A1(new_n1131), .A2(new_n886), .A3(G330), .A4(new_n893), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n915), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT120), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1133), .A2(new_n915), .A3(new_n1134), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1138), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n915), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1141), .A2(KEYINPUT120), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n1081), .A2(new_n1082), .A3(new_n1070), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1068), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n1074), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT116), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1146), .A2(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1093), .A2(KEYINPUT116), .A3(new_n1074), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1065), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1121), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n845), .A2(new_n201), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(new_n1016), .A2(G132), .B1(new_n769), .B2(G150), .ZN(new_n1153));
  INV_X1    g0953(.A(G128), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n1153), .B1(new_n777), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(G125), .ZN(new_n1156));
  OAI22_X1  g0956(.A1(new_n788), .A2(new_n1156), .B1(new_n782), .B2(new_n1106), .ZN(new_n1157));
  AOI211_X1 g0957(.A(new_n1155), .B(new_n1157), .C1(G137), .C2(new_n829), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT59), .ZN(new_n1159));
  AOI21_X1  g0959(.A(G41), .B1(new_n780), .B2(G159), .ZN(new_n1160));
  AOI21_X1  g0960(.A(G33), .B1(new_n794), .B2(G124), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(G97), .A2(new_n1016), .B1(new_n829), .B2(new_n316), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n1163), .B1(new_n838), .B2(new_n762), .ZN(new_n1164));
  NOR4_X1   g0964(.A1(new_n1164), .A2(G41), .A3(new_n273), .A4(new_n985), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n779), .A2(new_n202), .ZN(new_n1166));
  AOI211_X1 g0966(.A(new_n1018), .B(new_n1166), .C1(new_n778), .C2(G107), .ZN(new_n1167));
  OAI211_X1 g0967(.A(new_n1165), .B(new_n1167), .C1(new_n208), .C2(new_n788), .ZN(new_n1168));
  XNOR2_X1  g0968(.A(new_n1168), .B(KEYINPUT58), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n201), .B1(new_n280), .B2(G41), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1162), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(new_n1171), .B(KEYINPUT118), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n746), .B1(new_n1172), .B2(new_n804), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1152), .B(new_n1173), .C1(new_n1132), .C2(new_n751), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1151), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT119), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1133), .A2(new_n915), .A3(new_n1134), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1176), .B1(new_n1177), .B2(new_n1141), .ZN(new_n1178));
  NAND3_X1  g0978(.A1(new_n1137), .A2(KEYINPUT119), .A3(new_n1139), .ZN(new_n1179));
  AND2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1065), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1181), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n678), .A2(KEYINPUT57), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1180), .B1(new_n1184), .B2(new_n972), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1175), .A2(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(new_n1186), .ZN(G375));
  AND2_X1   g0987(.A1(new_n1069), .A2(new_n1073), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1188), .A2(new_n1065), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1189), .A2(KEYINPUT121), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT121), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1191), .A3(new_n1065), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n952), .ZN(new_n1194));
  NAND3_X1  g0994(.A1(new_n1193), .A2(new_n1194), .A3(new_n1075), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n901), .A2(new_n751), .ZN(new_n1196));
  OR2_X1    g0996(.A1(new_n1196), .A2(KEYINPUT122), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1196), .A2(KEYINPUT122), .ZN(new_n1198));
  OAI221_X1 g0998(.A(new_n282), .B1(new_n762), .B2(new_n451), .C1(new_n208), .C2(new_n766), .ZN(new_n1199));
  AOI211_X1 g0999(.A(new_n1014), .B(new_n1199), .C1(G107), .C2(new_n829), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n778), .A2(G283), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n990), .B1(new_n789), .B2(G294), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n783), .A2(G97), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n778), .A2(G137), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n829), .A2(G150), .ZN(new_n1206));
  OAI221_X1 g1006(.A(new_n273), .B1(new_n762), .B2(new_n1154), .C1(new_n766), .C2(new_n1106), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(G50), .B2(new_n769), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n1166), .B1(G159), .B2(new_n783), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1205), .A2(new_n1206), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n788), .A2(new_n835), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1204), .B1(new_n1210), .B2(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(new_n1212), .A2(new_n804), .B1(new_n203), .B2(new_n845), .ZN(new_n1213));
  NAND4_X1  g1013(.A1(new_n1197), .A2(new_n745), .A3(new_n1198), .A4(new_n1213), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n1188), .B2(new_n972), .ZN(new_n1215));
  INV_X1    g1015(.A(new_n1215), .ZN(new_n1216));
  NAND2_X1  g1016(.A1(new_n1195), .A2(new_n1216), .ZN(G381));
  INV_X1    g1017(.A(G378), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1186), .A2(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT123), .ZN(new_n1220));
  INV_X1    g1020(.A(G396), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n999), .A2(new_n1221), .A3(new_n1036), .A4(new_n848), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1219), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n974), .A2(new_n996), .A3(new_n1062), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1222), .A2(new_n1220), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1224), .A2(new_n1225), .A3(G381), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1223), .A2(new_n1226), .ZN(G407));
  OAI211_X1 g1027(.A(G407), .B(G213), .C1(G343), .C2(new_n1219), .ZN(G409));
  OAI21_X1  g1028(.A(G378), .B1(new_n1175), .B2(new_n1185), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n662), .A2(G213), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1140), .A2(new_n973), .A3(new_n1142), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1174), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT124), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n952), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1234), .A2(new_n1182), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT124), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1231), .A2(new_n1236), .A3(new_n1174), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1233), .A2(new_n1218), .A3(new_n1235), .A4(new_n1237), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1229), .A2(new_n1230), .A3(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1230), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1240), .A2(G2897), .ZN(new_n1241));
  XNOR2_X1  g1041(.A(new_n1241), .B(KEYINPUT125), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1239), .A2(new_n1243), .ZN(new_n1244));
  AND3_X1   g1044(.A1(new_n1188), .A2(KEYINPUT60), .A3(new_n1065), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1075), .A2(KEYINPUT60), .ZN(new_n1246));
  AOI211_X1 g1046(.A(new_n678), .B(new_n1245), .C1(new_n1193), .C2(new_n1246), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n848), .B1(new_n1247), .B2(new_n1215), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1245), .B1(new_n1193), .B2(new_n1246), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1249), .A2(new_n677), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1250), .A2(G384), .A3(new_n1216), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1244), .A2(new_n1252), .ZN(new_n1253));
  AND2_X1   g1053(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1239), .A2(new_n1254), .A3(new_n1243), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(KEYINPUT63), .A3(new_n1255), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(G393), .B(new_n1221), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(new_n1224), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1062), .B1(new_n974), .B2(new_n996), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT126), .ZN(new_n1261));
  NOR3_X1   g1061(.A1(new_n1259), .A2(new_n1260), .A3(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(G387), .A2(G390), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT126), .B1(new_n1263), .B2(new_n1224), .ZN(new_n1264));
  OAI21_X1  g1064(.A(new_n1258), .B1(new_n1262), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1261), .B1(new_n1259), .B2(new_n1260), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(new_n1257), .ZN(new_n1267));
  AOI21_X1  g1067(.A(KEYINPUT61), .B1(new_n1265), .B2(new_n1267), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1231), .A2(new_n1236), .A3(new_n1174), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1236), .B1(new_n1231), .B2(new_n1174), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  AOI21_X1  g1071(.A(G378), .B1(new_n1182), .B2(new_n1234), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1240), .B1(new_n1271), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1273), .A2(new_n1254), .A3(new_n1229), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT63), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1256), .A2(new_n1268), .A3(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1274), .A2(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT61), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  AOI211_X1 g1080(.A(new_n1252), .B(new_n1242), .C1(new_n1273), .C2(new_n1229), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1254), .B1(new_n1239), .B2(new_n1243), .ZN(new_n1282));
  NOR2_X1   g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT62), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1280), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1265), .A2(new_n1267), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1277), .B1(new_n1285), .B2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(new_n1219), .A2(new_n1229), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1254), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1286), .ZN(G402));
endmodule


