//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n720, new_n721, new_n722, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n202));
  NAND2_X1  g001(.A1(G43gat), .A2(G50gat), .ZN(new_n203));
  INV_X1    g002(.A(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(G43gat), .A2(G50gat), .ZN(new_n205));
  OAI21_X1  g004(.A(KEYINPUT15), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G29gat), .A2(G36gat), .ZN(new_n208));
  NOR3_X1   g007(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n209));
  OAI21_X1  g008(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT92), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  OAI211_X1 g011(.A(KEYINPUT92), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n214), .A2(KEYINPUT93), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT93), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n209), .B1(new_n215), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT94), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n208), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(new_n209), .ZN(new_n221));
  AND3_X1   g020(.A1(new_n212), .A2(new_n216), .A3(new_n213), .ZN(new_n222));
  AOI21_X1  g021(.A(new_n216), .B1(new_n212), .B2(new_n213), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n219), .B(new_n221), .C1(new_n222), .C2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(new_n224), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n207), .B1(new_n220), .B2(new_n225), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT95), .B(G50gat), .Z(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n228), .B2(G43gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n214), .A2(new_n221), .ZN(new_n230));
  NAND4_X1  g029(.A1(new_n229), .A2(new_n230), .A3(new_n206), .A4(new_n208), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n226), .A2(KEYINPUT17), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(G8gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(G1gat), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n238), .B2(G1gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n233), .B1(new_n237), .B2(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT97), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(G8gat), .B1(new_n235), .B2(new_n236), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n234), .B(KEYINPUT97), .C1(new_n238), .C2(G1gat), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n242), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT98), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n242), .A2(new_n243), .A3(KEYINPUT98), .A4(new_n244), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n240), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n232), .A2(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n231), .ZN(new_n251));
  OAI21_X1  g050(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(KEYINPUT94), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n253), .A2(new_n224), .A3(new_n208), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n251), .B1(new_n254), .B2(new_n207), .ZN(new_n255));
  OAI21_X1  g054(.A(KEYINPUT96), .B1(new_n255), .B2(KEYINPUT17), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n226), .A2(new_n231), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT96), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT17), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n250), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(new_n249), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n257), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n263), .A2(KEYINPUT18), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n202), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(new_n262), .B1(new_n255), .B2(KEYINPUT17), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n258), .B1(new_n257), .B2(new_n259), .ZN(new_n268));
  NOR3_X1   g067(.A1(new_n255), .A2(KEYINPUT96), .A3(KEYINPUT17), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n263), .A2(new_n264), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n270), .A2(KEYINPUT99), .A3(KEYINPUT18), .A4(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n266), .A2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n249), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  XOR2_X1   g074(.A(new_n264), .B(KEYINPUT13), .Z(new_n276));
  AND2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n270), .A2(new_n271), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT18), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G113gat), .B(G141gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(G197gat), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT11), .B(G169gat), .Z(new_n283));
  XNOR2_X1  g082(.A(new_n282), .B(new_n283), .ZN(new_n284));
  XNOR2_X1  g083(.A(KEYINPUT91), .B(KEYINPUT12), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n273), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n287), .B1(new_n273), .B2(new_n280), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  XNOR2_X1  g090(.A(G197gat), .B(G204gat), .ZN(new_n292));
  INV_X1    g091(.A(G211gat), .ZN(new_n293));
  INV_X1    g092(.A(G218gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n292), .B1(KEYINPUT22), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(G211gat), .B(G218gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n296), .B(new_n297), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n291), .B1(new_n298), .B2(KEYINPUT29), .ZN(new_n299));
  INV_X1    g098(.A(G141gat), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G148gat), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT73), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n300), .A2(KEYINPUT73), .A3(G148gat), .ZN(new_n304));
  INV_X1    g103(.A(G148gat), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(G141gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n303), .A2(new_n304), .A3(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G155gat), .A2(G162gat), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  INV_X1    g108(.A(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n308), .B1(new_n311), .B2(KEYINPUT2), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n307), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n301), .A2(new_n306), .B1(new_n314), .B2(KEYINPUT2), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n308), .A2(KEYINPUT72), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n314), .A2(G155gat), .A3(G162gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n316), .A2(new_n317), .A3(new_n311), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n313), .B1(new_n315), .B2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n299), .A2(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(G228gat), .ZN(new_n321));
  INV_X1    g120(.A(G233gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n320), .A2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT82), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n315), .A2(new_n318), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n326), .B1(new_n312), .B2(new_n307), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT29), .B1(new_n327), .B2(new_n291), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n298), .B1(new_n328), .B2(KEYINPUT81), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT29), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n330), .B1(new_n319), .B2(KEYINPUT3), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT81), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n325), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n298), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n335), .B1(new_n331), .B2(new_n332), .ZN(new_n336));
  OAI211_X1 g135(.A(new_n336), .B(KEYINPUT82), .C1(new_n332), .C2(new_n331), .ZN(new_n337));
  AOI21_X1  g136(.A(new_n324), .B1(new_n334), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n331), .A2(new_n298), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n323), .B1(new_n320), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(G22gat), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR3_X1   g140(.A1(new_n338), .A2(G22gat), .A3(new_n340), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n341), .B1(new_n342), .B2(KEYINPUT83), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344));
  OAI211_X1 g143(.A(new_n344), .B(G22gat), .C1(new_n338), .C2(new_n340), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n343), .A2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G78gat), .B(G106gat), .Z(new_n347));
  XNOR2_X1  g146(.A(new_n347), .B(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT80), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT79), .B(KEYINPUT31), .ZN(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n346), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g152(.A1(new_n338), .A2(new_n340), .ZN(new_n354));
  INV_X1    g153(.A(G22gat), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT85), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n352), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT84), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(KEYINPUT84), .B1(new_n338), .B2(new_n340), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n360), .A2(new_n361), .A3(G22gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n342), .A2(KEYINPUT85), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n362), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n353), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(KEYINPUT86), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT86), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n353), .A2(new_n364), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G15gat), .B(G43gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(G71gat), .B(G99gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT23), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT23), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n375), .B1(G169gat), .B2(G176gat), .ZN(new_n376));
  INV_X1    g175(.A(G169gat), .ZN(new_n377));
  INV_X1    g176(.A(G176gat), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n374), .B(new_n376), .C1(new_n377), .C2(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n380));
  NOR2_X1   g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g180(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(G183gat), .A2(G190gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n383), .B1(KEYINPUT64), .B2(KEYINPUT24), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT64), .A2(KEYINPUT24), .ZN(new_n385));
  OAI221_X1 g184(.A(new_n382), .B1(G183gat), .B2(G190gat), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n381), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n381), .A2(KEYINPUT65), .A3(new_n386), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n382), .B1(G183gat), .B2(G190gat), .ZN(new_n391));
  INV_X1    g190(.A(KEYINPUT24), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n391), .B1(new_n392), .B2(new_n383), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n380), .B1(new_n393), .B2(new_n379), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n389), .A2(new_n390), .A3(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n383), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n377), .A2(new_n378), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n397), .A2(KEYINPUT26), .A3(new_n373), .ZN(new_n398));
  AOI211_X1 g197(.A(new_n396), .B(new_n398), .C1(KEYINPUT26), .C2(new_n373), .ZN(new_n399));
  INV_X1    g198(.A(G183gat), .ZN(new_n400));
  OR2_X1    g199(.A1(new_n400), .A2(KEYINPUT66), .ZN(new_n401));
  AOI21_X1  g200(.A(G190gat), .B1(new_n401), .B2(KEYINPUT27), .ZN(new_n402));
  OR3_X1    g201(.A1(new_n400), .A2(KEYINPUT66), .A3(KEYINPUT27), .ZN(new_n403));
  AOI21_X1  g202(.A(KEYINPUT28), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XOR2_X1   g203(.A(KEYINPUT27), .B(G183gat), .Z(new_n405));
  INV_X1    g204(.A(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(G190gat), .ZN(new_n407));
  AND3_X1   g206(.A1(new_n406), .A2(KEYINPUT28), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n399), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n395), .A2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT68), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  XNOR2_X1  g211(.A(G113gat), .B(G120gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n413), .A2(KEYINPUT1), .ZN(new_n414));
  INV_X1    g213(.A(G127gat), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(G134gat), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(KEYINPUT67), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(G134gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(G127gat), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n416), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n416), .C1(new_n414), .C2(KEYINPUT67), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND3_X1  g222(.A1(new_n395), .A2(KEYINPUT68), .A3(new_n409), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n412), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n410), .A2(new_n411), .A3(new_n422), .A4(new_n421), .ZN(new_n426));
  NAND4_X1  g225(.A1(new_n425), .A2(G227gat), .A3(G233gat), .A4(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n372), .B1(new_n427), .B2(KEYINPUT32), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(KEYINPUT33), .B2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(new_n372), .ZN(new_n431));
  OR2_X1    g230(.A1(new_n431), .A2(KEYINPUT69), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(KEYINPUT69), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(KEYINPUT33), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n427), .A2(KEYINPUT32), .A3(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n430), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n425), .A2(new_n426), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT34), .ZN(new_n438));
  NAND2_X1  g237(.A1(G227gat), .A2(G233gat), .ZN(new_n439));
  AND3_X1   g238(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n438), .B1(new_n437), .B2(new_n439), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n430), .A2(new_n442), .A3(new_n435), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(KEYINPUT70), .A3(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT70), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n436), .A2(new_n447), .A3(new_n443), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n446), .A2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n423), .A2(new_n319), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(KEYINPUT4), .ZN(new_n451));
  INV_X1    g250(.A(KEYINPUT4), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n452), .B1(new_n423), .B2(new_n319), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT78), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(KEYINPUT78), .A3(new_n453), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n459));
  NAND2_X1  g258(.A1(G225gat), .A2(G233gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n421), .A2(KEYINPUT74), .A3(new_n422), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT74), .B1(new_n421), .B2(new_n422), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  XNOR2_X1  g264(.A(new_n319), .B(new_n291), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n461), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n458), .A2(new_n459), .A3(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n454), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n459), .B1(new_n469), .B2(new_n467), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n471), .B1(new_n465), .B2(new_n319), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT74), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n423), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(new_n471), .A3(new_n319), .A4(new_n462), .ZN(new_n475));
  INV_X1    g274(.A(new_n450), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n461), .B1(new_n472), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT77), .ZN(new_n479));
  AND3_X1   g278(.A1(new_n470), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n479), .B1(new_n470), .B2(new_n478), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n468), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(G1gat), .B(G29gat), .ZN(new_n483));
  XNOR2_X1  g282(.A(new_n483), .B(KEYINPUT0), .ZN(new_n484));
  XNOR2_X1  g283(.A(G57gat), .B(G85gat), .ZN(new_n485));
  XOR2_X1   g284(.A(new_n484), .B(new_n485), .Z(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n482), .A2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT6), .ZN(new_n489));
  OAI211_X1 g288(.A(new_n486), .B(new_n468), .C1(new_n480), .C2(new_n481), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n482), .A2(KEYINPUT6), .A3(new_n487), .ZN(new_n492));
  INV_X1    g291(.A(G226gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n493), .A2(new_n322), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n494), .A2(KEYINPUT29), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n495), .B1(new_n395), .B2(new_n409), .ZN(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n395), .B(new_n409), .C1(new_n493), .C2(new_n322), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n497), .A2(new_n335), .A3(new_n498), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n499), .A2(KEYINPUT71), .ZN(new_n500));
  INV_X1    g299(.A(new_n498), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n298), .B1(new_n501), .B2(new_n496), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(new_n499), .A3(KEYINPUT71), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n500), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g303(.A(G8gat), .B(G36gat), .ZN(new_n505));
  XNOR2_X1  g304(.A(G64gat), .B(G92gat), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n505), .B(new_n506), .Z(new_n507));
  OAI21_X1  g306(.A(KEYINPUT30), .B1(new_n504), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(new_n504), .ZN(new_n510));
  INV_X1    g309(.A(new_n507), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n509), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g311(.A1(new_n510), .A2(new_n511), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n508), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n491), .A2(new_n492), .B1(new_n512), .B2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT35), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n369), .A2(new_n449), .A3(new_n515), .A4(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT90), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n491), .A2(new_n492), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n512), .A2(new_n514), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n520), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(KEYINPUT90), .A3(new_n369), .A4(new_n449), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n519), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n444), .A2(new_n445), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n525), .B1(new_n366), .B2(new_n368), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n516), .B1(new_n526), .B2(new_n515), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT40), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n487), .B1(KEYINPUT87), .B2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n465), .A2(new_n466), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n460), .B1(new_n458), .B2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT39), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n532), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OR3_X1    g335(.A1(new_n472), .A2(new_n477), .A3(new_n461), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n456), .A2(new_n457), .B1(new_n465), .B2(new_n466), .ZN(new_n538));
  OAI211_X1 g337(.A(new_n537), .B(KEYINPUT39), .C1(new_n538), .C2(new_n460), .ZN(new_n539));
  NOR2_X1   g338(.A1(new_n530), .A2(KEYINPUT87), .ZN(new_n540));
  AND3_X1   g339(.A1(new_n536), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n536), .B2(new_n539), .ZN(new_n542));
  NOR2_X1   g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g342(.A1(new_n543), .A2(new_n488), .A3(new_n514), .A4(new_n512), .ZN(new_n544));
  XOR2_X1   g343(.A(KEYINPUT88), .B(KEYINPUT37), .Z(new_n545));
  AOI21_X1  g344(.A(new_n507), .B1(new_n504), .B2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT37), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n546), .B1(new_n547), .B2(new_n504), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n548), .A2(KEYINPUT38), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n502), .A2(new_n499), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT38), .B1(new_n550), .B2(KEYINPUT37), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n513), .B1(new_n546), .B2(new_n551), .ZN(new_n552));
  NAND4_X1  g351(.A1(new_n491), .A2(new_n549), .A3(new_n552), .A4(new_n492), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n369), .A2(new_n544), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT89), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n366), .A2(new_n368), .ZN(new_n557));
  INV_X1    g356(.A(new_n515), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT36), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n446), .A2(new_n559), .A3(new_n448), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n444), .A2(KEYINPUT36), .A3(new_n445), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n557), .A2(new_n558), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  NAND4_X1  g361(.A1(new_n369), .A2(new_n544), .A3(KEYINPUT89), .A4(new_n553), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  AOI21_X1  g363(.A(new_n290), .B1(new_n529), .B2(new_n564), .ZN(new_n565));
  OR2_X1    g364(.A1(G99gat), .A2(G106gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G99gat), .A2(G106gat), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G85gat), .A2(G92gat), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n569), .A2(KEYINPUT7), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT7), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n571), .A2(G85gat), .A3(G92gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n570), .A2(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(G85gat), .ZN(new_n574));
  INV_X1    g373(.A(G92gat), .ZN(new_n575));
  AOI22_X1  g374(.A1(KEYINPUT8), .A2(new_n567), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n568), .B1(new_n573), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n573), .A2(new_n576), .A3(new_n568), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  OAI211_X1 g379(.A(new_n232), .B(new_n580), .C1(new_n268), .C2(new_n269), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n573), .A2(new_n568), .A3(new_n576), .ZN(new_n582));
  NOR2_X1   g381(.A1(new_n582), .A2(new_n577), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n257), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g385(.A(G190gat), .B(G218gat), .Z(new_n587));
  NAND2_X1  g386(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n587), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n581), .A2(new_n589), .A3(new_n585), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n592));
  XNOR2_X1  g391(.A(G134gat), .B(G162gat), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n591), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n588), .A2(new_n594), .A3(new_n590), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT21), .ZN(new_n599));
  NAND2_X1  g398(.A1(G71gat), .A2(G78gat), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n604));
  AND2_X1   g403(.A1(G57gat), .A2(G64gat), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n600), .B(new_n603), .C1(new_n604), .C2(new_n605), .ZN(new_n606));
  NAND2_X1  g405(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g408(.A1(G71gat), .A2(G78gat), .ZN(new_n610));
  NOR2_X1   g409(.A1(G71gat), .A2(G78gat), .ZN(new_n611));
  OAI21_X1  g410(.A(new_n609), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  NAND3_X1  g411(.A1(KEYINPUT100), .A2(G57gat), .A3(G64gat), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n613), .B1(new_n610), .B2(KEYINPUT9), .ZN(new_n614));
  NOR3_X1   g413(.A1(new_n612), .A2(new_n614), .A3(KEYINPUT101), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT101), .ZN(new_n616));
  AOI22_X1  g415(.A1(new_n603), .A2(new_n600), .B1(new_n608), .B2(new_n607), .ZN(new_n617));
  AND2_X1   g416(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT9), .ZN(new_n619));
  AOI22_X1  g418(.A1(new_n618), .A2(G64gat), .B1(new_n600), .B2(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n616), .B1(new_n617), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n606), .B1(new_n615), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n249), .B1(new_n599), .B2(new_n622), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n623), .B(KEYINPUT104), .ZN(new_n624));
  XOR2_X1   g423(.A(G127gat), .B(G155gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT103), .ZN(new_n626));
  NAND2_X1  g425(.A1(G231gat), .A2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(KEYINPUT102), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n626), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n624), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n622), .A2(new_n599), .ZN(new_n631));
  XOR2_X1   g430(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(G183gat), .B(G211gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n630), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n630), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n622), .A2(new_n580), .ZN(new_n639));
  INV_X1    g438(.A(KEYINPUT10), .ZN(new_n640));
  OAI21_X1  g439(.A(KEYINPUT101), .B1(new_n612), .B2(new_n614), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n617), .A2(new_n616), .A3(new_n620), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n583), .A2(new_n643), .A3(new_n606), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  NAND4_X1  g444(.A1(new_n583), .A2(new_n643), .A3(KEYINPUT10), .A4(new_n606), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(G230gat), .A2(G233gat), .ZN(new_n648));
  XOR2_X1   g447(.A(new_n648), .B(KEYINPUT105), .Z(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g450(.A1(new_n639), .A2(new_n644), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n652), .B2(new_n650), .ZN(new_n653));
  XNOR2_X1  g452(.A(G120gat), .B(G148gat), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n654), .B(KEYINPUT106), .ZN(new_n655));
  XNOR2_X1  g454(.A(G176gat), .B(G204gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n653), .A2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n653), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n598), .A2(new_n638), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n565), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(new_n520), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n667), .B(new_n236), .ZN(G1324gat));
  INV_X1    g467(.A(KEYINPUT42), .ZN(new_n669));
  INV_X1    g468(.A(new_n521), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n565), .A2(new_n670), .A3(new_n665), .ZN(new_n671));
  XOR2_X1   g470(.A(KEYINPUT16), .B(G8gat), .Z(new_n672));
  INV_X1    g471(.A(new_n672), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n669), .B1(new_n671), .B2(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(new_n673), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(G8gat), .B2(new_n671), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n674), .B1(new_n676), .B2(new_n669), .ZN(G1325gat));
  AND2_X1   g476(.A1(new_n560), .A2(new_n561), .ZN(new_n678));
  INV_X1    g477(.A(new_n678), .ZN(new_n679));
  OAI21_X1  g478(.A(G15gat), .B1(new_n666), .B2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(new_n449), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n681), .A2(G15gat), .A3(new_n664), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n565), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(G1326gat));
  NOR2_X1   g483(.A1(new_n666), .A2(new_n369), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT43), .B(G22gat), .Z(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AND2_X1   g486(.A1(new_n596), .A2(new_n597), .ZN(new_n688));
  AND3_X1   g487(.A1(new_n556), .A2(new_n562), .A3(new_n563), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n527), .B1(new_n519), .B2(new_n523), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT44), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  OAI211_X1 g492(.A(KEYINPUT44), .B(new_n688), .C1(new_n689), .C2(new_n690), .ZN(new_n694));
  AND2_X1   g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n638), .B(KEYINPUT107), .Z(new_n696));
  XOR2_X1   g495(.A(new_n662), .B(KEYINPUT108), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NOR3_X1   g497(.A1(new_n696), .A2(new_n290), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n695), .A2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(G29gat), .B1(new_n700), .B2(new_n520), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT45), .ZN(new_n702));
  NOR3_X1   g501(.A1(new_n598), .A2(new_n638), .A3(new_n662), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n565), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n520), .A2(G29gat), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n702), .B1(new_n704), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g506(.A1(new_n565), .A2(KEYINPUT45), .A3(new_n703), .A4(new_n705), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n701), .A2(new_n707), .A3(new_n708), .ZN(G1328gat));
  OAI21_X1  g508(.A(G36gat), .B1(new_n700), .B2(new_n521), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n521), .A2(G36gat), .ZN(new_n711));
  INV_X1    g510(.A(new_n711), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT46), .B1(new_n704), .B2(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n704), .A2(KEYINPUT46), .A3(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n710), .A2(new_n713), .A3(new_n714), .ZN(G1329gat));
  NOR3_X1   g514(.A1(new_n704), .A2(G43gat), .A3(new_n681), .ZN(new_n716));
  NAND4_X1  g515(.A1(new_n693), .A2(new_n678), .A3(new_n694), .A4(new_n699), .ZN(new_n717));
  AOI21_X1  g516(.A(new_n716), .B1(G43gat), .B2(new_n717), .ZN(new_n718));
  XNOR2_X1  g517(.A(new_n718), .B(KEYINPUT47), .ZN(G1330gat));
  NOR3_X1   g518(.A1(new_n704), .A2(new_n228), .A3(new_n369), .ZN(new_n720));
  NAND4_X1  g519(.A1(new_n693), .A2(new_n557), .A3(new_n694), .A4(new_n699), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n720), .B1(new_n228), .B2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(KEYINPUT48), .ZN(G1331gat));
  NAND2_X1  g522(.A1(new_n598), .A2(new_n638), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n698), .A2(new_n290), .ZN(new_n725));
  AOI211_X1 g524(.A(new_n724), .B(new_n725), .C1(new_n529), .C2(new_n564), .ZN(new_n726));
  INV_X1    g525(.A(new_n520), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g528(.A(new_n521), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT109), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n726), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n732), .B(new_n733), .Z(G1333gat));
  AOI21_X1  g533(.A(new_n601), .B1(new_n726), .B2(new_n678), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n681), .A2(G71gat), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n735), .B1(new_n726), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n737), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g537(.A1(new_n726), .A2(new_n557), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G78gat), .ZN(G1335gat));
  INV_X1    g539(.A(new_n290), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n741), .A2(new_n638), .A3(new_n663), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n695), .A2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(G85gat), .B1(new_n743), .B2(new_n520), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n741), .A2(new_n638), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n688), .B(new_n745), .C1(new_n689), .C2(new_n690), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n520), .A2(G85gat), .A3(new_n663), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n749), .B(KEYINPUT110), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n748), .A2(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n744), .A2(new_n751), .ZN(G1336gat));
  NAND4_X1  g551(.A1(new_n748), .A2(new_n575), .A3(new_n670), .A4(new_n698), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n693), .A2(new_n670), .A3(new_n694), .A4(new_n742), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G92gat), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT52), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT52), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n753), .A2(new_n758), .A3(new_n755), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1337gat));
  XOR2_X1   g559(.A(KEYINPUT111), .B(G99gat), .Z(new_n761));
  NAND4_X1  g560(.A1(new_n748), .A2(new_n449), .A3(new_n662), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n743), .A2(new_n679), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n762), .B1(new_n763), .B2(new_n761), .ZN(G1338gat));
  INV_X1    g563(.A(KEYINPUT53), .ZN(new_n765));
  NOR3_X1   g564(.A1(new_n369), .A2(G106gat), .A3(new_n697), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n766), .B(KEYINPUT112), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n598), .B1(new_n529), .B2(new_n564), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(new_n768), .B2(new_n745), .ZN(new_n769));
  NOR2_X1   g568(.A1(new_n746), .A2(new_n747), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n767), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  NAND4_X1  g570(.A1(new_n693), .A2(new_n557), .A3(new_n694), .A4(new_n742), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n773), .A2(G106gat), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n772), .A2(KEYINPUT114), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n765), .B(new_n771), .C1(new_n774), .C2(new_n775), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n772), .A2(G106gat), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(new_n771), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n777), .B1(new_n779), .B2(KEYINPUT53), .ZN(new_n780));
  AOI211_X1 g579(.A(KEYINPUT113), .B(new_n765), .C1(new_n778), .C2(new_n771), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n776), .B1(new_n780), .B2(new_n781), .ZN(G1339gat));
  NOR2_X1   g581(.A1(new_n664), .A2(new_n741), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n645), .A2(new_n646), .A3(new_n649), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n651), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT115), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT115), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n651), .A2(new_n788), .A3(KEYINPUT54), .A4(new_n785), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n647), .A2(new_n790), .A3(new_n650), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n658), .ZN(new_n792));
  NAND4_X1  g591(.A1(new_n787), .A2(KEYINPUT55), .A3(new_n789), .A4(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT116), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n793), .A2(new_n794), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n791), .A2(new_n658), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n796), .B1(KEYINPUT115), .B2(new_n786), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n797), .A2(KEYINPUT116), .A3(KEYINPUT55), .A4(new_n789), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n789), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT55), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n659), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(new_n799), .B(new_n802), .C1(new_n288), .C2(new_n289), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n273), .A2(new_n280), .A3(new_n287), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n264), .B1(new_n270), .B2(new_n263), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n275), .A2(new_n276), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n284), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n804), .A2(new_n662), .A3(new_n807), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n688), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n804), .A2(new_n807), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n799), .A2(new_n802), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n598), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n784), .B1(new_n813), .B2(new_n696), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n814), .A2(new_n727), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(new_n526), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n670), .ZN(new_n817));
  AOI21_X1  g616(.A(G113gat), .B1(new_n817), .B2(new_n741), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n557), .A2(new_n681), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n814), .A2(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n727), .A2(new_n521), .ZN(new_n821));
  NOR2_X1   g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n741), .A2(G113gat), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n818), .B1(new_n822), .B2(new_n823), .ZN(G1340gat));
  AOI21_X1  g623(.A(G120gat), .B1(new_n817), .B2(new_n662), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n698), .A2(G120gat), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n822), .B2(new_n826), .ZN(G1341gat));
  NAND3_X1  g626(.A1(new_n817), .A2(new_n415), .A3(new_n638), .ZN(new_n828));
  INV_X1    g627(.A(new_n822), .ZN(new_n829));
  INV_X1    g628(.A(new_n696), .ZN(new_n830));
  OAI21_X1  g629(.A(G127gat), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n828), .A2(new_n831), .ZN(G1342gat));
  NOR4_X1   g631(.A1(new_n816), .A2(G134gat), .A3(new_n670), .A4(new_n598), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT56), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n418), .B1(new_n822), .B2(new_n688), .ZN(new_n835));
  XOR2_X1   g634(.A(new_n835), .B(KEYINPUT117), .Z(new_n836));
  NAND2_X1  g635(.A1(new_n834), .A2(new_n836), .ZN(G1343gat));
  NAND2_X1  g636(.A1(new_n679), .A2(new_n557), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n838), .B1(new_n815), .B2(KEYINPUT118), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n839), .B1(KEYINPUT118), .B2(new_n815), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n840), .A2(new_n670), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n741), .A2(new_n300), .ZN(new_n842));
  XNOR2_X1  g641(.A(new_n842), .B(KEYINPUT119), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT57), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n814), .A2(new_n845), .A3(new_n557), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n678), .A2(new_n821), .ZN(new_n847));
  INV_X1    g646(.A(new_n638), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n848), .B1(new_n809), .B2(new_n812), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n369), .B1(new_n849), .B2(new_n784), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n846), .B(new_n847), .C1(new_n845), .C2(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G141gat), .B1(new_n851), .B2(new_n290), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n844), .A2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT58), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n854), .B1(new_n852), .B2(KEYINPUT120), .ZN(new_n855));
  XNOR2_X1  g654(.A(new_n853), .B(new_n855), .ZN(G1344gat));
  NOR2_X1   g655(.A1(new_n305), .A2(KEYINPUT59), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n857), .B1(new_n851), .B2(new_n663), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT121), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n859), .B1(new_n850), .B2(KEYINPUT57), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n273), .A2(new_n280), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(new_n286), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n811), .B1(new_n862), .B2(new_n804), .ZN(new_n863));
  INV_X1    g662(.A(new_n808), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n598), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  OR3_X1    g664(.A1(new_n598), .A2(new_n810), .A3(new_n811), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n783), .B1(new_n867), .B2(new_n848), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT121), .B(new_n845), .C1(new_n868), .C2(new_n369), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n814), .A2(KEYINPUT57), .A3(new_n557), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n860), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n678), .A2(new_n663), .A3(new_n821), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(G148gat), .ZN(new_n874));
  AOI21_X1  g673(.A(KEYINPUT122), .B1(new_n871), .B2(new_n872), .ZN(new_n875));
  OAI211_X1 g674(.A(KEYINPUT123), .B(KEYINPUT59), .C1(new_n874), .C2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n872), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n880), .A2(G148gat), .A3(new_n873), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT123), .B1(new_n881), .B2(KEYINPUT59), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n858), .B1(new_n877), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n841), .A2(new_n305), .A3(new_n662), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n883), .A2(new_n884), .ZN(G1345gat));
  NOR3_X1   g684(.A1(new_n851), .A2(new_n309), .A3(new_n830), .ZN(new_n886));
  NOR3_X1   g685(.A1(new_n840), .A2(new_n670), .A3(new_n848), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n887), .A2(KEYINPUT124), .ZN(new_n888));
  AOI21_X1  g687(.A(G155gat), .B1(new_n887), .B2(KEYINPUT124), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n886), .B1(new_n888), .B2(new_n889), .ZN(G1346gat));
  OAI21_X1  g689(.A(G162gat), .B1(new_n851), .B2(new_n598), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n521), .A2(new_n310), .A3(new_n688), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n891), .B1(new_n840), .B2(new_n892), .ZN(G1347gat));
  NOR2_X1   g692(.A1(new_n727), .A2(new_n521), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n814), .A2(new_n819), .A3(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n895), .A2(new_n377), .A3(new_n290), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n814), .A2(new_n520), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n526), .A2(new_n670), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(new_n741), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n896), .B1(new_n901), .B2(new_n377), .ZN(G1348gat));
  OAI21_X1  g701(.A(G176gat), .B1(new_n895), .B2(new_n697), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n662), .A2(new_n378), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n903), .B1(new_n899), .B2(new_n904), .ZN(G1349gat));
  OAI21_X1  g704(.A(G183gat), .B1(new_n895), .B2(new_n830), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n638), .A2(new_n406), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n906), .B1(new_n899), .B2(new_n907), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g708(.A1(new_n900), .A2(new_n407), .A3(new_n688), .ZN(new_n910));
  OAI21_X1  g709(.A(G190gat), .B1(new_n895), .B2(new_n598), .ZN(new_n911));
  AND2_X1   g710(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n911), .A2(KEYINPUT61), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g713(.A(new_n914), .B(KEYINPUT125), .ZN(G1351gat));
  NOR2_X1   g714(.A1(new_n838), .A2(new_n521), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(new_n897), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g717(.A(G197gat), .B1(new_n918), .B2(new_n741), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n679), .A2(new_n894), .ZN(new_n920));
  XNOR2_X1  g719(.A(new_n920), .B(KEYINPUT126), .ZN(new_n921));
  AND2_X1   g720(.A1(new_n871), .A2(new_n921), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n741), .A2(G197gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(G1352gat));
  NOR3_X1   g723(.A1(new_n917), .A2(G204gat), .A3(new_n663), .ZN(new_n925));
  XNOR2_X1  g724(.A(KEYINPUT127), .B(KEYINPUT62), .ZN(new_n926));
  XNOR2_X1  g725(.A(new_n925), .B(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n698), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n928), .A2(G204gat), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n927), .A2(new_n929), .ZN(G1353gat));
  NAND3_X1  g729(.A1(new_n918), .A2(new_n293), .A3(new_n638), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n922), .A2(new_n638), .ZN(new_n932));
  AND3_X1   g731(.A1(new_n932), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n933));
  AOI21_X1  g732(.A(KEYINPUT63), .B1(new_n932), .B2(G211gat), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n933), .B2(new_n934), .ZN(G1354gat));
  NAND3_X1  g734(.A1(new_n918), .A2(new_n294), .A3(new_n688), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n922), .A2(new_n688), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n294), .ZN(G1355gat));
endmodule


