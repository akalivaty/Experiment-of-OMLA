//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 1 0 0 1 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 1 0 1 0 0 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n699, new_n700, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n727, new_n728, new_n729, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n769, new_n770, new_n771,
    new_n772, new_n773, new_n774, new_n775, new_n777, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n854, new_n855,
    new_n857, new_n858, new_n860, new_n861, new_n862, new_n863, new_n864,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n912, new_n913, new_n915, new_n916, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n958, new_n959;
  INV_X1    g000(.A(KEYINPUT95), .ZN(new_n202));
  NAND2_X1  g001(.A1(G228gat), .A2(G233gat), .ZN(new_n203));
  XOR2_X1   g002(.A(new_n203), .B(G22gat), .Z(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G148gat), .ZN(new_n206));
  INV_X1    g005(.A(G148gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n207), .A2(G141gat), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT81), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT2), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(G141gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n205), .A2(G148gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT81), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n209), .A2(new_n210), .A3(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G162gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n216), .A2(G155gat), .ZN(new_n217));
  INV_X1    g016(.A(G155gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G162gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT82), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT82), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(G141gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n223), .A3(G148gat), .ZN(new_n224));
  AOI21_X1  g023(.A(new_n220), .B1(new_n224), .B2(new_n211), .ZN(new_n225));
  AND2_X1   g024(.A1(KEYINPUT83), .A2(G162gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(KEYINPUT83), .A2(G162gat), .ZN(new_n227));
  NOR2_X1   g026(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(KEYINPUT2), .B1(new_n228), .B2(new_n218), .ZN(new_n229));
  AOI22_X1  g028(.A1(new_n215), .A2(new_n220), .B1(new_n225), .B2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT22), .ZN(new_n231));
  XOR2_X1   g030(.A(KEYINPUT77), .B(G211gat), .Z(new_n232));
  INV_X1    g031(.A(G218gat), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n232), .B2(new_n233), .ZN(new_n234));
  XNOR2_X1  g033(.A(G197gat), .B(G204gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G211gat), .B(G218gat), .ZN(new_n237));
  XNOR2_X1  g036(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT29), .ZN(new_n239));
  INV_X1    g038(.A(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n230), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(new_n238), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT29), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n230), .A2(new_n241), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n204), .B1(new_n242), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G78gat), .B(G106gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(G50gat), .ZN(new_n249));
  XNOR2_X1  g048(.A(KEYINPUT88), .B(KEYINPUT31), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n249), .B(new_n250), .ZN(new_n251));
  AND2_X1   g050(.A1(new_n251), .A2(KEYINPUT89), .ZN(new_n252));
  INV_X1    g051(.A(new_n246), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n214), .A2(new_n210), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n213), .B1(new_n211), .B2(new_n212), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n220), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n224), .A2(new_n211), .ZN(new_n257));
  INV_X1    g056(.A(new_n220), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n229), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n256), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n239), .B2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g060(.A(new_n204), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n253), .A2(new_n261), .A3(new_n262), .ZN(new_n263));
  AND3_X1   g062(.A1(new_n247), .A2(new_n252), .A3(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n251), .B(KEYINPUT89), .ZN(new_n265));
  AOI21_X1  g064(.A(new_n265), .B1(new_n247), .B2(new_n263), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT35), .ZN(new_n268));
  XNOR2_X1  g067(.A(G1gat), .B(G29gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n269), .B(KEYINPUT86), .ZN(new_n270));
  XNOR2_X1  g069(.A(G57gat), .B(G85gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(new_n270), .B(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(KEYINPUT85), .B(KEYINPUT0), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n271), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n270), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n273), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n274), .A2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT90), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n274), .A2(new_n278), .A3(KEYINPUT90), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(G225gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(G113gat), .A2(G120gat), .ZN(new_n289));
  INV_X1    g088(.A(G134gat), .ZN(new_n290));
  NOR2_X1   g089(.A1(new_n290), .A2(G127gat), .ZN(new_n291));
  AOI22_X1  g090(.A1(new_n288), .A2(new_n289), .B1(new_n291), .B2(KEYINPUT67), .ZN(new_n292));
  XNOR2_X1  g091(.A(G127gat), .B(G134gat), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT70), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT1), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI22_X1  g098(.A1(new_n286), .A2(new_n287), .B1(KEYINPUT70), .B2(KEYINPUT1), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT69), .ZN(new_n301));
  OAI211_X1 g100(.A(new_n299), .B(new_n300), .C1(new_n293), .C2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(G127gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(G134gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n290), .A2(G127gat), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n305), .A3(new_n301), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT68), .B(G120gat), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n306), .B1(new_n307), .B2(new_n286), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n296), .B1(new_n302), .B2(new_n308), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n260), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n287), .A2(KEYINPUT68), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT68), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(G120gat), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  AOI22_X1  g113(.A1(G113gat), .A2(new_n314), .B1(new_n293), .B2(new_n301), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n301), .B1(new_n304), .B2(new_n305), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n286), .A2(new_n287), .ZN(new_n317));
  NAND2_X1  g116(.A1(KEYINPUT70), .A2(KEYINPUT1), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n299), .A3(new_n318), .ZN(new_n319));
  NOR2_X1   g118(.A1(new_n316), .A2(new_n319), .ZN(new_n320));
  AOI22_X1  g119(.A1(new_n315), .A2(new_n320), .B1(new_n295), .B2(new_n292), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n230), .A2(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n285), .B1(new_n310), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n309), .B1(new_n230), .B2(new_n241), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n326));
  OAI21_X1  g125(.A(KEYINPUT84), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n321), .B1(new_n260), .B2(KEYINPUT3), .ZN(new_n328));
  INV_X1    g127(.A(KEYINPUT84), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n328), .A2(new_n329), .A3(new_n245), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n327), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  OAI21_X1  g131(.A(new_n332), .B1(new_n260), .B2(new_n309), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n230), .A2(new_n321), .A3(KEYINPUT4), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n333), .A2(new_n284), .A3(new_n334), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n324), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT5), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n333), .A2(new_n337), .A3(new_n334), .A4(new_n284), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n338), .B1(new_n327), .B2(new_n330), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n283), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n339), .A2(new_n279), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n342));
  AND4_X1   g141(.A1(new_n329), .A2(new_n342), .A3(new_n245), .A4(new_n309), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n329), .B1(new_n328), .B2(new_n245), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n335), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g144(.A1(new_n323), .A2(KEYINPUT5), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n341), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT6), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n340), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n279), .ZN(new_n351));
  INV_X1    g150(.A(new_n338), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n331), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n351), .B1(new_n347), .B2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT6), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  AND3_X1   g155(.A1(new_n267), .A2(new_n268), .A3(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT24), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n358), .A2(G183gat), .A3(G190gat), .ZN(new_n359));
  XNOR2_X1  g158(.A(G183gat), .B(G190gat), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n360), .B2(new_n358), .ZN(new_n361));
  NOR2_X1   g160(.A1(G169gat), .A2(G176gat), .ZN(new_n362));
  NAND2_X1  g161(.A1(G169gat), .A2(G176gat), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n362), .B1(KEYINPUT23), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(G169gat), .ZN(new_n365));
  INV_X1    g164(.A(G176gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT23), .ZN(new_n368));
  OAI21_X1  g167(.A(KEYINPUT25), .B1(new_n367), .B2(new_n368), .ZN(new_n369));
  NOR3_X1   g168(.A1(new_n361), .A2(new_n364), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(KEYINPUT23), .ZN(new_n371));
  AND2_X1   g170(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n372));
  NOR2_X1   g171(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n373));
  NOR3_X1   g172(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(KEYINPUT66), .B1(new_n374), .B2(new_n364), .ZN(new_n375));
  NOR2_X1   g174(.A1(new_n368), .A2(G169gat), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT65), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n377), .A2(new_n366), .ZN(new_n378));
  NAND2_X1  g177(.A1(KEYINPUT65), .A2(G176gat), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n376), .A2(new_n378), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT66), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n359), .ZN(new_n385));
  XOR2_X1   g184(.A(G183gat), .B(G190gat), .Z(new_n386));
  AOI21_X1  g185(.A(new_n385), .B1(new_n386), .B2(KEYINPUT24), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n375), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n370), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(KEYINPUT27), .B(G183gat), .ZN(new_n391));
  INV_X1    g190(.A(G190gat), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT28), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n391), .A2(KEYINPUT28), .A3(new_n392), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(new_n363), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n398), .A2(KEYINPUT26), .A3(new_n362), .ZN(new_n399));
  INV_X1    g198(.A(KEYINPUT26), .ZN(new_n400));
  INV_X1    g199(.A(G183gat), .ZN(new_n401));
  OAI22_X1  g200(.A1(new_n367), .A2(new_n400), .B1(new_n401), .B2(new_n392), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n399), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  OAI21_X1  g204(.A(new_n321), .B1(new_n390), .B2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n383), .B1(new_n380), .B2(new_n382), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n407), .A2(new_n361), .ZN(new_n408));
  AOI21_X1  g207(.A(KEYINPUT25), .B1(new_n408), .B2(new_n384), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n309), .B(new_n404), .C1(new_n409), .C2(new_n370), .ZN(new_n410));
  NAND2_X1  g209(.A1(G227gat), .A2(G233gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(KEYINPUT64), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n406), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT33), .ZN(new_n414));
  XOR2_X1   g213(.A(G15gat), .B(G43gat), .Z(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT72), .ZN(new_n416));
  XNOR2_X1  g215(.A(G71gat), .B(G99gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(new_n416), .B(new_n417), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n413), .B(KEYINPUT32), .C1(new_n414), .C2(new_n418), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n413), .B2(KEYINPUT32), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT71), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n413), .A2(new_n421), .A3(new_n414), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n420), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n421), .B1(new_n413), .B2(new_n414), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n419), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n406), .A2(new_n410), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT34), .ZN(new_n427));
  INV_X1    g226(.A(new_n412), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n426), .A2(new_n427), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(KEYINPUT73), .ZN(new_n430));
  AOI21_X1  g229(.A(new_n412), .B1(new_n406), .B2(new_n410), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(new_n432), .A3(new_n427), .ZN(new_n433));
  OAI211_X1 g232(.A(new_n430), .B(new_n433), .C1(new_n427), .C2(new_n431), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n425), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT76), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n413), .A2(new_n414), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(KEYINPUT71), .ZN(new_n438));
  NAND3_X1  g237(.A1(new_n438), .A2(new_n422), .A3(new_n420), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n427), .B1(new_n426), .B2(new_n428), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(KEYINPUT73), .B2(new_n429), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n439), .A2(new_n441), .A3(new_n419), .A4(new_n433), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n435), .A2(new_n436), .A3(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n425), .A2(KEYINPUT76), .A3(new_n434), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(G226gat), .A2(G233gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT78), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n244), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n390), .B2(new_n405), .ZN(new_n449));
  OAI211_X1 g248(.A(new_n404), .B(new_n447), .C1(new_n409), .C2(new_n370), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n449), .A2(new_n450), .A3(new_n243), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n243), .B1(new_n449), .B2(new_n450), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  XNOR2_X1  g253(.A(G8gat), .B(G36gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(G64gat), .B(G92gat), .ZN(new_n456));
  XOR2_X1   g255(.A(new_n455), .B(new_n456), .Z(new_n457));
  NAND4_X1  g256(.A1(new_n453), .A2(new_n454), .A3(KEYINPUT30), .A4(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n449), .A2(new_n450), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(new_n238), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n449), .A2(new_n450), .A3(new_n243), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n460), .A2(KEYINPUT30), .A3(new_n461), .A4(new_n457), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n453), .A2(new_n457), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT30), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n457), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(new_n451), .B2(new_n452), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT79), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT79), .ZN(new_n471));
  OAI211_X1 g270(.A(new_n471), .B(new_n468), .C1(new_n451), .C2(new_n452), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n464), .A2(new_n467), .A3(new_n473), .ZN(new_n474));
  AND3_X1   g273(.A1(new_n357), .A2(new_n445), .A3(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT87), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n353), .A2(new_n351), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n349), .B1(new_n477), .B2(new_n336), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n476), .B1(new_n478), .B2(new_n354), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n279), .B1(new_n336), .B2(new_n339), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n480), .A2(new_n348), .A3(KEYINPUT87), .A4(new_n349), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n479), .A2(new_n481), .A3(new_n355), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n482), .A2(new_n474), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n267), .A2(new_n435), .A3(new_n442), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT35), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  AND2_X1   g286(.A1(new_n435), .A2(new_n442), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n488), .A2(new_n482), .A3(new_n474), .A4(new_n267), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n489), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n475), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n435), .A2(KEYINPUT36), .A3(new_n442), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n492), .A2(KEYINPUT74), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT74), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n435), .A2(new_n442), .A3(new_n494), .A4(KEYINPUT36), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n497));
  NAND3_X1  g296(.A1(new_n443), .A2(new_n444), .A3(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT39), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n343), .A2(new_n344), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n333), .A2(new_n334), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n500), .B(new_n285), .C1(new_n501), .C2(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n310), .A2(new_n322), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n504), .B2(new_n284), .ZN(new_n505));
  AOI21_X1  g304(.A(new_n502), .B1(new_n327), .B2(new_n330), .ZN(new_n506));
  OAI21_X1  g305(.A(new_n505), .B1(new_n506), .B2(new_n284), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n281), .A2(new_n282), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n503), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(KEYINPUT91), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT40), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT91), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n510), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT92), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND4_X1  g315(.A1(new_n510), .A2(KEYINPUT92), .A3(new_n511), .A4(new_n513), .ZN(new_n517));
  NAND4_X1  g316(.A1(new_n503), .A2(new_n507), .A3(new_n508), .A4(KEYINPUT40), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n340), .ZN(new_n519));
  AOI22_X1  g318(.A1(new_n470), .A2(new_n472), .B1(new_n465), .B2(new_n466), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n519), .B1(new_n464), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n516), .A2(new_n517), .A3(new_n521), .ZN(new_n522));
  OR2_X1    g321(.A1(new_n264), .A2(new_n266), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT37), .ZN(new_n524));
  AOI21_X1  g323(.A(new_n457), .B1(new_n453), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT38), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT93), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n460), .A2(new_n527), .A3(new_n461), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n243), .A2(new_n527), .ZN(new_n529));
  AOI21_X1  g328(.A(new_n524), .B1(new_n452), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n525), .A2(new_n526), .A3(new_n531), .ZN(new_n532));
  AND3_X1   g331(.A1(new_n532), .A2(new_n350), .A3(new_n355), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n525), .B1(new_n524), .B2(new_n453), .ZN(new_n534));
  AOI22_X1  g333(.A1(new_n534), .A2(KEYINPUT38), .B1(new_n453), .B2(new_n457), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n523), .B1(new_n533), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n522), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n483), .A2(new_n523), .ZN(new_n538));
  AND3_X1   g337(.A1(new_n499), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n202), .B1(new_n491), .B2(new_n539), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n357), .A2(new_n445), .A3(new_n474), .ZN(new_n541));
  AND3_X1   g340(.A1(new_n489), .A2(KEYINPUT94), .A3(KEYINPUT35), .ZN(new_n542));
  AOI21_X1  g341(.A(KEYINPUT94), .B1(new_n489), .B2(KEYINPUT35), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AOI22_X1  g343(.A1(new_n522), .A2(new_n536), .B1(new_n483), .B2(new_n523), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n545), .A2(new_n499), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n544), .A2(KEYINPUT95), .A3(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT96), .B(G36gat), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g349(.A1(G29gat), .A2(G36gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(KEYINPUT14), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT15), .ZN(new_n553));
  OR3_X1    g352(.A1(new_n550), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G43gat), .B(G50gat), .ZN(new_n555));
  OR2_X1    g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n553), .B1(new_n550), .B2(new_n552), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n554), .A2(new_n557), .A3(new_n555), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n559), .B(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(G8gat), .ZN(new_n561));
  XNOR2_X1  g360(.A(G15gat), .B(G22gat), .ZN(new_n562));
  OR2_X1    g361(.A1(new_n562), .A2(G1gat), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n561), .B1(new_n563), .B2(KEYINPUT97), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT16), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n562), .B1(new_n565), .B2(G1gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n564), .B(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n560), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(G229gat), .A2(G233gat), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n559), .A2(new_n568), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT18), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(new_n559), .B(new_n568), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT98), .B(KEYINPUT13), .Z(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n571), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n576), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT99), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n576), .A2(KEYINPUT99), .A3(new_n578), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(new_n575), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(G197gat), .ZN(new_n586));
  XOR2_X1   g385(.A(KEYINPUT11), .B(G169gat), .Z(new_n587));
  XNOR2_X1  g386(.A(new_n586), .B(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(new_n588), .B(KEYINPUT12), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  AND2_X1   g389(.A1(new_n570), .A2(new_n572), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n591), .A2(KEYINPUT18), .A3(new_n571), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n584), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND3_X1  g392(.A1(new_n592), .A2(new_n575), .A3(new_n583), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n594), .A2(new_n589), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  AND3_X1   g395(.A1(new_n540), .A2(new_n547), .A3(new_n596), .ZN(new_n597));
  XOR2_X1   g396(.A(KEYINPUT101), .B(G57gat), .Z(new_n598));
  NAND2_X1  g397(.A1(new_n598), .A2(G64gat), .ZN(new_n599));
  INV_X1    g398(.A(G64gat), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n600), .A2(G57gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(G71gat), .ZN(new_n603));
  INV_X1    g402(.A(G78gat), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n603), .A2(new_n604), .A3(KEYINPUT9), .ZN(new_n605));
  AOI22_X1  g404(.A1(new_n599), .A2(new_n601), .B1(new_n602), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n607));
  XNOR2_X1  g406(.A(new_n606), .B(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n601), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n600), .A2(G57gat), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT9), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n602), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT100), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n604), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n612), .B1(new_n613), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g414(.A(new_n611), .B(new_n615), .C1(new_n613), .C2(new_n614), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n608), .A2(new_n616), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT21), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G231gat), .A2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n621), .B(new_n303), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n569), .B1(new_n617), .B2(new_n618), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G155gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(G183gat), .B(G211gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  OR2_X1    g427(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n624), .A2(new_n628), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g430(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n632));
  INV_X1    g431(.A(new_n559), .ZN(new_n633));
  NOR2_X1   g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  NAND2_X1  g433(.A1(G99gat), .A2(G106gat), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n634), .B1(KEYINPUT8), .B2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n636), .B(KEYINPUT104), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(G99gat), .B(G106gat), .Z(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  OAI21_X1  g441(.A(new_n632), .B1(new_n633), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n643), .B1(new_n560), .B2(new_n642), .ZN(new_n644));
  XOR2_X1   g443(.A(G190gat), .B(G218gat), .Z(new_n645));
  NAND2_X1  g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n646), .A2(KEYINPUT105), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT103), .B(G134gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(G162gat), .ZN(new_n649));
  AOI21_X1  g448(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n649), .B(new_n650), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g451(.A(new_n644), .B(new_n645), .ZN(new_n653));
  OR2_X1    g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n652), .A2(new_n653), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(new_n656), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n631), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g457(.A1(new_n617), .A2(new_n642), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n617), .A2(new_n642), .ZN(new_n660));
  OR3_X1    g459(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT10), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(KEYINPUT10), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(G230gat), .A2(G233gat), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n664), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n666), .B1(new_n659), .B2(new_n660), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  XNOR2_X1  g467(.A(G120gat), .B(G148gat), .ZN(new_n669));
  XNOR2_X1  g468(.A(G176gat), .B(G204gat), .ZN(new_n670));
  XOR2_X1   g469(.A(new_n669), .B(new_n670), .Z(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n665), .A2(new_n667), .A3(new_n671), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g474(.A1(new_n658), .A2(new_n675), .ZN(new_n676));
  OR2_X1    g475(.A1(new_n482), .A2(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n482), .A2(KEYINPUT106), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND3_X1  g479(.A1(new_n597), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g480(.A(new_n681), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g481(.A1(new_n597), .A2(new_n676), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n474), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n561), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  XNOR2_X1  g485(.A(KEYINPUT16), .B(G8gat), .ZN(new_n687));
  NOR3_X1   g486(.A1(new_n683), .A2(new_n474), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n689), .B1(KEYINPUT42), .B2(new_n688), .ZN(G1325gat));
  INV_X1    g489(.A(KEYINPUT107), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n499), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n496), .A2(KEYINPUT107), .A3(new_n498), .ZN(new_n693));
  AND2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g493(.A(G15gat), .B1(new_n683), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G15gat), .ZN(new_n696));
  NAND4_X1  g495(.A1(new_n597), .A2(new_n696), .A3(new_n445), .A4(new_n676), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1326gat));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n267), .ZN(new_n699));
  XOR2_X1   g498(.A(KEYINPUT43), .B(G22gat), .Z(new_n700));
  XNOR2_X1  g499(.A(new_n699), .B(new_n700), .ZN(G1327gat));
  NAND3_X1  g500(.A1(new_n540), .A2(new_n547), .A3(new_n656), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(KEYINPUT44), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT109), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n692), .A2(new_n545), .A3(new_n693), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n657), .B1(new_n705), .B2(new_n544), .ZN(new_n706));
  INV_X1    g505(.A(KEYINPUT44), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n704), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n703), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n702), .A2(new_n704), .A3(KEYINPUT44), .ZN(new_n710));
  AND2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n631), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n675), .A2(KEYINPUT108), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n712), .A2(new_n715), .A3(new_n596), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g516(.A(G29gat), .B1(new_n717), .B2(new_n679), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT45), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n631), .A2(new_n657), .A3(new_n675), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n597), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n680), .A2(new_n549), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n719), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  OR3_X1    g522(.A1(new_n721), .A2(new_n719), .A3(new_n722), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n718), .A2(new_n723), .A3(new_n724), .ZN(G1328gat));
  NAND2_X1  g524(.A1(new_n685), .A2(new_n548), .ZN(new_n726));
  OAI21_X1  g525(.A(KEYINPUT46), .B1(new_n721), .B2(new_n726), .ZN(new_n727));
  OR3_X1    g526(.A1(new_n721), .A2(KEYINPUT46), .A3(new_n726), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n717), .A2(new_n474), .ZN(new_n729));
  OAI211_X1 g528(.A(new_n727), .B(new_n728), .C1(new_n729), .C2(new_n548), .ZN(G1329gat));
  INV_X1    g529(.A(new_n694), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n709), .A2(new_n731), .A3(new_n710), .A4(new_n716), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(G43gat), .ZN(new_n733));
  INV_X1    g532(.A(new_n445), .ZN(new_n734));
  OR3_X1    g533(.A1(new_n721), .A2(G43gat), .A3(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n733), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g535(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n737));
  XNOR2_X1  g536(.A(new_n736), .B(new_n737), .ZN(G1330gat));
  NAND4_X1  g537(.A1(new_n709), .A2(new_n523), .A3(new_n710), .A4(new_n716), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NOR3_X1   g539(.A1(new_n721), .A2(G50gat), .A3(new_n267), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  NOR2_X1   g541(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT112), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n739), .A2(new_n745), .A3(G50gat), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n739), .B2(G50gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n746), .A2(new_n747), .A3(new_n741), .ZN(new_n748));
  XOR2_X1   g547(.A(KEYINPUT111), .B(KEYINPUT48), .Z(new_n749));
  OAI21_X1  g548(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(G1331gat));
  NOR3_X1   g549(.A1(new_n658), .A2(new_n715), .A3(new_n596), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT113), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n705), .A2(new_n544), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n751), .A2(new_n752), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n752), .B1(new_n751), .B2(new_n753), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n680), .ZN(new_n758));
  XOR2_X1   g557(.A(new_n758), .B(new_n598), .Z(G1332gat));
  INV_X1    g558(.A(KEYINPUT114), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(new_n755), .B2(new_n756), .ZN(new_n761));
  INV_X1    g560(.A(new_n756), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n762), .A2(KEYINPUT114), .A3(new_n754), .ZN(new_n763));
  AND2_X1   g562(.A1(new_n761), .A2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n685), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n765), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n766));
  XOR2_X1   g565(.A(KEYINPUT49), .B(G64gat), .Z(new_n767));
  OAI21_X1  g566(.A(new_n766), .B1(new_n765), .B2(new_n767), .ZN(G1333gat));
  NAND3_X1  g567(.A1(new_n761), .A2(new_n763), .A3(new_n731), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G71gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n757), .A2(new_n603), .A3(new_n445), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT50), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n770), .A2(KEYINPUT50), .A3(new_n771), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n774), .A2(new_n775), .ZN(G1334gat));
  NAND2_X1  g575(.A1(new_n764), .A2(new_n523), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g577(.A1(new_n631), .A2(new_n596), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n706), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT51), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT51), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n706), .A2(new_n782), .A3(new_n779), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n781), .A2(new_n783), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT115), .ZN(new_n785));
  INV_X1    g584(.A(new_n675), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n679), .A2(G85gat), .A3(new_n786), .ZN(new_n787));
  XNOR2_X1  g586(.A(new_n787), .B(KEYINPUT116), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n785), .A2(new_n788), .ZN(new_n789));
  NOR3_X1   g588(.A1(new_n631), .A2(new_n596), .A3(new_n786), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n711), .A2(new_n790), .ZN(new_n791));
  OAI21_X1  g590(.A(G85gat), .B1(new_n791), .B2(new_n679), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n789), .A2(new_n792), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n711), .A2(new_n685), .A3(new_n790), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(G92gat), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n715), .A2(G92gat), .A3(new_n474), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n784), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT117), .B1(KEYINPUT118), .B2(KEYINPUT51), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n706), .B2(new_n779), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT118), .B1(new_n780), .B2(KEYINPUT117), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n800), .B1(new_n801), .B2(new_n782), .ZN(new_n802));
  AOI22_X1  g601(.A1(new_n794), .A2(G92gat), .B1(new_n802), .B2(new_n796), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n798), .B1(new_n803), .B2(new_n804), .ZN(G1337gat));
  NOR3_X1   g604(.A1(new_n786), .A2(new_n734), .A3(G99gat), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n785), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(G99gat), .B1(new_n791), .B2(new_n694), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1338gat));
  NOR3_X1   g608(.A1(new_n715), .A2(G106gat), .A3(new_n267), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n781), .A2(new_n783), .A3(new_n810), .ZN(new_n811));
  XOR2_X1   g610(.A(KEYINPUT119), .B(KEYINPUT53), .Z(new_n812));
  NAND2_X1  g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n709), .A2(new_n523), .A3(new_n710), .A4(new_n790), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n813), .B1(new_n814), .B2(G106gat), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT120), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n815), .A2(new_n816), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT53), .ZN(new_n819));
  AOI22_X1  g618(.A1(new_n814), .A2(G106gat), .B1(new_n802), .B2(new_n810), .ZN(new_n820));
  OAI22_X1  g619(.A1(new_n817), .A2(new_n818), .B1(new_n819), .B2(new_n820), .ZN(G1339gat));
  NAND3_X1  g620(.A1(new_n661), .A2(new_n662), .A3(new_n666), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n665), .A2(KEYINPUT54), .A3(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n666), .B1(new_n661), .B2(new_n662), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n671), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n823), .A2(KEYINPUT55), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n674), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AND2_X1   g628(.A1(new_n823), .A2(new_n826), .ZN(new_n830));
  OAI211_X1 g629(.A(new_n829), .B(new_n596), .C1(KEYINPUT55), .C2(new_n830), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n591), .A2(new_n571), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n576), .A2(new_n578), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n588), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n675), .A2(new_n593), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n656), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n656), .B1(KEYINPUT55), .B2(new_n830), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n593), .A2(new_n834), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n837), .A2(new_n838), .A3(new_n828), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n712), .B1(new_n836), .B2(new_n839), .ZN(new_n840));
  INV_X1    g639(.A(new_n596), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n676), .A2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n679), .A2(new_n685), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n484), .ZN(new_n846));
  AND2_X1   g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n596), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n734), .A2(new_n523), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n843), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n844), .ZN(new_n851));
  NOR3_X1   g650(.A1(new_n851), .A2(new_n286), .A3(new_n841), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n848), .A2(new_n852), .ZN(G1340gat));
  NAND3_X1  g652(.A1(new_n847), .A2(new_n307), .A3(new_n675), .ZN(new_n854));
  OAI21_X1  g653(.A(G120gat), .B1(new_n851), .B2(new_n715), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n854), .A2(new_n855), .ZN(G1341gat));
  NAND3_X1  g655(.A1(new_n847), .A2(new_n303), .A3(new_n631), .ZN(new_n857));
  OAI21_X1  g656(.A(G127gat), .B1(new_n851), .B2(new_n712), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(G1342gat));
  NOR2_X1   g658(.A1(new_n657), .A2(G134gat), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n843), .A2(new_n846), .A3(new_n844), .A4(new_n860), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(KEYINPUT56), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n850), .A2(new_n656), .A3(new_n844), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(G134gat), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n865), .B1(new_n861), .B2(KEYINPUT56), .ZN(new_n866));
  AND3_X1   g665(.A1(new_n861), .A2(new_n865), .A3(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(KEYINPUT122), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  OAI211_X1 g669(.A(new_n864), .B(KEYINPUT122), .C1(new_n866), .C2(new_n867), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n870), .A2(new_n871), .ZN(G1343gat));
  AND2_X1   g671(.A1(new_n221), .A2(new_n223), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n694), .A2(new_n844), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n596), .A2(new_n674), .A3(new_n827), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n823), .A2(KEYINPUT124), .A3(new_n826), .ZN(new_n876));
  AOI21_X1  g675(.A(KEYINPUT124), .B1(new_n823), .B2(new_n826), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT55), .ZN(new_n878));
  OAI21_X1  g677(.A(new_n835), .B1(new_n875), .B2(new_n878), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n656), .B1(new_n879), .B2(KEYINPUT125), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT125), .ZN(new_n881));
  OAI211_X1 g680(.A(new_n881), .B(new_n835), .C1(new_n875), .C2(new_n878), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n839), .B1(new_n880), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n842), .B1(new_n883), .B2(new_n631), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n884), .A2(KEYINPUT57), .A3(new_n523), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n843), .A2(new_n523), .ZN(new_n886));
  XOR2_X1   g685(.A(KEYINPUT123), .B(KEYINPUT57), .Z(new_n887));
  NAND2_X1  g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n874), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n873), .B1(new_n889), .B2(new_n596), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n694), .A2(new_n523), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT126), .ZN(new_n892));
  OR2_X1    g691(.A1(new_n891), .A2(KEYINPUT126), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n845), .A2(new_n892), .A3(new_n893), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n894), .A2(G141gat), .A3(new_n841), .ZN(new_n895));
  OAI21_X1  g694(.A(KEYINPUT58), .B1(new_n890), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n894), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n897), .A2(new_n205), .A3(new_n596), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT58), .ZN(new_n899));
  AOI211_X1 g698(.A(new_n841), .B(new_n874), .C1(new_n885), .C2(new_n888), .ZN(new_n900));
  OAI211_X1 g699(.A(new_n898), .B(new_n899), .C1(new_n900), .C2(new_n873), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n896), .A2(new_n901), .ZN(G1344gat));
  AOI21_X1  g701(.A(KEYINPUT57), .B1(new_n884), .B2(new_n523), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n886), .A2(new_n887), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n694), .A2(new_n675), .A3(new_n844), .ZN(new_n906));
  OAI211_X1 g705(.A(KEYINPUT59), .B(G148gat), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT59), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n889), .A2(new_n908), .A3(new_n675), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n908), .B1(new_n897), .B2(new_n675), .ZN(new_n910));
  OAI211_X1 g709(.A(new_n907), .B(new_n909), .C1(G148gat), .C2(new_n910), .ZN(G1345gat));
  NAND3_X1  g710(.A1(new_n897), .A2(new_n218), .A3(new_n631), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n889), .A2(new_n631), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n913), .B2(new_n218), .ZN(G1346gat));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n656), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n657), .A2(new_n228), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n915), .A2(new_n228), .B1(new_n889), .B2(new_n916), .ZN(G1347gat));
  NOR2_X1   g716(.A1(new_n680), .A2(new_n474), .ZN(new_n918));
  INV_X1    g717(.A(new_n918), .ZN(new_n919));
  AOI211_X1 g718(.A(new_n484), .B(new_n919), .C1(new_n840), .C2(new_n842), .ZN(new_n920));
  AOI21_X1  g719(.A(G169gat), .B1(new_n920), .B2(new_n596), .ZN(new_n921));
  AND3_X1   g720(.A1(new_n843), .A2(new_n849), .A3(new_n918), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n841), .A2(new_n365), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(G1348gat));
  AOI21_X1  g723(.A(G176gat), .B1(new_n920), .B2(new_n675), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n715), .B1(new_n378), .B2(new_n379), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n922), .B2(new_n926), .ZN(G1349gat));
  NAND2_X1  g726(.A1(new_n922), .A2(new_n631), .ZN(new_n928));
  AND2_X1   g727(.A1(new_n631), .A2(new_n391), .ZN(new_n929));
  AOI22_X1  g728(.A1(new_n928), .A2(G183gat), .B1(new_n920), .B2(new_n929), .ZN(new_n930));
  XOR2_X1   g729(.A(new_n930), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g730(.A1(new_n920), .A2(new_n392), .A3(new_n656), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n922), .A2(new_n656), .ZN(new_n933));
  NOR2_X1   g732(.A1(KEYINPUT127), .A2(KEYINPUT61), .ZN(new_n934));
  AOI21_X1  g733(.A(new_n392), .B1(KEYINPUT127), .B2(KEYINPUT61), .ZN(new_n935));
  AND3_X1   g734(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n932), .B1(new_n936), .B2(new_n937), .ZN(G1351gat));
  NOR2_X1   g737(.A1(new_n731), .A2(new_n919), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n886), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(G197gat), .B1(new_n941), .B2(new_n596), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n905), .A2(new_n940), .ZN(new_n943));
  AND2_X1   g742(.A1(new_n596), .A2(G197gat), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n943), .B2(new_n944), .ZN(G1352gat));
  INV_X1    g744(.A(new_n941), .ZN(new_n946));
  INV_X1    g745(.A(G204gat), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n675), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g747(.A(KEYINPUT62), .B1(new_n946), .B2(new_n948), .ZN(new_n949));
  OR3_X1    g748(.A1(new_n946), .A2(KEYINPUT62), .A3(new_n948), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n905), .A2(new_n715), .A3(new_n940), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n949), .B(new_n950), .C1(new_n951), .C2(new_n947), .ZN(G1353gat));
  NAND3_X1  g751(.A1(new_n941), .A2(new_n232), .A3(new_n631), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n631), .B(new_n939), .C1(new_n903), .C2(new_n904), .ZN(new_n954));
  AND3_X1   g753(.A1(new_n954), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n955));
  AOI21_X1  g754(.A(KEYINPUT63), .B1(new_n954), .B2(G211gat), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(G1354gat));
  NAND3_X1  g756(.A1(new_n941), .A2(new_n233), .A3(new_n656), .ZN(new_n958));
  NOR3_X1   g757(.A1(new_n905), .A2(new_n657), .A3(new_n940), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n958), .B1(new_n959), .B2(new_n233), .ZN(G1355gat));
endmodule


