//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 0 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  INV_X1    g002(.A(G140), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G125), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(KEYINPUT16), .ZN(new_n191));
  INV_X1    g005(.A(G125), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G140), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(new_n193), .A3(KEYINPUT16), .ZN(new_n194));
  INV_X1    g008(.A(KEYINPUT82), .ZN(new_n195));
  AOI21_X1  g009(.A(new_n191), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NOR3_X1   g010(.A1(new_n190), .A2(KEYINPUT82), .A3(KEYINPUT16), .ZN(new_n197));
  OAI21_X1  g011(.A(new_n188), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(new_n197), .ZN(new_n199));
  XNOR2_X1  g013(.A(G125), .B(G140), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT82), .B1(new_n200), .B2(KEYINPUT16), .ZN(new_n201));
  OAI211_X1 g015(.A(G146), .B(new_n199), .C1(new_n201), .C2(new_n191), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n198), .A2(new_n202), .ZN(new_n203));
  AND2_X1   g017(.A1(KEYINPUT73), .A2(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(KEYINPUT73), .A2(G128), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT23), .A3(G119), .ZN(new_n207));
  INV_X1    g021(.A(G128), .ZN(new_n208));
  AOI21_X1  g022(.A(KEYINPUT23), .B1(new_n208), .B2(G119), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n208), .A2(G119), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n207), .A2(new_n211), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n210), .B1(new_n206), .B2(G119), .ZN(new_n213));
  XOR2_X1   g027(.A(KEYINPUT24), .B(G110), .Z(new_n214));
  AOI22_X1  g028(.A1(new_n212), .A2(G110), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n203), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT83), .ZN(new_n217));
  XNOR2_X1  g031(.A(new_n216), .B(new_n217), .ZN(new_n218));
  OAI22_X1  g032(.A1(new_n212), .A2(G110), .B1(new_n213), .B2(new_n214), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n188), .A2(KEYINPUT66), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT66), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(G146), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(new_n200), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n219), .A2(new_n225), .A3(new_n202), .ZN(new_n226));
  XNOR2_X1  g040(.A(new_n226), .B(KEYINPUT84), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n218), .A2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(G953), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT78), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(G953), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(KEYINPUT22), .B(G137), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n228), .A2(new_n237), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n218), .A2(new_n227), .A3(new_n236), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  OAI21_X1  g054(.A(new_n187), .B1(new_n240), .B2(G902), .ZN(new_n241));
  INV_X1    g055(.A(G902), .ZN(new_n242));
  NAND4_X1  g056(.A1(new_n238), .A2(KEYINPUT25), .A3(new_n242), .A4(new_n239), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  INV_X1    g058(.A(G217), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n245), .B1(G234), .B2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n240), .B(KEYINPUT85), .ZN(new_n248));
  INV_X1    g062(.A(new_n248), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n246), .A2(G902), .ZN(new_n250));
  INV_X1    g064(.A(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n247), .B1(new_n249), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(G472), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n220), .A2(new_n222), .A3(G143), .ZN(new_n254));
  INV_X1    g068(.A(G143), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT65), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n258), .A3(G146), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n254), .A2(new_n259), .A3(new_n260), .A4(G128), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n256), .A2(new_n258), .ZN(new_n262));
  AOI22_X1  g076(.A1(new_n255), .A2(new_n223), .B1(new_n262), .B2(new_n188), .ZN(new_n263));
  AOI21_X1  g077(.A(new_n206), .B1(new_n254), .B2(KEYINPUT1), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n261), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(G137), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(G134), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT72), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n269), .B1(G134), .B2(new_n266), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n267), .A2(new_n268), .ZN(new_n271));
  OAI21_X1  g085(.A(G131), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT70), .B1(new_n266), .B2(G134), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT70), .ZN(new_n274));
  INV_X1    g088(.A(G134), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(G137), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n273), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT69), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n278), .B1(new_n275), .B2(G137), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT11), .ZN(new_n280));
  INV_X1    g094(.A(G131), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT11), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n267), .A2(new_n278), .A3(new_n282), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n277), .A2(new_n280), .A3(new_n281), .A4(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT71), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n284), .A2(new_n285), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n265), .B(new_n272), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT77), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n282), .B1(new_n267), .B2(new_n278), .ZN(new_n290));
  AOI211_X1 g104(.A(KEYINPUT69), .B(KEYINPUT11), .C1(new_n266), .C2(G134), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND4_X1  g106(.A1(new_n292), .A2(KEYINPUT71), .A3(new_n281), .A4(new_n277), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n284), .A2(new_n285), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n292), .A2(new_n277), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n296), .A2(G131), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  AND2_X1   g112(.A1(KEYINPUT0), .A2(G128), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n254), .A2(new_n259), .A3(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT67), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n254), .A2(new_n259), .A3(KEYINPUT67), .A4(new_n299), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n257), .A2(G143), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n255), .A2(KEYINPUT65), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n188), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n306), .B1(new_n224), .B2(G143), .ZN(new_n307));
  NOR2_X1   g121(.A1(KEYINPUT0), .A2(G128), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n299), .A2(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n302), .A2(new_n303), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n298), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT2), .ZN(new_n312));
  INV_X1    g126(.A(G113), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(new_n313), .A3(KEYINPUT74), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT74), .ZN(new_n315));
  OAI21_X1  g129(.A(new_n315), .B1(KEYINPUT2), .B2(G113), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(KEYINPUT2), .A2(G113), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(G116), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G116), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n323), .A3(G119), .ZN(new_n324));
  INV_X1    g138(.A(G119), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G116), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n317), .A2(new_n324), .A3(new_n318), .A4(new_n326), .ZN(new_n329));
  AND3_X1   g143(.A1(new_n328), .A2(new_n329), .A3(KEYINPUT76), .ZN(new_n330));
  AOI21_X1  g144(.A(KEYINPUT76), .B1(new_n328), .B2(new_n329), .ZN(new_n331));
  NOR2_X1   g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT77), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n295), .A2(new_n333), .A3(new_n265), .A4(new_n272), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n289), .A2(new_n311), .A3(new_n332), .A4(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(new_n288), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n302), .A2(new_n303), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n307), .A2(new_n309), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT68), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g153(.A1(new_n293), .A2(new_n294), .B1(new_n296), .B2(G131), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n336), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n335), .B1(new_n343), .B2(new_n332), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n344), .A2(KEYINPUT28), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n338), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n332), .B(new_n288), .C1(new_n340), .C2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT28), .ZN(new_n348));
  AND3_X1   g162(.A1(new_n347), .A2(KEYINPUT79), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(KEYINPUT79), .B1(new_n347), .B2(new_n348), .ZN(new_n350));
  NOR2_X1   g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(G237), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n233), .A2(G210), .A3(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(new_n353), .B(KEYINPUT27), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT26), .B(G101), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n354), .B(new_n355), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n345), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  OR2_X1    g171(.A1(new_n330), .A2(new_n331), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n289), .A2(new_n311), .A3(KEYINPUT30), .A4(new_n334), .ZN(new_n359));
  XOR2_X1   g173(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n360));
  OAI211_X1 g174(.A(new_n358), .B(new_n359), .C1(new_n343), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(new_n335), .ZN(new_n362));
  INV_X1    g176(.A(new_n356), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT29), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n357), .A2(new_n364), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n334), .B1(new_n340), .B2(new_n346), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n265), .A2(new_n272), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n333), .B1(new_n368), .B2(new_n295), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n358), .B1(new_n367), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n348), .B1(new_n370), .B2(new_n335), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n332), .A2(new_n288), .ZN(new_n372));
  NOR2_X1   g186(.A1(new_n340), .A2(new_n346), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n348), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT79), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n347), .A2(KEYINPUT79), .A3(new_n348), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n371), .A2(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(new_n363), .A2(new_n365), .ZN(new_n380));
  AOI21_X1  g194(.A(G902), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n253), .B1(new_n366), .B2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n384));
  AOI211_X1 g198(.A(new_n384), .B(new_n253), .C1(new_n366), .C2(new_n381), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n361), .A2(new_n335), .A3(new_n356), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(KEYINPUT31), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n337), .A2(KEYINPUT68), .A3(new_n338), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n389), .A2(new_n339), .A3(new_n340), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n358), .B1(new_n390), .B2(new_n336), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n348), .B1(new_n391), .B2(new_n335), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n363), .B1(new_n392), .B2(new_n378), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT31), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n361), .A2(new_n394), .A3(new_n335), .A4(new_n356), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n388), .A2(new_n393), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n253), .A2(new_n242), .ZN(new_n397));
  XNOR2_X1  g211(.A(new_n397), .B(KEYINPUT80), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(KEYINPUT32), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT32), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n396), .A2(new_n401), .A3(new_n398), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n252), .B1(new_n386), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(KEYINPUT9), .B(G234), .ZN(new_n405));
  OAI21_X1  g219(.A(G221), .B1(new_n405), .B2(G902), .ZN(new_n406));
  INV_X1    g220(.A(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT88), .ZN(new_n409));
  INV_X1    g223(.A(G104), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT3), .B1(new_n410), .B2(G107), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT3), .ZN(new_n412));
  INV_X1    g226(.A(G107), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(new_n413), .A3(G104), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n410), .A2(G107), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(G101), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n415), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n410), .A2(G107), .ZN(new_n420));
  OAI21_X1  g234(.A(G101), .B1(new_n419), .B2(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n261), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n254), .A2(new_n259), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n260), .B1(new_n262), .B2(new_n188), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n424), .B1(new_n425), .B2(new_n208), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n423), .B1(new_n426), .B2(KEYINPUT87), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT87), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n424), .B(new_n428), .C1(new_n425), .C2(new_n208), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n409), .B(new_n422), .C1(new_n427), .C2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n208), .B1(new_n306), .B2(KEYINPUT1), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n254), .A2(new_n259), .ZN(new_n432));
  OAI21_X1  g246(.A(KEYINPUT87), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n433), .A2(new_n429), .A3(new_n261), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n418), .A2(new_n421), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT88), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n408), .B1(new_n430), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n411), .A2(new_n414), .A3(new_n415), .ZN(new_n438));
  OR2_X1    g252(.A1(new_n438), .A2(KEYINPUT86), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n417), .B1(new_n438), .B2(KEYINPUT86), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT4), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  AOI22_X1  g257(.A1(new_n439), .A2(new_n440), .B1(new_n417), .B2(new_n416), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n443), .B1(new_n444), .B2(new_n442), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n422), .A2(new_n408), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n445), .A2(new_n310), .B1(new_n265), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n437), .A2(new_n340), .A3(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT89), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n437), .A2(KEYINPUT89), .A3(new_n340), .A4(new_n447), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  OR2_X1    g266(.A1(new_n435), .A2(new_n265), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n430), .B2(new_n436), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n298), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT12), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n454), .A2(KEYINPUT12), .A3(new_n298), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n452), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n233), .A2(G227), .ZN(new_n461));
  XOR2_X1   g275(.A(G110), .B(G140), .Z(new_n462));
  XNOR2_X1  g276(.A(new_n461), .B(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n437), .A2(new_n447), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n298), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n450), .B2(new_n451), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT90), .ZN(new_n468));
  OAI21_X1  g282(.A(new_n466), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  AOI211_X1 g283(.A(KEYINPUT90), .B(new_n463), .C1(new_n450), .C2(new_n451), .ZN(new_n470));
  OAI211_X1 g284(.A(G469), .B(new_n464), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(G469), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n472), .A2(new_n242), .ZN(new_n473));
  INV_X1    g287(.A(new_n473), .ZN(new_n474));
  AND2_X1   g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n452), .A2(new_n466), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT91), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(new_n477), .A3(new_n463), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n450), .A2(new_n451), .B1(new_n465), .B2(new_n298), .ZN(new_n479));
  INV_X1    g293(.A(new_n463), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT91), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n467), .A2(new_n459), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n478), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(new_n472), .A3(new_n242), .ZN(new_n484));
  AOI21_X1  g298(.A(new_n407), .B1(new_n475), .B2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT17), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n233), .A2(G143), .A3(G214), .A4(new_n352), .ZN(new_n487));
  INV_X1    g301(.A(new_n262), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n230), .A2(new_n232), .A3(G214), .A4(new_n352), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI211_X1 g304(.A(new_n486), .B(new_n281), .C1(new_n487), .C2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(KEYINPUT95), .B1(new_n203), .B2(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n281), .B1(new_n487), .B2(new_n490), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT17), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT95), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n202), .A4(new_n198), .ZN(new_n496));
  INV_X1    g310(.A(new_n493), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n487), .A2(new_n281), .A3(new_n490), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n497), .A2(new_n486), .A3(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n492), .A2(new_n496), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n225), .B1(new_n188), .B2(new_n200), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n487), .A2(new_n490), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n503), .A2(new_n281), .ZN(new_n504));
  OAI221_X1 g318(.A(new_n501), .B1(new_n502), .B2(new_n504), .C1(new_n497), .C2(new_n503), .ZN(new_n505));
  XNOR2_X1  g319(.A(G113), .B(G122), .ZN(new_n506));
  XNOR2_X1  g320(.A(KEYINPUT94), .B(G104), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n506), .B(new_n507), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n505), .A3(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(new_n510), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n509), .B1(new_n500), .B2(new_n505), .ZN(new_n512));
  OAI21_X1  g326(.A(new_n242), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(G475), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT20), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT19), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n200), .B(new_n516), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n517), .A2(new_n223), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n196), .A2(new_n188), .A3(new_n197), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT93), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n497), .A2(new_n498), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n202), .B(new_n522), .C1(new_n223), .C2(new_n517), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n505), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(new_n508), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n526), .A2(new_n510), .ZN(new_n527));
  NOR2_X1   g341(.A1(G475), .A2(G902), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n515), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(new_n528), .ZN(new_n530));
  AOI211_X1 g344(.A(KEYINPUT20), .B(new_n530), .C1(new_n526), .C2(new_n510), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n514), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT98), .ZN(new_n534));
  AOI211_X1 g348(.A(new_n242), .B(new_n233), .C1(G234), .C2(G237), .ZN(new_n535));
  XOR2_X1   g349(.A(KEYINPUT21), .B(G898), .Z(new_n536));
  XNOR2_X1  g350(.A(new_n536), .B(KEYINPUT96), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G952), .ZN(new_n539));
  AOI211_X1 g353(.A(G953), .B(new_n539), .C1(G234), .C2(G237), .ZN(new_n540));
  INV_X1    g354(.A(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n538), .A2(new_n541), .ZN(new_n542));
  XOR2_X1   g356(.A(new_n542), .B(KEYINPUT97), .Z(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT75), .B(G116), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(G122), .ZN(new_n545));
  OR2_X1    g359(.A1(new_n320), .A2(G122), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n547), .A2(G107), .ZN(new_n548));
  INV_X1    g362(.A(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n544), .A2(KEYINPUT14), .A3(G122), .ZN(new_n550));
  OAI211_X1 g364(.A(G107), .B(new_n550), .C1(new_n547), .C2(KEYINPUT14), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n488), .A2(G128), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n206), .A2(G143), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(new_n275), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n275), .B1(new_n552), .B2(new_n553), .ZN(new_n556));
  OAI211_X1 g370(.A(new_n549), .B(new_n551), .C1(new_n555), .C2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(new_n547), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n558), .A2(new_n413), .ZN(new_n559));
  OAI21_X1  g373(.A(new_n554), .B1(new_n559), .B2(new_n548), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT13), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n552), .A2(new_n561), .B1(G143), .B2(new_n206), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n488), .A2(KEYINPUT13), .A3(G128), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n275), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n557), .B1(new_n560), .B2(new_n564), .ZN(new_n565));
  NOR3_X1   g379(.A1(new_n405), .A2(new_n245), .A3(G953), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI211_X1 g382(.A(new_n557), .B(new_n566), .C1(new_n560), .C2(new_n564), .ZN(new_n569));
  AOI21_X1  g383(.A(G902), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G478), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n570), .A2(KEYINPUT15), .A3(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(new_n571), .A2(KEYINPUT15), .ZN(new_n573));
  AOI211_X1 g387(.A(G902), .B(new_n573), .C1(new_n568), .C2(new_n569), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n572), .A2(new_n574), .ZN(new_n575));
  NAND4_X1  g389(.A1(new_n533), .A2(new_n534), .A3(new_n543), .A4(new_n575), .ZN(new_n576));
  OAI211_X1 g390(.A(new_n575), .B(new_n514), .C1(new_n529), .C2(new_n531), .ZN(new_n577));
  INV_X1    g391(.A(new_n543), .ZN(new_n578));
  OAI21_X1  g392(.A(KEYINPUT98), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n576), .A2(new_n579), .ZN(new_n580));
  OAI21_X1  g394(.A(G214), .B1(G237), .B2(G902), .ZN(new_n581));
  INV_X1    g395(.A(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n346), .A2(G125), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n265), .A2(G125), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(G224), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n586), .A2(G953), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT5), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n327), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n325), .A3(G116), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT92), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n313), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n592), .B1(new_n591), .B2(new_n590), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n435), .B(new_n329), .C1(new_n589), .C2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n329), .B1(new_n589), .B2(new_n593), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n422), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n594), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(G110), .B(G122), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT8), .ZN(new_n599));
  AOI22_X1  g413(.A1(new_n585), .A2(new_n587), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n358), .A2(new_n445), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n601), .A2(new_n594), .A3(new_n598), .ZN(new_n602));
  INV_X1    g416(.A(new_n587), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n583), .A2(KEYINPUT7), .A3(new_n603), .A4(new_n584), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n585), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n600), .A2(new_n602), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n607), .A2(new_n242), .ZN(new_n608));
  NOR2_X1   g422(.A1(new_n595), .A2(new_n422), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n609), .B1(new_n358), .B2(new_n445), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n598), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT6), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n614), .B1(new_n610), .B2(new_n598), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n585), .B(new_n587), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n611), .A2(new_n614), .A3(new_n612), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n616), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n608), .A2(new_n619), .ZN(new_n620));
  OAI21_X1  g434(.A(G210), .B1(G237), .B2(G902), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n608), .A2(new_n619), .A3(new_n621), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n582), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n404), .A2(new_n485), .A3(new_n580), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  AOI21_X1  g441(.A(new_n253), .B1(new_n396), .B2(new_n242), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT99), .ZN(new_n629));
  AND2_X1   g443(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n399), .B1(new_n628), .B2(new_n629), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n252), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n485), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n633), .B(KEYINPUT100), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n625), .A2(new_n543), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT101), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n571), .A2(G902), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT33), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n568), .A2(new_n638), .A3(new_n569), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n638), .B1(new_n568), .B2(new_n569), .ZN(new_n641));
  OAI211_X1 g455(.A(new_n636), .B(new_n637), .C1(new_n640), .C2(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n568), .A2(new_n569), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(KEYINPUT33), .ZN(new_n644));
  AOI211_X1 g458(.A(new_n571), .B(G902), .C1(new_n644), .C2(new_n639), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT101), .B1(new_n570), .B2(G478), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n642), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n532), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n635), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n634), .A2(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT102), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT34), .B(G104), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  NAND2_X1  g468(.A1(new_n527), .A2(new_n528), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT20), .ZN(new_n656));
  INV_X1    g470(.A(KEYINPUT103), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n527), .A2(new_n515), .A3(new_n528), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n656), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI22_X1  g473(.A1(new_n531), .A2(KEYINPUT103), .B1(new_n513), .B2(G475), .ZN(new_n660));
  OR2_X1    g474(.A1(new_n572), .A2(new_n574), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n635), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n634), .A2(new_n663), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT35), .B(G107), .Z(new_n665));
  XNOR2_X1  g479(.A(new_n664), .B(new_n665), .ZN(G9));
  NOR2_X1   g480(.A1(new_n630), .A2(new_n631), .ZN(new_n667));
  INV_X1    g481(.A(new_n625), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n237), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(KEYINPUT104), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n228), .B(new_n670), .ZN(new_n671));
  AOI22_X1  g485(.A1(new_n244), .A2(new_n246), .B1(new_n250), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g487(.A1(new_n485), .A2(new_n580), .A3(new_n667), .A4(new_n673), .ZN(new_n674));
  XOR2_X1   g488(.A(KEYINPUT37), .B(G110), .Z(new_n675));
  XNOR2_X1  g489(.A(new_n674), .B(new_n675), .ZN(G12));
  INV_X1    g490(.A(KEYINPUT106), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n370), .A2(new_n335), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(KEYINPUT28), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n351), .A3(new_n380), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n242), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n392), .A2(new_n378), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT29), .B1(new_n682), .B2(new_n356), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n681), .B1(new_n683), .B2(new_n364), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n384), .B1(new_n684), .B2(new_n253), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n382), .A2(KEYINPUT81), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n403), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(G900), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n540), .B1(new_n535), .B2(new_n688), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n659), .A2(new_n660), .A3(new_n661), .A4(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n687), .A2(new_n673), .A3(new_n693), .ZN(new_n694));
  AND3_X1   g508(.A1(new_n483), .A2(new_n472), .A3(new_n242), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n471), .A2(new_n474), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n406), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n677), .B1(new_n694), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n672), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n625), .ZN(new_n700));
  AOI21_X1  g514(.A(new_n700), .B1(new_n386), .B2(new_n403), .ZN(new_n701));
  NAND4_X1  g515(.A1(new_n701), .A2(new_n485), .A3(KEYINPUT106), .A4(new_n693), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G128), .ZN(G30));
  XOR2_X1   g518(.A(new_n689), .B(KEYINPUT39), .Z(new_n705));
  NAND2_X1  g519(.A1(new_n485), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(KEYINPUT40), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n362), .A2(new_n356), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n242), .B1(new_n678), .B2(new_n356), .ZN(new_n710));
  OAI21_X1  g524(.A(G472), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n699), .B1(new_n403), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n623), .A2(new_n624), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(KEYINPUT38), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n533), .A2(new_n575), .ZN(new_n715));
  AND4_X1   g529(.A1(new_n581), .A2(new_n712), .A3(new_n714), .A4(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT40), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n485), .A2(new_n717), .A3(new_n705), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n707), .A2(new_n716), .A3(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n262), .ZN(G45));
  OAI211_X1 g534(.A(new_n406), .B(new_n690), .C1(new_n695), .C2(new_n696), .ZN(new_n721));
  INV_X1    g535(.A(new_n649), .ZN(new_n722));
  NAND3_X1  g536(.A1(new_n687), .A2(new_n722), .A3(new_n673), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(new_n188), .ZN(G48));
  AOI21_X1  g539(.A(new_n472), .B1(new_n483), .B2(new_n242), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n695), .A2(new_n726), .A3(new_n407), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n404), .A3(new_n650), .ZN(new_n728));
  XOR2_X1   g542(.A(KEYINPUT41), .B(G113), .Z(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT107), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n727), .A2(new_n404), .A3(new_n663), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  AOI21_X1  g547(.A(new_n672), .B1(new_n576), .B2(new_n579), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n727), .A2(new_n625), .A3(new_n687), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  INV_X1    g550(.A(KEYINPUT108), .ZN(new_n737));
  OAI211_X1 g551(.A(new_n388), .B(new_n395), .C1(new_n356), .C2(new_n379), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n398), .ZN(new_n739));
  AOI21_X1  g553(.A(new_n628), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI22_X1  g554(.A1(new_n250), .A2(new_n248), .B1(new_n244), .B2(new_n246), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n738), .A2(KEYINPUT108), .A3(new_n398), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n740), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n715), .A2(new_n625), .A3(new_n543), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n745), .A2(new_n727), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G122), .ZN(G24));
  NAND2_X1  g561(.A1(new_n483), .A2(new_n242), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(G469), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n749), .A2(new_n406), .A3(new_n484), .A4(new_n625), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n649), .A2(new_n689), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(new_n740), .A3(new_n699), .A4(new_n742), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(new_n192), .ZN(G27));
  NAND3_X1  g568(.A1(new_n623), .A2(new_n581), .A3(new_n624), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT109), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n757), .B(new_n406), .C1(new_n695), .C2(new_n696), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n687), .A2(new_n741), .ZN(new_n759));
  NOR2_X1   g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(new_n751), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(new_n751), .ZN(new_n764));
  NOR4_X1   g578(.A1(new_n758), .A2(new_n759), .A3(new_n762), .A4(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(G131), .ZN(G33));
  NAND2_X1  g582(.A1(new_n760), .A2(new_n693), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n769), .B(G134), .ZN(G36));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n647), .A2(new_n532), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT43), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT111), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g589(.A(KEYINPUT111), .B(KEYINPUT43), .Z(new_n776));
  OAI21_X1  g590(.A(new_n776), .B1(new_n647), .B2(new_n532), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n778), .A2(new_n699), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n771), .B1(new_n779), .B2(new_n667), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n672), .B1(new_n775), .B2(new_n777), .ZN(new_n781));
  OAI211_X1 g595(.A(new_n781), .B(KEYINPUT44), .C1(new_n630), .C2(new_n631), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n757), .A3(new_n782), .ZN(new_n783));
  INV_X1    g597(.A(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n464), .B1(new_n469), .B2(new_n470), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT45), .ZN(new_n786));
  OR2_X1    g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n472), .B1(new_n785), .B2(new_n786), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n474), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT110), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n790), .A2(new_n791), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n473), .B1(new_n787), .B2(new_n788), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT110), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n795));
  AOI21_X1  g609(.A(new_n695), .B1(new_n794), .B2(KEYINPUT46), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n793), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n784), .A2(new_n797), .A3(new_n406), .A4(new_n705), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT112), .B(G137), .Z(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G39));
  XNOR2_X1  g614(.A(KEYINPUT113), .B(KEYINPUT47), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n801), .B1(new_n797), .B2(new_n406), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n406), .A3(new_n801), .ZN(new_n804));
  INV_X1    g618(.A(new_n687), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n805), .A2(new_n252), .A3(new_n751), .A4(new_n757), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n803), .A2(new_n804), .A3(new_n807), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G140), .ZN(G42));
  INV_X1    g623(.A(new_n714), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n727), .A2(new_n582), .A3(new_n810), .ZN(new_n811));
  OR2_X1    g625(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n778), .A2(new_n540), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n743), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n811), .A2(KEYINPUT117), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n812), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(KEYINPUT50), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT118), .ZN(new_n818));
  OR2_X1    g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n727), .A2(new_n757), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(new_n813), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n740), .A2(new_n699), .A3(new_n742), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n403), .A2(new_n741), .A3(new_n711), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n820), .A2(new_n541), .A3(new_n824), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n532), .A3(new_n648), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n695), .A2(new_n726), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n407), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n797), .A2(new_n406), .A3(new_n801), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n828), .B1(new_n829), .B2(new_n802), .ZN(new_n830));
  INV_X1    g644(.A(new_n757), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n813), .A2(new_n831), .A3(new_n743), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n823), .B(new_n826), .C1(new_n830), .C2(new_n832), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n817), .A2(new_n818), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n819), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n821), .A2(new_n759), .ZN(new_n838));
  XOR2_X1   g652(.A(new_n838), .B(KEYINPUT48), .Z(new_n839));
  INV_X1    g653(.A(new_n750), .ZN(new_n840));
  AOI211_X1 g654(.A(new_n539), .B(G953), .C1(new_n840), .C2(new_n814), .ZN(new_n841));
  OAI211_X1 g655(.A(new_n839), .B(new_n841), .C1(new_n649), .C2(new_n825), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n817), .A2(new_n836), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n842), .B1(new_n833), .B2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT116), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n659), .A2(new_n660), .A3(new_n575), .A4(new_n690), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n672), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n847), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n752), .B1(new_n805), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n697), .A2(new_n831), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n760), .A2(new_n693), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(KEYINPUT42), .B1(new_n760), .B2(new_n751), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n851), .B1(new_n852), .B2(new_n765), .ZN(new_n853));
  OAI22_X1  g667(.A1(new_n721), .A2(new_n723), .B1(new_n750), .B2(new_n752), .ZN(new_n854));
  INV_X1    g668(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n715), .A2(new_n625), .ZN(new_n856));
  INV_X1    g670(.A(new_n856), .ZN(new_n857));
  NAND4_X1  g671(.A1(new_n485), .A2(new_n690), .A3(new_n712), .A4(new_n857), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n855), .A2(new_n703), .A3(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT52), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n855), .A2(new_n703), .A3(KEYINPUT52), .A4(new_n858), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n853), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND2_X1   g677(.A1(new_n728), .A2(new_n746), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT114), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n865), .A3(new_n732), .A4(new_n735), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT115), .ZN(new_n867));
  OAI211_X1 g681(.A(new_n406), .B(new_n580), .C1(new_n695), .C2(new_n696), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n667), .A2(new_n673), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n687), .A2(new_n625), .A3(new_n741), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n868), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n577), .B1(new_n648), .B2(new_n533), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n635), .A2(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n485), .A2(new_n632), .A3(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n867), .B1(new_n871), .B2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n485), .A2(new_n632), .A3(new_n873), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n626), .A2(new_n674), .A3(new_n876), .A4(KEYINPUT115), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n875), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n735), .A2(new_n732), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n728), .A2(new_n746), .ZN(new_n880));
  OAI21_X1  g694(.A(KEYINPUT114), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n866), .A2(new_n878), .A3(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n882), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT53), .B1(new_n863), .B2(new_n882), .ZN(new_n884));
  OAI21_X1  g698(.A(KEYINPUT54), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT53), .ZN(new_n886));
  INV_X1    g700(.A(new_n853), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n854), .B1(new_n698), .B2(new_n702), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT52), .B1(new_n888), .B2(new_n858), .ZN(new_n889));
  INV_X1    g703(.A(new_n862), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n887), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n866), .A2(new_n878), .A3(new_n881), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n886), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT54), .ZN(new_n894));
  NOR3_X1   g708(.A1(new_n879), .A2(new_n880), .A3(new_n886), .ZN(new_n895));
  AND2_X1   g709(.A1(new_n895), .A2(new_n878), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n863), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n893), .A2(new_n894), .A3(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n837), .A2(new_n844), .A3(new_n885), .A4(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n539), .A2(new_n229), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n810), .A2(new_n406), .A3(new_n581), .A4(new_n772), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT49), .ZN(new_n903));
  NOR2_X1   g717(.A1(new_n827), .A2(new_n903), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n902), .A2(new_n904), .A3(new_n824), .ZN(new_n905));
  INV_X1    g719(.A(new_n827), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n905), .B1(KEYINPUT49), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n907), .ZN(G75));
  NOR2_X1   g722(.A1(new_n233), .A2(G952), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT119), .Z(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT56), .ZN(new_n912));
  INV_X1    g726(.A(new_n897), .ZN(new_n913));
  OAI21_X1  g727(.A(G902), .B1(new_n913), .B2(new_n884), .ZN(new_n914));
  INV_X1    g728(.A(G210), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n912), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n616), .A2(new_n618), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n617), .ZN(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT55), .Z(new_n919));
  INV_X1    g733(.A(new_n919), .ZN(new_n920));
  OR2_X1    g734(.A1(new_n916), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n916), .A2(new_n920), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n911), .B1(new_n921), .B2(new_n922), .ZN(G51));
  XNOR2_X1  g737(.A(new_n473), .B(KEYINPUT57), .ZN(new_n924));
  INV_X1    g738(.A(new_n898), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n894), .B1(new_n893), .B2(new_n897), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n924), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  XOR2_X1   g741(.A(new_n483), .B(KEYINPUT120), .Z(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  OR2_X1    g743(.A1(new_n914), .A2(new_n789), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n909), .B1(new_n929), .B2(new_n930), .ZN(G54));
  INV_X1    g745(.A(new_n527), .ZN(new_n932));
  NAND2_X1  g746(.A1(KEYINPUT58), .A2(G475), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n932), .B1(new_n914), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(new_n909), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n914), .A2(new_n932), .A3(new_n933), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n936), .A2(new_n937), .ZN(G60));
  NAND2_X1  g752(.A1(G478), .A2(G902), .ZN(new_n939));
  XOR2_X1   g753(.A(new_n939), .B(KEYINPUT59), .Z(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n885), .B2(new_n898), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n640), .A2(new_n641), .ZN(new_n942));
  INV_X1    g756(.A(new_n942), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n910), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n942), .A2(new_n940), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n925), .B2(new_n926), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g762(.A(KEYINPUT121), .B(new_n945), .C1(new_n925), .C2(new_n926), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n944), .B1(new_n948), .B2(new_n949), .ZN(G63));
  NOR2_X1   g764(.A1(new_n913), .A2(new_n884), .ZN(new_n951));
  NAND2_X1  g765(.A1(G217), .A2(G902), .ZN(new_n952));
  XOR2_X1   g766(.A(new_n952), .B(KEYINPUT122), .Z(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n249), .B1(new_n951), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n954), .B1(new_n893), .B2(new_n897), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n671), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n955), .A2(new_n957), .A3(new_n910), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n955), .A2(new_n957), .A3(KEYINPUT61), .A4(new_n910), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n960), .A2(new_n961), .ZN(G66));
  OAI21_X1  g776(.A(G953), .B1(new_n537), .B2(new_n586), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n892), .A2(KEYINPUT123), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT123), .ZN(new_n965));
  NAND4_X1  g779(.A1(new_n866), .A2(new_n878), .A3(new_n965), .A4(new_n881), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n233), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n963), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n917), .B1(G898), .B2(new_n233), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n969), .B(new_n970), .ZN(G69));
  OAI21_X1  g785(.A(new_n359), .B1(new_n343), .B2(new_n360), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(new_n517), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n888), .A2(new_n719), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n888), .A2(KEYINPUT62), .A3(new_n719), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OR4_X1    g792(.A1(new_n759), .A2(new_n706), .A3(new_n831), .A4(new_n872), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n798), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n978), .A2(new_n808), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n973), .B1(new_n981), .B2(new_n233), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n982), .A2(KEYINPUT124), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n783), .B1(new_n759), .B2(new_n856), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n985), .A2(new_n797), .A3(new_n406), .A4(new_n705), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n986), .A2(new_n767), .A3(new_n769), .A4(new_n888), .ZN(new_n987));
  NOR3_X1   g801(.A1(new_n829), .A2(new_n802), .A3(new_n806), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n233), .ZN(new_n990));
  OAI211_X1 g804(.A(new_n990), .B(new_n973), .C1(new_n688), .C2(new_n233), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n983), .A2(new_n984), .A3(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n233), .B1(G227), .B2(G900), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n993), .ZN(new_n995));
  NAND4_X1  g809(.A1(new_n983), .A2(new_n995), .A3(new_n984), .A4(new_n991), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n994), .A2(new_n996), .ZN(G72));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n998));
  XNOR2_X1  g812(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n999));
  NOR2_X1   g813(.A1(new_n253), .A2(new_n242), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n999), .B(new_n1000), .Z(new_n1001));
  INV_X1    g815(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(new_n981), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n967), .ZN(new_n1004));
  OAI21_X1  g818(.A(new_n998), .B1(new_n1004), .B2(new_n708), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n981), .B1(new_n964), .B2(new_n966), .ZN(new_n1006));
  OAI211_X1 g820(.A(KEYINPUT126), .B(new_n709), .C1(new_n1006), .C2(new_n1002), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  AOI21_X1  g822(.A(new_n1002), .B1(new_n967), .B2(new_n989), .ZN(new_n1009));
  NAND3_X1  g823(.A1(new_n361), .A2(new_n335), .A3(new_n363), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n935), .B1(new_n1009), .B2(new_n1010), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT127), .ZN(new_n1012));
  OR2_X1    g826(.A1(new_n883), .A2(new_n884), .ZN(new_n1013));
  AND3_X1   g827(.A1(new_n708), .A2(new_n1001), .A3(new_n1010), .ZN(new_n1014));
  AOI22_X1  g828(.A1(new_n1011), .A2(new_n1012), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI211_X1 g829(.A(KEYINPUT127), .B(new_n935), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1008), .A2(new_n1015), .A3(new_n1016), .ZN(G57));
endmodule


