

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772;

  NOR2_X1 U377 ( .A1(n445), .A2(n354), .ZN(n444) );
  AND2_X1 U378 ( .A1(n575), .A2(n587), .ZN(n353) );
  AND2_X1 U379 ( .A1(n441), .A2(n596), .ZN(n354) );
  NOR2_X1 U380 ( .A1(n587), .A2(n575), .ZN(n725) );
  NAND2_X2 U381 ( .A1(n383), .A2(n370), .ZN(n461) );
  NAND2_X2 U382 ( .A1(n609), .A2(n490), .ZN(n610) );
  NOR2_X2 U383 ( .A1(G902), .A2(n730), .ZN(n518) );
  XNOR2_X2 U384 ( .A(G146), .B(G125), .ZN(n540) );
  XNOR2_X2 U385 ( .A(n601), .B(n410), .ZN(n569) );
  XNOR2_X2 U386 ( .A(n610), .B(KEYINPUT0), .ZN(n617) );
  XNOR2_X2 U387 ( .A(n389), .B(n492), .ZN(n549) );
  XNOR2_X2 U388 ( .A(n502), .B(n501), .ZN(n591) );
  OR2_X1 U389 ( .A1(n657), .A2(n658), .ZN(n654) );
  INV_X2 U390 ( .A(G953), .ZN(n762) );
  AND2_X1 U391 ( .A1(n461), .A2(n462), .ZN(n393) );
  NOR2_X1 U392 ( .A1(n770), .A2(n626), .ZN(n627) );
  NOR2_X1 U393 ( .A1(n726), .A2(n712), .ZN(n428) );
  INV_X1 U394 ( .A(n617), .ZN(n420) );
  XNOR2_X1 U395 ( .A(n480), .B(n493), .ZN(n546) );
  XNOR2_X1 U396 ( .A(KEYINPUT86), .B(G119), .ZN(n481) );
  INV_X1 U397 ( .A(KEYINPUT22), .ZN(n454) );
  XNOR2_X1 U398 ( .A(n382), .B(n371), .ZN(n381) );
  NOR2_X1 U399 ( .A1(n444), .A2(n468), .ZN(n373) );
  NAND2_X1 U400 ( .A1(n396), .A2(n395), .ZN(n769) );
  AND2_X1 U401 ( .A1(n398), .A2(n397), .ZN(n396) );
  XNOR2_X1 U402 ( .A(n418), .B(n416), .ZN(n770) );
  NAND2_X1 U403 ( .A1(n360), .A2(n435), .ZN(n395) );
  INV_X1 U404 ( .A(n676), .ZN(n355) );
  XNOR2_X1 U405 ( .A(n662), .B(n443), .ZN(n633) );
  AND2_X1 U406 ( .A1(n618), .A2(n457), .ZN(n456) );
  OR2_X1 U407 ( .A1(n591), .A2(n504), .ZN(n506) );
  XNOR2_X1 U408 ( .A(n431), .B(n415), .ZN(n596) );
  XNOR2_X1 U409 ( .A(n533), .B(n534), .ZN(n657) );
  XOR2_X1 U410 ( .A(KEYINPUT13), .B(n567), .Z(n587) );
  NOR2_X1 U411 ( .A1(G902), .A2(n708), .ZN(n502) );
  XNOR2_X1 U412 ( .A(n413), .B(n412), .ZN(n567) );
  XNOR2_X1 U413 ( .A(n752), .B(n547), .ZN(n695) );
  XNOR2_X1 U414 ( .A(n432), .B(n517), .ZN(n730) );
  XNOR2_X1 U415 ( .A(n403), .B(n546), .ZN(n752) );
  XNOR2_X1 U416 ( .A(n545), .B(n544), .ZN(n403) );
  XNOR2_X1 U417 ( .A(n483), .B(n482), .ZN(n545) );
  INV_X1 U418 ( .A(n745), .ZN(n380) );
  XNOR2_X1 U419 ( .A(n484), .B(G104), .ZN(n483) );
  XNOR2_X1 U420 ( .A(n543), .B(KEYINPUT16), .ZN(n544) );
  XNOR2_X1 U421 ( .A(n500), .B(G472), .ZN(n501) );
  XNOR2_X1 U422 ( .A(n388), .B(KEYINPUT64), .ZN(n539) );
  XNOR2_X1 U423 ( .A(n481), .B(KEYINPUT3), .ZN(n480) );
  XOR2_X1 U424 ( .A(KEYINPUT70), .B(G122), .Z(n543) );
  NOR2_X1 U425 ( .A1(n704), .A2(n745), .ZN(n707) );
  NOR2_X1 U426 ( .A1(n740), .A2(n745), .ZN(n408) );
  XNOR2_X1 U427 ( .A(KEYINPUT65), .B(KEYINPUT75), .ZN(n492) );
  NAND2_X1 U428 ( .A1(n596), .A2(n414), .ZN(n628) );
  INV_X1 U429 ( .A(n654), .ZN(n414) );
  INV_X1 U430 ( .A(KEYINPUT77), .ZN(n452) );
  INV_X1 U431 ( .A(KEYINPUT94), .ZN(n427) );
  XNOR2_X1 U432 ( .A(KEYINPUT98), .B(n576), .ZN(n676) );
  NAND2_X1 U433 ( .A1(n505), .A2(n507), .ZN(n479) );
  XNOR2_X1 U434 ( .A(n529), .B(n409), .ZN(n535) );
  XNOR2_X1 U435 ( .A(n530), .B(KEYINPUT90), .ZN(n409) );
  XOR2_X1 U436 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n530) );
  XNOR2_X1 U437 ( .A(n539), .B(G137), .ZN(n387) );
  XNOR2_X1 U438 ( .A(n464), .B(n463), .ZN(n547) );
  XNOR2_X1 U439 ( .A(n539), .B(n361), .ZN(n463) );
  NOR2_X1 U440 ( .A1(n373), .A2(n433), .ZN(n372) );
  NOR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n503) );
  XNOR2_X1 U442 ( .A(n560), .B(n449), .ZN(n756) );
  INV_X1 U443 ( .A(n561), .ZN(n449) );
  AND2_X1 U444 ( .A1(n462), .A2(G210), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n613), .B(KEYINPUT68), .ZN(n614) );
  NAND2_X1 U446 ( .A1(n633), .A2(n402), .ZN(n593) );
  AND2_X1 U447 ( .A1(n353), .A2(n442), .ZN(n402) );
  INV_X1 U448 ( .A(n592), .ZN(n442) );
  INV_X1 U449 ( .A(KEYINPUT1), .ZN(n415) );
  INV_X1 U450 ( .A(n633), .ZN(n620) );
  XNOR2_X1 U451 ( .A(n528), .B(n527), .ZN(n743) );
  XNOR2_X1 U452 ( .A(n756), .B(n446), .ZN(n737) );
  XNOR2_X1 U453 ( .A(n448), .B(n447), .ZN(n446) );
  XNOR2_X1 U454 ( .A(n563), .B(n566), .ZN(n447) );
  XNOR2_X1 U455 ( .A(n564), .B(n364), .ZN(n448) );
  AND2_X1 U456 ( .A1(n462), .A2(G475), .ZN(n385) );
  NOR2_X1 U457 ( .A1(G952), .A2(n762), .ZN(n745) );
  NAND2_X1 U458 ( .A1(n589), .A2(n359), .ZN(n445) );
  AND2_X1 U459 ( .A1(n421), .A2(n450), .ZN(n589) );
  INV_X1 U460 ( .A(KEYINPUT4), .ZN(n388) );
  INV_X1 U461 ( .A(KEYINPUT38), .ZN(n410) );
  XNOR2_X1 U462 ( .A(G101), .B(G131), .ZN(n494) );
  XOR2_X1 U463 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n495) );
  XNOR2_X1 U464 ( .A(n425), .B(n424), .ZN(n488) );
  INV_X1 U465 ( .A(KEYINPUT99), .ZN(n424) );
  NAND2_X1 U466 ( .A1(n426), .A2(n355), .ZN(n425) );
  INV_X1 U467 ( .A(G134), .ZN(n390) );
  XNOR2_X1 U468 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n519) );
  NOR2_X1 U469 ( .A1(G953), .A2(G237), .ZN(n565) );
  XOR2_X1 U470 ( .A(G131), .B(G140), .Z(n561) );
  XNOR2_X1 U471 ( .A(n698), .B(n460), .ZN(n458) );
  INV_X1 U472 ( .A(KEYINPUT78), .ZN(n460) );
  INV_X1 U473 ( .A(n585), .ZN(n400) );
  INV_X1 U474 ( .A(n658), .ZN(n457) );
  NOR2_X1 U475 ( .A1(n608), .A2(n514), .ZN(n571) );
  NAND2_X1 U476 ( .A1(n479), .A2(n478), .ZN(n477) );
  NAND2_X1 U477 ( .A1(KEYINPUT106), .A2(KEYINPUT30), .ZN(n478) );
  NAND2_X1 U478 ( .A1(n476), .A2(n475), .ZN(n474) );
  NAND2_X1 U479 ( .A1(n505), .A2(KEYINPUT30), .ZN(n476) );
  NAND2_X1 U480 ( .A1(KEYINPUT106), .A2(n507), .ZN(n475) );
  XNOR2_X1 U481 ( .A(n401), .B(n559), .ZN(n586) );
  NOR2_X1 U482 ( .A1(n741), .A2(G902), .ZN(n401) );
  XNOR2_X1 U483 ( .A(G107), .B(G110), .ZN(n482) );
  XNOR2_X1 U484 ( .A(G119), .B(G137), .ZN(n522) );
  XNOR2_X1 U485 ( .A(n540), .B(KEYINPUT10), .ZN(n560) );
  XNOR2_X1 U486 ( .A(G140), .B(KEYINPUT89), .ZN(n524) );
  XNOR2_X1 U487 ( .A(G116), .B(G107), .ZN(n550) );
  XOR2_X1 U488 ( .A(KEYINPUT96), .B(G122), .Z(n551) );
  NAND2_X1 U489 ( .A1(n400), .A2(n436), .ZN(n435) );
  INV_X1 U490 ( .A(G475), .ZN(n412) );
  NOR2_X1 U491 ( .A1(n737), .A2(G902), .ZN(n413) );
  XNOR2_X1 U492 ( .A(n532), .B(n531), .ZN(n533) );
  INV_X1 U493 ( .A(KEYINPUT25), .ZN(n531) );
  INV_X1 U494 ( .A(KEYINPUT6), .ZN(n443) );
  NAND2_X1 U495 ( .A1(n384), .A2(n461), .ZN(n382) );
  AND2_X1 U496 ( .A1(n462), .A2(G472), .ZN(n384) );
  XNOR2_X1 U497 ( .A(n697), .B(n696), .ZN(n703) );
  XNOR2_X1 U498 ( .A(n599), .B(n411), .ZN(n602) );
  XNOR2_X1 U499 ( .A(n600), .B(KEYINPUT43), .ZN(n411) );
  XNOR2_X1 U500 ( .A(n417), .B(KEYINPUT35), .ZN(n416) );
  NAND2_X1 U501 ( .A1(n356), .A2(n394), .ZN(n418) );
  INV_X1 U502 ( .A(KEYINPUT73), .ZN(n417) );
  NAND2_X1 U503 ( .A1(n393), .A2(G217), .ZN(n742) );
  XNOR2_X1 U504 ( .A(n741), .B(KEYINPUT124), .ZN(n486) );
  XNOR2_X1 U505 ( .A(n737), .B(n736), .ZN(n738) );
  AND2_X1 U506 ( .A1(n465), .A2(n365), .ZN(n356) );
  AND2_X1 U507 ( .A1(n437), .A2(n353), .ZN(n357) );
  AND2_X1 U508 ( .A1(n357), .A2(n568), .ZN(n358) );
  AND2_X1 U509 ( .A1(n584), .A2(n583), .ZN(n359) );
  AND2_X1 U510 ( .A1(n438), .A2(n358), .ZN(n360) );
  XOR2_X1 U511 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n361) );
  XOR2_X1 U512 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n362) );
  AND2_X1 U513 ( .A1(G210), .A2(n548), .ZN(n363) );
  XNOR2_X1 U514 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n364) );
  AND2_X1 U515 ( .A1(n466), .A2(n616), .ZN(n365) );
  AND2_X1 U516 ( .A1(n436), .A2(n440), .ZN(n366) );
  AND2_X1 U517 ( .A1(n438), .A2(n437), .ZN(n367) );
  XOR2_X1 U518 ( .A(n590), .B(KEYINPUT36), .Z(n368) );
  XOR2_X1 U519 ( .A(KEYINPUT107), .B(KEYINPUT28), .Z(n369) );
  INV_X1 U520 ( .A(n568), .ZN(n440) );
  XNOR2_X1 U521 ( .A(KEYINPUT66), .B(n701), .ZN(n370) );
  XOR2_X1 U522 ( .A(n709), .B(KEYINPUT112), .Z(n371) );
  XNOR2_X1 U523 ( .A(G902), .B(KEYINPUT15), .ZN(n700) );
  INV_X1 U524 ( .A(n700), .ZN(n419) );
  NAND2_X1 U525 ( .A1(n374), .A2(n372), .ZN(n603) );
  NAND2_X1 U526 ( .A1(n377), .A2(n375), .ZN(n374) );
  NAND2_X1 U527 ( .A1(n434), .A2(n376), .ZN(n375) );
  NAND2_X1 U528 ( .A1(n444), .A2(n468), .ZN(n376) );
  NAND2_X1 U529 ( .A1(n378), .A2(n468), .ZN(n377) );
  INV_X1 U530 ( .A(n434), .ZN(n378) );
  XNOR2_X1 U531 ( .A(n379), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U532 ( .A1(n381), .A2(n380), .ZN(n379) );
  XNOR2_X1 U533 ( .A(n491), .B(n390), .ZN(n389) );
  XNOR2_X2 U534 ( .A(G128), .B(G143), .ZN(n491) );
  NAND2_X1 U535 ( .A1(n459), .A2(n458), .ZN(n383) );
  NAND2_X1 U536 ( .A1(n461), .A2(n385), .ZN(n739) );
  NAND2_X1 U537 ( .A1(n461), .A2(n386), .ZN(n405) );
  XNOR2_X2 U538 ( .A(n549), .B(n387), .ZN(n757) );
  INV_X1 U539 ( .A(n491), .ZN(n391) );
  XNOR2_X1 U540 ( .A(n428), .B(n427), .ZN(n426) );
  NAND2_X1 U541 ( .A1(n617), .A2(KEYINPUT34), .ZN(n466) );
  OR2_X1 U542 ( .A1(n617), .A2(KEYINPUT34), .ZN(n467) );
  XNOR2_X1 U543 ( .A(n391), .B(n492), .ZN(n392) );
  OR2_X1 U544 ( .A1(n682), .A2(n467), .ZN(n394) );
  XNOR2_X2 U545 ( .A(n615), .B(n614), .ZN(n682) );
  NAND2_X1 U546 ( .A1(n438), .A2(n357), .ZN(n399) );
  NAND2_X1 U547 ( .A1(n400), .A2(n366), .ZN(n397) );
  NAND2_X1 U548 ( .A1(n399), .A2(n440), .ZN(n398) );
  NAND2_X1 U549 ( .A1(n355), .A2(n721), .ZN(n423) );
  XNOR2_X1 U550 ( .A(n405), .B(n703), .ZN(n704) );
  XNOR2_X1 U551 ( .A(n594), .B(n579), .ZN(n605) );
  NOR2_X1 U552 ( .A1(n632), .A2(n633), .ZN(n634) );
  XNOR2_X1 U553 ( .A(n404), .B(KEYINPUT46), .ZN(n434) );
  NAND2_X1 U554 ( .A1(n585), .A2(n439), .ZN(n438) );
  NOR2_X1 U555 ( .A1(n537), .A2(n571), .ZN(n406) );
  NOR2_X2 U556 ( .A1(n769), .A2(n771), .ZN(n404) );
  NAND2_X1 U557 ( .A1(n470), .A2(n406), .ZN(n538) );
  BUF_X1 U558 ( .A(n431), .Z(n407) );
  XNOR2_X1 U559 ( .A(n408), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U560 ( .A(n455), .B(n454), .ZN(n623) );
  NOR2_X2 U561 ( .A1(n431), .A2(n654), .ZN(n630) );
  XOR2_X1 U562 ( .A(KEYINPUT42), .B(n574), .Z(n771) );
  NAND2_X1 U563 ( .A1(n746), .A2(n419), .ZN(n698) );
  XNOR2_X2 U564 ( .A(n638), .B(KEYINPUT45), .ZN(n746) );
  NAND2_X1 U565 ( .A1(n420), .A2(n667), .ZN(n629) );
  NAND2_X1 U566 ( .A1(n420), .A2(n456), .ZN(n455) );
  NAND2_X1 U567 ( .A1(n420), .A2(n630), .ZN(n631) );
  NAND2_X1 U568 ( .A1(n422), .A2(n451), .ZN(n421) );
  NAND2_X1 U569 ( .A1(n423), .A2(n452), .ZN(n422) );
  INV_X1 U570 ( .A(n580), .ZN(n577) );
  NAND2_X1 U571 ( .A1(n430), .A2(n429), .ZN(n580) );
  INV_X1 U572 ( .A(n407), .ZN(n429) );
  XNOR2_X1 U573 ( .A(n573), .B(n369), .ZN(n430) );
  XNOR2_X2 U574 ( .A(n518), .B(G469), .ZN(n431) );
  XNOR2_X1 U575 ( .A(n392), .B(n542), .ZN(n464) );
  XNOR2_X1 U576 ( .A(n432), .B(n499), .ZN(n708) );
  XNOR2_X2 U577 ( .A(n757), .B(G146), .ZN(n432) );
  INV_X1 U578 ( .A(n729), .ZN(n433) );
  NAND2_X1 U579 ( .A1(n367), .A2(n435), .ZN(n639) );
  NOR2_X1 U580 ( .A1(n569), .A2(n439), .ZN(n436) );
  NAND2_X1 U581 ( .A1(n569), .A2(n439), .ZN(n437) );
  INV_X1 U582 ( .A(KEYINPUT39), .ZN(n439) );
  XNOR2_X1 U583 ( .A(n628), .B(n611), .ZN(n612) );
  XNOR2_X2 U584 ( .A(n538), .B(KEYINPUT72), .ZN(n585) );
  XNOR2_X1 U585 ( .A(n603), .B(KEYINPUT80), .ZN(n646) );
  NOR2_X1 U586 ( .A1(n646), .A2(n645), .ZN(n647) );
  INV_X1 U587 ( .A(n506), .ZN(n473) );
  NAND2_X1 U588 ( .A1(n473), .A2(n477), .ZN(n472) );
  XNOR2_X1 U589 ( .A(n595), .B(n368), .ZN(n441) );
  INV_X1 U590 ( .A(n720), .ZN(n450) );
  INV_X1 U591 ( .A(KEYINPUT47), .ZN(n451) );
  NAND2_X1 U592 ( .A1(n578), .A2(n672), .ZN(n594) );
  XNOR2_X2 U593 ( .A(n453), .B(n363), .ZN(n578) );
  NAND2_X1 U594 ( .A1(n695), .A2(n700), .ZN(n453) );
  NAND2_X1 U595 ( .A1(n624), .A2(n623), .ZN(n625) );
  INV_X1 U596 ( .A(n699), .ZN(n459) );
  INV_X1 U597 ( .A(n702), .ZN(n462) );
  XNOR2_X1 U598 ( .A(n647), .B(KEYINPUT79), .ZN(n699) );
  NAND2_X1 U599 ( .A1(n682), .A2(KEYINPUT34), .ZN(n465) );
  XNOR2_X2 U600 ( .A(n625), .B(KEYINPUT32), .ZN(n767) );
  INV_X1 U601 ( .A(KEYINPUT48), .ZN(n468) );
  NAND2_X1 U602 ( .A1(n669), .A2(n577), .ZN(n574) );
  XNOR2_X2 U603 ( .A(n469), .B(n570), .ZN(n669) );
  NOR2_X2 U604 ( .A1(n677), .A2(n675), .ZN(n469) );
  NAND2_X1 U605 ( .A1(n673), .A2(n672), .ZN(n677) );
  NAND2_X1 U606 ( .A1(n472), .A2(n471), .ZN(n470) );
  NAND2_X1 U607 ( .A1(n506), .A2(n474), .ZN(n471) );
  XNOR2_X2 U608 ( .A(G101), .B(KEYINPUT85), .ZN(n484) );
  NOR2_X1 U609 ( .A1(n485), .A2(n745), .ZN(G63) );
  XNOR2_X1 U610 ( .A(n487), .B(n486), .ZN(n485) );
  NAND2_X1 U611 ( .A1(n393), .A2(G478), .ZN(n487) );
  AND2_X1 U612 ( .A1(n710), .A2(n488), .ZN(n489) );
  OR2_X1 U613 ( .A1(n608), .A2(n607), .ZN(n490) );
  XNOR2_X1 U614 ( .A(n541), .B(n540), .ZN(n542) );
  INV_X1 U615 ( .A(KEYINPUT100), .ZN(n611) );
  INV_X1 U616 ( .A(KEYINPUT19), .ZN(n579) );
  INV_X1 U617 ( .A(KEYINPUT59), .ZN(n736) );
  XNOR2_X1 U618 ( .A(n521), .B(n560), .ZN(n528) );
  XNOR2_X1 U619 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n568) );
  XNOR2_X1 U620 ( .A(n694), .B(n693), .ZN(G75) );
  XNOR2_X1 U621 ( .A(G116), .B(G113), .ZN(n493) );
  XNOR2_X1 U622 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U623 ( .A(n546), .B(n496), .Z(n498) );
  NAND2_X1 U624 ( .A1(n565), .A2(G210), .ZN(n497) );
  XNOR2_X1 U625 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U626 ( .A(KEYINPUT69), .B(KEYINPUT93), .ZN(n500) );
  XNOR2_X1 U627 ( .A(n503), .B(KEYINPUT71), .ZN(n548) );
  NAND2_X1 U628 ( .A1(G214), .A2(n548), .ZN(n672) );
  INV_X1 U629 ( .A(n672), .ZN(n504) );
  INV_X1 U630 ( .A(KEYINPUT106), .ZN(n505) );
  INV_X1 U631 ( .A(KEYINPUT30), .ZN(n507) );
  NAND2_X1 U632 ( .A1(G234), .A2(G237), .ZN(n508) );
  XNOR2_X1 U633 ( .A(n508), .B(KEYINPUT14), .ZN(n510) );
  NAND2_X1 U634 ( .A1(n510), .A2(G952), .ZN(n509) );
  XOR2_X1 U635 ( .A(KEYINPUT87), .B(n509), .Z(n688) );
  NOR2_X1 U636 ( .A1(G953), .A2(n688), .ZN(n608) );
  NAND2_X1 U637 ( .A1(G902), .A2(n510), .ZN(n511) );
  XOR2_X1 U638 ( .A(KEYINPUT88), .B(n511), .Z(n512) );
  NAND2_X1 U639 ( .A1(G953), .A2(n512), .ZN(n606) );
  NOR2_X1 U640 ( .A1(G900), .A2(n606), .ZN(n513) );
  XOR2_X1 U641 ( .A(KEYINPUT101), .B(n513), .Z(n514) );
  XNOR2_X1 U642 ( .A(n545), .B(n561), .ZN(n516) );
  AND2_X1 U643 ( .A1(G227), .A2(n762), .ZN(n515) );
  XNOR2_X1 U644 ( .A(n516), .B(n515), .ZN(n517) );
  NAND2_X1 U645 ( .A1(n762), .A2(G234), .ZN(n520) );
  XNOR2_X1 U646 ( .A(n520), .B(n519), .ZN(n554) );
  NAND2_X1 U647 ( .A1(G221), .A2(n554), .ZN(n521) );
  XOR2_X1 U648 ( .A(G110), .B(G128), .Z(n523) );
  XNOR2_X1 U649 ( .A(n523), .B(n522), .ZN(n526) );
  XNOR2_X1 U650 ( .A(n362), .B(n524), .ZN(n525) );
  XOR2_X1 U651 ( .A(n526), .B(n525), .Z(n527) );
  NOR2_X1 U652 ( .A1(G902), .A2(n743), .ZN(n534) );
  NAND2_X1 U653 ( .A1(G234), .A2(n700), .ZN(n529) );
  NAND2_X1 U654 ( .A1(G217), .A2(n535), .ZN(n532) );
  NAND2_X1 U655 ( .A1(G221), .A2(n535), .ZN(n536) );
  XNOR2_X1 U656 ( .A(KEYINPUT21), .B(n536), .ZN(n658) );
  XNOR2_X1 U657 ( .A(n630), .B(KEYINPUT105), .ZN(n537) );
  NAND2_X1 U658 ( .A1(G224), .A2(n762), .ZN(n541) );
  INV_X1 U659 ( .A(n578), .ZN(n601) );
  XNOR2_X1 U660 ( .A(KEYINPUT97), .B(G478), .ZN(n559) );
  INV_X1 U661 ( .A(n549), .ZN(n553) );
  XNOR2_X1 U662 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U663 ( .A(n553), .B(n552), .ZN(n558) );
  XOR2_X1 U664 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n556) );
  NAND2_X1 U665 ( .A1(G217), .A2(n554), .ZN(n555) );
  XNOR2_X1 U666 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U667 ( .A(n558), .B(n557), .ZN(n741) );
  INV_X1 U668 ( .A(n586), .ZN(n575) );
  XNOR2_X1 U669 ( .A(G113), .B(G104), .ZN(n562) );
  XNOR2_X1 U670 ( .A(n562), .B(KEYINPUT95), .ZN(n564) );
  XNOR2_X1 U671 ( .A(G143), .B(G122), .ZN(n563) );
  NAND2_X1 U672 ( .A1(G214), .A2(n565), .ZN(n566) );
  INV_X1 U673 ( .A(n569), .ZN(n673) );
  NOR2_X1 U674 ( .A1(n587), .A2(n586), .ZN(n618) );
  INV_X1 U675 ( .A(n618), .ZN(n675) );
  XNOR2_X1 U676 ( .A(KEYINPUT41), .B(KEYINPUT109), .ZN(n570) );
  NOR2_X1 U677 ( .A1(n571), .A2(n658), .ZN(n572) );
  NAND2_X1 U678 ( .A1(n657), .A2(n572), .ZN(n592) );
  NOR2_X1 U679 ( .A1(n592), .A2(n591), .ZN(n573) );
  NOR2_X1 U680 ( .A1(n353), .A2(n725), .ZN(n576) );
  NAND2_X1 U681 ( .A1(n355), .A2(KEYINPUT77), .ZN(n584) );
  NOR2_X1 U682 ( .A1(n580), .A2(n605), .ZN(n721) );
  OR2_X1 U683 ( .A1(n355), .A2(KEYINPUT77), .ZN(n581) );
  NAND2_X1 U684 ( .A1(n721), .A2(n581), .ZN(n582) );
  NAND2_X1 U685 ( .A1(KEYINPUT47), .A2(n582), .ZN(n583) );
  NAND2_X1 U686 ( .A1(n587), .A2(n586), .ZN(n604) );
  OR2_X1 U687 ( .A1(n601), .A2(n604), .ZN(n588) );
  NOR2_X1 U688 ( .A1(n585), .A2(n588), .ZN(n720) );
  INV_X1 U689 ( .A(n596), .ZN(n655) );
  XNOR2_X1 U690 ( .A(KEYINPUT83), .B(KEYINPUT110), .ZN(n590) );
  INV_X1 U691 ( .A(n591), .ZN(n662) );
  XNOR2_X1 U692 ( .A(KEYINPUT102), .B(n593), .ZN(n597) );
  NOR2_X1 U693 ( .A1(n594), .A2(n597), .ZN(n595) );
  XOR2_X1 U694 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n600) );
  NOR2_X1 U695 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U696 ( .A1(n598), .A2(n672), .ZN(n599) );
  NAND2_X1 U697 ( .A1(n602), .A2(n601), .ZN(n729) );
  INV_X1 U698 ( .A(n604), .ZN(n616) );
  INV_X1 U699 ( .A(n605), .ZN(n609) );
  NOR2_X1 U700 ( .A1(G898), .A2(n606), .ZN(n607) );
  NAND2_X1 U701 ( .A1(n612), .A2(n633), .ZN(n615) );
  XOR2_X1 U702 ( .A(KEYINPUT33), .B(KEYINPUT84), .Z(n613) );
  NAND2_X1 U703 ( .A1(n655), .A2(n623), .ZN(n632) );
  NOR2_X1 U704 ( .A1(n662), .A2(n632), .ZN(n619) );
  NAND2_X1 U705 ( .A1(n619), .A2(n657), .ZN(n716) );
  NAND2_X1 U706 ( .A1(n657), .A2(n620), .ZN(n621) );
  NOR2_X1 U707 ( .A1(n655), .A2(n621), .ZN(n622) );
  XNOR2_X1 U708 ( .A(KEYINPUT74), .B(n622), .ZN(n624) );
  NAND2_X1 U709 ( .A1(n716), .A2(n767), .ZN(n626) );
  XNOR2_X1 U710 ( .A(n627), .B(KEYINPUT44), .ZN(n637) );
  NOR2_X1 U711 ( .A1(n591), .A2(n628), .ZN(n667) );
  XNOR2_X1 U712 ( .A(n629), .B(KEYINPUT31), .ZN(n726) );
  NOR2_X1 U713 ( .A1(n662), .A2(n631), .ZN(n712) );
  XNOR2_X1 U714 ( .A(n634), .B(KEYINPUT82), .ZN(n636) );
  INV_X1 U715 ( .A(n657), .ZN(n635) );
  NAND2_X1 U716 ( .A1(n636), .A2(n635), .ZN(n710) );
  NAND2_X1 U717 ( .A1(n637), .A2(n489), .ZN(n638) );
  INV_X1 U718 ( .A(n725), .ZN(n640) );
  NOR2_X1 U719 ( .A1(n640), .A2(n639), .ZN(n641) );
  XNOR2_X1 U720 ( .A(n641), .B(KEYINPUT111), .ZN(n766) );
  NAND2_X1 U721 ( .A1(KEYINPUT2), .A2(n766), .ZN(n642) );
  XOR2_X1 U722 ( .A(KEYINPUT76), .B(n642), .Z(n643) );
  NAND2_X1 U723 ( .A1(n746), .A2(n643), .ZN(n644) );
  NOR2_X1 U724 ( .A1(n646), .A2(n644), .ZN(n702) );
  INV_X1 U725 ( .A(n766), .ZN(n645) );
  BUF_X1 U726 ( .A(n699), .Z(n761) );
  INV_X1 U727 ( .A(n746), .ZN(n648) );
  NOR2_X1 U728 ( .A1(n761), .A2(n648), .ZN(n649) );
  NOR2_X1 U729 ( .A1(KEYINPUT2), .A2(n649), .ZN(n650) );
  NOR2_X1 U730 ( .A1(n702), .A2(n650), .ZN(n653) );
  INV_X1 U731 ( .A(n669), .ZN(n651) );
  NOR2_X1 U732 ( .A1(n682), .A2(n651), .ZN(n652) );
  NOR2_X1 U733 ( .A1(n653), .A2(n652), .ZN(n691) );
  NAND2_X1 U734 ( .A1(n655), .A2(n654), .ZN(n656) );
  XOR2_X1 U735 ( .A(KEYINPUT50), .B(n656), .Z(n665) );
  XOR2_X1 U736 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n660) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  XNOR2_X1 U738 ( .A(n660), .B(n659), .ZN(n661) );
  NOR2_X1 U739 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U740 ( .A(KEYINPUT116), .B(n663), .Z(n664) );
  NOR2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U742 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U743 ( .A(KEYINPUT51), .B(n668), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n670), .A2(n669), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n671), .B(KEYINPUT117), .ZN(n684) );
  NOR2_X1 U746 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n680) );
  NOR2_X1 U748 ( .A1(n677), .A2(n676), .ZN(n678) );
  XNOR2_X1 U749 ( .A(n678), .B(KEYINPUT118), .ZN(n679) );
  NOR2_X1 U750 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U751 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U752 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U753 ( .A(n685), .B(KEYINPUT52), .Z(n686) );
  XNOR2_X1 U754 ( .A(KEYINPUT119), .B(n686), .ZN(n687) );
  NOR2_X1 U755 ( .A1(n688), .A2(n687), .ZN(n689) );
  NOR2_X1 U756 ( .A1(G953), .A2(n689), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n694) );
  INV_X1 U758 ( .A(KEYINPUT120), .ZN(n692) );
  XNOR2_X1 U759 ( .A(n692), .B(KEYINPUT53), .ZN(n693) );
  XOR2_X1 U760 ( .A(KEYINPUT121), .B(KEYINPUT54), .Z(n697) );
  XNOR2_X1 U761 ( .A(n695), .B(KEYINPUT55), .ZN(n696) );
  NAND2_X1 U762 ( .A1(n419), .A2(KEYINPUT2), .ZN(n701) );
  XOR2_X1 U763 ( .A(KEYINPUT81), .B(KEYINPUT122), .Z(n705) );
  XNOR2_X1 U764 ( .A(n705), .B(KEYINPUT56), .ZN(n706) );
  XNOR2_X1 U765 ( .A(n707), .B(n706), .ZN(G51) );
  XNOR2_X1 U766 ( .A(n708), .B(KEYINPUT62), .ZN(n709) );
  XNOR2_X1 U767 ( .A(G101), .B(n710), .ZN(G3) );
  NAND2_X1 U768 ( .A1(n712), .A2(n353), .ZN(n711) );
  XNOR2_X1 U769 ( .A(n711), .B(G104), .ZN(G6) );
  XOR2_X1 U770 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n714) );
  NAND2_X1 U771 ( .A1(n712), .A2(n725), .ZN(n713) );
  XNOR2_X1 U772 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U773 ( .A(G107), .B(n715), .ZN(G9) );
  XNOR2_X1 U774 ( .A(G110), .B(n716), .ZN(G12) );
  XOR2_X1 U775 ( .A(KEYINPUT113), .B(KEYINPUT29), .Z(n718) );
  NAND2_X1 U776 ( .A1(n721), .A2(n725), .ZN(n717) );
  XNOR2_X1 U777 ( .A(n718), .B(n717), .ZN(n719) );
  XOR2_X1 U778 ( .A(G128), .B(n719), .Z(G30) );
  XOR2_X1 U779 ( .A(G143), .B(n720), .Z(G45) );
  NAND2_X1 U780 ( .A1(n721), .A2(n353), .ZN(n722) );
  XNOR2_X1 U781 ( .A(n722), .B(KEYINPUT114), .ZN(n723) );
  XNOR2_X1 U782 ( .A(G146), .B(n723), .ZN(G48) );
  NAND2_X1 U783 ( .A1(n726), .A2(n353), .ZN(n724) );
  XNOR2_X1 U784 ( .A(n724), .B(G113), .ZN(G15) );
  NAND2_X1 U785 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U786 ( .A(n727), .B(G116), .ZN(G18) );
  XNOR2_X1 U787 ( .A(G125), .B(n354), .ZN(n728) );
  XNOR2_X1 U788 ( .A(n728), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U789 ( .A(G140), .B(n729), .ZN(G42) );
  XNOR2_X1 U790 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n732) );
  XNOR2_X1 U791 ( .A(n730), .B(KEYINPUT57), .ZN(n731) );
  XNOR2_X1 U792 ( .A(n732), .B(n731), .ZN(n734) );
  NAND2_X1 U793 ( .A1(n393), .A2(G469), .ZN(n733) );
  XNOR2_X1 U794 ( .A(n734), .B(n733), .ZN(n735) );
  NOR2_X1 U795 ( .A1(n745), .A2(n735), .ZN(G54) );
  XNOR2_X1 U796 ( .A(n739), .B(n738), .ZN(n740) );
  XNOR2_X1 U797 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U798 ( .A1(n745), .A2(n744), .ZN(G66) );
  NAND2_X1 U799 ( .A1(n762), .A2(n746), .ZN(n750) );
  NAND2_X1 U800 ( .A1(G953), .A2(G224), .ZN(n747) );
  XNOR2_X1 U801 ( .A(KEYINPUT61), .B(n747), .ZN(n748) );
  NAND2_X1 U802 ( .A1(n748), .A2(G898), .ZN(n749) );
  NAND2_X1 U803 ( .A1(n750), .A2(n749), .ZN(n754) );
  NOR2_X1 U804 ( .A1(G898), .A2(n762), .ZN(n751) );
  NOR2_X1 U805 ( .A1(n752), .A2(n751), .ZN(n753) );
  XNOR2_X1 U806 ( .A(n754), .B(n753), .ZN(n755) );
  XOR2_X1 U807 ( .A(KEYINPUT125), .B(n755), .Z(G69) );
  XOR2_X1 U808 ( .A(n757), .B(n756), .Z(n760) );
  XNOR2_X1 U809 ( .A(G227), .B(n760), .ZN(n758) );
  NAND2_X1 U810 ( .A1(G900), .A2(n758), .ZN(n759) );
  NAND2_X1 U811 ( .A1(n759), .A2(G953), .ZN(n765) );
  XNOR2_X1 U812 ( .A(n761), .B(n760), .ZN(n763) );
  NAND2_X1 U813 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U814 ( .A1(n765), .A2(n764), .ZN(G72) );
  XNOR2_X1 U815 ( .A(G134), .B(n766), .ZN(G36) );
  XNOR2_X1 U816 ( .A(n767), .B(G119), .ZN(n768) );
  XNOR2_X1 U817 ( .A(n768), .B(KEYINPUT126), .ZN(G21) );
  XOR2_X1 U818 ( .A(n769), .B(G131), .Z(G33) );
  XOR2_X1 U819 ( .A(n770), .B(G122), .Z(G24) );
  XNOR2_X1 U820 ( .A(G137), .B(KEYINPUT127), .ZN(n772) );
  XNOR2_X1 U821 ( .A(n772), .B(n771), .ZN(G39) );
endmodule

