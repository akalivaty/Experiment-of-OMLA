//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1 0 1 1 0 1 1 0 0 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 0 1 1 0 0 1 1 0 1 1 1 1 0 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:22 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n605, new_n606, new_n607, new_n608,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n618, new_n619, new_n620, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n627, new_n628, new_n629, new_n630, new_n631,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n887, new_n888, new_n889, new_n890, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951;
  XNOR2_X1  g000(.A(G125), .B(G140), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT76), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n190));
  INV_X1    g004(.A(G146), .ZN(new_n191));
  AND3_X1   g005(.A1(new_n189), .A2(new_n190), .A3(new_n191), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n190), .B1(new_n189), .B2(new_n191), .ZN(new_n193));
  OAI22_X1  g007(.A1(new_n192), .A2(new_n193), .B1(new_n191), .B2(new_n187), .ZN(new_n194));
  INV_X1    g008(.A(G237), .ZN(new_n195));
  INV_X1    g009(.A(G953), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(new_n196), .A3(G214), .ZN(new_n197));
  XNOR2_X1  g011(.A(new_n197), .B(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT18), .A2(G131), .ZN(new_n199));
  XOR2_X1   g013(.A(new_n198), .B(new_n199), .Z(new_n200));
  NAND2_X1  g014(.A1(new_n194), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G125), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n202), .A2(KEYINPUT16), .A3(G140), .ZN(new_n203));
  AOI21_X1  g017(.A(new_n203), .B1(new_n187), .B2(KEYINPUT16), .ZN(new_n204));
  XNOR2_X1  g018(.A(new_n204), .B(new_n191), .ZN(new_n205));
  INV_X1    g019(.A(new_n198), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n206), .A2(KEYINPUT17), .A3(G131), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(G131), .ZN(new_n208));
  INV_X1    g022(.A(G131), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n198), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  OAI211_X1 g025(.A(new_n205), .B(new_n207), .C1(new_n211), .C2(KEYINPUT17), .ZN(new_n212));
  XNOR2_X1  g026(.A(G113), .B(G122), .ZN(new_n213));
  INV_X1    g027(.A(G104), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n213), .B(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(KEYINPUT89), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n201), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  AOI22_X1  g031(.A1(new_n208), .A2(new_n210), .B1(G146), .B2(new_n204), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT19), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n187), .A2(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n220), .B1(new_n189), .B2(new_n219), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n221), .A2(new_n191), .ZN(new_n222));
  AOI22_X1  g036(.A1(new_n194), .A2(new_n200), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n217), .B1(new_n215), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G475), .ZN(new_n225));
  INV_X1    g039(.A(G902), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT20), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  XNOR2_X1  g043(.A(G128), .B(G143), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(KEYINPUT13), .ZN(new_n231));
  INV_X1    g045(.A(G143), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(G128), .ZN(new_n233));
  OAI211_X1 g047(.A(new_n231), .B(G134), .C1(KEYINPUT13), .C2(new_n233), .ZN(new_n234));
  XOR2_X1   g048(.A(G116), .B(G122), .Z(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G107), .ZN(new_n236));
  XNOR2_X1  g050(.A(G116), .B(G122), .ZN(new_n237));
  INV_X1    g051(.A(G107), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(G134), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n234), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n230), .B(new_n241), .ZN(new_n244));
  INV_X1    g058(.A(G116), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT14), .A3(G122), .ZN(new_n246));
  OAI211_X1 g060(.A(G107), .B(new_n246), .C1(new_n235), .C2(KEYINPUT14), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n244), .A2(new_n239), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  XOR2_X1   g063(.A(KEYINPUT9), .B(G234), .Z(new_n250));
  NAND3_X1  g064(.A1(new_n250), .A2(G217), .A3(new_n196), .ZN(new_n251));
  XNOR2_X1  g065(.A(new_n249), .B(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(new_n226), .ZN(new_n253));
  INV_X1    g067(.A(G478), .ZN(new_n254));
  NOR2_X1   g068(.A1(new_n254), .A2(KEYINPUT15), .ZN(new_n255));
  XOR2_X1   g069(.A(new_n253), .B(new_n255), .Z(new_n256));
  INV_X1    g070(.A(new_n217), .ZN(new_n257));
  AOI21_X1  g071(.A(new_n215), .B1(new_n201), .B2(new_n212), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n226), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(G475), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n224), .A2(KEYINPUT20), .A3(new_n225), .A4(new_n226), .ZN(new_n261));
  NAND4_X1  g075(.A1(new_n229), .A2(new_n256), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G952), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n263), .A2(G953), .ZN(new_n264));
  NAND2_X1  g078(.A1(G234), .A2(G237), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  XOR2_X1   g080(.A(KEYINPUT21), .B(G898), .Z(new_n267));
  NAND3_X1  g081(.A1(new_n265), .A2(G902), .A3(G953), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n262), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT90), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n271), .B(new_n272), .ZN(new_n273));
  OAI21_X1  g087(.A(G214), .B1(G237), .B2(G902), .ZN(new_n274));
  XOR2_X1   g088(.A(new_n274), .B(KEYINPUT83), .Z(new_n275));
  OAI21_X1  g089(.A(KEYINPUT3), .B1(new_n214), .B2(G107), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT3), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(new_n238), .A3(G104), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n214), .A2(G107), .ZN(new_n279));
  AND3_X1   g093(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT80), .B(G101), .Z(new_n281));
  NAND2_X1  g095(.A1(new_n238), .A2(G104), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(new_n282), .ZN(new_n283));
  AOI22_X1  g097(.A1(new_n280), .A2(new_n281), .B1(G101), .B2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT67), .B1(new_n245), .B2(G119), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT67), .ZN(new_n286));
  INV_X1    g100(.A(G119), .ZN(new_n287));
  NAND3_X1  g101(.A1(new_n286), .A2(new_n287), .A3(G116), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n245), .A2(G119), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT2), .B(G113), .ZN(new_n291));
  OR2_X1    g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n287), .A3(G116), .ZN(new_n294));
  OAI211_X1 g108(.A(G113), .B(new_n294), .C1(new_n290), .C2(new_n293), .ZN(new_n295));
  NAND3_X1  g109(.A1(new_n284), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n281), .A2(new_n279), .A3(new_n278), .A4(new_n276), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(G101), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n297), .A2(new_n299), .A3(KEYINPUT4), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT4), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n301), .A3(G101), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n290), .A2(new_n291), .ZN(new_n304));
  AND2_X1   g118(.A1(new_n292), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n296), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT84), .ZN(new_n307));
  XOR2_X1   g121(.A(G110), .B(G122), .Z(new_n308));
  AND2_X1   g122(.A1(new_n308), .A2(KEYINPUT85), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT84), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n310), .B(new_n296), .C1(new_n303), .C2(new_n305), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n307), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT6), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OR2_X1    g128(.A1(new_n306), .A2(new_n308), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n307), .A2(new_n311), .A3(KEYINPUT6), .A4(new_n309), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n315), .A3(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n191), .A2(G143), .ZN(new_n318));
  AND3_X1   g132(.A1(new_n232), .A2(KEYINPUT64), .A3(G146), .ZN(new_n319));
  AOI21_X1  g133(.A(KEYINPUT64), .B1(new_n232), .B2(G146), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT0), .A2(G128), .ZN(new_n322));
  OR2_X1    g136(.A1(KEYINPUT0), .A2(G128), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n321), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n232), .A2(G146), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT65), .B1(new_n191), .B2(G143), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT65), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n327), .A2(new_n232), .A3(G146), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n329), .A2(KEYINPUT0), .A3(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n324), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(G125), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT86), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT1), .B1(new_n232), .B2(G146), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n334), .A2(KEYINPUT66), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n318), .A2(new_n336), .A3(KEYINPUT1), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(G128), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G128), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT1), .ZN(new_n340));
  AOI22_X1  g154(.A1(new_n338), .A2(new_n321), .B1(new_n329), .B2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n202), .ZN(new_n342));
  AND3_X1   g156(.A1(new_n332), .A2(new_n333), .A3(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n333), .B1(new_n332), .B2(new_n342), .ZN(new_n344));
  INV_X1    g158(.A(G224), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n345), .A2(G953), .ZN(new_n346));
  INV_X1    g160(.A(new_n346), .ZN(new_n347));
  OR3_X1    g161(.A1(new_n343), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  OAI21_X1  g162(.A(new_n347), .B1(new_n343), .B2(new_n344), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(G902), .B1(new_n317), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n332), .B1(new_n342), .B2(KEYINPUT87), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(KEYINPUT7), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(new_n353), .ZN(new_n355));
  OAI211_X1 g169(.A(new_n332), .B(new_n342), .C1(KEYINPUT87), .C2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n295), .A2(new_n292), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n283), .A2(G101), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n297), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  AND2_X1   g174(.A1(new_n360), .A2(new_n296), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n308), .B(KEYINPUT8), .ZN(new_n362));
  OAI211_X1 g176(.A(new_n354), .B(new_n356), .C1(new_n361), .C2(new_n362), .ZN(new_n363));
  OR2_X1    g177(.A1(new_n363), .A2(KEYINPUT88), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n363), .A2(KEYINPUT88), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n364), .A2(new_n315), .A3(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n351), .A2(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(G210), .B1(G237), .B2(G902), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n351), .A2(new_n368), .A3(new_n366), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n275), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(G221), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n373), .B1(new_n250), .B2(new_n226), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G469), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT1), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n377), .B1(G143), .B2(new_n191), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n339), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n334), .A2(KEYINPUT81), .ZN(new_n381));
  AOI21_X1  g195(.A(new_n329), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n377), .A2(G128), .ZN(new_n383));
  AOI211_X1 g197(.A(new_n383), .B(new_n325), .C1(new_n326), .C2(new_n328), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n284), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT10), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT11), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n388), .B1(new_n241), .B2(G137), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n241), .A2(G137), .ZN(new_n390));
  INV_X1    g204(.A(G137), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(KEYINPUT11), .A3(G134), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n389), .A2(new_n390), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G131), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n389), .A2(new_n392), .A3(new_n209), .A4(new_n390), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n338), .A2(new_n321), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n329), .A2(new_n340), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT10), .A3(new_n284), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n300), .A2(new_n330), .A3(new_n324), .A4(new_n302), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n387), .A2(new_n397), .A3(new_n401), .A4(new_n402), .ZN(new_n403));
  XNOR2_X1  g217(.A(G110), .B(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n196), .A2(G227), .ZN(new_n405));
  XNOR2_X1  g219(.A(new_n404), .B(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n387), .A2(new_n402), .A3(new_n401), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(new_n396), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  INV_X1    g225(.A(KEYINPUT12), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n341), .A2(new_n359), .ZN(new_n413));
  AND3_X1   g227(.A1(new_n413), .A2(new_n385), .A3(KEYINPUT82), .ZN(new_n414));
  OAI21_X1  g228(.A(new_n396), .B1(new_n413), .B2(KEYINPUT82), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n412), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR2_X1   g230(.A1(new_n400), .A2(new_n284), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT82), .ZN(new_n418));
  AOI21_X1  g232(.A(new_n397), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n413), .A2(new_n385), .A3(KEYINPUT82), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n419), .A2(KEYINPUT12), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n416), .A2(new_n421), .ZN(new_n422));
  AND2_X1   g236(.A1(new_n422), .A2(new_n403), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n411), .B1(new_n423), .B2(new_n406), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n376), .B1(new_n424), .B2(new_n226), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n407), .B1(new_n421), .B2(new_n416), .ZN(new_n426));
  AOI21_X1  g240(.A(new_n406), .B1(new_n410), .B2(new_n403), .ZN(new_n427));
  NOR2_X1   g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NOR3_X1   g242(.A1(new_n428), .A2(G469), .A3(G902), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n375), .B1(new_n425), .B2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n273), .A2(new_n372), .A3(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  INV_X1    g247(.A(KEYINPUT68), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n391), .A2(G134), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n241), .A2(G137), .ZN(new_n436));
  OAI21_X1  g250(.A(G131), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n395), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n434), .B1(new_n341), .B2(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n396), .A2(new_n324), .A3(new_n330), .ZN(new_n440));
  AND2_X1   g254(.A1(new_n395), .A2(new_n437), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT64), .ZN(new_n442));
  OAI21_X1  g256(.A(new_n442), .B1(new_n191), .B2(G143), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n232), .A2(KEYINPUT64), .A3(G146), .ZN(new_n444));
  AOI21_X1  g258(.A(new_n325), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n339), .B1(new_n378), .B2(new_n336), .ZN(new_n446));
  AOI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n335), .ZN(new_n447));
  OAI211_X1 g261(.A(KEYINPUT68), .B(new_n441), .C1(new_n447), .C2(new_n384), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n439), .A2(new_n305), .A3(new_n440), .A4(new_n448), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n439), .A2(new_n440), .A3(new_n448), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(KEYINPUT30), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n441), .B1(new_n447), .B2(new_n384), .ZN(new_n452));
  INV_X1    g266(.A(KEYINPUT30), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n452), .A2(new_n453), .A3(new_n440), .ZN(new_n454));
  INV_X1    g268(.A(new_n454), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n451), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(new_n305), .ZN(new_n457));
  AOI21_X1  g271(.A(KEYINPUT69), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n454), .B1(KEYINPUT30), .B2(new_n450), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT69), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n459), .A2(new_n460), .A3(new_n305), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n449), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n463));
  XNOR2_X1  g277(.A(new_n463), .B(G101), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n195), .A2(new_n196), .A3(G210), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n464), .B(new_n465), .Z(new_n466));
  NAND3_X1  g280(.A1(new_n462), .A2(KEYINPUT73), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT73), .ZN(new_n468));
  INV_X1    g282(.A(new_n449), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n456), .A2(KEYINPUT69), .A3(new_n457), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n460), .B1(new_n459), .B2(new_n305), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n469), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n466), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n468), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n396), .A2(new_n330), .A3(new_n324), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n438), .B1(new_n398), .B2(new_n399), .ZN(new_n476));
  NOR3_X1   g290(.A1(new_n475), .A2(new_n476), .A3(new_n457), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n477), .A2(KEYINPUT28), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n457), .B1(new_n475), .B2(new_n476), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n449), .A2(new_n479), .ZN(new_n480));
  XOR2_X1   g294(.A(KEYINPUT71), .B(KEYINPUT28), .Z(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT72), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n480), .A2(KEYINPUT72), .A3(new_n482), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n478), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT29), .B1(new_n487), .B2(new_n473), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n467), .A2(new_n474), .A3(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n450), .A2(new_n457), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n491), .A2(KEYINPUT74), .A3(new_n449), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT74), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n450), .A2(new_n493), .A3(new_n457), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n492), .A2(KEYINPUT28), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n478), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n495), .A2(KEYINPUT29), .A3(new_n496), .A4(new_n473), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n226), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT75), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n497), .A2(KEYINPUT75), .A3(new_n226), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g316(.A(G472), .B1(new_n490), .B2(new_n502), .ZN(new_n503));
  NOR2_X1   g317(.A1(G472), .A2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n469), .A2(new_n466), .ZN(new_n507));
  OAI211_X1 g321(.A(new_n506), .B(new_n507), .C1(new_n458), .C2(new_n461), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n509));
  INV_X1    g323(.A(new_n507), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n510), .B1(new_n470), .B2(new_n471), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT70), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n511), .A2(new_n512), .A3(new_n506), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n509), .A2(new_n513), .ZN(new_n514));
  OAI21_X1  g328(.A(new_n507), .B1(new_n458), .B2(new_n461), .ZN(new_n515));
  AOI21_X1  g329(.A(KEYINPUT72), .B1(new_n480), .B2(new_n482), .ZN(new_n516));
  AOI211_X1 g330(.A(new_n484), .B(new_n481), .C1(new_n449), .C2(new_n479), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n496), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g332(.A1(new_n515), .A2(KEYINPUT31), .B1(new_n466), .B2(new_n518), .ZN(new_n519));
  AOI211_X1 g333(.A(KEYINPUT32), .B(new_n505), .C1(new_n514), .C2(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(KEYINPUT32), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n508), .A2(KEYINPUT70), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n512), .B1(new_n511), .B2(new_n506), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n519), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(new_n504), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n503), .B1(new_n520), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n192), .A2(new_n193), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n287), .A2(G128), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n339), .A2(G119), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT24), .B(G110), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT23), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n339), .A2(KEYINPUT23), .A3(G119), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(new_n528), .A3(new_n535), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n532), .B1(new_n536), .B2(G110), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n204), .A2(G146), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  OR2_X1    g353(.A1(new_n527), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n536), .A2(G110), .ZN(new_n541));
  NOR2_X1   g355(.A1(new_n530), .A2(new_n531), .ZN(new_n542));
  NOR3_X1   g356(.A1(new_n205), .A2(new_n541), .A3(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT22), .B(G137), .ZN(new_n545));
  XNOR2_X1  g359(.A(new_n545), .B(KEYINPUT78), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n196), .A2(G221), .A3(G234), .ZN(new_n547));
  XNOR2_X1  g361(.A(new_n546), .B(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n540), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n548), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n527), .A2(new_n539), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n550), .B1(new_n551), .B2(new_n543), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n549), .A2(new_n226), .A3(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(G217), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(G234), .B2(new_n226), .ZN(new_n555));
  NOR2_X1   g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(KEYINPUT25), .ZN(new_n557));
  XNOR2_X1  g371(.A(new_n553), .B(new_n557), .ZN(new_n558));
  AOI21_X1  g372(.A(new_n556), .B1(new_n558), .B2(new_n555), .ZN(new_n559));
  AND3_X1   g373(.A1(new_n526), .A2(KEYINPUT79), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(KEYINPUT79), .B1(new_n526), .B2(new_n559), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n433), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  XOR2_X1   g376(.A(new_n562), .B(new_n281), .Z(G3));
  INV_X1    g377(.A(new_n371), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n368), .B1(new_n351), .B2(new_n366), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n269), .B(new_n274), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n251), .A2(KEYINPUT92), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(KEYINPUT33), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n568), .A2(KEYINPUT91), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n252), .A2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT33), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n569), .B1(KEYINPUT91), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n252), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  INV_X1    g389(.A(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n576), .A2(G478), .A3(new_n226), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n253), .A2(new_n254), .ZN(new_n578));
  XNOR2_X1  g392(.A(new_n578), .B(KEYINPUT93), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n229), .A2(new_n260), .A3(new_n261), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  OAI21_X1  g396(.A(KEYINPUT94), .B1(new_n566), .B2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n274), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n584), .B1(new_n370), .B2(new_n371), .ZN(new_n585));
  INV_X1    g399(.A(new_n582), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n585), .A2(new_n586), .A3(new_n587), .A4(new_n269), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI22_X1  g403(.A1(new_n511), .A2(new_n506), .B1(new_n487), .B2(new_n473), .ZN(new_n590));
  AOI21_X1  g404(.A(new_n590), .B1(new_n513), .B2(new_n509), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n591), .A2(new_n505), .ZN(new_n592));
  INV_X1    g406(.A(G472), .ZN(new_n593));
  AOI21_X1  g407(.A(new_n593), .B1(new_n524), .B2(new_n226), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n559), .B(new_n375), .C1(new_n425), .C2(new_n429), .ZN(new_n595));
  NOR3_X1   g409(.A1(new_n592), .A2(new_n594), .A3(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT34), .B(G104), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(KEYINPUT95), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n597), .B(new_n599), .ZN(G6));
  AND3_X1   g414(.A1(new_n229), .A2(new_n260), .A3(new_n261), .ZN(new_n601));
  INV_X1    g415(.A(new_n256), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n566), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT35), .B(G107), .ZN(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(new_n607));
  XNOR2_X1  g421(.A(KEYINPUT96), .B(KEYINPUT97), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(G9));
  OAI21_X1  g423(.A(G472), .B1(new_n591), .B2(G902), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n591), .B2(new_n505), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n558), .A2(new_n555), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n551), .A2(new_n543), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n550), .A2(KEYINPUT36), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n615), .A2(G902), .A3(new_n555), .ZN(new_n616));
  OR2_X1    g430(.A1(new_n612), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n617), .ZN(new_n618));
  NOR3_X1   g432(.A1(new_n432), .A2(new_n611), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(KEYINPUT37), .ZN(new_n620));
  XNOR2_X1  g434(.A(new_n620), .B(G110), .ZN(G12));
  XOR2_X1   g435(.A(new_n266), .B(KEYINPUT98), .Z(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(G900), .B2(new_n268), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n603), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n370), .A2(new_n371), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n627), .A2(new_n274), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n628), .A2(new_n430), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n526), .A2(new_n617), .A3(new_n626), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT99), .B(G128), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G30));
  AND2_X1   g446(.A1(new_n492), .A2(new_n494), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n511), .B1(new_n633), .B2(new_n466), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n634), .A2(G472), .ZN(new_n635));
  NAND2_X1  g449(.A1(G472), .A2(G902), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n635), .A2(KEYINPUT100), .A3(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT100), .ZN(new_n638));
  OAI211_X1 g452(.A(new_n638), .B(G472), .C1(new_n634), .C2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n637), .A2(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n640), .B1(new_n520), .B2(new_n525), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT38), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n627), .B(new_n643), .ZN(new_n644));
  NOR3_X1   g458(.A1(new_n642), .A2(new_n584), .A3(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n581), .A2(new_n602), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g461(.A(new_n624), .B(KEYINPUT39), .Z(new_n648));
  NOR2_X1   g462(.A1(new_n430), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(KEYINPUT40), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n645), .A2(new_n618), .A3(new_n647), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(G143), .ZN(G45));
  NOR2_X1   g466(.A1(new_n582), .A2(new_n625), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n526), .A2(new_n617), .A3(new_n629), .A4(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G146), .ZN(G48));
  INV_X1    g469(.A(KEYINPUT101), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n656), .B1(new_n428), .B2(G902), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n422), .A2(new_n408), .ZN(new_n658));
  INV_X1    g472(.A(new_n427), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n660), .A2(KEYINPUT101), .A3(new_n226), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n657), .A2(new_n661), .A3(G469), .ZN(new_n662));
  NOR2_X1   g476(.A1(new_n428), .A2(G902), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT102), .B1(new_n663), .B2(new_n376), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n657), .A2(new_n661), .A3(KEYINPUT102), .A4(G469), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n374), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  NAND4_X1  g481(.A1(new_n589), .A2(new_n526), .A3(new_n559), .A4(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT41), .B(G113), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n668), .B(new_n669), .ZN(G15));
  NAND4_X1  g484(.A1(new_n526), .A2(new_n604), .A3(new_n559), .A4(new_n667), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G116), .ZN(G18));
  NAND2_X1  g486(.A1(new_n665), .A2(new_n666), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n673), .A2(new_n585), .A3(new_n375), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n526), .A2(new_n674), .A3(new_n273), .A4(new_n617), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G119), .ZN(G21));
  INV_X1    g490(.A(KEYINPUT104), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n504), .B(KEYINPUT103), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n473), .B1(new_n495), .B2(new_n496), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n680), .B1(new_n509), .B2(new_n513), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n515), .A2(KEYINPUT31), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n594), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g498(.A1(new_n684), .A2(new_n559), .A3(new_n269), .A4(new_n647), .ZN(new_n685));
  INV_X1    g499(.A(new_n674), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n677), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  INV_X1    g501(.A(new_n559), .ZN(new_n688));
  NOR4_X1   g502(.A1(new_n594), .A2(new_n683), .A3(new_n688), .A4(new_n646), .ZN(new_n689));
  NAND4_X1  g503(.A1(new_n689), .A2(KEYINPUT104), .A3(new_n269), .A4(new_n674), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G122), .ZN(G24));
  NAND4_X1  g506(.A1(new_n674), .A2(new_n684), .A3(new_n617), .A4(new_n653), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G125), .ZN(G27));
  AND2_X1   g508(.A1(new_n500), .A2(new_n501), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n593), .B1(new_n695), .B2(new_n489), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT32), .B1(new_n591), .B2(new_n505), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n524), .A2(new_n521), .A3(new_n504), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n699), .A2(new_n688), .ZN(new_n700));
  INV_X1    g514(.A(new_n653), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n370), .A2(new_n371), .A3(new_n274), .ZN(new_n702));
  NOR3_X1   g516(.A1(new_n701), .A2(new_n430), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n700), .A2(KEYINPUT42), .A3(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT42), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n701), .A2(new_n702), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n431), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n526), .A2(new_n559), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n705), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n704), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  AOI21_X1  g525(.A(new_n702), .B1(new_n626), .B2(KEYINPUT105), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n626), .A2(KEYINPUT105), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n700), .A2(new_n431), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G134), .ZN(G36));
  NAND2_X1  g529(.A1(new_n601), .A2(new_n580), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT43), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n716), .B(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n611), .A2(new_n718), .A3(new_n617), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT106), .ZN(new_n722));
  INV_X1    g536(.A(new_n702), .ZN(new_n723));
  OAI21_X1  g537(.A(new_n723), .B1(new_n719), .B2(new_n720), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n424), .B(KEYINPUT45), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n726), .A2(G469), .ZN(new_n727));
  NAND2_X1  g541(.A1(G469), .A2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT46), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n429), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n727), .A2(KEYINPUT46), .A3(new_n728), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n375), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n734), .A2(new_n648), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n725), .A2(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G137), .ZN(G39));
  INV_X1    g551(.A(KEYINPUT47), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n734), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n733), .A2(KEYINPUT47), .A3(new_n375), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n741), .A2(new_n699), .A3(new_n688), .A4(new_n706), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G140), .ZN(G42));
  NOR2_X1   g557(.A1(new_n617), .A2(new_n625), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n641), .A2(new_n629), .A3(new_n647), .A4(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n630), .A2(new_n654), .A3(new_n745), .A4(new_n693), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n697), .A2(new_n698), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n618), .B1(new_n749), .B2(new_n503), .ZN(new_n750));
  OAI211_X1 g564(.A(new_n750), .B(new_n629), .C1(new_n626), .C2(new_n653), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n751), .A2(KEYINPUT52), .A3(new_n693), .A4(new_n745), .ZN(new_n752));
  AND3_X1   g566(.A1(new_n748), .A2(new_n752), .A3(KEYINPUT111), .ZN(new_n753));
  AOI21_X1  g567(.A(KEYINPUT111), .B1(new_n748), .B2(new_n752), .ZN(new_n754));
  NOR2_X1   g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  OR3_X1    g569(.A1(new_n432), .A2(new_n611), .A3(new_n618), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n691), .A2(new_n562), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n703), .A2(new_n684), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n702), .A2(new_n262), .A3(new_n625), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n526), .B(new_n431), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  AND2_X1   g575(.A1(new_n759), .A2(new_n760), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n758), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n617), .A2(new_n763), .B1(new_n704), .B2(new_n709), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n586), .A2(KEYINPUT108), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n603), .A2(KEYINPUT109), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT108), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n582), .A2(new_n767), .ZN(new_n768));
  OR3_X1    g582(.A1(new_n581), .A2(KEYINPUT109), .A3(new_n256), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n765), .A2(new_n766), .A3(new_n768), .A4(new_n769), .ZN(new_n770));
  NAND4_X1  g584(.A1(new_n596), .A2(new_n770), .A3(new_n269), .A4(new_n372), .ZN(new_n771));
  AND4_X1   g585(.A1(new_n668), .A2(new_n771), .A3(new_n671), .A4(new_n675), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n757), .A2(new_n764), .A3(new_n714), .A4(new_n772), .ZN(new_n773));
  OAI21_X1  g587(.A(KEYINPUT53), .B1(new_n755), .B2(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT79), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n708), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n526), .A2(KEYINPUT79), .A3(new_n559), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n619), .B1(new_n778), .B2(new_n433), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n772), .A3(new_n691), .A4(new_n714), .ZN(new_n780));
  INV_X1    g594(.A(new_n764), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n748), .A2(new_n752), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n782), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(KEYINPUT54), .B1(new_n774), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT113), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n788), .B(KEYINPUT54), .C1(new_n774), .C2(new_n785), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n787), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT114), .B(KEYINPUT51), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n716), .A2(new_n717), .ZN(new_n792));
  AOI21_X1  g606(.A(KEYINPUT43), .B1(new_n601), .B2(new_n580), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(KEYINPUT115), .B1(new_n794), .B2(new_n623), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT115), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n718), .A2(new_n796), .A3(new_n622), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  AND3_X1   g612(.A1(new_n798), .A2(new_n559), .A3(new_n684), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n644), .A2(new_n584), .A3(new_n667), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(KEYINPUT118), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n799), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n799), .A2(new_n801), .A3(KEYINPUT50), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n798), .A2(new_n667), .A3(new_n723), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n808), .A2(new_n617), .A3(new_n684), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n641), .A2(new_n266), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n559), .A3(new_n667), .A4(new_n723), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n811), .A2(new_n581), .A3(new_n580), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n806), .A2(new_n809), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(new_n673), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n815), .A2(KEYINPUT116), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(KEYINPUT116), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n816), .A2(new_n374), .A3(new_n817), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n739), .A2(new_n740), .A3(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n819), .A2(new_n723), .A3(new_n799), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT117), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(KEYINPUT117), .A3(new_n723), .A4(new_n799), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g638(.A(new_n791), .B1(new_n814), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n812), .B1(new_n804), .B2(new_n805), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n809), .A4(new_n820), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n825), .A2(new_n264), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n807), .A2(new_n708), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n829), .B(KEYINPUT48), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n811), .A2(new_n582), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n828), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT111), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n784), .A2(new_n833), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n748), .A2(new_n752), .A3(KEYINPUT111), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT53), .B1(new_n836), .B2(new_n782), .ZN(new_n837));
  INV_X1    g651(.A(new_n784), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n773), .A2(new_n783), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g653(.A(KEYINPUT54), .B1(new_n837), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT112), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n783), .B1(new_n755), .B2(new_n773), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n782), .A2(KEYINPUT53), .A3(new_n784), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n844), .A2(new_n845), .A3(KEYINPUT54), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n799), .A2(new_n674), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n790), .A2(new_n832), .A3(new_n847), .A4(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n263), .A2(new_n196), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NOR3_X1   g665(.A1(new_n688), .A2(new_n374), .A3(new_n275), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT107), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n815), .A2(KEYINPUT49), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n716), .B1(new_n852), .B2(new_n853), .ZN(new_n856));
  AND4_X1   g670(.A1(new_n644), .A2(new_n854), .A3(new_n855), .A4(new_n856), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n857), .B(new_n642), .C1(KEYINPUT49), .C2(new_n815), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n851), .A2(new_n858), .ZN(G75));
  AOI21_X1  g673(.A(new_n783), .B1(new_n836), .B2(new_n782), .ZN(new_n860));
  NOR3_X1   g674(.A1(new_n773), .A2(KEYINPUT53), .A3(new_n838), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n860), .A2(new_n861), .A3(new_n226), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n862), .A2(G210), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT56), .ZN(new_n864));
  XOR2_X1   g678(.A(new_n317), .B(new_n350), .Z(new_n865));
  XNOR2_X1  g679(.A(new_n865), .B(KEYINPUT55), .ZN(new_n866));
  AND3_X1   g680(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n866), .B1(new_n863), .B2(new_n864), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n196), .A2(G952), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G51));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n860), .A2(new_n861), .A3(new_n871), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n872), .A2(new_n786), .ZN(new_n873));
  XOR2_X1   g687(.A(new_n728), .B(KEYINPUT57), .Z(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(KEYINPUT119), .B(new_n660), .C1(new_n873), .C2(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT119), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n871), .B1(new_n860), .B2(new_n861), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n774), .A2(KEYINPUT54), .A3(new_n785), .ZN(new_n879));
  AOI21_X1  g693(.A(new_n875), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n877), .B1(new_n880), .B2(new_n428), .ZN(new_n881));
  XOR2_X1   g695(.A(new_n727), .B(KEYINPUT120), .Z(new_n882));
  NAND2_X1  g696(.A1(new_n862), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n876), .A2(new_n881), .A3(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n869), .ZN(new_n885));
  AND2_X1   g699(.A1(new_n884), .A2(new_n885), .ZN(G54));
  NAND3_X1  g700(.A1(new_n862), .A2(KEYINPUT58), .A3(G475), .ZN(new_n887));
  INV_X1    g701(.A(new_n224), .ZN(new_n888));
  AND2_X1   g702(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n887), .A2(new_n888), .ZN(new_n890));
  NOR3_X1   g704(.A1(new_n889), .A2(new_n890), .A3(new_n869), .ZN(G60));
  NAND2_X1  g705(.A1(new_n878), .A2(new_n788), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n786), .A2(KEYINPUT113), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n845), .B1(new_n844), .B2(KEYINPUT54), .ZN(new_n894));
  AOI211_X1 g708(.A(KEYINPUT112), .B(new_n871), .C1(new_n842), .C2(new_n843), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n892), .B(new_n893), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  XNOR2_X1  g710(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n254), .A2(new_n226), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n897), .B(new_n898), .Z(new_n899));
  AOI21_X1  g713(.A(new_n576), .B1(new_n896), .B2(new_n899), .ZN(new_n900));
  INV_X1    g714(.A(new_n899), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n873), .A2(new_n575), .A3(new_n901), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n900), .A2(new_n869), .A3(new_n902), .ZN(G63));
  NAND2_X1  g717(.A1(G217), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT60), .Z(new_n905));
  NAND3_X1  g719(.A1(new_n774), .A2(new_n785), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n549), .A2(new_n552), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n869), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n860), .A2(new_n861), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n615), .B(KEYINPUT123), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n909), .A2(KEYINPUT124), .A3(new_n905), .A4(new_n910), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n774), .A2(new_n785), .A3(new_n905), .A4(new_n910), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT124), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n908), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g729(.A1(new_n915), .A2(KEYINPUT122), .A3(KEYINPUT61), .ZN(new_n916));
  AOI21_X1  g730(.A(KEYINPUT61), .B1(new_n915), .B2(KEYINPUT122), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n916), .A2(new_n917), .ZN(G66));
  AOI21_X1  g732(.A(new_n196), .B1(new_n267), .B2(G224), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n757), .A2(new_n772), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n919), .B1(new_n920), .B2(new_n196), .ZN(new_n921));
  INV_X1    g735(.A(G898), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n317), .B1(new_n922), .B2(G953), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n921), .B(new_n923), .ZN(G69));
  XNOR2_X1  g738(.A(new_n459), .B(KEYINPUT125), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(new_n221), .ZN(new_n926));
  NAND2_X1  g740(.A1(G900), .A2(G953), .ZN(new_n927));
  NOR3_X1   g741(.A1(new_n708), .A2(new_n628), .A3(new_n646), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n735), .B1(new_n725), .B2(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n714), .A2(new_n693), .A3(new_n751), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n929), .A2(new_n710), .A3(new_n742), .A4(new_n930), .ZN(new_n931));
  OAI211_X1 g745(.A(new_n926), .B(new_n927), .C1(new_n931), .C2(G953), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n651), .A2(new_n693), .A3(new_n751), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT62), .Z(new_n934));
  OAI21_X1  g748(.A(new_n649), .B1(new_n770), .B2(KEYINPUT126), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(KEYINPUT126), .B2(new_n770), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n936), .A2(new_n778), .A3(new_n723), .ZN(new_n937));
  NAND4_X1  g751(.A1(new_n934), .A2(new_n736), .A3(new_n742), .A4(new_n937), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n938), .A2(new_n196), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n932), .B1(new_n939), .B2(new_n926), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n196), .B1(G227), .B2(G900), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT127), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n932), .B2(new_n942), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n940), .B(new_n943), .Z(G72));
  XOR2_X1   g758(.A(new_n636), .B(KEYINPUT63), .Z(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n938), .B2(new_n920), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n946), .A2(new_n473), .A3(new_n462), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n945), .B1(new_n931), .B2(new_n920), .ZN(new_n948));
  NAND3_X1  g762(.A1(new_n948), .A2(new_n466), .A3(new_n472), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n467), .A2(new_n474), .A3(new_n515), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n844), .A2(new_n945), .A3(new_n950), .ZN(new_n951));
  AND4_X1   g765(.A1(new_n885), .A2(new_n947), .A3(new_n949), .A4(new_n951), .ZN(G57));
endmodule


