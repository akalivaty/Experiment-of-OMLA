//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 0 1 1 1 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:14 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n763, new_n764,
    new_n765, new_n766, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n955,
    new_n956, new_n957, new_n958, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(G107), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G104), .ZN(new_n191));
  INV_X1    g005(.A(G104), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G107), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G101), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT3), .B1(new_n192), .B2(G107), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n197), .A2(new_n190), .A3(G104), .ZN(new_n198));
  INV_X1    g012(.A(G101), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .A4(new_n193), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n200), .A2(KEYINPUT81), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(KEYINPUT81), .ZN(new_n202));
  OAI21_X1  g016(.A(new_n195), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G113), .ZN(new_n204));
  INV_X1    g018(.A(G116), .ZN(new_n205));
  NOR2_X1   g019(.A1(new_n205), .A2(G119), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT5), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n204), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT67), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n209), .B1(new_n205), .B2(G119), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT67), .A3(G116), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n205), .A2(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n210), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n208), .B1(new_n214), .B2(new_n207), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n204), .A2(KEYINPUT2), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT2), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G113), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  NAND4_X1  g033(.A1(new_n219), .A2(new_n210), .A3(new_n212), .A4(new_n213), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n215), .A2(new_n220), .ZN(new_n221));
  NOR2_X1   g035(.A1(new_n203), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT2), .B(G113), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT69), .ZN(new_n226));
  OAI211_X1 g040(.A(new_n225), .B(new_n226), .C1(new_n214), .C2(new_n223), .ZN(new_n227));
  INV_X1    g041(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g042(.A(new_n226), .B1(new_n220), .B2(new_n225), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n224), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n225), .B1(new_n214), .B2(new_n223), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n231), .A2(KEYINPUT69), .ZN(new_n232));
  INV_X1    g046(.A(new_n224), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n232), .A2(new_n233), .A3(new_n227), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n230), .A2(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n196), .A2(new_n198), .A3(new_n193), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G101), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT82), .ZN(new_n238));
  OAI21_X1  g052(.A(KEYINPUT4), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT4), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n236), .A2(KEYINPUT82), .A3(new_n240), .A4(G101), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n198), .A2(new_n193), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT81), .ZN(new_n244));
  NAND4_X1  g058(.A1(new_n243), .A2(new_n244), .A3(new_n199), .A4(new_n196), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n200), .A2(KEYINPUT81), .ZN(new_n246));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n237), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n222), .B1(new_n235), .B2(new_n248), .ZN(new_n249));
  XNOR2_X1  g063(.A(G110), .B(G122), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n250), .ZN(new_n252));
  AOI22_X1  g066(.A1(new_n230), .A2(new_n234), .B1(new_n242), .B2(new_n247), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n252), .B1(new_n253), .B2(new_n222), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n251), .A2(KEYINPUT6), .A3(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G146), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G143), .ZN(new_n257));
  INV_X1    g071(.A(G143), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n257), .A2(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(KEYINPUT0), .A2(G128), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT64), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT0), .ZN(new_n263));
  INV_X1    g077(.A(G128), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n262), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  OAI21_X1  g079(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n260), .A2(new_n261), .A3(new_n265), .A4(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT65), .ZN(new_n268));
  XNOR2_X1  g082(.A(G143), .B(G146), .ZN(new_n269));
  INV_X1    g083(.A(new_n261), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(new_n266), .ZN(new_n273));
  NOR3_X1   g087(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND4_X1  g089(.A1(new_n275), .A2(new_n268), .A3(new_n260), .A4(new_n261), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n272), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G125), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n257), .A2(KEYINPUT1), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n260), .A2(new_n279), .A3(G128), .ZN(new_n280));
  OAI211_X1 g094(.A(new_n257), .B(new_n259), .C1(KEYINPUT1), .C2(new_n264), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n278), .B1(G125), .B2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(G224), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n284), .A2(G953), .ZN(new_n285));
  XOR2_X1   g099(.A(new_n283), .B(new_n285), .Z(new_n286));
  INV_X1    g100(.A(KEYINPUT85), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n228), .A2(new_n229), .A3(new_n224), .ZN(new_n288));
  AOI21_X1  g102(.A(new_n233), .B1(new_n232), .B2(new_n227), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n248), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n222), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n250), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT6), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n287), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NOR4_X1   g108(.A1(new_n249), .A2(KEYINPUT85), .A3(KEYINPUT6), .A4(new_n250), .ZN(new_n295));
  OAI211_X1 g109(.A(new_n255), .B(new_n286), .C1(new_n294), .C2(new_n295), .ZN(new_n296));
  OR2_X1    g110(.A1(new_n285), .A2(KEYINPUT87), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT7), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n298), .B1(new_n285), .B2(KEYINPUT87), .ZN(new_n299));
  AND3_X1   g113(.A1(new_n283), .A2(new_n297), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(KEYINPUT86), .A2(KEYINPUT7), .ZN(new_n301));
  INV_X1    g115(.A(KEYINPUT86), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n285), .B1(new_n302), .B2(new_n298), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n283), .B1(new_n301), .B2(new_n303), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n250), .B(KEYINPUT8), .Z(new_n305));
  NAND2_X1  g119(.A1(new_n203), .A2(new_n221), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n305), .B1(new_n291), .B2(new_n306), .ZN(new_n307));
  NOR3_X1   g121(.A1(new_n300), .A2(new_n304), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g122(.A(G902), .B1(new_n308), .B2(new_n251), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n189), .B1(new_n296), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n296), .A2(new_n309), .A3(new_n189), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n188), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT9), .B(G234), .ZN(new_n314));
  OAI21_X1  g128(.A(G221), .B1(new_n314), .B2(G902), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT11), .ZN(new_n317));
  INV_X1    g131(.A(G134), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n317), .B1(new_n318), .B2(G137), .ZN(new_n319));
  INV_X1    g133(.A(G137), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n320), .A2(KEYINPUT11), .A3(G134), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n318), .A2(G137), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G131), .ZN(new_n324));
  INV_X1    g138(.A(G131), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n319), .A2(new_n321), .A3(new_n325), .A4(new_n322), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n203), .A2(new_n282), .ZN(new_n328));
  INV_X1    g142(.A(new_n282), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n245), .A2(new_n246), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n329), .B1(new_n330), .B2(new_n195), .ZN(new_n331));
  OAI211_X1 g145(.A(KEYINPUT12), .B(new_n327), .C1(new_n328), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(KEYINPUT83), .ZN(new_n333));
  INV_X1    g147(.A(new_n327), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n203), .A2(new_n282), .ZN(new_n335));
  AOI22_X1  g149(.A1(new_n245), .A2(new_n246), .B1(G101), .B2(new_n194), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n329), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n334), .B1(new_n335), .B2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT83), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT12), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n327), .B1(new_n328), .B2(new_n331), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT12), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n333), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  AND3_X1   g158(.A1(new_n272), .A2(KEYINPUT70), .A3(new_n276), .ZN(new_n345));
  AOI21_X1  g159(.A(KEYINPUT70), .B1(new_n272), .B2(new_n276), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(new_n248), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT10), .ZN(new_n349));
  OAI21_X1  g163(.A(new_n349), .B1(new_n203), .B2(new_n282), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n280), .A2(KEYINPUT71), .A3(new_n281), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT71), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n282), .A2(new_n352), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n336), .A2(KEYINPUT10), .A3(new_n351), .A4(new_n353), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n348), .A2(new_n334), .A3(new_n350), .A4(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n344), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(G953), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n357), .A2(G227), .ZN(new_n358));
  XNOR2_X1  g172(.A(new_n358), .B(KEYINPUT80), .ZN(new_n359));
  XNOR2_X1  g173(.A(G110), .B(G140), .ZN(new_n360));
  XNOR2_X1  g174(.A(new_n359), .B(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n355), .A2(new_n362), .ZN(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n277), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n272), .A2(new_n276), .A3(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g182(.A(new_n200), .B(new_n244), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n369), .A2(new_n237), .B1(new_n239), .B2(new_n241), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n350), .B(new_n354), .C1(new_n368), .C2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(KEYINPUT84), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NAND4_X1  g187(.A1(new_n348), .A2(KEYINPUT84), .A3(new_n350), .A4(new_n354), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n327), .ZN(new_n375));
  AOI22_X1  g189(.A1(new_n356), .A2(new_n361), .B1(new_n364), .B2(new_n375), .ZN(new_n376));
  OAI21_X1  g190(.A(G469), .B1(new_n376), .B2(G902), .ZN(new_n377));
  INV_X1    g191(.A(G469), .ZN(new_n378));
  INV_X1    g192(.A(G902), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n362), .B1(new_n375), .B2(new_n355), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n339), .B1(new_n338), .B2(KEYINPUT12), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n338), .A2(KEYINPUT12), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n363), .B1(new_n383), .B2(new_n340), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n378), .B(new_n379), .C1(new_n380), .C2(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n316), .B1(new_n377), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(G475), .ZN(new_n387));
  INV_X1    g201(.A(G237), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n388), .A2(new_n357), .A3(G214), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n389), .A2(KEYINPUT88), .A3(new_n258), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n258), .A2(KEYINPUT88), .ZN(new_n391));
  NOR2_X1   g205(.A1(G237), .A2(G953), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(G214), .A3(new_n392), .ZN(new_n393));
  AOI21_X1  g207(.A(new_n325), .B1(new_n390), .B2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT17), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n325), .A3(new_n393), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT16), .ZN(new_n399));
  INV_X1    g213(.A(G140), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(new_n400), .A3(G125), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(G125), .ZN(new_n402));
  INV_X1    g216(.A(G125), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G140), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n402), .A2(new_n404), .ZN(new_n405));
  OAI211_X1 g219(.A(G146), .B(new_n401), .C1(new_n405), .C2(new_n399), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n401), .B1(new_n405), .B2(new_n399), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n407), .A2(new_n256), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n390), .A2(new_n393), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n409), .A2(KEYINPUT17), .A3(G131), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n398), .A2(new_n406), .A3(new_n408), .A4(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n409), .A2(KEYINPUT18), .A3(G131), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n405), .B(G146), .ZN(new_n413));
  NAND2_X1  g227(.A1(KEYINPUT18), .A2(G131), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n390), .A2(new_n414), .A3(new_n393), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n411), .A2(new_n416), .ZN(new_n417));
  XOR2_X1   g231(.A(G113), .B(G122), .Z(new_n418));
  XOR2_X1   g232(.A(KEYINPUT89), .B(G104), .Z(new_n419));
  XOR2_X1   g233(.A(new_n418), .B(new_n419), .Z(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n417), .A2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT91), .ZN(new_n423));
  AND3_X1   g237(.A1(new_n390), .A2(new_n325), .A3(new_n393), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n424), .A2(new_n394), .A3(KEYINPUT17), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n410), .A2(new_n406), .A3(new_n408), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n416), .B(new_n420), .C1(new_n425), .C2(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n422), .A2(new_n423), .A3(new_n427), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n420), .B1(new_n411), .B2(new_n416), .ZN(new_n429));
  AOI21_X1  g243(.A(G902), .B1(new_n429), .B2(KEYINPUT91), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n387), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  NOR2_X1   g245(.A1(G475), .A2(G902), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n402), .A2(new_n404), .A3(KEYINPUT19), .ZN(new_n433));
  AOI21_X1  g247(.A(KEYINPUT19), .B1(new_n402), .B2(new_n404), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n256), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  OAI211_X1 g249(.A(new_n406), .B(new_n435), .C1(new_n424), .C2(new_n394), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n416), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n421), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n438), .A2(new_n427), .A3(KEYINPUT90), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT90), .B1(new_n438), .B2(new_n427), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n432), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n441), .A2(KEYINPUT20), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n438), .A2(new_n427), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT20), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n443), .A2(new_n444), .A3(new_n432), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n431), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  INV_X1    g260(.A(G478), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT15), .ZN(new_n448));
  INV_X1    g262(.A(G122), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(G116), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n190), .B1(new_n450), .B2(KEYINPUT14), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n205), .A2(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n451), .A2(new_n453), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n264), .A2(G143), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT92), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n456), .B(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n258), .A2(G128), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n318), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n457), .A2(new_n258), .A3(G128), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n264), .B2(G143), .ZN(new_n462));
  OAI21_X1  g276(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n463), .A2(G134), .ZN(new_n464));
  OAI211_X1 g278(.A(new_n454), .B(new_n455), .C1(new_n460), .C2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n466));
  XNOR2_X1  g280(.A(new_n459), .B(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n461), .A2(new_n462), .ZN(new_n468));
  OAI21_X1  g282(.A(G134), .B1(new_n467), .B2(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n458), .A2(new_n318), .A3(new_n459), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n453), .B(G107), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G217), .ZN(new_n473));
  NOR3_X1   g287(.A1(new_n314), .A2(new_n473), .A3(G953), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n465), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n474), .B1(new_n465), .B2(new_n472), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n379), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n448), .B1(new_n478), .B2(KEYINPUT93), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(KEYINPUT93), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n465), .A2(new_n472), .ZN(new_n481));
  INV_X1    g295(.A(new_n474), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(G902), .B1(new_n483), .B2(new_n475), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT93), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n480), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n479), .B1(new_n487), .B2(new_n448), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n446), .A2(new_n488), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n357), .A2(G952), .ZN(new_n490));
  NAND2_X1  g304(.A1(G234), .A2(G237), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g306(.A(KEYINPUT21), .B(G898), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n379), .B1(G234), .B2(G237), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(G953), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g309(.A(new_n489), .B1(new_n492), .B2(new_n495), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n313), .A2(new_n386), .A3(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT29), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n366), .A2(new_n327), .A3(new_n367), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n318), .A2(G137), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n320), .A2(G134), .ZN(new_n501));
  OAI21_X1  g315(.A(G131), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n326), .A2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(new_n503), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n353), .A2(new_n504), .A3(new_n351), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n499), .A2(KEYINPUT30), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n277), .A2(new_n327), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT66), .B1(new_n282), .B2(new_n503), .ZN(new_n508));
  INV_X1    g322(.A(KEYINPUT66), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n329), .A2(new_n509), .A3(new_n504), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT30), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n506), .A2(new_n235), .A3(new_n513), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n499), .A2(new_n234), .A3(new_n230), .A4(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n392), .A2(G210), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(KEYINPUT27), .ZN(new_n518));
  XNOR2_X1  g332(.A(KEYINPUT26), .B(G101), .ZN(new_n519));
  XNOR2_X1  g333(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n516), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n511), .A2(new_n235), .ZN(new_n523));
  INV_X1    g337(.A(KEYINPUT73), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n511), .A2(new_n235), .A3(KEYINPUT73), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n515), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n527), .A2(KEYINPUT28), .ZN(new_n528));
  NOR3_X1   g342(.A1(new_n345), .A2(new_n346), .A3(new_n334), .ZN(new_n529));
  INV_X1    g343(.A(new_n505), .ZN(new_n530));
  OAI21_X1  g344(.A(KEYINPUT74), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n235), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT74), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n499), .A2(new_n533), .A3(new_n505), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT28), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n528), .A2(new_n537), .ZN(new_n538));
  OAI211_X1 g352(.A(new_n498), .B(new_n522), .C1(new_n538), .C2(new_n521), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n499), .A2(new_n505), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n235), .B1(new_n540), .B2(KEYINPUT74), .ZN(new_n541));
  AOI21_X1  g355(.A(KEYINPUT28), .B1(new_n541), .B2(new_n534), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n235), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n536), .B1(new_n543), .B2(new_n515), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n521), .A2(new_n498), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n539), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(G472), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT32), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT31), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT72), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n515), .A2(new_n552), .A3(new_n520), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(new_n514), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n552), .B1(new_n515), .B2(new_n520), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n515), .A2(new_n520), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n557), .A2(KEYINPUT72), .ZN(new_n558));
  NAND4_X1  g372(.A1(new_n558), .A2(KEYINPUT31), .A3(new_n514), .A4(new_n553), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n556), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n530), .B1(new_n347), .B2(new_n327), .ZN(new_n561));
  AOI22_X1  g375(.A1(new_n532), .A2(new_n561), .B1(new_n523), .B2(new_n524), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n536), .B1(new_n562), .B2(new_n526), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n521), .B1(new_n563), .B2(new_n542), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(G472), .A2(G902), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n550), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g381(.A(new_n566), .ZN(new_n568));
  AOI211_X1 g382(.A(KEYINPUT32), .B(new_n568), .C1(new_n560), .C2(new_n564), .ZN(new_n569));
  OAI21_X1  g383(.A(new_n549), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n264), .A2(KEYINPUT23), .A3(G119), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n571), .B(KEYINPUT75), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT23), .B1(new_n264), .B2(G119), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(KEYINPUT76), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n211), .A2(G128), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n575), .A2(new_n576), .A3(KEYINPUT23), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n264), .A2(G119), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G110), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n572), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n575), .A2(new_n578), .ZN(new_n582));
  XNOR2_X1  g396(.A(KEYINPUT24), .B(G110), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g398(.A1(new_n581), .A2(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n405), .A2(G146), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n585), .A2(new_n406), .A3(new_n587), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n582), .A2(new_n583), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n408), .B2(new_n406), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n572), .A2(new_n579), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(G110), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n588), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g408(.A(KEYINPUT22), .B(G137), .ZN(new_n595));
  NAND3_X1  g409(.A1(new_n357), .A2(G221), .A3(G234), .ZN(new_n596));
  XNOR2_X1  g410(.A(new_n595), .B(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(KEYINPUT77), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n594), .A2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n588), .A2(new_n593), .A3(new_n597), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n473), .B1(G234), .B2(new_n379), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n602), .A2(G902), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(KEYINPUT78), .ZN(new_n605));
  INV_X1    g419(.A(new_n602), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n600), .A2(new_n379), .A3(new_n601), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n606), .B1(new_n607), .B2(KEYINPUT25), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT25), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n600), .A2(new_n601), .A3(new_n609), .A4(new_n379), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n608), .A2(new_n610), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n605), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT79), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n497), .A2(new_n570), .A3(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(G101), .ZN(G3));
  AOI22_X1  g429(.A1(new_n538), .A2(new_n521), .B1(new_n556), .B2(new_n559), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n616), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n565), .A2(new_n566), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n620), .A2(new_n613), .A3(new_n386), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n495), .A2(new_n492), .ZN(new_n622));
  AND3_X1   g436(.A1(new_n296), .A2(new_n309), .A3(new_n189), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n187), .B(new_n622), .C1(new_n623), .C2(new_n310), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n483), .A2(new_n475), .ZN(new_n625));
  OAI21_X1  g439(.A(KEYINPUT33), .B1(new_n474), .B2(KEYINPUT94), .ZN(new_n626));
  OR2_X1    g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n626), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n447), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(G478), .A2(G902), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n478), .B2(G478), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  NOR3_X1   g447(.A1(new_n624), .A2(new_n446), .A3(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n621), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(KEYINPUT95), .B(KEYINPUT34), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n636), .B(new_n637), .ZN(G6));
  XNOR2_X1  g452(.A(new_n441), .B(KEYINPUT20), .ZN(new_n639));
  INV_X1    g453(.A(new_n431), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n485), .B1(new_n625), .B2(new_n379), .ZN(new_n641));
  AOI211_X1 g455(.A(KEYINPUT93), .B(G902), .C1(new_n483), .C2(new_n475), .ZN(new_n642));
  OAI21_X1  g456(.A(new_n448), .B1(new_n641), .B2(new_n642), .ZN(new_n643));
  INV_X1    g457(.A(new_n479), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n639), .A2(new_n640), .A3(new_n645), .ZN(new_n646));
  AND3_X1   g460(.A1(new_n313), .A2(new_n622), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n621), .A2(new_n647), .ZN(new_n648));
  XOR2_X1   g462(.A(KEYINPUT35), .B(G107), .Z(new_n649));
  XNOR2_X1  g463(.A(new_n648), .B(new_n649), .ZN(G9));
  INV_X1    g464(.A(KEYINPUT97), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n594), .B1(KEYINPUT36), .B2(new_n599), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT36), .ZN(new_n653));
  NAND4_X1  g467(.A1(new_n588), .A2(new_n598), .A3(new_n593), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n652), .A2(new_n603), .A3(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(new_n655), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n656), .B1(new_n608), .B2(new_n610), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT96), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n659));
  AOI211_X1 g473(.A(new_n659), .B(new_n656), .C1(new_n608), .C2(new_n610), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n651), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n611), .A2(new_n655), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n659), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n657), .A2(KEYINPUT96), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n663), .A2(KEYINPUT97), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n661), .A2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n497), .A2(new_n620), .A3(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT37), .B(G110), .Z(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G12));
  NAND2_X1  g483(.A1(G469), .A2(G902), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n356), .A2(new_n361), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n364), .A2(new_n375), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n671), .A2(G469), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n385), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n315), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n187), .B1(new_n623), .B2(new_n310), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g491(.A1(new_n357), .A2(G900), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n494), .A2(new_n678), .ZN(new_n679));
  OR2_X1    g493(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(KEYINPUT98), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n680), .A2(new_n492), .A3(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n639), .A2(new_n640), .A3(new_n645), .A4(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n683), .B1(new_n661), .B2(new_n665), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n677), .A2(new_n570), .A3(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n685), .A2(KEYINPUT99), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n677), .A2(new_n570), .A3(new_n684), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  NOR2_X1   g504(.A1(new_n623), .A2(new_n310), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n558), .A2(new_n514), .A3(new_n553), .ZN(new_n694));
  INV_X1    g508(.A(new_n515), .ZN(new_n695));
  AOI22_X1  g509(.A1(new_n499), .A2(new_n505), .B1(new_n234), .B2(new_n230), .ZN(new_n696));
  OAI21_X1  g510(.A(new_n521), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g512(.A(G472), .B1(new_n698), .B2(G902), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(new_n567), .B2(new_n569), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n663), .A2(new_n664), .ZN(new_n702));
  INV_X1    g516(.A(new_n446), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n703), .A2(new_n187), .A3(new_n645), .ZN(new_n704));
  NOR4_X1   g518(.A1(new_n693), .A2(new_n701), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n682), .B(KEYINPUT39), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n386), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n708));
  OR2_X1    g522(.A1(new_n707), .A2(KEYINPUT40), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n705), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT101), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  AND2_X1   g526(.A1(new_n570), .A2(new_n666), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n703), .A2(new_n632), .A3(new_n682), .ZN(new_n714));
  INV_X1    g528(.A(new_n714), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n313), .A2(new_n386), .A3(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n713), .A2(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G146), .ZN(G48));
  OAI21_X1  g533(.A(new_n379), .B1(new_n380), .B2(new_n384), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n720), .A2(G469), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(new_n315), .A3(new_n385), .ZN(new_n722));
  NAND4_X1  g536(.A1(new_n634), .A2(new_n570), .A3(new_n613), .A4(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(KEYINPUT41), .B(G113), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n723), .B(new_n724), .ZN(G15));
  NAND4_X1  g539(.A1(new_n647), .A2(new_n570), .A3(new_n613), .A4(new_n722), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(G116), .ZN(G18));
  NAND3_X1  g541(.A1(new_n721), .A2(new_n315), .A3(new_n385), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n676), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n570), .A2(new_n729), .A3(new_n496), .A4(new_n666), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G119), .ZN(G21));
  INV_X1    g545(.A(KEYINPUT102), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n732), .B1(new_n542), .B2(new_n544), .ZN(new_n733));
  OAI21_X1  g547(.A(KEYINPUT28), .B1(new_n695), .B2(new_n696), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n537), .A2(KEYINPUT102), .A3(new_n734), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n733), .A2(new_n735), .A3(new_n521), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n568), .B1(new_n736), .B2(new_n560), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n560), .B2(new_n564), .ZN(new_n738));
  INV_X1    g552(.A(G472), .ZN(new_n739));
  OAI22_X1  g553(.A1(new_n737), .A2(KEYINPUT103), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT103), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n741), .B(new_n568), .C1(new_n736), .C2(new_n560), .ZN(new_n742));
  NOR2_X1   g556(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(new_n612), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT104), .ZN(new_n745));
  OAI21_X1  g559(.A(new_n745), .B1(new_n446), .B2(new_n488), .ZN(new_n746));
  INV_X1    g560(.A(new_n445), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n747), .B1(new_n441), .B2(KEYINPUT20), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n645), .B(KEYINPUT104), .C1(new_n748), .C2(new_n431), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n746), .A2(new_n749), .ZN(new_n750));
  OR3_X1    g564(.A1(new_n624), .A2(new_n728), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n744), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(new_n449), .ZN(G24));
  NAND2_X1  g567(.A1(new_n537), .A2(new_n734), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n520), .B1(new_n754), .B2(new_n732), .ZN(new_n755));
  AOI22_X1  g569(.A1(new_n755), .A2(new_n735), .B1(new_n556), .B2(new_n559), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n741), .B1(new_n756), .B2(new_n568), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n617), .A3(new_n702), .A4(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n722), .A2(new_n313), .A3(new_n715), .ZN(new_n760));
  OAI21_X1  g574(.A(KEYINPUT105), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NOR3_X1   g575(.A1(new_n728), .A2(new_n676), .A3(new_n714), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT105), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n743), .A2(new_n762), .A3(new_n763), .A4(new_n702), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(KEYINPUT106), .B(G125), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n765), .B(new_n766), .ZN(G27));
  OAI21_X1  g581(.A(KEYINPUT32), .B1(new_n616), .B2(new_n568), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n565), .A2(new_n550), .A3(new_n566), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n770), .A2(KEYINPUT107), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT107), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n768), .A2(new_n769), .A3(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n771), .A2(new_n549), .A3(new_n773), .ZN(new_n774));
  NOR3_X1   g588(.A1(new_n623), .A2(new_n310), .A3(new_n188), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NOR3_X1   g590(.A1(new_n776), .A2(new_n675), .A3(new_n714), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n774), .A2(KEYINPUT42), .A3(new_n612), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n386), .A2(new_n775), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n779), .A2(new_n570), .A3(new_n613), .A4(new_n715), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT42), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n778), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  AND2_X1   g598(.A1(new_n570), .A2(new_n613), .ZN(new_n785));
  INV_X1    g599(.A(new_n683), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(KEYINPUT108), .A3(new_n786), .A4(new_n779), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n779), .A2(new_n570), .A3(new_n613), .A4(new_n786), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT108), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n790), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n791), .B(G134), .ZN(G36));
  XNOR2_X1  g606(.A(new_n775), .B(KEYINPUT110), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n633), .A2(new_n703), .ZN(new_n794));
  XOR2_X1   g608(.A(new_n794), .B(KEYINPUT43), .Z(new_n795));
  AOI21_X1  g609(.A(new_n795), .B1(new_n663), .B2(new_n664), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n619), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(KEYINPUT44), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT44), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n799), .A3(new_n619), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  OR2_X1    g615(.A1(new_n376), .A2(KEYINPUT45), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n376), .A2(KEYINPUT45), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(G469), .A3(new_n803), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n804), .A2(new_n670), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT46), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n807), .B(KEYINPUT109), .ZN(new_n808));
  INV_X1    g622(.A(new_n385), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n805), .B2(new_n806), .ZN(new_n810));
  AOI21_X1  g624(.A(new_n316), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n801), .A2(new_n706), .A3(new_n811), .ZN(new_n812));
  XNOR2_X1  g626(.A(new_n812), .B(G137), .ZN(G39));
  XOR2_X1   g627(.A(new_n811), .B(KEYINPUT47), .Z(new_n814));
  OR4_X1    g628(.A1(new_n570), .A2(new_n776), .A3(new_n613), .A4(new_n714), .ZN(new_n815));
  OR2_X1    g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  NAND2_X1  g631(.A1(new_n721), .A2(new_n385), .ZN(new_n818));
  XOR2_X1   g632(.A(new_n818), .B(KEYINPUT49), .Z(new_n819));
  NAND3_X1  g633(.A1(new_n612), .A2(new_n187), .A3(new_n315), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n794), .B1(new_n820), .B2(KEYINPUT111), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n821), .B1(KEYINPUT111), .B2(new_n820), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n819), .A2(new_n693), .A3(new_n701), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g637(.A1(new_n795), .A2(new_n492), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n824), .A2(new_n612), .A3(new_n743), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT116), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT50), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n187), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g642(.A1(new_n693), .A2(new_n722), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n825), .A2(new_n829), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n826), .A2(new_n827), .ZN(new_n831));
  XNOR2_X1  g645(.A(new_n830), .B(new_n831), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n721), .A2(new_n316), .A3(new_n385), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n814), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n825), .A2(new_n793), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(new_n832), .B1(new_n834), .B2(new_n836), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n776), .A2(new_n728), .ZN(new_n838));
  INV_X1    g652(.A(new_n492), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n613), .A2(new_n701), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n840), .A2(new_n446), .A3(new_n633), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n824), .A2(new_n838), .ZN(new_n844));
  INV_X1    g658(.A(new_n759), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n842), .A2(new_n843), .A3(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n837), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g662(.A1(new_n848), .A2(KEYINPUT51), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT52), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n676), .A2(new_n750), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n657), .A2(new_n682), .ZN(new_n852));
  AND3_X1   g666(.A1(new_n674), .A2(new_n315), .A3(new_n852), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n700), .A2(new_n851), .A3(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n570), .A2(new_n666), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n854), .B1(new_n855), .B2(new_n716), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n856), .B1(new_n688), .B2(new_n686), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n850), .B1(new_n857), .B2(new_n765), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n674), .A2(new_n315), .A3(new_n852), .ZN(new_n859));
  AOI21_X1  g673(.A(new_n859), .B1(new_n770), .B2(new_n699), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n713), .A2(new_n717), .B1(new_n860), .B2(new_n851), .ZN(new_n861));
  AND4_X1   g675(.A1(new_n850), .A2(new_n689), .A3(new_n765), .A4(new_n861), .ZN(new_n862));
  OAI21_X1  g676(.A(KEYINPUT114), .B1(new_n858), .B2(new_n862), .ZN(new_n863));
  AND4_X1   g677(.A1(new_n640), .A2(new_n639), .A3(new_n488), .A4(new_n682), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n779), .A2(new_n570), .A3(new_n666), .A4(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT112), .ZN(new_n866));
  OR2_X1    g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n865), .A2(new_n866), .ZN(new_n868));
  AOI22_X1  g682(.A1(new_n867), .A2(new_n868), .B1(new_n845), .B2(new_n777), .ZN(new_n869));
  AOI22_X1  g683(.A1(new_n778), .A2(new_n782), .B1(new_n787), .B2(new_n790), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n726), .A2(new_n614), .A3(new_n667), .A4(new_n723), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n489), .B1(new_n446), .B2(new_n632), .ZN(new_n872));
  NOR2_X1   g686(.A1(new_n624), .A2(new_n872), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n620), .A2(new_n873), .A3(new_n613), .A4(new_n386), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n874), .B(new_n730), .C1(new_n744), .C2(new_n751), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n871), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g690(.A1(new_n869), .A2(new_n870), .A3(new_n876), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n689), .A2(new_n765), .A3(new_n861), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n878), .A2(KEYINPUT52), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n857), .A2(new_n850), .A3(new_n765), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT114), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n863), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT53), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g699(.A(KEYINPUT115), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  AND4_X1   g702(.A1(new_n880), .A2(new_n876), .A3(new_n870), .A4(new_n869), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n689), .A2(new_n765), .ZN(new_n890));
  OR2_X1    g704(.A1(new_n890), .A2(KEYINPUT113), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n890), .A2(KEYINPUT113), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n856), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI211_X1 g707(.A(new_n889), .B(KEYINPUT53), .C1(new_n893), .C2(new_n850), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n883), .A2(KEYINPUT115), .A3(new_n884), .ZN(new_n895));
  NAND4_X1  g709(.A1(new_n887), .A2(new_n888), .A3(new_n894), .A4(new_n895), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n893), .A2(new_n850), .ZN(new_n897));
  AOI21_X1  g711(.A(KEYINPUT53), .B1(new_n897), .B2(new_n889), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n883), .A2(new_n884), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n896), .B1(new_n900), .B2(new_n888), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n774), .A2(new_n612), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n844), .A2(new_n902), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT48), .Z(new_n904));
  NAND3_X1  g718(.A1(new_n840), .A2(new_n703), .A3(new_n632), .ZN(new_n905));
  INV_X1    g719(.A(new_n729), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n905), .B(new_n490), .C1(new_n906), .C2(new_n825), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n904), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n847), .A2(KEYINPUT118), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n909), .A2(KEYINPUT51), .A3(new_n910), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n908), .B1(new_n837), .B2(new_n911), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n849), .A2(new_n901), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g727(.A1(G952), .A2(G953), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n823), .B1(new_n913), .B2(new_n914), .ZN(G75));
  NOR2_X1   g729(.A1(new_n357), .A2(G952), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n255), .B1(new_n294), .B2(new_n295), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(new_n286), .ZN(new_n918));
  XNOR2_X1  g732(.A(new_n918), .B(KEYINPUT55), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n895), .A2(new_n894), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT115), .B1(new_n883), .B2(new_n884), .ZN(new_n921));
  OAI211_X1 g735(.A(G210), .B(G902), .C1(new_n920), .C2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n919), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n919), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT119), .ZN(new_n926));
  INV_X1    g740(.A(KEYINPUT119), .ZN(new_n927));
  NAND4_X1  g741(.A1(new_n922), .A2(new_n927), .A3(new_n923), .A4(new_n919), .ZN(new_n928));
  AOI211_X1 g742(.A(new_n916), .B(new_n924), .C1(new_n926), .C2(new_n928), .ZN(G51));
  INV_X1    g743(.A(new_n804), .ZN(new_n930));
  OAI211_X1 g744(.A(G902), .B(new_n930), .C1(new_n920), .C2(new_n921), .ZN(new_n931));
  INV_X1    g745(.A(new_n931), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n380), .A2(new_n384), .ZN(new_n933));
  OAI21_X1  g747(.A(KEYINPUT54), .B1(new_n920), .B2(new_n921), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(new_n896), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n670), .B(KEYINPUT57), .Z(new_n936));
  AOI21_X1  g750(.A(new_n933), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n932), .B1(new_n937), .B2(KEYINPUT120), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT120), .ZN(new_n939));
  INV_X1    g753(.A(new_n936), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n940), .B1(new_n934), .B2(new_n896), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n933), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n916), .B1(new_n938), .B2(new_n942), .ZN(G54));
  INV_X1    g757(.A(new_n920), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n379), .B1(new_n944), .B2(new_n887), .ZN(new_n945));
  AND2_X1   g759(.A1(KEYINPUT58), .A2(G475), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g761(.A1(new_n439), .A2(new_n440), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(KEYINPUT121), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  AOI21_X1  g764(.A(new_n916), .B1(new_n947), .B2(new_n949), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT121), .ZN(new_n952));
  NAND4_X1  g766(.A1(new_n945), .A2(new_n952), .A3(new_n948), .A4(new_n946), .ZN(new_n953));
  AND3_X1   g767(.A1(new_n950), .A2(new_n951), .A3(new_n953), .ZN(G60));
  AND2_X1   g768(.A1(new_n627), .A2(new_n628), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n630), .B(KEYINPUT59), .ZN(new_n956));
  AND3_X1   g770(.A1(new_n935), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n955), .B1(new_n901), .B2(new_n956), .ZN(new_n958));
  NOR3_X1   g772(.A1(new_n957), .A2(new_n958), .A3(new_n916), .ZN(G63));
  XNOR2_X1  g773(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n473), .A2(new_n379), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n962), .B1(new_n920), .B2(new_n921), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n652), .A2(new_n654), .ZN(new_n964));
  OR2_X1    g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n916), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n600), .A2(new_n601), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n963), .A2(new_n967), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n965), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g783(.A(KEYINPUT61), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g785(.A1(new_n965), .A2(KEYINPUT61), .A3(new_n966), .A4(new_n968), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n493), .B2(new_n284), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n876), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n917), .B1(G898), .B2(new_n357), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  AOI21_X1  g791(.A(new_n357), .B1(G227), .B2(G900), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n506), .A2(new_n513), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n433), .A2(new_n434), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n980), .B(new_n981), .ZN(new_n982));
  XNOR2_X1  g796(.A(KEYINPUT124), .B(G900), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n979), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  XOR2_X1   g798(.A(new_n984), .B(KEYINPUT125), .Z(new_n985));
  AOI22_X1  g799(.A1(new_n891), .A2(new_n892), .B1(new_n713), .B2(new_n717), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n811), .A2(new_n706), .A3(new_n902), .A4(new_n851), .ZN(new_n987));
  AND3_X1   g801(.A1(new_n812), .A2(new_n870), .A3(new_n987), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n816), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n678), .B1(new_n989), .B2(new_n357), .ZN(new_n990));
  INV_X1    g804(.A(new_n982), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n979), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n986), .A2(new_n711), .ZN(new_n993));
  OR2_X1    g807(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(KEYINPUT62), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n776), .A2(new_n872), .ZN(new_n996));
  NAND4_X1  g810(.A1(new_n785), .A2(new_n386), .A3(new_n706), .A4(new_n996), .ZN(new_n997));
  XOR2_X1   g811(.A(new_n997), .B(KEYINPUT123), .Z(new_n998));
  AND2_X1   g812(.A1(new_n812), .A2(new_n998), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n994), .A2(new_n816), .A3(new_n995), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n982), .B1(new_n1000), .B2(new_n357), .ZN(new_n1001));
  OAI21_X1  g815(.A(new_n985), .B1(new_n992), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g816(.A(KEYINPUT126), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  OAI211_X1 g818(.A(KEYINPUT126), .B(new_n985), .C1(new_n992), .C2(new_n1001), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(G72));
  NAND2_X1  g820(.A1(G472), .A2(G902), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1007), .B(KEYINPUT63), .Z(new_n1008));
  INV_X1    g822(.A(new_n876), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1008), .B1(new_n1000), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n1010), .A2(new_n520), .A3(new_n516), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n1008), .B1(new_n989), .B2(new_n1009), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1012), .A2(new_n515), .A3(new_n521), .A4(new_n514), .ZN(new_n1013));
  INV_X1    g827(.A(new_n900), .ZN(new_n1014));
  INV_X1    g828(.A(new_n1008), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1015), .B1(new_n694), .B2(new_n522), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT127), .Z(new_n1017));
  AOI21_X1  g831(.A(new_n916), .B1(new_n1014), .B2(new_n1017), .ZN(new_n1018));
  AND3_X1   g832(.A1(new_n1011), .A2(new_n1013), .A3(new_n1018), .ZN(G57));
endmodule


