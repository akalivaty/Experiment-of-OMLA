

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585;

  XOR2_X2 U322 ( .A(n310), .B(n338), .Z(n311) );
  XNOR2_X2 U323 ( .A(KEYINPUT79), .B(n559), .ZN(n570) );
  XNOR2_X2 U324 ( .A(n420), .B(n419), .ZN(n559) );
  NOR2_X1 U325 ( .A1(n427), .A2(n426), .ZN(n428) );
  XNOR2_X1 U326 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U327 ( .A(n401), .B(n400), .Z(n556) );
  XOR2_X1 U328 ( .A(n383), .B(n382), .Z(n562) );
  XNOR2_X1 U329 ( .A(KEYINPUT55), .B(KEYINPUT120), .ZN(n290) );
  XOR2_X1 U330 ( .A(G92GAT), .B(G85GAT), .Z(n291) );
  XNOR2_X1 U331 ( .A(n389), .B(n388), .ZN(n391) );
  INV_X1 U332 ( .A(KEYINPUT24), .ZN(n304) );
  XNOR2_X1 U333 ( .A(n391), .B(n443), .ZN(n392) );
  XNOR2_X1 U334 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n432) );
  NOR2_X1 U335 ( .A1(n535), .A2(n455), .ZN(n456) );
  INV_X1 U336 ( .A(KEYINPUT54), .ZN(n447) );
  XNOR2_X1 U337 ( .A(n433), .B(n432), .ZN(n532) );
  XNOR2_X1 U338 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U339 ( .A(n448), .B(n447), .ZN(n449) );
  OR2_X1 U340 ( .A1(n411), .A2(KEYINPUT75), .ZN(n412) );
  XNOR2_X1 U341 ( .A(n479), .B(n290), .ZN(n480) );
  XNOR2_X1 U342 ( .A(n450), .B(KEYINPUT124), .ZN(n583) );
  NOR2_X1 U343 ( .A1(n565), .A2(n545), .ZN(n543) );
  XOR2_X1 U344 ( .A(n328), .B(n327), .Z(n535) );
  INV_X1 U345 ( .A(G29GAT), .ZN(n474) );
  XNOR2_X1 U346 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n452) );
  XNOR2_X1 U347 ( .A(n482), .B(n481), .ZN(n483) );
  XNOR2_X1 U348 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U349 ( .A(n453), .B(n452), .ZN(G1355GAT) );
  XNOR2_X1 U350 ( .A(n484), .B(n483), .ZN(G1349GAT) );
  XNOR2_X1 U351 ( .A(n477), .B(n476), .ZN(G1328GAT) );
  XOR2_X1 U352 ( .A(KEYINPUT21), .B(KEYINPUT89), .Z(n293) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(KEYINPUT88), .ZN(n292) );
  XNOR2_X1 U354 ( .A(n293), .B(n292), .ZN(n438) );
  XOR2_X1 U355 ( .A(KEYINPUT22), .B(KEYINPUT87), .Z(n295) );
  XNOR2_X1 U356 ( .A(G211GAT), .B(G204GAT), .ZN(n294) );
  XNOR2_X1 U357 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U358 ( .A(KEYINPUT23), .B(G106GAT), .Z(n297) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G78GAT), .Z(n352) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .Z(n397) );
  XNOR2_X1 U361 ( .A(n352), .B(n397), .ZN(n296) );
  XNOR2_X1 U362 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U363 ( .A(n299), .B(n298), .Z(n301) );
  NAND2_X1 U364 ( .A1(G228GAT), .A2(G233GAT), .ZN(n300) );
  XNOR2_X1 U365 ( .A(n301), .B(n300), .ZN(n307) );
  XOR2_X1 U366 ( .A(G162GAT), .B(KEYINPUT74), .Z(n303) );
  XNOR2_X1 U367 ( .A(G50GAT), .B(G218GAT), .ZN(n302) );
  XNOR2_X1 U368 ( .A(n303), .B(n302), .ZN(n414) );
  XNOR2_X1 U369 ( .A(n414), .B(KEYINPUT86), .ZN(n305) );
  XNOR2_X1 U370 ( .A(n438), .B(n308), .ZN(n310) );
  XOR2_X1 U371 ( .A(G141GAT), .B(KEYINPUT3), .Z(n309) );
  XOR2_X1 U372 ( .A(KEYINPUT2), .B(n309), .Z(n338) );
  XOR2_X1 U373 ( .A(G15GAT), .B(G127GAT), .Z(n389) );
  XOR2_X1 U374 ( .A(G120GAT), .B(KEYINPUT0), .Z(n313) );
  XNOR2_X1 U375 ( .A(G113GAT), .B(G134GAT), .ZN(n312) );
  XNOR2_X1 U376 ( .A(n313), .B(n312), .ZN(n339) );
  XOR2_X1 U377 ( .A(n389), .B(n339), .Z(n315) );
  NAND2_X1 U378 ( .A1(G227GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U379 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U380 ( .A(n316), .B(G176GAT), .Z(n320) );
  XOR2_X1 U381 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n318) );
  XNOR2_X1 U382 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n317) );
  XNOR2_X1 U383 ( .A(n318), .B(n317), .ZN(n442) );
  XNOR2_X1 U384 ( .A(n442), .B(KEYINPUT85), .ZN(n319) );
  XNOR2_X1 U385 ( .A(n320), .B(n319), .ZN(n328) );
  XOR2_X1 U386 ( .A(G71GAT), .B(G190GAT), .Z(n322) );
  XNOR2_X1 U387 ( .A(G43GAT), .B(G99GAT), .ZN(n321) );
  XNOR2_X1 U388 ( .A(n322), .B(n321), .ZN(n326) );
  XOR2_X1 U389 ( .A(KEYINPUT84), .B(KEYINPUT83), .Z(n324) );
  XNOR2_X1 U390 ( .A(G183GAT), .B(KEYINPUT20), .ZN(n323) );
  XNOR2_X1 U391 ( .A(n324), .B(n323), .ZN(n325) );
  XOR2_X1 U392 ( .A(n326), .B(n325), .Z(n327) );
  NOR2_X1 U393 ( .A1(n311), .A2(n535), .ZN(n329) );
  XNOR2_X1 U394 ( .A(n329), .B(KEYINPUT26), .ZN(n548) );
  XOR2_X1 U395 ( .A(KEYINPUT4), .B(KEYINPUT6), .Z(n331) );
  XNOR2_X1 U396 ( .A(G1GAT), .B(G57GAT), .ZN(n330) );
  XNOR2_X1 U397 ( .A(n331), .B(n330), .ZN(n347) );
  XOR2_X1 U398 ( .A(G155GAT), .B(G148GAT), .Z(n333) );
  XNOR2_X1 U399 ( .A(G29GAT), .B(G127GAT), .ZN(n332) );
  XNOR2_X1 U400 ( .A(n333), .B(n332), .ZN(n335) );
  XOR2_X1 U401 ( .A(G162GAT), .B(G85GAT), .Z(n334) );
  XNOR2_X1 U402 ( .A(n335), .B(n334), .ZN(n343) );
  XNOR2_X1 U403 ( .A(KEYINPUT5), .B(KEYINPUT1), .ZN(n336) );
  XNOR2_X1 U404 ( .A(n336), .B(KEYINPUT91), .ZN(n337) );
  XOR2_X1 U405 ( .A(n337), .B(KEYINPUT90), .Z(n341) );
  XNOR2_X1 U406 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U408 ( .A(n343), .B(n342), .ZN(n345) );
  NAND2_X1 U409 ( .A1(G225GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U410 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U411 ( .A(n347), .B(n346), .ZN(n522) );
  XNOR2_X1 U412 ( .A(G99GAT), .B(G106GAT), .ZN(n348) );
  XNOR2_X1 U413 ( .A(n291), .B(n348), .ZN(n407) );
  XOR2_X1 U414 ( .A(n407), .B(KEYINPUT32), .Z(n350) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U416 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U417 ( .A(n351), .B(KEYINPUT70), .Z(n354) );
  XNOR2_X1 U418 ( .A(G120GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U419 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U420 ( .A(KEYINPUT71), .B(KEYINPUT31), .Z(n356) );
  XNOR2_X1 U421 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n355) );
  XNOR2_X1 U422 ( .A(n356), .B(n355), .ZN(n357) );
  XNOR2_X1 U423 ( .A(n358), .B(n357), .ZN(n363) );
  XOR2_X1 U424 ( .A(G64GAT), .B(KEYINPUT13), .Z(n360) );
  XNOR2_X1 U425 ( .A(G71GAT), .B(G57GAT), .ZN(n359) );
  XNOR2_X1 U426 ( .A(n360), .B(n359), .ZN(n393) );
  XNOR2_X1 U427 ( .A(G176GAT), .B(G204GAT), .ZN(n361) );
  XNOR2_X1 U428 ( .A(n361), .B(KEYINPUT73), .ZN(n436) );
  XOR2_X1 U429 ( .A(n393), .B(n436), .Z(n362) );
  XNOR2_X1 U430 ( .A(n363), .B(n362), .ZN(n578) );
  XNOR2_X1 U431 ( .A(KEYINPUT41), .B(KEYINPUT64), .ZN(n364) );
  XNOR2_X1 U432 ( .A(n578), .B(n364), .ZN(n552) );
  XOR2_X1 U433 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n366) );
  XNOR2_X1 U434 ( .A(G22GAT), .B(G141GAT), .ZN(n365) );
  XNOR2_X1 U435 ( .A(n366), .B(n365), .ZN(n383) );
  XOR2_X1 U436 ( .A(G1GAT), .B(G8GAT), .Z(n368) );
  XNOR2_X1 U437 ( .A(KEYINPUT30), .B(KEYINPUT66), .ZN(n367) );
  XNOR2_X1 U438 ( .A(n368), .B(n367), .ZN(n376) );
  NAND2_X1 U439 ( .A1(G229GAT), .A2(G233GAT), .ZN(n374) );
  XOR2_X1 U440 ( .A(G197GAT), .B(G113GAT), .Z(n370) );
  XNOR2_X1 U441 ( .A(G169GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U442 ( .A(n370), .B(n369), .ZN(n372) );
  XOR2_X1 U443 ( .A(G50GAT), .B(G36GAT), .Z(n371) );
  XNOR2_X1 U444 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U445 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U446 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U447 ( .A(n377), .B(KEYINPUT67), .Z(n381) );
  XOR2_X1 U448 ( .A(G29GAT), .B(G43GAT), .Z(n379) );
  XNOR2_X1 U449 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n378) );
  XNOR2_X1 U450 ( .A(n379), .B(n378), .ZN(n408) );
  XNOR2_X1 U451 ( .A(n408), .B(KEYINPUT68), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n382) );
  NAND2_X1 U453 ( .A1(n552), .A2(n562), .ZN(n385) );
  XNOR2_X1 U454 ( .A(KEYINPUT46), .B(KEYINPUT112), .ZN(n384) );
  XNOR2_X1 U455 ( .A(n385), .B(n384), .ZN(n402) );
  XOR2_X1 U456 ( .A(KEYINPUT82), .B(KEYINPUT80), .Z(n387) );
  XNOR2_X1 U457 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n386) );
  XNOR2_X1 U458 ( .A(n387), .B(n386), .ZN(n401) );
  AND2_X1 U459 ( .A1(G231GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U460 ( .A(G8GAT), .B(G183GAT), .ZN(n390) );
  XNOR2_X1 U461 ( .A(n390), .B(G211GAT), .ZN(n443) );
  XOR2_X1 U462 ( .A(n392), .B(KEYINPUT12), .Z(n395) );
  XNOR2_X1 U463 ( .A(n393), .B(KEYINPUT81), .ZN(n394) );
  XNOR2_X1 U464 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U465 ( .A(n397), .B(n396), .Z(n399) );
  XNOR2_X1 U466 ( .A(G1GAT), .B(G78GAT), .ZN(n398) );
  XNOR2_X1 U467 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U468 ( .A(n556), .B(KEYINPUT111), .ZN(n565) );
  NAND2_X1 U469 ( .A1(n402), .A2(n565), .ZN(n421) );
  XOR2_X1 U470 ( .A(KEYINPUT65), .B(KEYINPUT9), .Z(n404) );
  NAND2_X1 U471 ( .A1(G232GAT), .A2(G233GAT), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n406) );
  XNOR2_X1 U473 ( .A(G36GAT), .B(G190GAT), .ZN(n405) );
  XNOR2_X1 U474 ( .A(n405), .B(KEYINPUT77), .ZN(n441) );
  XOR2_X1 U475 ( .A(n406), .B(n441), .Z(n410) );
  XNOR2_X1 U476 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U477 ( .A(n410), .B(n409), .ZN(n411) );
  NAND2_X1 U478 ( .A1(n411), .A2(KEYINPUT75), .ZN(n413) );
  NAND2_X1 U479 ( .A1(n413), .A2(n412), .ZN(n416) );
  XOR2_X1 U480 ( .A(n414), .B(KEYINPUT10), .Z(n415) );
  XNOR2_X1 U481 ( .A(n416), .B(n415), .ZN(n420) );
  XOR2_X1 U482 ( .A(KEYINPUT76), .B(KEYINPUT78), .Z(n418) );
  XNOR2_X1 U483 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n417) );
  XNOR2_X1 U484 ( .A(n418), .B(n417), .ZN(n419) );
  NOR2_X1 U485 ( .A1(n421), .A2(n559), .ZN(n422) );
  XNOR2_X1 U486 ( .A(KEYINPUT47), .B(n422), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n570), .B(KEYINPUT99), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n423), .B(KEYINPUT36), .ZN(n471) );
  NAND2_X1 U489 ( .A1(n556), .A2(n471), .ZN(n425) );
  XOR2_X1 U490 ( .A(KEYINPUT45), .B(KEYINPUT113), .Z(n424) );
  XNOR2_X1 U491 ( .A(n425), .B(n424), .ZN(n427) );
  INV_X1 U492 ( .A(n578), .ZN(n426) );
  XNOR2_X1 U493 ( .A(n428), .B(KEYINPUT114), .ZN(n429) );
  INV_X1 U494 ( .A(n562), .ZN(n573) );
  NAND2_X1 U495 ( .A1(n429), .A2(n573), .ZN(n430) );
  NAND2_X1 U496 ( .A1(n431), .A2(n430), .ZN(n433) );
  XOR2_X1 U497 ( .A(G92GAT), .B(G64GAT), .Z(n435) );
  NAND2_X1 U498 ( .A1(G226GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U499 ( .A(n435), .B(n434), .ZN(n437) );
  XOR2_X1 U500 ( .A(n437), .B(n436), .Z(n440) );
  XNOR2_X1 U501 ( .A(n438), .B(G218GAT), .ZN(n439) );
  XNOR2_X1 U502 ( .A(n440), .B(n439), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n444) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n458) );
  NOR2_X1 U506 ( .A1(n532), .A2(n458), .ZN(n448) );
  NOR2_X1 U507 ( .A1(n522), .A2(n449), .ZN(n478) );
  NAND2_X1 U508 ( .A1(n548), .A2(n478), .ZN(n450) );
  INV_X1 U509 ( .A(n583), .ZN(n451) );
  NAND2_X1 U510 ( .A1(n451), .A2(n471), .ZN(n453) );
  XOR2_X1 U511 ( .A(KEYINPUT27), .B(n458), .Z(n457) );
  NAND2_X1 U512 ( .A1(n522), .A2(n457), .ZN(n533) );
  XOR2_X2 U513 ( .A(KEYINPUT28), .B(n311), .Z(n537) );
  NOR2_X1 U514 ( .A1(n533), .A2(n537), .ZN(n454) );
  XOR2_X1 U515 ( .A(KEYINPUT92), .B(n454), .Z(n455) );
  XNOR2_X1 U516 ( .A(n456), .B(KEYINPUT93), .ZN(n467) );
  NAND2_X1 U517 ( .A1(n457), .A2(n548), .ZN(n463) );
  INV_X1 U518 ( .A(n458), .ZN(n524) );
  NAND2_X1 U519 ( .A1(n524), .A2(n535), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n459), .A2(n311), .ZN(n460) );
  XNOR2_X1 U521 ( .A(n460), .B(KEYINPUT94), .ZN(n461) );
  XOR2_X1 U522 ( .A(KEYINPUT25), .B(n461), .Z(n462) );
  NAND2_X1 U523 ( .A1(n463), .A2(n462), .ZN(n465) );
  INV_X1 U524 ( .A(n522), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n465), .A2(n464), .ZN(n466) );
  NAND2_X1 U526 ( .A1(n467), .A2(n466), .ZN(n486) );
  INV_X1 U527 ( .A(n556), .ZN(n582) );
  NAND2_X1 U528 ( .A1(n486), .A2(n582), .ZN(n469) );
  INV_X1 U529 ( .A(KEYINPUT100), .ZN(n468) );
  XNOR2_X1 U530 ( .A(n469), .B(n468), .ZN(n470) );
  AND2_X1 U531 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n472), .B(KEYINPUT37), .ZN(n521) );
  NAND2_X1 U533 ( .A1(n562), .A2(n578), .ZN(n488) );
  NOR2_X1 U534 ( .A1(n521), .A2(n488), .ZN(n473) );
  XNOR2_X2 U535 ( .A(n473), .B(KEYINPUT38), .ZN(n506) );
  AND2_X1 U536 ( .A1(n506), .A2(n522), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT39), .B(KEYINPUT101), .ZN(n475) );
  NAND2_X1 U538 ( .A1(n478), .A2(n311), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n480), .A2(n535), .ZN(n569) );
  INV_X1 U540 ( .A(n569), .ZN(n563) );
  NAND2_X1 U541 ( .A1(n563), .A2(n552), .ZN(n484) );
  XOR2_X1 U542 ( .A(KEYINPUT57), .B(KEYINPUT56), .Z(n482) );
  XOR2_X1 U543 ( .A(G176GAT), .B(KEYINPUT121), .Z(n481) );
  XOR2_X1 U544 ( .A(KEYINPUT34), .B(KEYINPUT96), .Z(n491) );
  NAND2_X1 U545 ( .A1(n570), .A2(n556), .ZN(n485) );
  XOR2_X1 U546 ( .A(KEYINPUT16), .B(n485), .Z(n487) );
  NAND2_X1 U547 ( .A1(n487), .A2(n486), .ZN(n509) );
  NOR2_X1 U548 ( .A1(n488), .A2(n509), .ZN(n489) );
  XOR2_X1 U549 ( .A(KEYINPUT95), .B(n489), .Z(n497) );
  NAND2_X1 U550 ( .A1(n497), .A2(n522), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U552 ( .A(G1GAT), .B(n492), .Z(G1324GAT) );
  NAND2_X1 U553 ( .A1(n497), .A2(n524), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT97), .B(KEYINPUT35), .Z(n495) );
  NAND2_X1 U556 ( .A1(n497), .A2(n535), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n495), .B(n494), .ZN(n496) );
  XOR2_X1 U558 ( .A(G15GAT), .B(n496), .Z(G1326GAT) );
  NAND2_X1 U559 ( .A1(n537), .A2(n497), .ZN(n498) );
  XNOR2_X1 U560 ( .A(n498), .B(KEYINPUT98), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G22GAT), .B(n499), .ZN(G1327GAT) );
  NAND2_X1 U562 ( .A1(n506), .A2(n524), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(KEYINPUT102), .ZN(n501) );
  XNOR2_X1 U564 ( .A(G36GAT), .B(n501), .ZN(G1329GAT) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(KEYINPUT104), .ZN(n505) );
  XOR2_X1 U566 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n503) );
  NAND2_X1 U567 ( .A1(n506), .A2(n535), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(G1330GAT) );
  XOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT105), .Z(n508) );
  NAND2_X1 U571 ( .A1(n537), .A2(n506), .ZN(n507) );
  XNOR2_X1 U572 ( .A(n508), .B(n507), .ZN(G1331GAT) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n511) );
  NAND2_X1 U574 ( .A1(n552), .A2(n573), .ZN(n520) );
  NOR2_X1 U575 ( .A1(n520), .A2(n509), .ZN(n516) );
  NAND2_X1 U576 ( .A1(n516), .A2(n522), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n511), .B(n510), .ZN(n512) );
  XOR2_X1 U578 ( .A(G57GAT), .B(n512), .Z(G1332GAT) );
  XOR2_X1 U579 ( .A(G64GAT), .B(KEYINPUT107), .Z(n514) );
  NAND2_X1 U580 ( .A1(n516), .A2(n524), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n516), .A2(n535), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n515), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U585 ( .A1(n516), .A2(n537), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n519) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n519), .ZN(G1335GAT) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n529) );
  NAND2_X1 U589 ( .A1(n529), .A2(n522), .ZN(n523) );
  XNOR2_X1 U590 ( .A(G85GAT), .B(n523), .ZN(G1336GAT) );
  XOR2_X1 U591 ( .A(G92GAT), .B(KEYINPUT109), .Z(n526) );
  NAND2_X1 U592 ( .A1(n529), .A2(n524), .ZN(n525) );
  XNOR2_X1 U593 ( .A(n526), .B(n525), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n529), .A2(n535), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n527), .B(KEYINPUT110), .ZN(n528) );
  XNOR2_X1 U596 ( .A(G99GAT), .B(n528), .ZN(G1338GAT) );
  NAND2_X1 U597 ( .A1(n537), .A2(n529), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n530), .B(KEYINPUT44), .ZN(n531) );
  XNOR2_X1 U599 ( .A(G106GAT), .B(n531), .ZN(G1339GAT) );
  XOR2_X1 U600 ( .A(G113GAT), .B(KEYINPUT117), .Z(n539) );
  NOR2_X1 U601 ( .A1(n533), .A2(n532), .ZN(n534) );
  XNOR2_X1 U602 ( .A(n534), .B(KEYINPUT116), .ZN(n549) );
  NAND2_X1 U603 ( .A1(n549), .A2(n535), .ZN(n536) );
  NOR2_X1 U604 ( .A1(n537), .A2(n536), .ZN(n542) );
  NAND2_X1 U605 ( .A1(n542), .A2(n562), .ZN(n538) );
  XNOR2_X1 U606 ( .A(n539), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U607 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U608 ( .A1(n542), .A2(n552), .ZN(n540) );
  XNOR2_X1 U609 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  INV_X1 U610 ( .A(n542), .ZN(n545) );
  XOR2_X1 U611 ( .A(KEYINPUT50), .B(n543), .Z(n544) );
  XNOR2_X1 U612 ( .A(G127GAT), .B(n544), .ZN(G1342GAT) );
  NOR2_X1 U613 ( .A1(n570), .A2(n545), .ZN(n547) );
  XNOR2_X1 U614 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U617 ( .A(KEYINPUT118), .B(n550), .Z(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n562), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n551), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U620 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  NAND2_X1 U621 ( .A1(n552), .A2(n560), .ZN(n553) );
  XNOR2_X1 U622 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(G148GAT), .B(n555), .ZN(G1345GAT) );
  XOR2_X1 U624 ( .A(G155GAT), .B(KEYINPUT119), .Z(n558) );
  NAND2_X1 U625 ( .A1(n556), .A2(n560), .ZN(n557) );
  XNOR2_X1 U626 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NAND2_X1 U627 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(n561), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  NOR2_X1 U631 ( .A1(n565), .A2(n569), .ZN(n566) );
  XOR2_X1 U632 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n568) );
  XNOR2_X1 U634 ( .A(G190GAT), .B(KEYINPUT123), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n572) );
  NOR2_X1 U636 ( .A1(n570), .A2(n569), .ZN(n571) );
  XOR2_X1 U637 ( .A(n572), .B(n571), .Z(G1351GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n583), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT60), .B(KEYINPUT125), .Z(n575) );
  XNOR2_X1 U640 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1352GAT) );
  XNOR2_X1 U643 ( .A(KEYINPUT61), .B(KEYINPUT126), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n578), .A2(n583), .ZN(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(G204GAT), .B(n581), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n583), .A2(n582), .ZN(n585) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n584) );
  XNOR2_X1 U649 ( .A(n585), .B(n584), .ZN(G1354GAT) );
endmodule

