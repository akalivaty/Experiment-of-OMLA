//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:21:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n589, new_n590, new_n591, new_n592, new_n593, new_n594, new_n595,
    new_n596, new_n597, new_n599, new_n600, new_n601, new_n602, new_n603,
    new_n604, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n694, new_n695, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n864, new_n865, new_n866, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n888, new_n889, new_n890, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924;
  INV_X1    g000(.A(G125), .ZN(new_n187));
  NOR3_X1   g001(.A1(new_n187), .A2(KEYINPUT16), .A3(G140), .ZN(new_n188));
  XNOR2_X1  g002(.A(G125), .B(G140), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n188), .B1(new_n189), .B2(KEYINPUT16), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n190), .B(G146), .ZN(new_n191));
  INV_X1    g005(.A(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G119), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT73), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(KEYINPUT23), .ZN(new_n196));
  INV_X1    g010(.A(G119), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G128), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT23), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n193), .A2(new_n194), .A3(new_n199), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n196), .A2(new_n198), .A3(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(G110), .ZN(new_n202));
  AND2_X1   g016(.A1(new_n198), .A2(new_n193), .ZN(new_n203));
  XOR2_X1   g017(.A(KEYINPUT24), .B(G110), .Z(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n191), .A2(new_n202), .A3(new_n205), .ZN(new_n206));
  OAI22_X1  g020(.A1(new_n201), .A2(G110), .B1(new_n203), .B2(new_n204), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n190), .A2(G146), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n189), .A2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n207), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n206), .A2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(G953), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(G221), .A3(G234), .ZN(new_n214));
  XNOR2_X1  g028(.A(new_n214), .B(KEYINPUT22), .ZN(new_n215));
  XNOR2_X1  g029(.A(new_n215), .B(G137), .ZN(new_n216));
  XNOR2_X1  g030(.A(new_n212), .B(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G902), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XOR2_X1   g033(.A(new_n219), .B(KEYINPUT25), .Z(new_n220));
  INV_X1    g034(.A(G217), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n221), .B1(G234), .B2(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n222), .A2(G902), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n217), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT32), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT68), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT11), .ZN(new_n230));
  INV_X1    g044(.A(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n230), .B1(new_n231), .B2(G137), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n231), .A2(G137), .ZN(new_n233));
  INV_X1    g047(.A(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n234), .A2(KEYINPUT11), .A3(G134), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(G131), .ZN(new_n237));
  INV_X1    g051(.A(G131), .ZN(new_n238));
  NAND4_X1  g052(.A1(new_n232), .A2(new_n235), .A3(new_n238), .A4(new_n233), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n209), .A2(G143), .ZN(new_n243));
  INV_X1    g057(.A(G143), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G146), .ZN(new_n245));
  AND3_X1   g059(.A1(new_n242), .A2(new_n243), .A3(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT64), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT0), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n247), .A2(new_n248), .A3(new_n192), .ZN(new_n249));
  OAI21_X1  g063(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n250));
  NAND3_X1  g064(.A1(new_n249), .A2(new_n241), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(G143), .B(G146), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n246), .B1(new_n252), .B2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n234), .A2(G134), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n238), .B1(new_n233), .B2(new_n256), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n244), .A2(G128), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n209), .A2(G143), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT1), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(G128), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n209), .A2(new_n258), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n192), .A2(KEYINPUT1), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n253), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(new_n257), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  AOI22_X1  g079(.A1(new_n240), .A2(new_n255), .B1(new_n265), .B2(new_n239), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT66), .A2(G116), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT66), .A2(G116), .ZN(new_n268));
  OAI21_X1  g082(.A(G119), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G116), .ZN(new_n270));
  OR3_X1    g084(.A1(new_n270), .A2(KEYINPUT65), .A3(G119), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT65), .B1(new_n270), .B2(G119), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XNOR2_X1  g087(.A(KEYINPUT2), .B(G113), .ZN(new_n274));
  AND2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n273), .A2(new_n274), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n229), .B1(new_n266), .B2(new_n277), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n273), .B(new_n274), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n253), .A2(new_n242), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n280), .B1(new_n251), .B2(new_n253), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n281), .B1(new_n237), .B2(new_n239), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n233), .A2(new_n256), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(G131), .ZN(new_n284));
  AND3_X1   g098(.A1(new_n263), .A2(new_n243), .A3(new_n245), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n192), .A2(new_n209), .A3(G143), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n286), .B1(new_n263), .B2(new_n245), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n284), .B(new_n239), .C1(new_n285), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n279), .B(KEYINPUT68), .C1(new_n282), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n255), .A2(new_n240), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n262), .A2(new_n264), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT67), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n292), .A2(new_n293), .A3(new_n239), .A4(new_n284), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(KEYINPUT67), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n277), .A2(new_n291), .A3(new_n294), .A4(new_n295), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n278), .A2(new_n290), .A3(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n297), .A2(KEYINPUT28), .ZN(new_n298));
  INV_X1    g112(.A(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT28), .ZN(new_n301));
  INV_X1    g115(.A(new_n266), .ZN(new_n302));
  OAI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n279), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n297), .A2(KEYINPUT69), .A3(KEYINPUT28), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n300), .A2(new_n303), .A3(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(G101), .ZN(new_n307));
  NOR2_X1   g121(.A1(G237), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(G210), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n307), .B(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT31), .ZN(new_n313));
  INV_X1    g127(.A(new_n296), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n291), .A2(new_n295), .A3(new_n294), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT30), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT30), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n266), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n314), .B1(new_n319), .B2(new_n279), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n313), .B1(new_n320), .B2(new_n310), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n277), .B1(new_n316), .B2(new_n318), .ZN(new_n322));
  NOR4_X1   g136(.A1(new_n322), .A2(KEYINPUT31), .A3(new_n311), .A4(new_n314), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n312), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g139(.A1(G472), .A2(G902), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n228), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  AOI211_X1 g142(.A(KEYINPUT70), .B(new_n328), .C1(new_n312), .C2(new_n324), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n227), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n328), .B1(new_n312), .B2(new_n324), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT32), .ZN(new_n332));
  AOI21_X1  g146(.A(KEYINPUT71), .B1(new_n315), .B2(new_n279), .ZN(new_n333));
  XNOR2_X1  g147(.A(new_n333), .B(new_n296), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n303), .B1(new_n334), .B2(new_n301), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n310), .A2(KEYINPUT29), .ZN(new_n336));
  NOR3_X1   g150(.A1(new_n322), .A2(new_n310), .A3(new_n314), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n337), .B1(new_n305), .B2(new_n310), .ZN(new_n338));
  OAI221_X1 g152(.A(new_n218), .B1(new_n335), .B2(new_n336), .C1(new_n338), .C2(KEYINPUT29), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G472), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n330), .A2(new_n332), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT72), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n330), .A2(new_n340), .A3(KEYINPUT72), .A4(new_n332), .ZN(new_n344));
  AOI21_X1  g158(.A(new_n226), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  AND2_X1   g159(.A1(KEYINPUT3), .A2(G107), .ZN(new_n346));
  NOR2_X1   g160(.A1(KEYINPUT3), .A2(G107), .ZN(new_n347));
  AOI21_X1  g161(.A(new_n346), .B1(G104), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT76), .ZN(new_n349));
  XNOR2_X1  g163(.A(KEYINPUT75), .B(G104), .ZN(new_n350));
  OAI211_X1 g164(.A(new_n348), .B(new_n349), .C1(new_n350), .C2(new_n347), .ZN(new_n351));
  INV_X1    g165(.A(G104), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n352), .A2(KEYINPUT75), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT75), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G104), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n347), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT3), .ZN(new_n357));
  INV_X1    g171(.A(G107), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n357), .A2(new_n358), .A3(G104), .ZN(new_n359));
  NAND2_X1  g173(.A1(KEYINPUT3), .A2(G107), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  OAI21_X1  g175(.A(KEYINPUT76), .B1(new_n356), .B2(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n351), .A2(new_n362), .A3(G101), .ZN(new_n363));
  INV_X1    g177(.A(G101), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n348), .B(new_n364), .C1(new_n350), .C2(new_n347), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n363), .A2(KEYINPUT4), .A3(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT4), .ZN(new_n367));
  NAND4_X1  g181(.A1(new_n351), .A2(new_n362), .A3(new_n367), .A4(G101), .ZN(new_n368));
  AND2_X1   g182(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n368), .A2(KEYINPUT77), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n279), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT80), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT78), .ZN(new_n373));
  NOR3_X1   g187(.A1(new_n356), .A2(new_n361), .A3(G101), .ZN(new_n374));
  AOI21_X1  g188(.A(G107), .B1(new_n353), .B2(new_n355), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n352), .A2(new_n358), .ZN(new_n376));
  NOR3_X1   g190(.A1(new_n375), .A2(new_n364), .A3(new_n376), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n373), .B1(new_n374), .B2(new_n377), .ZN(new_n378));
  INV_X1    g192(.A(new_n376), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n379), .B(G101), .C1(new_n350), .C2(G107), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n365), .A2(KEYINPUT78), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(new_n276), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT5), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n384), .A2(new_n197), .A3(G116), .ZN(new_n385));
  OAI211_X1 g199(.A(G113), .B(new_n385), .C1(new_n273), .C2(new_n384), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n382), .A2(new_n383), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n368), .B(KEYINPUT77), .ZN(new_n388));
  INV_X1    g202(.A(KEYINPUT80), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n388), .A2(new_n389), .A3(new_n279), .A4(new_n366), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n372), .A2(new_n387), .A3(new_n390), .ZN(new_n391));
  XOR2_X1   g205(.A(G110), .B(G122), .Z(new_n392));
  NAND2_X1  g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(new_n392), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n372), .A2(new_n390), .A3(new_n394), .A4(new_n387), .ZN(new_n395));
  NAND3_X1  g209(.A1(new_n393), .A2(KEYINPUT6), .A3(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT6), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n391), .A2(new_n397), .A3(new_n392), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n281), .A2(G125), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n399), .B1(G125), .B2(new_n292), .ZN(new_n400));
  INV_X1    g214(.A(G224), .ZN(new_n401));
  NOR2_X1   g215(.A1(new_n401), .A2(G953), .ZN(new_n402));
  XNOR2_X1  g216(.A(new_n402), .B(KEYINPUT81), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n400), .B(new_n403), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n396), .A2(new_n398), .A3(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(G210), .B1(G237), .B2(G902), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT7), .B1(new_n401), .B2(G953), .ZN(new_n407));
  XNOR2_X1  g221(.A(new_n400), .B(new_n407), .ZN(new_n408));
  XOR2_X1   g222(.A(new_n392), .B(KEYINPUT8), .Z(new_n409));
  NAND2_X1  g223(.A1(new_n383), .A2(new_n386), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n365), .A2(new_n380), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n410), .B(new_n411), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n409), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g227(.A(G902), .B1(new_n395), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  AOI21_X1  g230(.A(new_n406), .B1(new_n405), .B2(new_n414), .ZN(new_n417));
  NOR2_X1   g231(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G469), .ZN(new_n419));
  XOR2_X1   g233(.A(G110), .B(G140), .Z(new_n420));
  XNOR2_X1  g234(.A(new_n420), .B(KEYINPUT74), .ZN(new_n421));
  INV_X1    g235(.A(G227), .ZN(new_n422));
  NOR2_X1   g236(.A1(new_n422), .A2(G953), .ZN(new_n423));
  XOR2_X1   g237(.A(new_n421), .B(new_n423), .Z(new_n424));
  OAI211_X1 g238(.A(new_n255), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n425));
  INV_X1    g239(.A(new_n292), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n411), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT10), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n426), .B1(new_n378), .B2(new_n381), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(new_n428), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n432));
  AND3_X1   g246(.A1(new_n425), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n432), .B1(new_n425), .B2(new_n431), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n240), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n240), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n425), .A2(new_n431), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n424), .B1(new_n435), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n424), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n292), .B1(new_n365), .B2(new_n380), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n240), .B1(new_n427), .B2(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n439), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n419), .B(new_n218), .C1(new_n438), .C2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n424), .ZN(new_n445));
  INV_X1    g259(.A(new_n437), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n445), .B1(new_n446), .B2(new_n442), .ZN(new_n447));
  INV_X1    g261(.A(new_n435), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n447), .B(G469), .C1(new_n448), .C2(new_n439), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n419), .A2(new_n218), .ZN(new_n450));
  INV_X1    g264(.A(new_n450), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n444), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT9), .B(G234), .Z(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G221), .B1(new_n454), .B2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G214), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NOR3_X1   g272(.A1(new_n418), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  XOR2_X1   g273(.A(KEYINPUT89), .B(KEYINPUT13), .Z(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(G128), .A3(new_n244), .ZN(new_n461));
  XOR2_X1   g275(.A(G128), .B(G143), .Z(new_n462));
  OAI211_X1 g276(.A(new_n461), .B(G134), .C1(new_n462), .C2(new_n460), .ZN(new_n463));
  OAI21_X1  g277(.A(G122), .B1(new_n267), .B2(new_n268), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n270), .A2(G122), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n358), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n358), .A3(new_n465), .ZN(new_n467));
  INV_X1    g281(.A(new_n467), .ZN(new_n468));
  OAI221_X1 g282(.A(new_n463), .B1(G134), .B2(new_n462), .C1(new_n466), .C2(new_n468), .ZN(new_n469));
  OR2_X1    g283(.A1(new_n464), .A2(KEYINPUT14), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n270), .A2(G122), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n471), .B1(new_n464), .B2(KEYINPUT14), .ZN(new_n472));
  AND3_X1   g286(.A1(new_n470), .A2(KEYINPUT90), .A3(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G107), .B1(new_n472), .B2(KEYINPUT90), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n462), .B(new_n231), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n469), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n454), .A2(new_n221), .A3(G953), .ZN(new_n478));
  XOR2_X1   g292(.A(new_n477), .B(new_n478), .Z(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(new_n218), .ZN(new_n480));
  INV_X1    g294(.A(G478), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n481), .A2(KEYINPUT15), .ZN(new_n482));
  XNOR2_X1  g296(.A(new_n480), .B(new_n482), .ZN(new_n483));
  XOR2_X1   g297(.A(KEYINPUT87), .B(G475), .Z(new_n484));
  NAND3_X1  g298(.A1(new_n308), .A2(G143), .A3(G214), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  AOI21_X1  g300(.A(G143), .B1(new_n308), .B2(G214), .ZN(new_n487));
  OAI21_X1  g301(.A(G131), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT17), .ZN(new_n489));
  INV_X1    g303(.A(G237), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n213), .A3(G214), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(new_n244), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n492), .A2(new_n238), .A3(new_n485), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n488), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT85), .ZN(new_n495));
  OR2_X1    g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n495), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n492), .A2(new_n485), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n499), .A2(KEYINPUT17), .A3(G131), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(KEYINPUT84), .ZN(new_n501));
  INV_X1    g315(.A(new_n191), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n498), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XOR2_X1   g317(.A(G113), .B(G122), .Z(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(KEYINPUT83), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n352), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n499), .A2(KEYINPUT18), .A3(G131), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n189), .B(new_n209), .ZN(new_n508));
  NAND2_X1  g322(.A1(KEYINPUT18), .A2(G131), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n492), .A2(new_n485), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n507), .A2(new_n508), .A3(new_n510), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n503), .A2(new_n506), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT86), .ZN(new_n513));
  INV_X1    g327(.A(new_n511), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n191), .B1(new_n496), .B2(new_n497), .ZN(new_n515));
  AOI21_X1  g329(.A(new_n514), .B1(new_n515), .B2(new_n501), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT86), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n516), .A2(new_n517), .A3(new_n506), .ZN(new_n518));
  AND2_X1   g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n516), .ZN(new_n520));
  INV_X1    g334(.A(new_n506), .ZN(new_n521));
  NAND3_X1  g335(.A1(new_n520), .A2(KEYINPUT88), .A3(new_n521), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT88), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n516), .B2(new_n506), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n522), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n218), .B1(new_n519), .B2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n483), .B1(new_n484), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n488), .A2(new_n493), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n189), .B(KEYINPUT19), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI211_X1 g344(.A(new_n208), .B(new_n528), .C1(new_n530), .C2(G146), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n511), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n513), .A2(new_n518), .B1(new_n521), .B2(new_n532), .ZN(new_n533));
  NOR4_X1   g347(.A1(new_n533), .A2(KEYINPUT20), .A3(G475), .A4(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n513), .A2(new_n518), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n521), .A2(new_n532), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  INV_X1    g352(.A(G475), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n538), .A2(new_n539), .A3(new_n218), .ZN(new_n540));
  XNOR2_X1  g354(.A(KEYINPUT82), .B(KEYINPUT20), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n535), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(G952), .ZN(new_n544));
  AOI211_X1 g358(.A(G953), .B(new_n544), .C1(G234), .C2(G237), .ZN(new_n545));
  XNOR2_X1  g359(.A(KEYINPUT21), .B(G898), .ZN(new_n546));
  XNOR2_X1  g360(.A(new_n546), .B(KEYINPUT91), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  AOI211_X1 g362(.A(new_n218), .B(new_n213), .C1(G234), .C2(G237), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n545), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n527), .A2(new_n543), .A3(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(new_n459), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n345), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(new_n554), .B(G101), .ZN(G3));
  OR2_X1    g369(.A1(new_n327), .A2(new_n329), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n223), .A2(new_n225), .A3(new_n455), .ZN(new_n557));
  INV_X1    g371(.A(new_n325), .ZN(new_n558));
  OAI21_X1  g372(.A(G472), .B1(new_n558), .B2(G902), .ZN(new_n559));
  AND4_X1   g373(.A1(new_n556), .A2(new_n557), .A3(new_n452), .A4(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n560), .B(KEYINPUT92), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n457), .B(new_n551), .C1(new_n416), .C2(new_n417), .ZN(new_n562));
  NAND2_X1  g376(.A1(new_n526), .A2(new_n484), .ZN(new_n563));
  INV_X1    g377(.A(new_n541), .ZN(new_n564));
  AOI21_X1  g378(.A(G475), .B1(new_n536), .B2(new_n537), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n564), .B1(new_n565), .B2(new_n218), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n563), .B1(new_n566), .B2(new_n534), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n479), .B(KEYINPUT33), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n568), .A2(G478), .A3(new_n218), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT93), .B(G478), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n480), .A2(new_n570), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n567), .A2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n562), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n561), .A2(new_n574), .ZN(new_n575));
  XOR2_X1   g389(.A(KEYINPUT34), .B(G104), .Z(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(G6));
  NOR3_X1   g391(.A1(new_n533), .A2(G475), .A3(G902), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(new_n564), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n542), .A3(KEYINPUT94), .ZN(new_n580));
  OR3_X1    g394(.A1(new_n540), .A2(KEYINPUT94), .A3(new_n541), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n563), .A2(new_n483), .ZN(new_n583));
  OR2_X1    g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(new_n562), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n561), .A2(new_n585), .ZN(new_n586));
  XOR2_X1   g400(.A(KEYINPUT35), .B(G107), .Z(new_n587));
  XNOR2_X1  g401(.A(new_n586), .B(new_n587), .ZN(G9));
  AND2_X1   g402(.A1(new_n556), .A2(new_n559), .ZN(new_n589));
  INV_X1    g403(.A(new_n216), .ZN(new_n590));
  NOR2_X1   g404(.A1(new_n590), .A2(KEYINPUT36), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(new_n212), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n224), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n223), .A2(new_n593), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n459), .A2(new_n552), .A3(new_n589), .A4(new_n594), .ZN(new_n595));
  XNOR2_X1  g409(.A(new_n595), .B(KEYINPUT95), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT37), .B(G110), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n596), .B(new_n597), .ZN(G12));
  INV_X1    g412(.A(new_n594), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n599), .B1(new_n343), .B2(new_n344), .ZN(new_n600));
  INV_X1    g414(.A(G900), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n545), .B1(new_n549), .B2(new_n601), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n584), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n600), .A2(new_n459), .A3(new_n603), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n604), .B(G128), .ZN(G30));
  NAND2_X1  g419(.A1(new_n405), .A2(new_n414), .ZN(new_n606));
  INV_X1    g420(.A(new_n406), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n608), .A2(new_n415), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT38), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n567), .A2(new_n457), .A3(new_n483), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n334), .A2(new_n311), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n218), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n320), .A2(new_n311), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n330), .A2(new_n332), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT96), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND4_X1  g434(.A1(new_n330), .A2(KEYINPUT96), .A3(new_n332), .A4(new_n617), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n602), .B(KEYINPUT39), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n456), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(KEYINPUT40), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n613), .A2(new_n599), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G143), .ZN(G45));
  NAND2_X1  g441(.A1(new_n343), .A2(new_n344), .ZN(new_n628));
  INV_X1    g442(.A(new_n602), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n567), .A2(new_n572), .A3(new_n629), .ZN(new_n630));
  INV_X1    g444(.A(new_n630), .ZN(new_n631));
  NAND4_X1  g445(.A1(new_n628), .A2(new_n459), .A3(new_n594), .A4(new_n631), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT97), .B(G146), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G48));
  OAI21_X1  g448(.A(new_n218), .B1(new_n438), .B2(new_n443), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n635), .A2(G469), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n636), .A2(new_n455), .A3(new_n444), .ZN(new_n637));
  INV_X1    g451(.A(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n636), .A2(KEYINPUT98), .A3(new_n455), .A4(new_n444), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(KEYINPUT99), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT99), .ZN(new_n643));
  NAND3_X1  g457(.A1(new_n639), .A2(new_n643), .A3(new_n640), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n345), .A3(new_n574), .ZN(new_n646));
  XNOR2_X1  g460(.A(KEYINPUT41), .B(G113), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G15));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n345), .A3(new_n585), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(G116), .ZN(G18));
  AOI21_X1  g464(.A(new_n458), .B1(new_n608), .B2(new_n415), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n641), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n600), .A2(new_n552), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G119), .ZN(G21));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n559), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n226), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n335), .A2(new_n311), .ZN(new_n659));
  INV_X1    g473(.A(new_n324), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n326), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI211_X1 g475(.A(KEYINPUT100), .B(G472), .C1(new_n558), .C2(G902), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n657), .A2(new_n658), .A3(new_n661), .A4(new_n662), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n663), .A2(new_n550), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n612), .A2(new_n418), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n645), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(G122), .ZN(G24));
  NAND4_X1  g482(.A1(new_n657), .A2(new_n594), .A3(new_n661), .A4(new_n662), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n641), .A2(new_n669), .A3(new_n652), .A4(new_n630), .ZN(new_n670));
  XNOR2_X1  g484(.A(new_n670), .B(new_n187), .ZN(G27));
  INV_X1    g485(.A(new_n455), .ZN(new_n672));
  AND2_X1   g486(.A1(new_n444), .A2(new_n451), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT102), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n449), .A2(new_n674), .ZN(new_n675));
  NAND3_X1  g489(.A1(new_n435), .A2(new_n437), .A3(new_n424), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n676), .A2(KEYINPUT102), .A3(G469), .A4(new_n447), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n673), .A2(KEYINPUT103), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  NAND4_X1  g492(.A1(new_n675), .A2(new_n444), .A3(new_n451), .A4(new_n677), .ZN(new_n679));
  INV_X1    g493(.A(KEYINPUT103), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(new_n672), .B1(new_n678), .B2(new_n681), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n630), .A2(new_n458), .A3(new_n609), .ZN(new_n683));
  AND2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT42), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n684), .A2(new_n345), .A3(new_n685), .ZN(new_n686));
  AOI22_X1  g500(.A1(new_n339), .A2(G472), .B1(KEYINPUT32), .B2(new_n331), .ZN(new_n687));
  OR2_X1    g501(.A1(new_n331), .A2(KEYINPUT32), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n226), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n682), .A2(new_n683), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(KEYINPUT42), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n686), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n238), .ZN(G33));
  NOR2_X1   g507(.A1(new_n609), .A2(new_n458), .ZN(new_n694));
  NAND4_X1  g508(.A1(new_n345), .A2(new_n603), .A3(new_n694), .A4(new_n682), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G134), .ZN(G36));
  NAND2_X1  g510(.A1(new_n418), .A2(new_n457), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n676), .A2(new_n447), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(G469), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n700), .A2(KEYINPUT46), .A3(new_n451), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT46), .ZN(new_n702));
  OAI211_X1 g516(.A(new_n702), .B(G469), .C1(new_n699), .C2(G902), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n701), .A2(new_n444), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n455), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n623), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT44), .ZN(new_n707));
  INV_X1    g521(.A(KEYINPUT43), .ZN(new_n708));
  INV_X1    g522(.A(new_n572), .ZN(new_n709));
  OAI21_X1  g523(.A(new_n708), .B1(new_n709), .B2(new_n567), .ZN(new_n710));
  INV_X1    g524(.A(new_n567), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n711), .A2(KEYINPUT43), .A3(new_n572), .ZN(new_n712));
  AOI21_X1  g526(.A(new_n589), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n594), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n706), .B1(new_n707), .B2(new_n714), .ZN(new_n715));
  AOI211_X1 g529(.A(new_n697), .B(new_n715), .C1(new_n707), .C2(new_n714), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT104), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(new_n234), .ZN(G39));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT47), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  AND2_X1   g535(.A1(new_n705), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n719), .A2(new_n720), .ZN(new_n723));
  AOI21_X1  g537(.A(new_n721), .B1(new_n705), .B2(new_n723), .ZN(new_n724));
  NOR2_X1   g538(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n628), .A2(new_n658), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n725), .A2(new_n683), .A3(new_n726), .ZN(new_n727));
  OR2_X1    g541(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n730), .B(G140), .ZN(G42));
  NAND2_X1  g545(.A1(new_n636), .A2(new_n444), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n622), .B1(KEYINPUT49), .B2(new_n732), .ZN(new_n733));
  NAND4_X1  g547(.A1(new_n711), .A2(new_n557), .A3(new_n457), .A4(new_n572), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT107), .Z(new_n735));
  NOR2_X1   g549(.A1(new_n732), .A2(KEYINPUT49), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(KEYINPUT108), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n733), .A2(new_n735), .A3(new_n611), .A4(new_n737), .ZN(new_n738));
  INV_X1    g552(.A(new_n725), .ZN(new_n739));
  XOR2_X1   g553(.A(new_n732), .B(KEYINPUT114), .Z(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n672), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n545), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n743), .B(new_n663), .C1(new_n710), .C2(new_n712), .ZN(new_n744));
  AND3_X1   g558(.A1(new_n742), .A2(new_n694), .A3(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(new_n641), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n610), .A2(new_n457), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n744), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  XOR2_X1   g562(.A(new_n748), .B(KEYINPUT50), .Z(new_n749));
  NOR2_X1   g563(.A1(new_n641), .A2(new_n697), .ZN(new_n750));
  AOI21_X1  g564(.A(new_n743), .B1(new_n712), .B2(new_n710), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n752), .A2(new_n669), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(KEYINPUT115), .ZN(new_n754));
  INV_X1    g568(.A(new_n622), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n658), .A3(new_n750), .A4(new_n545), .ZN(new_n756));
  OR3_X1    g570(.A1(new_n756), .A2(new_n567), .A3(new_n572), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n749), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n745), .A2(new_n758), .ZN(new_n759));
  OAI211_X1 g573(.A(G952), .B(new_n213), .C1(new_n759), .C2(KEYINPUT51), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n742), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n739), .A2(KEYINPUT116), .A3(new_n741), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n762), .A2(new_n694), .A3(new_n744), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n764), .A2(KEYINPUT51), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n765), .A2(new_n758), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n760), .A2(new_n766), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n609), .A2(new_n455), .A3(new_n452), .A4(new_n457), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n768), .B(new_n599), .C1(new_n343), .C2(new_n344), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n670), .B1(new_n769), .B2(new_n603), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n612), .A2(new_n418), .A3(new_n602), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n622), .A2(new_n599), .A3(new_n682), .A4(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n770), .A2(KEYINPUT52), .A3(new_n632), .A4(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n669), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n653), .A2(new_n631), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n604), .A2(new_n632), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(KEYINPUT52), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT111), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n773), .A2(new_n778), .A3(new_n779), .ZN(new_n780));
  OR3_X1    g594(.A1(new_n776), .A2(new_n779), .A3(new_n777), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n543), .A2(new_n483), .A3(new_n563), .ZN(new_n783));
  OAI21_X1  g597(.A(KEYINPUT109), .B1(new_n562), .B2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n583), .B1(new_n542), .B2(new_n535), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT109), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n785), .A2(new_n651), .A3(new_n786), .A4(new_n551), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n784), .A2(new_n787), .A3(new_n560), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n788), .A2(new_n595), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT110), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI22_X1  g605(.A1(new_n345), .A2(new_n553), .B1(new_n574), .B2(new_n560), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n788), .A2(new_n595), .A3(KEYINPUT110), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n791), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n646), .A2(new_n649), .A3(new_n666), .A4(new_n654), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n695), .A2(new_n686), .A3(new_n691), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  NOR3_X1   g612(.A1(new_n582), .A2(new_n456), .A3(new_n602), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n600), .A2(new_n527), .A3(new_n694), .A4(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n684), .A2(new_n774), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n796), .A2(new_n798), .A3(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n782), .A2(new_n804), .A3(KEYINPUT53), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n773), .A2(new_n778), .ZN(new_n806));
  OR2_X1    g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n805), .B1(KEYINPUT53), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT54), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n744), .A2(new_n653), .ZN(new_n810));
  AND2_X1   g624(.A1(new_n646), .A2(new_n666), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n649), .A2(new_n654), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n811), .A2(new_n812), .A3(KEYINPUT112), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n795), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT53), .A3(new_n815), .ZN(new_n816));
  OR3_X1    g630(.A1(new_n794), .A2(new_n797), .A3(new_n802), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  AND2_X1   g632(.A1(new_n780), .A2(new_n781), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT113), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT113), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n794), .A2(new_n797), .A3(new_n802), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n822), .A2(KEYINPUT53), .A3(new_n815), .A4(new_n813), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n821), .B1(new_n823), .B2(new_n782), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT54), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n826));
  OAI21_X1  g640(.A(new_n826), .B1(new_n804), .B2(new_n806), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n820), .A2(new_n824), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n767), .A2(new_n809), .A3(new_n810), .A4(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n756), .A2(new_n573), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n750), .A2(new_n751), .A3(new_n689), .ZN(new_n831));
  XOR2_X1   g645(.A(new_n831), .B(KEYINPUT48), .Z(new_n832));
  NOR3_X1   g646(.A1(new_n829), .A2(new_n830), .A3(new_n832), .ZN(new_n833));
  NOR2_X1   g647(.A1(G952), .A2(G953), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(KEYINPUT117), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n738), .B1(new_n833), .B2(new_n835), .ZN(G75));
  NAND3_X1  g650(.A1(new_n820), .A2(new_n827), .A3(new_n824), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(G210), .A3(G902), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT56), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n396), .A2(new_n398), .ZN(new_n841));
  XNOR2_X1  g655(.A(new_n841), .B(new_n404), .ZN(new_n842));
  XNOR2_X1  g656(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n843));
  XOR2_X1   g657(.A(new_n842), .B(new_n843), .Z(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n213), .A2(G952), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(new_n844), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n838), .A2(new_n839), .A3(new_n848), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n845), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n845), .A2(KEYINPUT119), .A3(new_n847), .A4(new_n849), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(G51));
  NAND2_X1  g668(.A1(new_n837), .A2(KEYINPUT54), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n855), .A2(new_n828), .ZN(new_n856));
  XOR2_X1   g670(.A(KEYINPUT120), .B(KEYINPUT57), .Z(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n450), .ZN(new_n858));
  OR2_X1    g672(.A1(new_n857), .A2(new_n450), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  OAI21_X1  g674(.A(new_n860), .B1(new_n438), .B2(new_n443), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n837), .A2(G469), .A3(G902), .A4(new_n699), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n846), .B1(new_n861), .B2(new_n862), .ZN(G54));
  NAND4_X1  g677(.A1(new_n837), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT121), .ZN(new_n865));
  OR3_X1    g679(.A1(new_n864), .A2(new_n865), .A3(new_n533), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n846), .B1(new_n864), .B2(new_n533), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n865), .B1(new_n864), .B2(new_n533), .ZN(new_n868));
  AND3_X1   g682(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G60));
  NAND2_X1  g683(.A1(G478), .A2(G902), .ZN(new_n870));
  XOR2_X1   g684(.A(new_n870), .B(KEYINPUT59), .Z(new_n871));
  AOI21_X1  g685(.A(new_n871), .B1(new_n809), .B2(new_n828), .ZN(new_n872));
  OAI21_X1  g686(.A(new_n847), .B1(new_n872), .B2(new_n568), .ZN(new_n873));
  INV_X1    g687(.A(new_n871), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n568), .A2(new_n874), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n873), .B1(new_n856), .B2(new_n875), .ZN(G63));
  NAND2_X1  g690(.A1(G217), .A2(G902), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT122), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT60), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n837), .A2(new_n592), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n847), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n217), .B1(new_n837), .B2(new_n879), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT123), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT61), .ZN(new_n884));
  OAI22_X1  g698(.A1(new_n881), .A2(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  XNOR2_X1  g700(.A(new_n885), .B(new_n886), .ZN(G66));
  OAI21_X1  g701(.A(G953), .B1(new_n548), .B2(new_n401), .ZN(new_n888));
  OAI21_X1  g702(.A(new_n888), .B1(new_n796), .B2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n841), .B1(G898), .B2(new_n213), .ZN(new_n890));
  XNOR2_X1  g704(.A(new_n889), .B(new_n890), .ZN(G69));
  AOI21_X1  g705(.A(new_n716), .B1(new_n728), .B2(new_n729), .ZN(new_n892));
  AND2_X1   g706(.A1(new_n770), .A2(new_n632), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n706), .A2(new_n665), .A3(new_n689), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n892), .A2(new_n893), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n798), .A2(new_n213), .ZN(new_n896));
  OAI22_X1  g710(.A1(new_n895), .A2(new_n896), .B1(new_n422), .B2(new_n213), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n319), .B(new_n530), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  OAI21_X1  g714(.A(G900), .B1(new_n899), .B2(G227), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n901), .A2(G953), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n893), .A2(new_n626), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT62), .Z(new_n904));
  NAND2_X1  g718(.A1(new_n783), .A2(new_n573), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n345), .A2(new_n624), .A3(new_n694), .A4(new_n905), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n904), .A2(new_n892), .A3(new_n906), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n907), .A2(new_n213), .A3(new_n898), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n900), .A2(new_n902), .A3(new_n908), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n909), .B(KEYINPUT124), .Z(G72));
  NOR2_X1   g724(.A1(new_n616), .A2(new_n337), .ZN(new_n911));
  XOR2_X1   g725(.A(KEYINPUT125), .B(KEYINPUT63), .Z(new_n912));
  NAND2_X1  g726(.A1(G472), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n912), .B(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n915), .B(KEYINPUT126), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n808), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g731(.A(new_n917), .B(KEYINPUT127), .ZN(new_n918));
  INV_X1    g732(.A(new_n796), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n914), .B1(new_n907), .B2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n616), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n796), .A2(new_n798), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n914), .B1(new_n895), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n846), .B1(new_n923), .B2(new_n337), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n918), .A2(new_n921), .A3(new_n924), .ZN(G57));
endmodule


