//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 1 0 1 0 1 0 0 0 0 1 0 1 1 0 0 1 1 1 0 0 0 1 0 1 1 1 1 0 0 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:31 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n774, new_n775, new_n776, new_n777, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n793, new_n794,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n991, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  INV_X1    g000(.A(KEYINPUT11), .ZN(new_n187));
  INV_X1    g001(.A(G134), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G137), .ZN(new_n189));
  INV_X1    g003(.A(G137), .ZN(new_n190));
  NAND3_X1  g004(.A1(new_n190), .A2(KEYINPUT11), .A3(G134), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n188), .A2(G137), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(G131), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  NAND4_X1  g009(.A1(new_n189), .A2(new_n191), .A3(new_n195), .A4(new_n192), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(KEYINPUT80), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT80), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n207), .B(KEYINPUT1), .C1(new_n202), .C2(G146), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n206), .A2(G128), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n201), .A2(new_n203), .ZN(new_n210));
  AOI21_X1  g024(.A(new_n204), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G107), .ZN(new_n213));
  INV_X1    g027(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g028(.A1(new_n212), .A2(G107), .ZN(new_n215));
  OAI21_X1  g029(.A(G101), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT3), .ZN(new_n218));
  INV_X1    g032(.A(G107), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G104), .ZN(new_n220));
  INV_X1    g034(.A(G101), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n217), .A2(new_n220), .A3(new_n221), .A4(new_n213), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n216), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g037(.A(KEYINPUT81), .B1(new_n211), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n208), .A2(G128), .ZN(new_n225));
  AOI21_X1  g039(.A(new_n207), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n226));
  OAI21_X1  g040(.A(new_n210), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n199), .A2(new_n201), .A3(new_n203), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT81), .ZN(new_n230));
  INV_X1    g044(.A(new_n223), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(KEYINPUT10), .B1(new_n224), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n217), .A2(new_n220), .A3(new_n213), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G101), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n235), .A2(KEYINPUT4), .A3(new_n222), .ZN(new_n236));
  XNOR2_X1  g050(.A(KEYINPUT0), .B(G128), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n210), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G143), .B(G146), .ZN(new_n239));
  NAND2_X1  g053(.A1(KEYINPUT0), .A2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n238), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT4), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n234), .A2(new_n243), .A3(G101), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n242), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT1), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n246), .B1(G143), .B2(new_n200), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n210), .B1(new_n247), .B2(new_n198), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(new_n228), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n231), .A2(new_n249), .A3(KEYINPUT10), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n197), .B1(new_n233), .B2(new_n251), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT10), .ZN(new_n253));
  NOR3_X1   g067(.A1(new_n211), .A2(KEYINPUT81), .A3(new_n223), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n230), .B1(new_n229), .B2(new_n231), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n197), .ZN(new_n257));
  INV_X1    g071(.A(new_n251), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT82), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n252), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  XNOR2_X1  g075(.A(G110), .B(G140), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(G227), .ZN(new_n264));
  XOR2_X1   g078(.A(new_n262), .B(new_n264), .Z(new_n265));
  OAI211_X1 g079(.A(KEYINPUT82), .B(new_n197), .C1(new_n233), .C2(new_n251), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n261), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  OAI22_X1  g081(.A1(new_n254), .A2(new_n255), .B1(new_n249), .B2(new_n231), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n268), .A2(KEYINPUT12), .A3(new_n197), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT12), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n231), .A2(new_n249), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n271), .B1(new_n224), .B2(new_n232), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(new_n257), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n269), .A2(new_n273), .A3(KEYINPUT83), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n233), .A2(new_n251), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n265), .B1(new_n275), .B2(new_n257), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT83), .B1(new_n269), .B2(new_n273), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n267), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G469), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT70), .B(G902), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n279), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT84), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n281), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT83), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT12), .B1(new_n268), .B2(new_n197), .ZN(new_n287));
  NOR3_X1   g101(.A1(new_n272), .A2(new_n270), .A3(new_n257), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n274), .A3(new_n276), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n285), .B1(new_n290), .B2(new_n267), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT84), .A3(new_n280), .ZN(new_n292));
  INV_X1    g106(.A(G902), .ZN(new_n293));
  AOI22_X1  g107(.A1(new_n269), .A2(new_n273), .B1(new_n275), .B2(new_n257), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT79), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n265), .B1(new_n294), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n265), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n294), .B2(KEYINPUT79), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n261), .A2(new_n266), .ZN(new_n299));
  OAI211_X1 g113(.A(new_n293), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n300));
  AOI22_X1  g114(.A1(new_n284), .A2(new_n292), .B1(G469), .B2(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(KEYINPUT9), .B(G234), .ZN(new_n302));
  OAI21_X1  g116(.A(G221), .B1(new_n302), .B2(G902), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(G475), .A2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(KEYINPUT75), .A2(G125), .ZN(new_n307));
  INV_X1    g121(.A(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(KEYINPUT75), .A2(G125), .A3(G140), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT16), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(G125), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT16), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT76), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT90), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G143), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n202), .A2(KEYINPUT90), .ZN(new_n320));
  NOR2_X1   g134(.A1(G237), .A2(G953), .ZN(new_n321));
  AOI22_X1  g135(.A1(new_n319), .A2(new_n320), .B1(new_n321), .B2(G214), .ZN(new_n322));
  INV_X1    g136(.A(G237), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n323), .A2(new_n263), .A3(G214), .ZN(new_n324));
  NOR2_X1   g138(.A1(new_n318), .A2(G143), .ZN(new_n325));
  NOR2_X1   g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  OAI21_X1  g140(.A(G131), .B1(new_n322), .B2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(G214), .A3(new_n321), .ZN(new_n328));
  INV_X1    g142(.A(new_n324), .ZN(new_n329));
  XNOR2_X1  g143(.A(KEYINPUT90), .B(G143), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n195), .B(new_n328), .C1(new_n329), .C2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n200), .B1(new_n311), .B2(new_n314), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n309), .A2(KEYINPUT19), .A3(new_n310), .ZN(new_n336));
  INV_X1    g150(.A(G125), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G140), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT19), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n312), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AND2_X1   g154(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n200), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n317), .A2(new_n332), .A3(new_n335), .A4(new_n342), .ZN(new_n343));
  OAI211_X1 g157(.A(KEYINPUT18), .B(G131), .C1(new_n322), .C2(new_n326), .ZN(new_n344));
  NAND2_X1  g158(.A1(KEYINPUT18), .A2(G131), .ZN(new_n345));
  OAI211_X1 g159(.A(new_n328), .B(new_n345), .C1(new_n329), .C2(new_n330), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n309), .A2(G146), .A3(new_n310), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n312), .A2(new_n338), .A3(new_n200), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n344), .A2(new_n346), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n343), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G113), .B(G122), .ZN(new_n352));
  XNOR2_X1  g166(.A(new_n352), .B(new_n212), .ZN(new_n353));
  INV_X1    g167(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n351), .A2(new_n354), .ZN(new_n355));
  INV_X1    g169(.A(KEYINPUT17), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n327), .A2(new_n356), .A3(new_n331), .ZN(new_n357));
  OAI211_X1 g171(.A(KEYINPUT17), .B(G131), .C1(new_n322), .C2(new_n326), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n311), .A2(new_n200), .A3(new_n314), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n316), .A3(new_n359), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n353), .B(new_n350), .C1(new_n357), .C2(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n306), .B1(new_n355), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT20), .ZN(new_n363));
  OAI21_X1  g177(.A(KEYINPUT91), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n361), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n353), .B1(new_n343), .B2(new_n350), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n305), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT91), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT20), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n362), .A2(new_n363), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n364), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n357), .A2(new_n360), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n353), .B1(new_n372), .B2(new_n350), .ZN(new_n373));
  OAI21_X1  g187(.A(new_n293), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G475), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n371), .A2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G122), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(G116), .ZN(new_n379));
  INV_X1    g193(.A(G116), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G122), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n379), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT92), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(G116), .B(G122), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT92), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n219), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n382), .A2(new_n383), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n385), .A2(KEYINPUT92), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n388), .A2(new_n389), .A3(G107), .ZN(new_n390));
  AOI21_X1  g204(.A(KEYINPUT13), .B1(new_n198), .B2(G143), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n188), .ZN(new_n392));
  XNOR2_X1  g206(.A(G128), .B(G143), .ZN(new_n393));
  OR2_X1    g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n393), .ZN(new_n395));
  AOI22_X1  g209(.A1(new_n387), .A2(new_n390), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n380), .A2(KEYINPUT14), .A3(G122), .ZN(new_n397));
  OAI211_X1 g211(.A(G107), .B(new_n397), .C1(new_n382), .C2(KEYINPUT14), .ZN(new_n398));
  OR2_X1    g212(.A1(new_n393), .A2(G134), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n393), .A2(G134), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n402));
  NOR2_X1   g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g217(.A(KEYINPUT93), .B1(new_n396), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n394), .A2(new_n395), .ZN(new_n405));
  INV_X1    g219(.A(new_n390), .ZN(new_n406));
  OAI21_X1  g220(.A(new_n405), .B1(new_n406), .B2(new_n402), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT93), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n387), .A2(new_n398), .A3(new_n399), .A4(new_n400), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n407), .A2(new_n408), .A3(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(G217), .ZN(new_n411));
  NOR3_X1   g225(.A1(new_n302), .A2(new_n411), .A3(G953), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n404), .A2(new_n410), .A3(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT94), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n407), .A2(new_n409), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(KEYINPUT93), .A3(new_n412), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n414), .A2(new_n415), .A3(new_n281), .A4(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G478), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n419), .A2(KEYINPUT15), .ZN(new_n420));
  AND2_X1   g234(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n414), .A2(new_n281), .A3(new_n417), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(KEYINPUT94), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n418), .ZN(new_n424));
  INV_X1    g238(.A(new_n420), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n421), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  AOI211_X1 g240(.A(new_n263), .B(new_n281), .C1(G234), .C2(G237), .ZN(new_n427));
  XNOR2_X1  g241(.A(KEYINPUT21), .B(G898), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G952), .ZN(new_n430));
  AOI211_X1 g244(.A(G953), .B(new_n430), .C1(G234), .C2(G237), .ZN(new_n431));
  NOR2_X1   g245(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n432), .B(KEYINPUT95), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n377), .A2(new_n426), .A3(new_n433), .ZN(new_n434));
  OAI21_X1  g248(.A(G210), .B1(G237), .B2(G902), .ZN(new_n435));
  INV_X1    g249(.A(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(G119), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G116), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n380), .A2(G119), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n438), .A2(new_n439), .A3(KEYINPUT5), .ZN(new_n440));
  OR3_X1    g254(.A1(new_n380), .A2(KEYINPUT5), .A3(G119), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n440), .A2(new_n441), .A3(G113), .ZN(new_n442));
  NAND2_X1  g256(.A1(KEYINPUT2), .A2(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT66), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT66), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n445), .A2(KEYINPUT2), .A3(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OR2_X1    g261(.A1(KEYINPUT2), .A2(G113), .ZN(new_n448));
  XNOR2_X1  g262(.A(G116), .B(G119), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n450), .A3(new_n216), .A4(new_n222), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n236), .A2(new_n244), .ZN(new_n452));
  AND3_X1   g266(.A1(new_n447), .A2(new_n448), .A3(new_n449), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n449), .B1(new_n447), .B2(new_n448), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g269(.A(new_n451), .B1(new_n452), .B2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G110), .B(G122), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n451), .B(new_n457), .C1(new_n452), .C2(new_n455), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT6), .ZN(new_n461));
  NOR2_X1   g275(.A1(new_n461), .A2(KEYINPUT86), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n459), .A2(new_n460), .A3(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n456), .B(new_n458), .C1(KEYINPUT86), .C2(new_n461), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n238), .A2(new_n241), .A3(G125), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n198), .B1(new_n201), .B2(KEYINPUT1), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n228), .B(new_n337), .C1(new_n467), .C2(new_n239), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT87), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g284(.A1(new_n248), .A2(KEYINPUT87), .A3(new_n337), .A4(new_n228), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n466), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n263), .A2(G224), .ZN(new_n473));
  XNOR2_X1  g287(.A(new_n472), .B(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n463), .A2(new_n464), .A3(new_n474), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n457), .B(KEYINPUT8), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n442), .A2(new_n450), .B1(new_n216), .B2(new_n222), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n477), .B1(new_n478), .B2(new_n451), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n442), .A2(new_n450), .ZN(new_n480));
  NAND3_X1  g294(.A1(new_n480), .A2(new_n478), .A3(new_n223), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  OAI21_X1  g296(.A(new_n476), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n470), .A2(new_n471), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n473), .A2(KEYINPUT7), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n465), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(new_n460), .A3(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n466), .B1(new_n484), .B2(KEYINPUT89), .ZN(new_n489));
  INV_X1    g303(.A(KEYINPUT89), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n470), .A2(new_n490), .A3(new_n471), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n486), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n293), .B1(new_n488), .B2(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n436), .B1(new_n475), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n460), .A2(new_n487), .ZN(new_n495));
  INV_X1    g309(.A(new_n476), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n451), .A2(new_n478), .ZN(new_n497));
  INV_X1    g311(.A(new_n477), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n496), .B1(new_n499), .B2(new_n481), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(new_n492), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n463), .A2(new_n464), .A3(new_n474), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n503), .A2(new_n435), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n494), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(G214), .B1(G237), .B2(G902), .ZN(new_n507));
  XOR2_X1   g321(.A(new_n507), .B(KEYINPUT85), .Z(new_n508));
  INV_X1    g322(.A(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n506), .A2(new_n509), .ZN(new_n510));
  NOR4_X1   g324(.A1(new_n301), .A2(new_n304), .A3(new_n434), .A4(new_n510), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n321), .A2(G210), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT27), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT26), .B(G101), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n197), .A2(new_n242), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n188), .A2(G137), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n190), .A2(G134), .ZN(new_n519));
  OAI21_X1  g333(.A(G131), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n196), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n249), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n517), .A2(new_n522), .A3(new_n455), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT65), .ZN(new_n525));
  AOI22_X1  g339(.A1(new_n197), .A2(new_n242), .B1(new_n521), .B2(new_n249), .ZN(new_n526));
  XOR2_X1   g340(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(new_n454), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(new_n450), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n526), .A2(KEYINPUT30), .ZN(new_n531));
  INV_X1    g345(.A(new_n527), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n205), .A2(G128), .B1(new_n201), .B2(new_n203), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n533), .A2(new_n204), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n196), .A2(new_n520), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  AOI22_X1  g350(.A1(new_n194), .A2(new_n196), .B1(new_n238), .B2(new_n241), .ZN(new_n537));
  OAI211_X1 g351(.A(KEYINPUT65), .B(new_n532), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND4_X1  g352(.A1(new_n528), .A2(new_n530), .A3(new_n531), .A4(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT67), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n527), .B1(new_n517), .B2(new_n522), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n541), .A2(KEYINPUT65), .B1(KEYINPUT30), .B2(new_n526), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT67), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n542), .A2(new_n543), .A3(new_n530), .A4(new_n528), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n516), .B(new_n524), .C1(new_n540), .C2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT28), .ZN(new_n546));
  OAI21_X1  g360(.A(new_n530), .B1(new_n536), .B2(new_n537), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n546), .B1(new_n547), .B2(new_n523), .ZN(new_n548));
  OAI21_X1  g362(.A(KEYINPUT68), .B1(new_n536), .B2(new_n537), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT68), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n517), .A2(new_n522), .A3(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n549), .A2(new_n551), .A3(new_n455), .ZN(new_n552));
  AOI21_X1  g366(.A(new_n548), .B1(new_n546), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n516), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n512), .B1(new_n545), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g370(.A1(new_n554), .A2(new_n512), .ZN(new_n557));
  AOI21_X1  g371(.A(KEYINPUT69), .B1(new_n553), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n552), .A2(new_n546), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n455), .B1(new_n517), .B2(new_n522), .ZN(new_n560));
  OAI21_X1  g374(.A(KEYINPUT28), .B1(new_n524), .B2(new_n560), .ZN(new_n561));
  AND4_X1   g375(.A1(KEYINPUT69), .A2(new_n559), .A3(new_n561), .A4(new_n557), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n281), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT71), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT71), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n565), .B(new_n281), .C1(new_n558), .C2(new_n562), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n556), .A2(new_n564), .A3(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n567), .A2(G472), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT31), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n540), .A2(new_n544), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n523), .A2(new_n516), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n569), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  AOI211_X1 g387(.A(KEYINPUT31), .B(new_n571), .C1(new_n540), .C2(new_n544), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n553), .A2(new_n516), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n573), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  NOR2_X1   g390(.A1(G472), .A2(G902), .ZN(new_n577));
  INV_X1    g391(.A(new_n577), .ZN(new_n578));
  NOR3_X1   g392(.A1(new_n576), .A2(KEYINPUT32), .A3(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT32), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n570), .A2(new_n572), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(KEYINPUT31), .ZN(new_n582));
  INV_X1    g396(.A(new_n575), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n570), .A2(new_n569), .A3(new_n572), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n580), .B1(new_n585), .B2(new_n577), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n568), .B1(new_n579), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT72), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n437), .A2(G128), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n198), .A2(G119), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT73), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n590), .A2(new_n591), .A3(KEYINPUT73), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  XNOR2_X1  g410(.A(KEYINPUT24), .B(G110), .ZN(new_n597));
  OR2_X1    g411(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g412(.A1(new_n590), .A2(KEYINPUT23), .ZN(new_n599));
  AOI21_X1  g413(.A(KEYINPUT74), .B1(new_n198), .B2(G119), .ZN(new_n600));
  OR2_X1    g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n599), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G110), .ZN(new_n604));
  INV_X1    g418(.A(new_n359), .ZN(new_n605));
  OAI211_X1 g419(.A(new_n598), .B(new_n604), .C1(new_n333), .C2(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n348), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n596), .A2(new_n597), .ZN(new_n609));
  INV_X1    g423(.A(G110), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n601), .A2(new_n602), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n608), .B1(new_n609), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n333), .A2(new_n334), .ZN(new_n613));
  AOI211_X1 g427(.A(KEYINPUT76), .B(new_n200), .C1(new_n311), .C2(new_n314), .ZN(new_n614));
  NOR2_X1   g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT77), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g432(.A1(new_n612), .A2(new_n615), .A3(KEYINPUT77), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n607), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n263), .A2(G221), .A3(G234), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(KEYINPUT78), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT22), .B(G137), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n620), .B(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n411), .B1(new_n281), .B2(G234), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n626), .A2(G902), .ZN(new_n627));
  INV_X1    g441(.A(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT25), .ZN(new_n630));
  OAI21_X1  g444(.A(new_n630), .B1(new_n625), .B2(new_n285), .ZN(new_n631));
  INV_X1    g445(.A(new_n624), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n620), .B(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n633), .A2(KEYINPUT25), .A3(new_n281), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  AOI21_X1  g449(.A(new_n629), .B1(new_n635), .B2(new_n626), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT32), .B1(new_n576), .B2(new_n578), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n585), .A2(new_n580), .A3(new_n577), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n639), .A2(KEYINPUT72), .A3(new_n568), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n511), .A2(new_n589), .A3(new_n636), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(G101), .ZN(G3));
  NAND2_X1  g456(.A1(new_n300), .A2(G469), .ZN(new_n643));
  AND4_X1   g457(.A1(KEYINPUT84), .A2(new_n279), .A3(new_n280), .A4(new_n281), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT84), .B1(new_n291), .B2(new_n280), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n303), .ZN(new_n647));
  OAI21_X1  g461(.A(G472), .B1(new_n576), .B2(new_n285), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n636), .B(new_n648), .C1(new_n578), .C2(new_n576), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT96), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n284), .A2(new_n292), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n304), .B1(new_n651), .B2(new_n643), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT96), .ZN(new_n653));
  INV_X1    g467(.A(G472), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n654), .B1(new_n585), .B2(new_n281), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n577), .B2(new_n585), .ZN(new_n656));
  NAND4_X1  g470(.A1(new_n652), .A2(new_n653), .A3(new_n656), .A4(new_n636), .ZN(new_n657));
  AND2_X1   g471(.A1(new_n650), .A2(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(KEYINPUT97), .ZN(new_n659));
  OAI211_X1 g473(.A(new_n659), .B(new_n436), .C1(new_n475), .C2(new_n493), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n507), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n475), .A2(new_n493), .A3(new_n436), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n435), .B1(new_n503), .B2(new_n504), .ZN(new_n663));
  NOR2_X1   g477(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n661), .B1(new_n664), .B2(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n422), .A2(new_n419), .ZN(new_n666));
  AOI21_X1  g480(.A(KEYINPUT33), .B1(new_n414), .B2(new_n417), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n416), .A2(KEYINPUT98), .A3(new_n413), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n413), .A2(KEYINPUT98), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n407), .A2(new_n409), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n668), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n667), .B1(KEYINPUT33), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n281), .A2(G478), .ZN(new_n673));
  OAI21_X1  g487(.A(new_n666), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n376), .A2(new_n674), .A3(new_n433), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n658), .A2(new_n665), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT34), .B(G104), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n677), .B(new_n678), .ZN(G6));
  AOI22_X1  g493(.A1(new_n327), .A2(new_n331), .B1(new_n341), .B2(new_n200), .ZN(new_n680));
  AND2_X1   g494(.A1(new_n346), .A2(new_n349), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n615), .A2(new_n680), .B1(new_n344), .B2(new_n681), .ZN(new_n682));
  OAI21_X1  g496(.A(new_n361), .B1(new_n682), .B2(new_n353), .ZN(new_n683));
  AOI211_X1 g497(.A(KEYINPUT91), .B(new_n363), .C1(new_n683), .C2(new_n305), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n368), .B1(new_n367), .B2(KEYINPUT20), .ZN(new_n685));
  OAI21_X1  g499(.A(KEYINPUT99), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT99), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n364), .A2(new_n687), .A3(new_n369), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  AOI21_X1  g503(.A(new_n426), .B1(new_n689), .B2(new_n370), .ZN(new_n690));
  XOR2_X1   g504(.A(new_n433), .B(KEYINPUT100), .Z(new_n691));
  NAND4_X1  g505(.A1(new_n665), .A2(new_n690), .A3(new_n375), .A4(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n658), .A2(new_n693), .ZN(new_n694));
  XOR2_X1   g508(.A(KEYINPUT35), .B(G107), .Z(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NAND2_X1  g510(.A1(new_n635), .A2(new_n626), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n632), .A2(KEYINPUT36), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n620), .B(new_n698), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n699), .A2(new_n627), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n511), .A2(new_n656), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(KEYINPUT101), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT37), .B(G110), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G12));
  INV_X1    g519(.A(G900), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n431), .B1(new_n427), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n707), .B1(new_n374), .B2(G475), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n665), .A2(new_n690), .A3(new_n708), .ZN(new_n709));
  NOR3_X1   g523(.A1(new_n301), .A2(new_n709), .A3(new_n304), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n710), .A2(new_n589), .A3(new_n640), .A4(new_n701), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G128), .ZN(G30));
  AOI21_X1  g526(.A(new_n554), .B1(new_n570), .B2(new_n523), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n524), .A2(new_n560), .ZN(new_n714));
  AOI21_X1  g528(.A(G902), .B1(new_n714), .B2(new_n554), .ZN(new_n715));
  INV_X1    g529(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(G472), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n639), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n697), .A3(new_n700), .ZN(new_n719));
  INV_X1    g533(.A(new_n507), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT102), .B(KEYINPUT38), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n506), .B(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n426), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n376), .ZN(new_n725));
  NOR4_X1   g539(.A1(new_n719), .A2(new_n720), .A3(new_n723), .A4(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(new_n707), .B(KEYINPUT39), .Z(new_n727));
  NAND2_X1  g541(.A1(new_n652), .A2(new_n727), .ZN(new_n728));
  OR2_X1    g542(.A1(new_n728), .A2(KEYINPUT40), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(KEYINPUT40), .ZN(new_n730));
  NAND3_X1  g544(.A1(new_n726), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G143), .ZN(G45));
  AND3_X1   g546(.A1(new_n639), .A2(KEYINPUT72), .A3(new_n568), .ZN(new_n733));
  AOI21_X1  g547(.A(KEYINPUT72), .B1(new_n639), .B2(new_n568), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g549(.A(new_n507), .B(new_n660), .C1(new_n506), .C2(new_n659), .ZN(new_n736));
  INV_X1    g550(.A(new_n707), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n376), .A2(new_n674), .A3(new_n737), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(KEYINPUT103), .ZN(new_n740));
  INV_X1    g554(.A(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n735), .A2(new_n741), .A3(new_n652), .A4(new_n701), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G146), .ZN(G48));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  OR2_X1    g558(.A1(new_n291), .A2(new_n280), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n651), .A2(new_n303), .A3(new_n665), .A4(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n675), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n735), .A2(new_n744), .A3(new_n636), .A4(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n589), .A2(new_n636), .A3(new_n640), .ZN(new_n749));
  INV_X1    g563(.A(new_n746), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n676), .ZN(new_n751));
  OAI21_X1  g565(.A(KEYINPUT104), .B1(new_n749), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n748), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  OAI211_X1 g569(.A(new_n303), .B(new_n745), .C1(new_n644), .C2(new_n645), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n756), .A2(new_n692), .ZN(new_n757));
  NAND4_X1  g571(.A1(new_n589), .A2(new_n757), .A3(new_n636), .A4(new_n640), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G116), .ZN(G18));
  NOR2_X1   g573(.A1(new_n746), .A2(new_n434), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n760), .A2(new_n589), .A3(new_n640), .A4(new_n701), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(G119), .ZN(G21));
  INV_X1    g576(.A(new_n636), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n573), .A2(new_n574), .ZN(new_n764));
  OR2_X1    g578(.A1(new_n553), .A2(KEYINPUT105), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n553), .A2(KEYINPUT105), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n765), .A2(new_n554), .A3(new_n766), .ZN(new_n767));
  AOI21_X1  g581(.A(new_n578), .B1(new_n764), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g582(.A1(new_n763), .A2(new_n655), .A3(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(new_n756), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n725), .A2(new_n736), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n691), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G122), .ZN(G24));
  NOR2_X1   g587(.A1(new_n655), .A2(new_n768), .ZN(new_n774));
  INV_X1    g588(.A(new_n738), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n774), .A2(new_n701), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n776), .A2(new_n746), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(new_n337), .ZN(G27));
  OAI21_X1  g592(.A(KEYINPUT106), .B1(new_n301), .B2(new_n304), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n646), .A2(new_n780), .A3(new_n303), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n664), .A2(new_n507), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n749), .A2(new_n784), .ZN(new_n785));
  NOR2_X1   g599(.A1(new_n738), .A2(KEYINPUT42), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n782), .B1(new_n647), .B2(KEYINPUT106), .ZN(new_n787));
  AOI21_X1  g601(.A(new_n763), .B1(new_n639), .B2(new_n568), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n787), .A2(new_n775), .A3(new_n788), .A4(new_n781), .ZN(new_n789));
  AOI22_X1  g603(.A1(new_n785), .A2(new_n786), .B1(new_n789), .B2(KEYINPUT42), .ZN(new_n790));
  XNOR2_X1  g604(.A(KEYINPUT107), .B(G131), .ZN(new_n791));
  XNOR2_X1  g605(.A(new_n790), .B(new_n791), .ZN(G33));
  NAND2_X1  g606(.A1(new_n690), .A2(new_n708), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n749), .A2(new_n784), .A3(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n188), .ZN(G36));
  NOR2_X1   g609(.A1(new_n298), .A2(new_n299), .ZN(new_n796));
  INV_X1    g610(.A(new_n296), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT45), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n800), .A2(new_n280), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  AOI22_X1  g616(.A1(new_n801), .A2(new_n802), .B1(G469), .B2(G902), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n803), .A2(KEYINPUT46), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n651), .B1(new_n803), .B2(KEYINPUT46), .ZN(new_n805));
  OAI211_X1 g619(.A(new_n303), .B(new_n727), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  INV_X1    g620(.A(new_n806), .ZN(new_n807));
  XNOR2_X1  g621(.A(new_n782), .B(KEYINPUT109), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n377), .A2(new_n674), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT108), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(KEYINPUT43), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n813), .B1(new_n810), .B2(new_n814), .ZN(new_n815));
  INV_X1    g629(.A(new_n656), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n816), .A3(new_n701), .ZN(new_n817));
  OR2_X1    g631(.A1(new_n817), .A2(KEYINPUT44), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(KEYINPUT44), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n809), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n807), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G137), .ZN(G39));
  OR4_X1    g636(.A1(new_n636), .A2(new_n735), .A3(new_n738), .A4(new_n782), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n303), .B1(new_n804), .B2(new_n805), .ZN(new_n824));
  INV_X1    g638(.A(KEYINPUT47), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OAI211_X1 g640(.A(KEYINPUT47), .B(new_n303), .C1(new_n804), .C2(new_n805), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n823), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  XNOR2_X1  g642(.A(new_n828), .B(new_n308), .ZN(G42));
  NOR4_X1   g643(.A1(new_n763), .A2(new_n810), .A3(new_n304), .A4(new_n508), .ZN(new_n830));
  INV_X1    g644(.A(new_n830), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n831), .A2(KEYINPUT110), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n722), .B1(new_n831), .B2(KEYINPUT110), .ZN(new_n833));
  INV_X1    g647(.A(new_n718), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n651), .A2(new_n745), .ZN(new_n835));
  XOR2_X1   g649(.A(new_n835), .B(KEYINPUT49), .Z(new_n836));
  NAND4_X1  g650(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n430), .A2(new_n263), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT51), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n827), .ZN(new_n840));
  INV_X1    g654(.A(new_n835), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n840), .B1(new_n304), .B2(new_n841), .ZN(new_n842));
  AND2_X1   g656(.A1(new_n815), .A2(new_n431), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n769), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n844), .A2(new_n809), .ZN(new_n845));
  XOR2_X1   g659(.A(new_n845), .B(KEYINPUT117), .Z(new_n846));
  NOR2_X1   g660(.A1(new_n842), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n756), .A2(new_n782), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n843), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g663(.A(new_n849), .B(KEYINPUT119), .Z(new_n850));
  NAND3_X1  g664(.A1(new_n850), .A2(new_n701), .A3(new_n774), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT118), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n770), .A2(new_n720), .A3(new_n723), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n852), .B1(new_n844), .B2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(KEYINPUT50), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n834), .A2(new_n848), .A3(new_n636), .A4(new_n431), .ZN(new_n856));
  OR3_X1    g670(.A1(new_n856), .A2(new_n376), .A3(new_n674), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n851), .A2(new_n855), .A3(new_n857), .ZN(new_n858));
  OAI21_X1  g672(.A(new_n839), .B1(new_n847), .B2(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(new_n858), .ZN(new_n860));
  OAI211_X1 g674(.A(new_n860), .B(KEYINPUT51), .C1(new_n842), .C2(new_n846), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n430), .A2(G953), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n376), .A2(new_n674), .ZN(new_n863));
  OAI221_X1 g677(.A(new_n862), .B1(new_n856), .B2(new_n863), .C1(new_n746), .C2(new_n844), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n850), .A2(new_n788), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT48), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(KEYINPUT48), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n859), .A2(new_n861), .A3(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n777), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n589), .A2(new_n640), .A3(new_n652), .A4(new_n701), .ZN(new_n871));
  OAI211_X1 g685(.A(new_n711), .B(new_n870), .C1(new_n871), .C2(new_n740), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n652), .A2(new_n737), .A3(new_n771), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n719), .A2(new_n873), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT114), .B1(new_n872), .B2(new_n874), .ZN(new_n875));
  AND3_X1   g689(.A1(new_n589), .A2(new_n640), .A3(new_n701), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n777), .B1(new_n876), .B2(new_n710), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT114), .ZN(new_n878));
  INV_X1    g692(.A(new_n874), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n877), .A2(new_n878), .A3(new_n742), .A4(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n880), .A3(KEYINPUT52), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n689), .A2(new_n370), .ZN(new_n882));
  INV_X1    g696(.A(new_n708), .ZN(new_n883));
  NOR4_X1   g697(.A1(new_n882), .A2(new_n782), .A3(new_n724), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n871), .A2(new_n885), .B1(new_n784), .B2(new_n776), .ZN(new_n886));
  OAI21_X1  g700(.A(KEYINPUT111), .B1(new_n794), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g701(.A1(new_n779), .A2(new_n781), .A3(new_n783), .ZN(new_n888));
  INV_X1    g702(.A(new_n793), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n888), .A2(new_n636), .A3(new_n735), .A4(new_n889), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT111), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n784), .A2(new_n776), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n735), .A2(new_n652), .A3(new_n701), .A4(new_n884), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n376), .A2(new_n426), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(new_n376), .B2(new_n674), .ZN(new_n897));
  INV_X1    g711(.A(new_n691), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n897), .A2(new_n510), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n650), .A2(new_n657), .A3(new_n899), .ZN(new_n900));
  AND3_X1   g714(.A1(new_n900), .A2(new_n641), .A3(new_n702), .ZN(new_n901));
  AND3_X1   g715(.A1(new_n761), .A2(new_n758), .A3(new_n772), .ZN(new_n902));
  AND3_X1   g716(.A1(new_n901), .A2(new_n753), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n881), .A2(new_n790), .A3(new_n895), .A4(new_n903), .ZN(new_n904));
  AOI21_X1  g718(.A(KEYINPUT52), .B1(new_n875), .B2(new_n880), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT53), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT112), .ZN(new_n907));
  AND2_X1   g721(.A1(new_n887), .A2(new_n894), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n790), .A2(new_n753), .A3(new_n902), .A4(new_n901), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n907), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  NAND4_X1  g724(.A1(new_n903), .A2(new_n895), .A3(KEYINPUT112), .A4(new_n790), .ZN(new_n911));
  OAI211_X1 g725(.A(KEYINPUT113), .B(KEYINPUT52), .C1(new_n872), .C2(new_n874), .ZN(new_n912));
  XOR2_X1   g726(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n913));
  NAND4_X1  g727(.A1(new_n877), .A2(new_n742), .A3(new_n879), .A4(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n915), .A2(KEYINPUT53), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n910), .A2(new_n911), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n906), .A2(new_n917), .A3(KEYINPUT54), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT53), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n904), .B2(new_n905), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT54), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n753), .A2(new_n902), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT116), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n753), .A2(new_n902), .A3(KEYINPUT116), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n915), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n790), .A2(KEYINPUT53), .A3(new_n901), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n908), .A2(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n926), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n920), .A2(new_n921), .A3(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT115), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n918), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n906), .A2(new_n917), .A3(KEYINPUT115), .A4(KEYINPUT54), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n869), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n838), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g750(.A(KEYINPUT120), .B(new_n869), .C1(new_n932), .C2(new_n933), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n837), .B1(new_n936), .B2(new_n937), .ZN(G75));
  INV_X1    g752(.A(KEYINPUT56), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n281), .B1(new_n920), .B2(new_n929), .ZN(new_n940));
  INV_X1    g754(.A(new_n940), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n939), .B1(new_n941), .B2(new_n435), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n463), .A2(new_n464), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n474), .ZN(new_n944));
  NOR2_X1   g758(.A1(new_n944), .A2(new_n475), .ZN(new_n945));
  XOR2_X1   g759(.A(new_n945), .B(KEYINPUT55), .Z(new_n946));
  AND2_X1   g760(.A1(new_n942), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n942), .A2(new_n946), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n263), .A2(G952), .ZN(new_n949));
  NOR3_X1   g763(.A1(new_n947), .A2(new_n948), .A3(new_n949), .ZN(G51));
  NAND2_X1  g764(.A1(new_n920), .A2(new_n929), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n951), .A2(KEYINPUT54), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n930), .ZN(new_n953));
  NAND2_X1  g767(.A1(G469), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT57), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n279), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n940), .A2(new_n802), .A3(new_n801), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n949), .B1(new_n957), .B2(new_n958), .ZN(G54));
  INV_X1    g773(.A(new_n683), .ZN(new_n960));
  NAND2_X1  g774(.A1(KEYINPUT58), .A2(G475), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n960), .B1(new_n941), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n949), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n940), .A2(KEYINPUT58), .A3(G475), .A4(new_n683), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n963), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT121), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT121), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n962), .A2(new_n967), .A3(new_n963), .A4(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n968), .ZN(G60));
  XOR2_X1   g783(.A(new_n672), .B(KEYINPUT122), .Z(new_n970));
  NAND2_X1  g784(.A1(G478), .A2(G902), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n971), .B(KEYINPUT59), .Z(new_n972));
  NOR2_X1   g786(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n953), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(new_n963), .ZN(new_n975));
  INV_X1    g789(.A(new_n972), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n932), .A2(new_n933), .A3(new_n976), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n975), .B1(new_n970), .B2(new_n977), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT60), .Z(new_n980));
  NAND3_X1  g794(.A1(new_n951), .A2(new_n699), .A3(new_n980), .ZN(new_n981));
  AND2_X1   g795(.A1(new_n951), .A2(new_n980), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n963), .B(new_n981), .C1(new_n982), .C2(new_n633), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G66));
  INV_X1    g799(.A(new_n428), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n263), .B1(new_n986), .B2(G224), .ZN(new_n987));
  INV_X1    g801(.A(new_n903), .ZN(new_n988));
  AOI21_X1  g802(.A(new_n987), .B1(new_n988), .B2(new_n263), .ZN(new_n989));
  INV_X1    g803(.A(G898), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n943), .B1(new_n990), .B2(G953), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n989), .B(new_n991), .ZN(G69));
  AND2_X1   g806(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n993));
  NOR2_X1   g807(.A1(new_n872), .A2(KEYINPUT123), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n788), .A2(new_n771), .ZN(new_n996));
  OR3_X1    g810(.A1(new_n806), .A2(KEYINPUT124), .A3(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(KEYINPUT124), .B1(new_n806), .B2(new_n996), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n995), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n821), .ZN(new_n1000));
  NOR2_X1   g814(.A1(new_n1000), .A2(new_n828), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n790), .A2(new_n890), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n999), .A2(new_n1001), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1003), .A2(KEYINPUT125), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  NAND4_X1  g819(.A1(new_n999), .A2(new_n1005), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1004), .A2(new_n263), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n542), .A2(new_n528), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(new_n341), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1009), .B1(G900), .B2(G953), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NOR4_X1   g825(.A1(new_n749), .A2(new_n728), .A3(new_n782), .A4(new_n897), .ZN(new_n1012));
  NOR3_X1   g826(.A1(new_n1000), .A2(new_n828), .A3(new_n1012), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n731), .B1(new_n993), .B2(new_n994), .ZN(new_n1014));
  OR2_X1    g828(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1014), .A2(KEYINPUT62), .ZN(new_n1016));
  AND3_X1   g830(.A1(new_n1013), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1009), .B1(new_n1017), .B2(G953), .ZN(new_n1018));
  NAND2_X1  g832(.A1(new_n1011), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n263), .B1(G227), .B2(G900), .ZN(new_n1020));
  XNOR2_X1  g834(.A(new_n1019), .B(new_n1020), .ZN(G72));
  INV_X1    g835(.A(new_n713), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1013), .A2(new_n1015), .A3(new_n903), .A4(new_n1016), .ZN(new_n1023));
  XNOR2_X1  g837(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1024));
  NOR2_X1   g838(.A1(new_n654), .A2(new_n293), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1024), .B(new_n1025), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n1022), .B1(new_n1023), .B2(new_n1026), .ZN(new_n1027));
  XNOR2_X1  g841(.A(new_n1027), .B(KEYINPUT127), .ZN(new_n1028));
  INV_X1    g842(.A(new_n545), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1004), .A2(new_n903), .A3(new_n1006), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n1026), .ZN(new_n1031));
  AND3_X1   g845(.A1(new_n1022), .A2(new_n1029), .A3(new_n1026), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n906), .A2(new_n917), .A3(new_n1032), .ZN(new_n1033));
  NOR4_X1   g847(.A1(new_n1028), .A2(new_n949), .A3(new_n1031), .A4(new_n1033), .ZN(G57));
endmodule


