//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 1 1 0 1 1 1 1 0 0 0 0 0 0 0 0 0 0 0 0 1 0 0 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 1 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n447, new_n449, new_n450, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n560, new_n561, new_n563, new_n564, new_n565, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n640, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201, new_n1202;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT64), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XNOR2_X1  g017(.A(new_n442), .B(KEYINPUT65), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  INV_X1    g023(.A(G567), .ZN(new_n449));
  NOR2_X1   g024(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT66), .Z(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G219), .A2(G220), .A3(G218), .A4(G221), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n454), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n454), .A2(new_n458), .B1(new_n449), .B2(new_n455), .ZN(new_n459));
  XOR2_X1   g034(.A(new_n459), .B(KEYINPUT67), .Z(G319));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  AOI21_X1  g040(.A(KEYINPUT68), .B1(new_n465), .B2(G2105), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  AOI211_X1 g043(.A(new_n467), .B(new_n468), .C1(new_n463), .C2(new_n464), .ZN(new_n469));
  OR2_X1    g044(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  AND3_X1   g045(.A1(new_n468), .A2(G101), .A3(G2104), .ZN(new_n471));
  OAI211_X1 g046(.A(G137), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(KEYINPUT69), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT3), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n476), .A2(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND4_X1  g054(.A1(new_n478), .A2(new_n479), .A3(G137), .A4(new_n468), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n471), .B1(new_n473), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n470), .A2(new_n481), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(G160));
  OAI21_X1  g058(.A(G2104), .B1(new_n468), .B2(G112), .ZN(new_n484));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AOI21_X1  g060(.A(new_n484), .B1(new_n485), .B2(new_n468), .ZN(new_n486));
  AOI21_X1  g061(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n487));
  INV_X1    g062(.A(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  OR3_X1    g064(.A1(new_n488), .A2(KEYINPUT70), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT70), .B1(new_n488), .B2(new_n489), .ZN(new_n491));
  AND2_X1   g066(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n478), .A2(G2105), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  AOI211_X1 g069(.A(new_n486), .B(new_n492), .C1(G124), .C2(new_n494), .ZN(G162));
  OAI211_X1 g070(.A(KEYINPUT4), .B(G138), .C1(new_n461), .C2(new_n462), .ZN(new_n496));
  NAND2_X1  g071(.A1(G102), .A2(G2104), .ZN(new_n497));
  AOI21_X1  g072(.A(G2105), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g073(.A(KEYINPUT4), .B1(new_n487), .B2(G138), .ZN(new_n499));
  OAI21_X1  g074(.A(G126), .B1(new_n461), .B2(new_n462), .ZN(new_n500));
  NAND2_X1  g075(.A1(G114), .A2(G2104), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n468), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n498), .A2(new_n499), .A3(new_n502), .ZN(G164));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(G50), .A3(G543), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT71), .ZN(new_n506));
  XNOR2_X1  g081(.A(new_n505), .B(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(KEYINPUT72), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(G543), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  INV_X1    g088(.A(G651), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AND3_X1   g090(.A1(KEYINPUT72), .A2(KEYINPUT5), .A3(G543), .ZN(new_n516));
  AOI21_X1  g091(.A(G543), .B1(KEYINPUT72), .B2(KEYINPUT5), .ZN(new_n517));
  NOR2_X1   g092(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT6), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n520), .A2(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n518), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n507), .A2(new_n515), .A3(new_n524), .ZN(G303));
  INV_X1    g100(.A(G303), .ZN(G166));
  NAND2_X1  g101(.A1(G63), .A2(G651), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n522), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n529), .A2(new_n512), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n520), .A2(G651), .ZN(new_n531));
  NOR2_X1   g106(.A1(new_n514), .A2(KEYINPUT6), .ZN(new_n532));
  OAI21_X1  g107(.A(KEYINPUT73), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT73), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n519), .A2(new_n521), .A3(new_n534), .ZN(new_n535));
  NAND4_X1  g110(.A1(new_n533), .A2(G51), .A3(G543), .A4(new_n535), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  AND3_X1   g113(.A1(new_n530), .A2(new_n536), .A3(new_n538), .ZN(G168));
  NAND2_X1  g114(.A1(new_n523), .A2(G90), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n533), .A2(G52), .A3(G543), .A4(new_n535), .ZN(new_n541));
  INV_X1    g116(.A(G64), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n542), .B1(new_n510), .B2(new_n511), .ZN(new_n543));
  INV_X1    g118(.A(G77), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n544), .A2(new_n509), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND3_X1  g121(.A1(new_n540), .A2(new_n541), .A3(new_n546), .ZN(G301));
  INV_X1    g122(.A(G301), .ZN(G171));
  NAND4_X1  g123(.A1(new_n533), .A2(G43), .A3(G543), .A4(new_n535), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n550), .B1(new_n510), .B2(new_n511), .ZN(new_n551));
  AND2_X1   g126(.A1(G68), .A2(G543), .ZN(new_n552));
  OAI21_X1  g127(.A(G651), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT74), .B(G81), .ZN(new_n554));
  NAND3_X1  g129(.A1(new_n512), .A2(new_n504), .A3(new_n554), .ZN(new_n555));
  AND3_X1   g130(.A1(new_n549), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G860), .ZN(G153));
  AND3_X1   g132(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n558), .A2(G36), .ZN(G176));
  NAND2_X1  g134(.A1(G1), .A2(G3), .ZN(new_n560));
  XNOR2_X1  g135(.A(new_n560), .B(KEYINPUT8), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n558), .A2(new_n561), .ZN(G188));
  AND3_X1   g137(.A1(new_n519), .A2(new_n521), .A3(new_n534), .ZN(new_n563));
  AOI21_X1  g138(.A(new_n534), .B1(new_n519), .B2(new_n521), .ZN(new_n564));
  NOR2_X1   g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n565), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n566));
  NAND4_X1  g141(.A1(new_n533), .A2(G53), .A3(G543), .A4(new_n535), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT9), .ZN(new_n568));
  NAND2_X1  g143(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n523), .A2(G91), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n518), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND4_X1  g149(.A1(new_n566), .A2(new_n569), .A3(new_n570), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT75), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n567), .A2(new_n568), .B1(new_n573), .B2(G651), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n577), .A2(new_n578), .A3(new_n570), .A4(new_n566), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G299));
  NAND3_X1  g155(.A1(new_n530), .A2(new_n536), .A3(new_n538), .ZN(G286));
  NOR3_X1   g156(.A1(new_n563), .A2(new_n564), .A3(new_n509), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n582), .A2(KEYINPUT76), .A3(G49), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND3_X1  g159(.A1(new_n533), .A2(G543), .A3(new_n535), .ZN(new_n585));
  INV_X1    g160(.A(G49), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n584), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  AOI22_X1  g162(.A1(new_n583), .A2(new_n587), .B1(G87), .B2(new_n523), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n589));
  AND3_X1   g164(.A1(new_n588), .A2(KEYINPUT77), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(KEYINPUT77), .B1(new_n588), .B2(new_n589), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G288));
  NAND2_X1  g168(.A1(new_n523), .A2(G86), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT78), .ZN(new_n595));
  NAND2_X1  g170(.A1(G48), .A2(G543), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n522), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n504), .A2(KEYINPUT78), .A3(G48), .A4(G543), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n512), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n600));
  OAI211_X1 g175(.A(new_n594), .B(new_n599), .C1(new_n514), .C2(new_n600), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT79), .ZN(new_n602));
  XNOR2_X1  g177(.A(new_n601), .B(new_n602), .ZN(G305));
  INV_X1    g178(.A(G60), .ZN(new_n604));
  INV_X1    g179(.A(G72), .ZN(new_n605));
  OAI22_X1  g180(.A1(new_n518), .A2(new_n604), .B1(new_n605), .B2(new_n509), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n606), .A2(KEYINPUT80), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT80), .ZN(new_n608));
  OAI221_X1 g183(.A(new_n608), .B1(new_n605), .B2(new_n509), .C1(new_n518), .C2(new_n604), .ZN(new_n609));
  NAND3_X1  g184(.A1(new_n607), .A2(G651), .A3(new_n609), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n533), .A2(G47), .A3(G543), .A4(new_n535), .ZN(new_n611));
  INV_X1    g186(.A(KEYINPUT81), .ZN(new_n612));
  NAND3_X1  g187(.A1(new_n512), .A2(G85), .A3(new_n504), .ZN(new_n613));
  AND3_X1   g188(.A1(new_n611), .A2(new_n612), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n612), .B1(new_n611), .B2(new_n613), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n610), .B1(new_n614), .B2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT82), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  OAI211_X1 g193(.A(new_n610), .B(KEYINPUT82), .C1(new_n614), .C2(new_n615), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n618), .A2(new_n619), .ZN(G290));
  NAND2_X1  g195(.A1(G301), .A2(G868), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n622));
  INV_X1    g197(.A(G79), .ZN(new_n623));
  INV_X1    g198(.A(G66), .ZN(new_n624));
  OAI221_X1 g199(.A(new_n622), .B1(new_n623), .B2(new_n509), .C1(new_n518), .C2(new_n624), .ZN(new_n625));
  AOI21_X1  g200(.A(new_n624), .B1(new_n510), .B2(new_n511), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n623), .A2(new_n509), .ZN(new_n627));
  OAI21_X1  g202(.A(KEYINPUT83), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g203(.A1(new_n625), .A2(G651), .A3(new_n628), .ZN(new_n629));
  NAND3_X1  g204(.A1(new_n523), .A2(KEYINPUT10), .A3(G92), .ZN(new_n630));
  INV_X1    g205(.A(KEYINPUT10), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n512), .A2(new_n504), .ZN(new_n632));
  INV_X1    g207(.A(G92), .ZN(new_n633));
  OAI21_X1  g208(.A(new_n631), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n630), .A2(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n582), .A2(G54), .ZN(new_n636));
  AND3_X1   g211(.A1(new_n629), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n621), .B1(new_n637), .B2(G868), .ZN(G284));
  XOR2_X1   g213(.A(G284), .B(KEYINPUT84), .Z(G321));
  INV_X1    g214(.A(G868), .ZN(new_n640));
  MUX2_X1   g215(.A(G286), .B(G299), .S(new_n640), .Z(G297));
  XOR2_X1   g216(.A(G297), .B(KEYINPUT85), .Z(G280));
  INV_X1    g217(.A(G559), .ZN(new_n643));
  OAI21_X1  g218(.A(new_n637), .B1(new_n643), .B2(G860), .ZN(G148));
  NAND3_X1  g219(.A1(new_n549), .A2(new_n553), .A3(new_n555), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n645), .A2(new_n640), .ZN(new_n646));
  INV_X1    g221(.A(new_n637), .ZN(new_n647));
  NOR2_X1   g222(.A1(new_n647), .A2(G559), .ZN(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n648), .B2(new_n640), .ZN(G323));
  XNOR2_X1  g224(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g225(.A1(new_n487), .A2(G2104), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT12), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT86), .Z(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT13), .ZN(new_n654));
  NOR2_X1   g229(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n655));
  AND2_X1   g230(.A1(KEYINPUT87), .A2(G2100), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n487), .A2(G135), .ZN(new_n658));
  NOR2_X1   g233(.A1(G99), .A2(G2105), .ZN(new_n659));
  OAI21_X1  g234(.A(G2104), .B1(new_n468), .B2(G111), .ZN(new_n660));
  INV_X1    g235(.A(G123), .ZN(new_n661));
  OAI221_X1 g236(.A(new_n658), .B1(new_n659), .B2(new_n660), .C1(new_n661), .C2(new_n493), .ZN(new_n662));
  XOR2_X1   g237(.A(new_n662), .B(G2096), .Z(new_n663));
  OAI211_X1 g238(.A(new_n657), .B(new_n663), .C1(new_n655), .C2(new_n654), .ZN(G156));
  XNOR2_X1  g239(.A(KEYINPUT15), .B(G2435), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT89), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(G2438), .ZN(new_n667));
  XNOR2_X1  g242(.A(G2427), .B(G2430), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n669), .A2(KEYINPUT14), .ZN(new_n670));
  XNOR2_X1  g245(.A(G2451), .B(G2454), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G2443), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2446), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  XNOR2_X1  g249(.A(KEYINPUT88), .B(KEYINPUT16), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n674), .B(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1341), .B(G1348), .ZN(new_n677));
  OR2_X1    g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n676), .A2(new_n677), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n678), .A2(G14), .A3(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT90), .ZN(G401));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  INV_X1    g257(.A(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G2067), .B(G2678), .Z(new_n684));
  OR2_X1    g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT17), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT18), .ZN(new_n688));
  NAND2_X1  g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g264(.A(G2072), .B(G2078), .Z(new_n690));
  AOI21_X1  g265(.A(new_n690), .B1(new_n685), .B2(KEYINPUT18), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n689), .B(new_n691), .ZN(new_n692));
  XNOR2_X1  g267(.A(G2096), .B(G2100), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(G227));
  XNOR2_X1  g269(.A(G1971), .B(G1976), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT91), .ZN(new_n696));
  XOR2_X1   g271(.A(new_n696), .B(KEYINPUT19), .Z(new_n697));
  XOR2_X1   g272(.A(G1956), .B(G2474), .Z(new_n698));
  XOR2_X1   g273(.A(G1961), .B(G1966), .Z(new_n699));
  AND2_X1   g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n701), .B(KEYINPUT20), .ZN(new_n702));
  NOR2_X1   g277(.A1(new_n698), .A2(new_n699), .ZN(new_n703));
  OR3_X1    g278(.A1(new_n697), .A2(new_n700), .A3(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n697), .A2(new_n703), .ZN(new_n705));
  NAND3_X1  g280(.A1(new_n702), .A2(new_n704), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(G1991), .B(G1996), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1981), .B(G1986), .ZN(new_n709));
  XNOR2_X1  g284(.A(new_n708), .B(new_n709), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(G229));
  NOR2_X1   g287(.A1(G5), .A2(G16), .ZN(new_n713));
  AOI21_X1  g288(.A(new_n713), .B1(G171), .B2(G16), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n714), .A2(G1961), .ZN(new_n715));
  INV_X1    g290(.A(G29), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(G35), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G162), .B2(new_n716), .ZN(new_n718));
  XOR2_X1   g293(.A(new_n718), .B(KEYINPUT29), .Z(new_n719));
  INV_X1    g294(.A(new_n719), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT28), .ZN(new_n721));
  INV_X1    g296(.A(G26), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n721), .B1(new_n722), .B2(G29), .ZN(new_n723));
  NOR2_X1   g298(.A1(new_n722), .A2(G29), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n487), .A2(G140), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT97), .Z(new_n726));
  NAND2_X1  g301(.A1(new_n494), .A2(G128), .ZN(new_n727));
  NOR2_X1   g302(.A1(G104), .A2(G2105), .ZN(new_n728));
  OAI21_X1  g303(.A(G2104), .B1(new_n468), .B2(G116), .ZN(new_n729));
  OAI211_X1 g304(.A(new_n726), .B(new_n727), .C1(new_n728), .C2(new_n729), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n724), .B1(new_n730), .B2(G29), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n723), .B1(new_n731), .B2(new_n721), .ZN(new_n732));
  AOI22_X1  g307(.A1(new_n720), .A2(G2090), .B1(G2067), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n716), .A2(G27), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G164), .B2(new_n716), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G2078), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n716), .A2(G33), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT25), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n487), .A2(G139), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n478), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n741));
  OAI211_X1 g316(.A(new_n739), .B(new_n740), .C1(new_n741), .C2(new_n468), .ZN(new_n742));
  AOI21_X1  g317(.A(new_n737), .B1(new_n742), .B2(G29), .ZN(new_n743));
  INV_X1    g318(.A(new_n743), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n744), .A2(G2072), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT31), .B(G11), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n744), .A2(G2072), .ZN(new_n747));
  XOR2_X1   g322(.A(KEYINPUT30), .B(G28), .Z(new_n748));
  MUX2_X1   g323(.A(new_n748), .B(new_n662), .S(G29), .Z(new_n749));
  NAND4_X1  g324(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G2090), .ZN(new_n751));
  AOI211_X1 g326(.A(new_n736), .B(new_n750), .C1(new_n719), .C2(new_n751), .ZN(new_n752));
  OR2_X1    g327(.A1(new_n732), .A2(G2067), .ZN(new_n753));
  AND2_X1   g328(.A1(KEYINPUT24), .A2(G34), .ZN(new_n754));
  NOR2_X1   g329(.A1(KEYINPUT24), .A2(G34), .ZN(new_n755));
  NOR3_X1   g330(.A1(new_n754), .A2(new_n755), .A3(G29), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(new_n482), .B2(G29), .ZN(new_n757));
  INV_X1    g332(.A(G2084), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G1961), .B2(new_n714), .ZN(new_n760));
  NOR2_X1   g335(.A1(G16), .A2(G19), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n556), .B2(G16), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(G1341), .Z(new_n763));
  NAND2_X1  g338(.A1(new_n716), .A2(G32), .ZN(new_n764));
  AND3_X1   g339(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT26), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n487), .A2(G141), .ZN(new_n767));
  INV_X1    g342(.A(G129), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n766), .B(new_n767), .C1(new_n768), .C2(new_n493), .ZN(new_n769));
  NAND3_X1  g344(.A1(new_n468), .A2(G105), .A3(G2104), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT99), .Z(new_n771));
  NOR2_X1   g346(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n764), .B1(new_n772), .B2(new_n716), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT100), .Z(new_n774));
  XOR2_X1   g349(.A(KEYINPUT27), .B(G1996), .Z(new_n775));
  OAI21_X1  g350(.A(new_n763), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n760), .B(new_n776), .C1(new_n775), .C2(new_n774), .ZN(new_n777));
  NAND4_X1  g352(.A1(new_n733), .A2(new_n752), .A3(new_n753), .A4(new_n777), .ZN(new_n778));
  INV_X1    g353(.A(G16), .ZN(new_n779));
  AND3_X1   g354(.A1(new_n779), .A2(KEYINPUT23), .A3(G20), .ZN(new_n780));
  AOI21_X1  g355(.A(KEYINPUT23), .B1(new_n779), .B2(G20), .ZN(new_n781));
  AOI211_X1 g356(.A(new_n780), .B(new_n781), .C1(G299), .C2(G16), .ZN(new_n782));
  INV_X1    g357(.A(G1956), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g359(.A1(new_n757), .A2(new_n758), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT98), .Z(new_n786));
  OAI21_X1  g361(.A(KEYINPUT101), .B1(G16), .B2(G21), .ZN(new_n787));
  NOR2_X1   g362(.A1(G286), .A2(new_n779), .ZN(new_n788));
  MUX2_X1   g363(.A(new_n787), .B(KEYINPUT101), .S(new_n788), .Z(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G1966), .ZN(new_n790));
  OAI21_X1  g365(.A(KEYINPUT96), .B1(G4), .B2(G16), .ZN(new_n791));
  OR3_X1    g366(.A1(KEYINPUT96), .A2(G4), .A3(G16), .ZN(new_n792));
  OAI211_X1 g367(.A(new_n791), .B(new_n792), .C1(new_n647), .C2(new_n779), .ZN(new_n793));
  XNOR2_X1  g368(.A(new_n793), .B(G1348), .ZN(new_n794));
  NAND3_X1  g369(.A1(new_n786), .A2(new_n790), .A3(new_n794), .ZN(new_n795));
  NOR3_X1   g370(.A1(new_n778), .A2(new_n784), .A3(new_n795), .ZN(new_n796));
  AND2_X1   g371(.A1(new_n779), .A2(G23), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n588), .A2(new_n589), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n797), .B1(new_n798), .B2(G16), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT33), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(G1976), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n779), .A2(G22), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G166), .B2(new_n779), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n803), .A2(G1971), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n779), .A2(G6), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(G305), .B2(G16), .ZN(new_n806));
  XNOR2_X1  g381(.A(KEYINPUT32), .B(G1981), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(KEYINPUT94), .ZN(new_n808));
  AND2_X1   g383(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n806), .A2(new_n808), .ZN(new_n810));
  AND2_X1   g385(.A1(new_n803), .A2(G1971), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n809), .A2(new_n810), .A3(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n800), .A2(G1976), .ZN(new_n813));
  NAND4_X1  g388(.A1(new_n801), .A2(new_n804), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT34), .ZN(new_n815));
  MUX2_X1   g390(.A(G24), .B(G290), .S(G16), .Z(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(G1986), .Z(new_n817));
  AOI22_X1  g392(.A1(new_n494), .A2(G119), .B1(G131), .B2(new_n487), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n468), .A2(G107), .ZN(new_n819));
  OR3_X1    g394(.A1(KEYINPUT92), .A2(G95), .A3(G2105), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT92), .B1(G95), .B2(G2105), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n820), .A2(G2104), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n818), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  MUX2_X1   g398(.A(G25), .B(new_n823), .S(G29), .Z(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT35), .B(G1991), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT93), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n824), .B(new_n826), .ZN(new_n827));
  OAI211_X1 g402(.A(new_n817), .B(new_n827), .C1(new_n814), .C2(KEYINPUT34), .ZN(new_n828));
  INV_X1    g403(.A(KEYINPUT95), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AND2_X1   g405(.A1(new_n812), .A2(new_n813), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT34), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n831), .A2(new_n832), .A3(new_n804), .A4(new_n801), .ZN(new_n833));
  NAND4_X1  g408(.A1(new_n833), .A2(KEYINPUT95), .A3(new_n817), .A4(new_n827), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n815), .B1(new_n830), .B2(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(KEYINPUT36), .ZN(new_n836));
  NOR2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AOI211_X1 g412(.A(KEYINPUT36), .B(new_n815), .C1(new_n830), .C2(new_n834), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n715), .B(new_n796), .C1(new_n837), .C2(new_n838), .ZN(G150));
  INV_X1    g414(.A(G150), .ZN(G311));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n510), .B2(new_n511), .ZN(new_n842));
  INV_X1    g417(.A(G80), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n843), .A2(new_n509), .ZN(new_n844));
  OAI21_X1  g419(.A(G651), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(KEYINPUT102), .B(G93), .Z(new_n846));
  NAND3_X1  g421(.A1(new_n846), .A2(new_n512), .A3(new_n504), .ZN(new_n847));
  INV_X1    g422(.A(G55), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n845), .B(new_n847), .C1(new_n585), .C2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n849), .A2(G860), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT37), .Z(new_n851));
  NAND2_X1  g426(.A1(new_n637), .A2(G559), .ZN(new_n852));
  XOR2_X1   g427(.A(new_n852), .B(KEYINPUT39), .Z(new_n853));
  XNOR2_X1  g428(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n853), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n556), .A2(new_n849), .ZN(new_n856));
  OAI22_X1  g431(.A1(new_n518), .A2(new_n841), .B1(new_n843), .B2(new_n509), .ZN(new_n857));
  AOI22_X1  g432(.A1(new_n857), .A2(G651), .B1(new_n523), .B2(new_n846), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n582), .A2(G55), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n645), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n855), .B(new_n862), .ZN(new_n863));
  OAI21_X1  g438(.A(new_n851), .B1(new_n863), .B2(G860), .ZN(G145));
  OAI211_X1 g439(.A(G138), .B(new_n468), .C1(new_n461), .C2(new_n462), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT4), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  INV_X1    g442(.A(G126), .ZN(new_n868));
  AOI21_X1  g443(.A(new_n868), .B1(new_n476), .B2(new_n477), .ZN(new_n869));
  INV_X1    g444(.A(new_n501), .ZN(new_n870));
  OAI21_X1  g445(.A(G2105), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n497), .ZN(new_n872));
  INV_X1    g447(.A(G138), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n873), .B1(new_n476), .B2(new_n477), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n872), .B1(new_n874), .B2(KEYINPUT4), .ZN(new_n875));
  OAI211_X1 g450(.A(new_n867), .B(new_n871), .C1(new_n875), .C2(G2105), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n772), .B(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(new_n730), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n742), .A2(KEYINPUT104), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n742), .B(KEYINPUT104), .Z(new_n881));
  OAI21_X1  g456(.A(new_n880), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n487), .A2(G142), .ZN(new_n883));
  NOR2_X1   g458(.A1(G106), .A2(G2105), .ZN(new_n884));
  OAI21_X1  g459(.A(G2104), .B1(new_n468), .B2(G118), .ZN(new_n885));
  INV_X1    g460(.A(G130), .ZN(new_n886));
  OAI221_X1 g461(.A(new_n883), .B1(new_n884), .B2(new_n885), .C1(new_n886), .C2(new_n493), .ZN(new_n887));
  XNOR2_X1  g462(.A(new_n652), .B(new_n887), .ZN(new_n888));
  XNOR2_X1  g463(.A(new_n888), .B(new_n823), .ZN(new_n889));
  XNOR2_X1  g464(.A(KEYINPUT105), .B(KEYINPUT106), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n889), .B(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n882), .B(new_n891), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n482), .B(new_n662), .ZN(new_n893));
  XOR2_X1   g468(.A(new_n893), .B(G162), .Z(new_n894));
  INV_X1    g469(.A(new_n894), .ZN(new_n895));
  OR2_X1    g470(.A1(new_n892), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n892), .A2(new_n895), .ZN(new_n897));
  INV_X1    g472(.A(G37), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n849), .A2(new_n640), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n618), .A2(new_n798), .A3(new_n619), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n798), .B1(new_n618), .B2(new_n619), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n902), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n798), .ZN(new_n906));
  NAND2_X1  g481(.A1(G290), .A2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n618), .A2(new_n798), .A3(new_n619), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(KEYINPUT107), .A3(new_n908), .ZN(new_n909));
  XNOR2_X1  g484(.A(G305), .B(G303), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  XNOR2_X1  g486(.A(G305), .B(G166), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n912), .A2(KEYINPUT107), .A3(new_n907), .A4(new_n908), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(new_n914), .B(KEYINPUT42), .ZN(new_n915));
  INV_X1    g490(.A(KEYINPUT41), .ZN(new_n916));
  AND3_X1   g491(.A1(new_n576), .A2(new_n579), .A3(new_n637), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n637), .B1(new_n576), .B2(new_n579), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(G299), .A2(new_n647), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n576), .A2(new_n637), .A3(new_n579), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n920), .A2(KEYINPUT41), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n919), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n648), .B(new_n862), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NOR2_X1   g500(.A1(new_n917), .A2(new_n918), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n925), .B1(new_n926), .B2(new_n924), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n915), .B(new_n927), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n901), .B1(new_n928), .B2(new_n640), .ZN(G295));
  OAI21_X1  g504(.A(new_n901), .B1(new_n928), .B2(new_n640), .ZN(G331));
  AND2_X1   g505(.A1(new_n919), .A2(new_n922), .ZN(new_n931));
  NAND2_X1  g506(.A1(G168), .A2(G301), .ZN(new_n932));
  NAND4_X1  g507(.A1(G286), .A2(new_n541), .A3(new_n546), .A4(new_n540), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n861), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT109), .ZN(new_n936));
  NAND4_X1  g511(.A1(new_n932), .A2(new_n933), .A3(new_n856), .A4(new_n860), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n862), .A2(KEYINPUT109), .A3(new_n932), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n935), .A2(new_n937), .ZN(new_n942));
  INV_X1    g517(.A(new_n942), .ZN(new_n943));
  AOI22_X1  g518(.A1(new_n931), .A2(new_n941), .B1(new_n926), .B2(new_n943), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n944), .A2(KEYINPUT110), .A3(new_n911), .A4(new_n913), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n943), .A2(new_n926), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n947), .B1(new_n923), .B2(new_n940), .ZN(new_n948));
  OAI21_X1  g523(.A(new_n946), .B1(new_n914), .B2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n914), .A2(new_n948), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n945), .A2(new_n949), .A3(new_n898), .A4(new_n950), .ZN(new_n951));
  AND3_X1   g526(.A1(new_n951), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n952));
  AOI21_X1  g527(.A(KEYINPUT111), .B1(new_n951), .B2(KEYINPUT43), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n940), .A2(new_n926), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT112), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n919), .A2(new_n922), .A3(new_n942), .ZN(new_n957));
  NAND3_X1  g532(.A1(new_n940), .A2(KEYINPUT112), .A3(new_n926), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n959), .A2(new_n914), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n945), .A2(new_n960), .A3(new_n949), .A4(new_n898), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n961), .A2(KEYINPUT43), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n952), .A2(new_n953), .A3(new_n962), .ZN(new_n963));
  XNOR2_X1  g538(.A(KEYINPUT108), .B(KEYINPUT44), .ZN(new_n964));
  OAI21_X1  g539(.A(KEYINPUT113), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  OR2_X1    g540(.A1(new_n951), .A2(KEYINPUT43), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n967), .B1(new_n961), .B2(KEYINPUT43), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n966), .A2(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT114), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n966), .A2(new_n968), .A3(KEYINPUT114), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n953), .ZN(new_n974));
  INV_X1    g549(.A(new_n962), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n951), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n974), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT113), .ZN(new_n978));
  INV_X1    g553(.A(new_n964), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n977), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n965), .A2(new_n973), .A3(new_n980), .ZN(G397));
  INV_X1    g556(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g557(.A(new_n982), .B1(G164), .B2(G1384), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n481), .B(G40), .C1(new_n466), .C2(new_n469), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1996), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n987), .A2(new_n769), .A3(new_n771), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(KEYINPUT115), .ZN(new_n989));
  AND2_X1   g564(.A1(new_n988), .A2(KEYINPUT115), .ZN(new_n990));
  INV_X1    g565(.A(G2067), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n730), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g567(.A(new_n992), .B1(new_n986), .B2(new_n772), .ZN(new_n993));
  AOI211_X1 g568(.A(new_n989), .B(new_n990), .C1(new_n985), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n985), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n823), .B(new_n825), .Z(new_n996));
  OAI21_X1  g571(.A(new_n994), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NOR3_X1   g572(.A1(G290), .A2(new_n995), .A3(G1986), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n998), .B(KEYINPUT48), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NOR2_X1   g575(.A1(new_n823), .A2(new_n825), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n994), .A2(new_n1001), .ZN(new_n1002));
  OR2_X1    g577(.A1(new_n730), .A2(G2067), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n995), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n995), .B1(new_n992), .B2(new_n772), .ZN(new_n1005));
  INV_X1    g580(.A(new_n987), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n1006), .A2(KEYINPUT46), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n1005), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  XOR2_X1   g584(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n1010));
  XNOR2_X1  g585(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  NOR3_X1   g586(.A1(new_n1000), .A2(new_n1004), .A3(new_n1011), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT126), .ZN(new_n1013));
  XNOR2_X1  g588(.A(G290), .B(G1986), .ZN(new_n1014));
  AOI21_X1  g589(.A(new_n997), .B1(new_n985), .B2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT121), .ZN(new_n1016));
  NOR3_X1   g591(.A1(G164), .A2(new_n982), .A3(G1384), .ZN(new_n1017));
  INV_X1    g592(.A(G1384), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT45), .B1(new_n876), .B2(new_n1018), .ZN(new_n1019));
  NOR3_X1   g594(.A1(new_n1017), .A2(new_n1019), .A3(new_n984), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1016), .B1(new_n1020), .B2(G1966), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT50), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n876), .A2(new_n1022), .A3(new_n1018), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT117), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n876), .A2(KEYINPUT117), .A3(new_n1022), .A4(new_n1018), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1022), .B1(new_n876), .B2(new_n1018), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1028), .A2(new_n984), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n1027), .A2(new_n758), .A3(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n984), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n876), .A2(KEYINPUT45), .A3(new_n1018), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1031), .A2(new_n983), .A3(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G1966), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(KEYINPUT121), .A3(new_n1034), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n1021), .A2(new_n1030), .A3(new_n1035), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(G8), .ZN(new_n1038));
  NOR2_X1   g613(.A1(G168), .A2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(KEYINPUT51), .B1(new_n1039), .B2(KEYINPUT122), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1037), .A2(new_n1040), .A3(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT116), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1044), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n984), .B1(new_n983), .B2(KEYINPUT116), .ZN(new_n1046));
  INV_X1    g621(.A(G2078), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1045), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n1049));
  NOR2_X1   g624(.A1(new_n498), .A2(new_n502), .ZN(new_n1050));
  AOI21_X1  g625(.A(G1384), .B1(new_n1050), .B2(new_n867), .ZN(new_n1051));
  AOI21_X1  g626(.A(KEYINPUT117), .B1(new_n1051), .B2(new_n1022), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1026), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1029), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  XOR2_X1   g629(.A(KEYINPUT123), .B(G1961), .Z(new_n1055));
  AOI22_X1  g630(.A1(new_n1048), .A2(new_n1049), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n1020), .A2(KEYINPUT53), .A3(new_n1047), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1058), .A2(KEYINPUT62), .A3(G171), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1036), .A2(G8), .A3(G286), .ZN(new_n1060));
  OAI211_X1 g635(.A(G8), .B(new_n1041), .C1(new_n1036), .C2(G286), .ZN(new_n1061));
  NAND4_X1  g636(.A1(new_n1043), .A2(new_n1059), .A3(new_n1060), .A4(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT125), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT55), .ZN(new_n1064));
  NOR3_X1   g639(.A1(G166), .A2(new_n1064), .A3(new_n1038), .ZN(new_n1065));
  AOI21_X1  g640(.A(KEYINPUT55), .B1(G303), .B2(G8), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1054), .A2(G2090), .ZN(new_n1068));
  AOI21_X1  g643(.A(G1971), .B1(new_n1045), .B2(new_n1046), .ZN(new_n1069));
  OAI211_X1 g644(.A(new_n1067), .B(G8), .C1(new_n1068), .C2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n588), .A2(G1976), .A3(new_n589), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT118), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND4_X1  g648(.A1(new_n588), .A2(KEYINPUT118), .A3(G1976), .A4(new_n589), .ZN(new_n1074));
  AND2_X1   g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n876), .A2(new_n1018), .ZN(new_n1077));
  NOR2_X1   g652(.A1(new_n984), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1038), .ZN(new_n1079));
  INV_X1    g654(.A(G1976), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1080), .B1(new_n590), .B2(new_n591), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1075), .A2(new_n1076), .A3(new_n1079), .A4(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n1073), .A2(new_n1079), .A3(new_n1074), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(KEYINPUT52), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT49), .ZN(new_n1085));
  AND2_X1   g660(.A1(new_n601), .A2(G1981), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n601), .A2(G1981), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OR2_X1    g663(.A1(new_n601), .A2(G1981), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n601), .A2(G1981), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1089), .A2(KEYINPUT49), .A3(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1079), .A2(new_n1088), .A3(new_n1091), .ZN(new_n1092));
  AND4_X1   g667(.A1(new_n1070), .A2(new_n1082), .A3(new_n1084), .A4(new_n1092), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1067), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1028), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1095), .A2(new_n1031), .A3(new_n1023), .ZN(new_n1096));
  NOR2_X1   g671(.A1(new_n1096), .A2(G2090), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1069), .A2(new_n1097), .ZN(new_n1098));
  OAI21_X1  g673(.A(new_n1094), .B1(new_n1098), .B2(new_n1038), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1063), .B1(new_n1093), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1070), .A2(new_n1082), .A3(new_n1084), .A4(new_n1092), .ZN(new_n1101));
  OR2_X1    g676(.A1(new_n1069), .A2(new_n1097), .ZN(new_n1102));
  AOI21_X1  g677(.A(new_n1067), .B1(new_n1102), .B2(G8), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1101), .A2(KEYINPUT125), .A3(new_n1103), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n1062), .B1(new_n1100), .B2(new_n1104), .ZN(new_n1105));
  XNOR2_X1  g680(.A(new_n575), .B(KEYINPUT57), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1106), .ZN(new_n1107));
  XNOR2_X1  g682(.A(KEYINPUT56), .B(G2072), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1045), .A2(new_n1046), .A3(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1096), .A2(new_n783), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1107), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1348), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1054), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1078), .A2(new_n991), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n647), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1109), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1111), .B1(new_n1115), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g692(.A(G1348), .B1(new_n1027), .B2(new_n1029), .ZN(new_n1118));
  INV_X1    g693(.A(new_n1114), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1118), .A2(new_n637), .A3(new_n1119), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT60), .B1(new_n1115), .B2(new_n1120), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT61), .ZN(new_n1122));
  AND3_X1   g697(.A1(new_n1109), .A2(new_n1107), .A3(new_n1110), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1122), .B1(new_n1123), .B2(new_n1111), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1125), .A2(new_n1106), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1126), .A2(KEYINPUT61), .A3(new_n1116), .ZN(new_n1127));
  NOR2_X1   g702(.A1(new_n647), .A2(KEYINPUT60), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1113), .A2(new_n1114), .A3(new_n1128), .ZN(new_n1129));
  NAND4_X1  g704(.A1(new_n1121), .A2(new_n1124), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  NOR2_X1   g705(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1131));
  AND2_X1   g706(.A1(KEYINPUT58), .A2(G1341), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n1078), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  AOI21_X1  g708(.A(KEYINPUT116), .B1(new_n983), .B2(new_n1032), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n1031), .B1(new_n1019), .B2(new_n1044), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1133), .B1(new_n1136), .B2(new_n986), .ZN(new_n1137));
  OAI21_X1  g712(.A(KEYINPUT59), .B1(new_n1137), .B2(new_n645), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n1139));
  NOR3_X1   g714(.A1(new_n1134), .A2(new_n1135), .A3(G1996), .ZN(new_n1140));
  OAI211_X1 g715(.A(new_n1139), .B(new_n556), .C1(new_n1140), .C2(new_n1133), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1138), .A2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(new_n1142), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1117), .B1(new_n1130), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(KEYINPUT54), .B1(new_n1058), .B2(G171), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n465), .A2(G2105), .ZN(new_n1147));
  AND3_X1   g722(.A1(new_n481), .A2(KEYINPUT53), .A3(new_n1047), .ZN(new_n1148));
  NAND4_X1  g723(.A1(new_n1146), .A2(G40), .A3(new_n1147), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g724(.A(G301), .B1(new_n1056), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1145), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1058), .A2(G171), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1056), .A2(G301), .A3(new_n1149), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(KEYINPUT124), .A3(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT54), .ZN(new_n1156));
  OR2_X1    g731(.A1(new_n1154), .A2(KEYINPUT124), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1155), .A2(new_n1156), .A3(new_n1157), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1144), .A2(new_n1152), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1043), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1153), .B1(new_n1160), .B2(KEYINPUT62), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g737(.A(new_n1105), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  NAND3_X1  g738(.A1(new_n1092), .A2(new_n592), .A3(new_n1080), .ZN(new_n1164));
  AND3_X1   g739(.A1(new_n1164), .A2(KEYINPUT120), .A3(new_n1089), .ZN(new_n1165));
  AOI21_X1  g740(.A(KEYINPUT120), .B1(new_n1164), .B2(new_n1089), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1167));
  INV_X1    g742(.A(new_n1167), .ZN(new_n1168));
  NOR2_X1   g743(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1169));
  NOR4_X1   g744(.A1(new_n1165), .A2(new_n1166), .A3(new_n1168), .A4(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(KEYINPUT63), .ZN(new_n1171));
  AND2_X1   g746(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1172));
  NAND4_X1  g747(.A1(new_n1172), .A2(new_n1099), .A3(new_n1070), .A4(new_n1082), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1036), .A2(G8), .A3(G168), .ZN(new_n1174));
  OAI21_X1  g749(.A(new_n1171), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  INV_X1    g750(.A(new_n1174), .ZN(new_n1176));
  OAI21_X1  g751(.A(G8), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1177));
  AOI21_X1  g752(.A(new_n1171), .B1(new_n1177), .B2(new_n1094), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1093), .A2(new_n1176), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1170), .B1(new_n1175), .B2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1172), .A2(new_n1082), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n1180), .B1(new_n1070), .B2(new_n1181), .ZN(new_n1182));
  OAI211_X1 g757(.A(new_n1013), .B(new_n1015), .C1(new_n1163), .C2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1181), .A2(new_n1070), .ZN(new_n1185));
  AOI211_X1 g760(.A(new_n1185), .B(new_n1170), .C1(new_n1175), .C2(new_n1179), .ZN(new_n1186));
  INV_X1    g761(.A(new_n1129), .ZN(new_n1187));
  NAND3_X1  g762(.A1(new_n1113), .A2(new_n647), .A3(new_n1114), .ZN(new_n1188));
  OAI21_X1  g763(.A(new_n637), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1189));
  NAND2_X1  g764(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  AOI21_X1  g765(.A(new_n1187), .B1(new_n1190), .B2(KEYINPUT60), .ZN(new_n1191));
  NAND4_X1  g766(.A1(new_n1191), .A2(new_n1142), .A3(new_n1127), .A4(new_n1124), .ZN(new_n1192));
  AOI21_X1  g767(.A(new_n1151), .B1(new_n1192), .B2(new_n1117), .ZN(new_n1193));
  AOI21_X1  g768(.A(new_n1161), .B1(new_n1193), .B2(new_n1158), .ZN(new_n1194));
  OAI21_X1  g769(.A(new_n1186), .B1(new_n1194), .B2(new_n1105), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1013), .B1(new_n1195), .B2(new_n1015), .ZN(new_n1196));
  OAI21_X1  g771(.A(new_n1012), .B1(new_n1184), .B2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g772(.A(G227), .ZN(new_n1199));
  AND3_X1   g773(.A1(new_n899), .A2(new_n680), .A3(new_n1199), .ZN(new_n1200));
  INV_X1    g774(.A(G319), .ZN(new_n1201));
  NOR2_X1   g775(.A1(G229), .A2(new_n1201), .ZN(new_n1202));
  NAND3_X1  g776(.A1(new_n1200), .A2(new_n1202), .A3(new_n977), .ZN(G225));
  INV_X1    g777(.A(G225), .ZN(G308));
endmodule


