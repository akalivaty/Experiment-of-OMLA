//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 0 0 1 0 1 1 1 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 1 0 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:07 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1259, new_n1260,
    new_n1261, new_n1262, new_n1263, new_n1265, new_n1266, new_n1267,
    new_n1268, new_n1269, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1346, new_n1347,
    new_n1348, new_n1349, new_n1350, new_n1351, new_n1352;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  XNOR2_X1  g0012(.A(KEYINPUT64), .B(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G238), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G77), .B2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G58), .A2(G232), .ZN(new_n219));
  NAND4_X1  g0019(.A1(new_n216), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n209), .B1(new_n215), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n207), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(new_n201), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n212), .B1(KEYINPUT1), .B2(new_n221), .C1(new_n224), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n221), .ZN(G361));
  XNOR2_X1  g0028(.A(G238), .B(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G232), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(new_n233), .B(new_n236), .Z(G358));
  XOR2_X1   g0037(.A(G87), .B(G97), .Z(new_n238));
  XNOR2_X1  g0038(.A(G107), .B(G116), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(KEYINPUT65), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n202), .A2(G68), .ZN(new_n242));
  INV_X1    g0042(.A(G68), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n243), .A2(G50), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G58), .B(G77), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n241), .B(new_n247), .ZN(G351));
  INV_X1    g0048(.A(KEYINPUT3), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT3), .A2(G33), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G223), .A3(G1698), .ZN(new_n254));
  INV_X1    g0054(.A(G77), .ZN(new_n255));
  INV_X1    g0055(.A(G1698), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n253), .A2(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G222), .ZN(new_n258));
  OAI221_X1 g0058(.A(new_n254), .B1(new_n255), .B2(new_n253), .C1(new_n257), .C2(new_n258), .ZN(new_n259));
  AOI21_X1  g0059(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G274), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n263));
  NOR3_X1   g0063(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(G41), .ZN(new_n266));
  OAI211_X1 g0066(.A(G1), .B(G13), .C1(new_n250), .C2(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT66), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT66), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n267), .A2(new_n270), .A3(new_n263), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G226), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n261), .A2(new_n265), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n274), .A2(G200), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n261), .A2(G190), .A3(new_n265), .A4(new_n273), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n202), .B1(new_n206), .B2(G20), .ZN(new_n277));
  XNOR2_X1  g0077(.A(new_n277), .B(KEYINPUT68), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n279));
  NAND3_X1  g0079(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(new_n222), .A3(new_n280), .ZN(new_n281));
  OAI22_X1  g0081(.A1(new_n278), .A2(new_n281), .B1(G50), .B2(new_n279), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n280), .A2(new_n222), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n207), .A2(G33), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT67), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n207), .A2(KEYINPUT67), .A3(G33), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n286), .A2(new_n289), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(G20), .A2(G33), .ZN(new_n292));
  AOI22_X1  g0092(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n284), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n282), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT9), .ZN(new_n296));
  AND3_X1   g0096(.A1(new_n275), .A2(new_n276), .A3(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT10), .ZN(new_n298));
  INV_X1    g0098(.A(KEYINPUT9), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n299), .B1(new_n282), .B2(new_n294), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n300), .B(KEYINPUT70), .ZN(new_n301));
  NAND3_X1  g0101(.A1(new_n297), .A2(new_n298), .A3(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n275), .A2(new_n276), .A3(new_n296), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT70), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n300), .B(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(KEYINPUT10), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n302), .A2(new_n306), .ZN(new_n307));
  OR2_X1    g0107(.A1(new_n274), .A2(G179), .ZN(new_n308));
  INV_X1    g0108(.A(new_n295), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n274), .A2(new_n310), .ZN(new_n311));
  AND3_X1   g0111(.A1(new_n308), .A2(new_n309), .A3(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n206), .A2(G20), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(G77), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n281), .A2(new_n316), .B1(G77), .B2(new_n279), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n286), .A2(new_n292), .B1(G20), .B2(G77), .ZN(new_n318));
  XNOR2_X1  g0118(.A(KEYINPUT15), .B(G87), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n318), .B1(new_n287), .B2(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n320), .B2(new_n283), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n253), .A2(G238), .A3(G1698), .ZN(new_n322));
  INV_X1    g0122(.A(G107), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n322), .B1(new_n323), .B2(new_n253), .C1(new_n257), .C2(new_n230), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n260), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n272), .A2(G244), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n325), .A2(new_n265), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n327), .A2(KEYINPUT69), .ZN(new_n328));
  INV_X1    g0128(.A(KEYINPUT69), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n325), .A2(new_n329), .A3(new_n265), .A4(new_n326), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G179), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n321), .B1(new_n331), .B2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n328), .A2(new_n310), .A3(new_n330), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G200), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n321), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G190), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n328), .B2(new_n330), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n314), .A2(new_n336), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G226), .A2(G1698), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n230), .B2(G1698), .ZN(new_n344));
  AOI22_X1  g0144(.A1(new_n344), .A2(new_n253), .B1(G33), .B2(G97), .ZN(new_n345));
  OAI21_X1  g0145(.A(new_n265), .B1(new_n345), .B2(new_n267), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n214), .B1(new_n269), .B2(new_n271), .ZN(new_n347));
  OAI21_X1  g0147(.A(KEYINPUT13), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n253), .ZN(new_n349));
  NAND2_X1  g0149(.A1(G33), .A2(G97), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n264), .B1(new_n351), .B2(new_n260), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT13), .ZN(new_n353));
  INV_X1    g0153(.A(new_n271), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n270), .B1(new_n267), .B2(new_n263), .ZN(new_n355));
  OAI21_X1  g0155(.A(G238), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n352), .A2(new_n353), .A3(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n348), .A2(KEYINPUT71), .A3(new_n357), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT71), .ZN(new_n359));
  OAI211_X1 g0159(.A(new_n359), .B(KEYINPUT13), .C1(new_n346), .C2(new_n347), .ZN(new_n360));
  AND2_X1   g0160(.A1(KEYINPUT73), .A2(G169), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n358), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(KEYINPUT14), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT14), .ZN(new_n364));
  NAND4_X1  g0164(.A1(new_n358), .A2(new_n364), .A3(new_n360), .A4(new_n361), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n348), .A2(G179), .A3(new_n357), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n289), .A2(G77), .A3(new_n290), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n213), .A2(G20), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n292), .A2(G50), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n368), .A2(new_n369), .A3(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT72), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n371), .A2(new_n372), .A3(new_n283), .ZN(new_n373));
  INV_X1    g0173(.A(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n372), .B1(new_n371), .B2(new_n283), .ZN(new_n375));
  OAI21_X1  g0175(.A(KEYINPUT11), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n371), .A2(new_n283), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT72), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT11), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n378), .A2(new_n379), .A3(new_n373), .ZN(new_n380));
  INV_X1    g0180(.A(new_n281), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n381), .A2(G68), .A3(new_n315), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT12), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n279), .B2(G68), .ZN(new_n384));
  INV_X1    g0184(.A(G13), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n385), .A2(G1), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n213), .A2(KEYINPUT12), .A3(G20), .A4(new_n386), .ZN(new_n387));
  AND3_X1   g0187(.A1(new_n382), .A2(new_n384), .A3(new_n387), .ZN(new_n388));
  AND3_X1   g0188(.A1(new_n376), .A2(new_n380), .A3(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n367), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n358), .A2(G200), .A3(new_n360), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n348), .A2(G190), .A3(new_n357), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(G58), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n225), .B1(new_n213), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n292), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n251), .A2(new_n207), .A3(new_n252), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT74), .ZN(new_n401));
  AND2_X1   g0201(.A1(KEYINPUT3), .A2(G33), .ZN(new_n402));
  NOR2_X1   g0202(.A1(KEYINPUT3), .A2(G33), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n401), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n251), .A2(KEYINPUT74), .A3(new_n252), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n405), .A3(new_n207), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n400), .B1(new_n406), .B2(new_n399), .ZN(new_n407));
  OAI211_X1 g0207(.A(KEYINPUT16), .B(new_n397), .C1(new_n407), .C2(new_n243), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT16), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n396), .A2(G20), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n292), .A2(G159), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n398), .A2(new_n399), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n402), .A2(new_n403), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n414), .A2(KEYINPUT7), .A3(new_n207), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n213), .B1(new_n413), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n409), .B1(new_n412), .B2(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n408), .A2(new_n417), .A3(new_n283), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n285), .B1(new_n206), .B2(G20), .ZN(new_n419));
  INV_X1    g0219(.A(new_n279), .ZN(new_n420));
  AOI22_X1  g0220(.A1(new_n419), .A2(new_n381), .B1(new_n420), .B2(new_n285), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n418), .A2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n265), .B1(new_n230), .B2(new_n268), .ZN(new_n423));
  INV_X1    g0223(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n253), .A2(G223), .A3(new_n256), .ZN(new_n425));
  NAND2_X1  g0225(.A1(G33), .A2(G87), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  OAI211_X1 g0227(.A(G226), .B(G1698), .C1(new_n402), .C2(new_n403), .ZN(new_n428));
  INV_X1    g0228(.A(KEYINPUT75), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  NAND4_X1  g0230(.A1(new_n253), .A2(KEYINPUT75), .A3(G226), .A4(G1698), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n427), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI211_X1 g0232(.A(new_n424), .B(G179), .C1(new_n267), .C2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n427), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n430), .A2(new_n431), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n267), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g0236(.A(G169), .B1(new_n436), .B2(new_n423), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n422), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n439), .A2(KEYINPUT18), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT18), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n422), .A2(new_n438), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n424), .B(G190), .C1(new_n267), .C2(new_n432), .ZN(new_n444));
  OAI21_X1  g0244(.A(G200), .B1(new_n436), .B2(new_n423), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n446), .A2(KEYINPUT17), .A3(new_n418), .A4(new_n421), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n418), .A2(new_n444), .A3(new_n421), .A4(new_n445), .ZN(new_n448));
  INV_X1    g0248(.A(KEYINPUT17), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  NOR2_X1   g0251(.A1(new_n443), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n342), .A2(new_n391), .A3(new_n394), .A4(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n292), .A2(G77), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT6), .ZN(new_n455));
  INV_X1    g0255(.A(G97), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n455), .A2(new_n456), .A3(G107), .ZN(new_n457));
  XNOR2_X1  g0257(.A(G97), .B(G107), .ZN(new_n458));
  AOI21_X1  g0258(.A(new_n457), .B1(new_n455), .B2(new_n458), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n454), .B1(new_n459), .B2(new_n207), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n323), .B1(new_n413), .B2(new_n415), .ZN(new_n461));
  OAI21_X1  g0261(.A(new_n283), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n420), .A2(new_n456), .ZN(new_n463));
  OR3_X1    g0263(.A1(new_n250), .A2(KEYINPUT76), .A3(G1), .ZN(new_n464));
  OAI21_X1  g0264(.A(KEYINPUT76), .B1(new_n250), .B2(G1), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g0266(.A1(new_n466), .A2(new_n281), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(G97), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n462), .A2(new_n463), .A3(new_n468), .ZN(new_n469));
  XNOR2_X1  g0269(.A(KEYINPUT5), .B(G41), .ZN(new_n470));
  INV_X1    g0270(.A(G45), .ZN(new_n471));
  NOR2_X1   g0271(.A1(new_n471), .A2(G1), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n470), .A2(new_n267), .A3(G274), .A4(new_n472), .ZN(new_n473));
  AND2_X1   g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  NOR2_X1   g0274(.A1(KEYINPUT5), .A2(G41), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n472), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n267), .ZN(new_n477));
  INV_X1    g0277(.A(G257), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n473), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  OAI211_X1 g0279(.A(G244), .B(new_n256), .C1(new_n402), .C2(new_n403), .ZN(new_n480));
  INV_X1    g0280(.A(KEYINPUT4), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n253), .A2(KEYINPUT4), .A3(G244), .A4(new_n256), .ZN(new_n483));
  NAND2_X1  g0283(.A1(G33), .A2(G283), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n253), .A2(G250), .A3(G1698), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n482), .A2(new_n483), .A3(new_n484), .A4(new_n485), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n479), .B1(new_n486), .B2(new_n260), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n469), .B1(G190), .B2(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(new_n479), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n486), .A2(KEYINPUT77), .A3(new_n260), .ZN(new_n490));
  AOI21_X1  g0290(.A(KEYINPUT77), .B1(new_n486), .B2(new_n260), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n489), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(G200), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n488), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(new_n332), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n495));
  OR2_X1    g0295(.A1(new_n487), .A2(G169), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(new_n496), .A3(new_n469), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n494), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n214), .A2(new_n256), .ZN(new_n499));
  INV_X1    g0299(.A(G244), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G1698), .ZN(new_n501));
  OAI211_X1 g0301(.A(new_n499), .B(new_n501), .C1(new_n402), .C2(new_n403), .ZN(new_n502));
  NAND2_X1  g0302(.A1(G33), .A2(G116), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT78), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n502), .A2(KEYINPUT78), .A3(new_n503), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n267), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n267), .A2(G274), .A3(new_n472), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n206), .A2(G45), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n267), .A2(G250), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NOR3_X1   g0312(.A1(new_n508), .A2(G179), .A3(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n507), .ZN(new_n514));
  AOI21_X1  g0314(.A(KEYINPUT78), .B1(new_n502), .B2(new_n503), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n260), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g0316(.A(new_n512), .ZN(new_n517));
  AOI21_X1  g0317(.A(G169), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  OAI21_X1  g0318(.A(KEYINPUT79), .B1(new_n513), .B2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT81), .ZN(new_n520));
  INV_X1    g0320(.A(new_n319), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n521), .A2(new_n279), .ZN(new_n522));
  NAND3_X1  g0322(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n523), .A2(new_n207), .ZN(new_n524));
  INV_X1    g0324(.A(G87), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n525), .A2(new_n456), .A3(new_n323), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT80), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n524), .A2(KEYINPUT80), .A3(new_n526), .ZN(new_n530));
  OAI211_X1 g0330(.A(new_n207), .B(G68), .C1(new_n402), .C2(new_n403), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n532), .B1(new_n287), .B2(new_n456), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n529), .A2(new_n530), .A3(new_n531), .A4(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n522), .B1(new_n534), .B2(new_n283), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n467), .A2(new_n521), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n520), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT80), .B1(new_n524), .B2(new_n526), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n283), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n522), .ZN(new_n541));
  AND4_X1   g0341(.A1(new_n520), .A2(new_n540), .A3(new_n541), .A4(new_n536), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n516), .A2(new_n332), .A3(new_n517), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT79), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n508), .A2(new_n512), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n544), .B(new_n545), .C1(new_n546), .C2(G169), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n519), .A2(new_n543), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n516), .A2(G190), .A3(new_n517), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n467), .A2(G87), .ZN(new_n550));
  AND3_X1   g0350(.A1(new_n540), .A2(new_n541), .A3(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(new_n549), .B(new_n551), .C1(new_n546), .C2(new_n337), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n484), .B(new_n207), .C1(G33), .C2(new_n456), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT83), .ZN(new_n555));
  INV_X1    g0355(.A(G116), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G20), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n283), .A2(new_n555), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(new_n555), .B1(new_n283), .B2(new_n557), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n554), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  INV_X1    g0360(.A(KEYINPUT20), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  OAI211_X1 g0362(.A(KEYINPUT20), .B(new_n554), .C1(new_n558), .C2(new_n559), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n420), .A2(new_n556), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n467), .A2(G116), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n564), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(G303), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n267), .B1(new_n414), .B2(new_n568), .ZN(new_n569));
  NOR2_X1   g0369(.A1(G257), .A2(G1698), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n256), .A2(G264), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n253), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n569), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n476), .A2(G270), .A3(new_n267), .ZN(new_n574));
  INV_X1    g0374(.A(KEYINPUT82), .ZN(new_n575));
  AND3_X1   g0375(.A1(new_n574), .A2(new_n473), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g0376(.A(new_n575), .B1(new_n574), .B2(new_n473), .ZN(new_n577));
  OAI21_X1  g0377(.A(new_n573), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n567), .A2(KEYINPUT21), .A3(G169), .A4(new_n578), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n381), .A2(new_n464), .A3(new_n465), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n565), .B1(new_n580), .B2(new_n556), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n562), .B2(new_n563), .ZN(new_n582));
  OAI211_X1 g0382(.A(G190), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n583));
  INV_X1    g0383(.A(new_n578), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n337), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n578), .A2(G169), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n586), .B1(new_n587), .B2(new_n582), .ZN(new_n588));
  OAI211_X1 g0388(.A(G179), .B(new_n573), .C1(new_n576), .C2(new_n577), .ZN(new_n589));
  INV_X1    g0389(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n567), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n579), .A2(new_n585), .A3(new_n588), .A4(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n503), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n207), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n323), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n253), .A2(new_n207), .A3(G87), .ZN(new_n599));
  AND2_X1   g0399(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n599), .A2(KEYINPUT22), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(KEYINPUT24), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n284), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  OAI211_X1 g0404(.A(KEYINPUT24), .B(new_n598), .C1(new_n600), .C2(new_n601), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n420), .A2(new_n323), .ZN(new_n606));
  XOR2_X1   g0406(.A(new_n606), .B(KEYINPUT25), .Z(new_n607));
  INV_X1    g0407(.A(KEYINPUT84), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n467), .A2(G107), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n607), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n580), .A2(new_n323), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n606), .B(KEYINPUT25), .ZN(new_n612));
  OAI21_X1  g0412(.A(KEYINPUT84), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  AOI22_X1  g0413(.A1(new_n604), .A2(new_n605), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n476), .A2(G264), .A3(new_n267), .ZN(new_n615));
  NOR2_X1   g0415(.A1(G250), .A2(G1698), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n616), .B1(new_n478), .B2(G1698), .ZN(new_n617));
  AOI22_X1  g0417(.A1(new_n617), .A2(new_n253), .B1(G33), .B2(G294), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n260), .B1(new_n618), .B2(KEYINPUT85), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n617), .A2(new_n253), .ZN(new_n620));
  NAND2_X1  g0420(.A1(G33), .A2(G294), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(KEYINPUT85), .A3(new_n621), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n473), .B(new_n615), .C1(new_n619), .C2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(KEYINPUT86), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n620), .A2(new_n621), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT85), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n618), .A2(KEYINPUT85), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n627), .A2(new_n628), .A3(new_n260), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT86), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n473), .A4(new_n615), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n624), .A2(new_n631), .A3(G169), .ZN(new_n632));
  INV_X1    g0432(.A(new_n615), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n267), .B1(new_n625), .B2(new_n626), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n634), .B2(new_n628), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n635), .A2(G179), .A3(new_n473), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n614), .B1(new_n632), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(G190), .B1(new_n624), .B2(new_n631), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n623), .A2(new_n337), .ZN(new_n640));
  INV_X1    g0440(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n614), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n593), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NOR4_X1   g0443(.A1(new_n453), .A2(new_n498), .A3(new_n553), .A4(new_n643), .ZN(G372));
  NAND2_X1  g0444(.A1(new_n512), .A2(KEYINPUT87), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT87), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n509), .A2(new_n511), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n310), .B1(new_n648), .B2(new_n508), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n535), .A2(new_n536), .ZN(new_n650));
  NAND3_X1  g0450(.A1(new_n649), .A2(new_n544), .A3(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(G200), .B1(new_n648), .B2(new_n508), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n652), .A2(new_n549), .A3(new_n551), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n642), .A2(new_n497), .A3(new_n494), .A4(new_n653), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n579), .A2(new_n588), .A3(new_n591), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n637), .A2(new_n655), .ZN(new_n656));
  OAI21_X1  g0456(.A(new_n651), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n651), .A2(new_n653), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n495), .A2(new_n496), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT88), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n495), .A2(KEYINPUT88), .A3(new_n496), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n659), .A2(new_n662), .A3(new_n469), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT89), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n548), .A2(new_n552), .ZN(new_n668));
  AND3_X1   g0468(.A1(new_n495), .A2(new_n496), .A3(new_n469), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n668), .A2(KEYINPUT26), .A3(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(KEYINPUT89), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n664), .A2(new_n671), .A3(new_n665), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n667), .A2(new_n670), .A3(new_n672), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n453), .B1(new_n658), .B2(new_n673), .ZN(new_n674));
  XOR2_X1   g0474(.A(new_n674), .B(KEYINPUT90), .Z(new_n675));
  INV_X1    g0475(.A(new_n443), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n336), .A2(new_n394), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n677), .A2(new_n391), .ZN(new_n678));
  OAI21_X1  g0478(.A(new_n676), .B1(new_n678), .B2(new_n451), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n307), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(new_n313), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n675), .A2(new_n682), .ZN(G369));
  NAND2_X1  g0483(.A1(new_n604), .A2(new_n605), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n610), .A2(new_n613), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n624), .A2(new_n631), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(new_n339), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n686), .B1(new_n688), .B2(new_n640), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n637), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n386), .A2(new_n207), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(KEYINPUT27), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n692), .A2(new_n693), .A3(G213), .ZN(new_n694));
  INV_X1    g0494(.A(G343), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n690), .B1(new_n614), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n698), .B1(new_n638), .B2(new_n697), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n582), .A2(new_n697), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n655), .A2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n701), .B1(new_n592), .B2(new_n700), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n702), .A2(G330), .ZN(new_n703));
  INV_X1    g0503(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n699), .A2(new_n704), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n655), .A2(new_n697), .ZN(new_n706));
  AOI22_X1  g0506(.A1(new_n690), .A2(new_n706), .B1(new_n637), .B2(new_n697), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n705), .A2(new_n707), .ZN(G399));
  NAND3_X1  g0508(.A1(new_n210), .A2(KEYINPUT91), .A3(new_n266), .ZN(new_n709));
  INV_X1    g0509(.A(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(KEYINPUT91), .B1(new_n210), .B2(new_n266), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n526), .A2(G116), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NOR3_X1   g0514(.A1(new_n712), .A2(new_n206), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(new_n226), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n715), .B1(new_n716), .B2(new_n712), .ZN(new_n717));
  XNOR2_X1  g0517(.A(KEYINPUT92), .B(KEYINPUT28), .ZN(new_n718));
  XNOR2_X1  g0518(.A(new_n717), .B(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n696), .B1(new_n673), .B2(new_n658), .ZN(new_n720));
  OAI21_X1  g0520(.A(KEYINPUT93), .B1(new_n720), .B2(KEYINPUT29), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n672), .A2(new_n670), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n671), .B1(new_n664), .B2(new_n665), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n658), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n697), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT93), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT29), .ZN(new_n727));
  NAND3_X1  g0527(.A1(new_n725), .A2(new_n726), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT94), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n548), .A2(new_n669), .A3(new_n552), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n730), .A2(new_n665), .ZN(new_n731));
  INV_X1    g0531(.A(new_n469), .ZN(new_n732));
  AOI21_X1  g0532(.A(new_n732), .B1(new_n660), .B2(new_n661), .ZN(new_n733));
  NAND4_X1  g0533(.A1(new_n733), .A2(KEYINPUT26), .A3(new_n659), .A4(new_n663), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n697), .B1(new_n735), .B2(new_n657), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n729), .B1(new_n736), .B2(new_n727), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n731), .A2(new_n734), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n696), .B1(new_n658), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g0539(.A1(new_n739), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n740));
  AOI22_X1  g0540(.A1(new_n721), .A2(new_n728), .B1(new_n737), .B2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(G330), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n553), .A2(new_n498), .A3(new_n696), .ZN(new_n743));
  NOR3_X1   g0543(.A1(new_n689), .A2(new_n592), .A3(new_n637), .ZN(new_n744));
  INV_X1    g0544(.A(KEYINPUT30), .ZN(new_n745));
  NAND3_X1  g0545(.A1(new_n546), .A2(new_n635), .A3(new_n487), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n745), .B1(new_n746), .B2(new_n589), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n615), .B1(new_n619), .B2(new_n622), .ZN(new_n748));
  NOR3_X1   g0548(.A1(new_n748), .A2(new_n512), .A3(new_n508), .ZN(new_n749));
  NAND4_X1  g0549(.A1(new_n749), .A2(KEYINPUT30), .A3(new_n590), .A4(new_n487), .ZN(new_n750));
  AND2_X1   g0550(.A1(new_n645), .A2(new_n647), .ZN(new_n751));
  AOI21_X1  g0551(.A(G179), .B1(new_n751), .B2(new_n516), .ZN(new_n752));
  NAND4_X1  g0552(.A1(new_n492), .A2(new_n752), .A3(new_n623), .A4(new_n578), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n747), .A2(new_n750), .A3(new_n753), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(new_n696), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n743), .A2(new_n744), .B1(new_n756), .B2(KEYINPUT31), .ZN(new_n757));
  INV_X1    g0557(.A(KEYINPUT31), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n742), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n741), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n719), .B1(new_n761), .B2(G1), .ZN(G364));
  NOR2_X1   g0562(.A1(new_n385), .A2(G20), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n206), .B1(new_n763), .B2(G45), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n712), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n704), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g0567(.A(new_n767), .B1(G330), .B2(new_n702), .ZN(new_n768));
  INV_X1    g0568(.A(new_n766), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n210), .A2(new_n253), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n770), .B1(KEYINPUT95), .B2(G355), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n771), .B1(KEYINPUT95), .B2(G355), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n247), .A2(new_n471), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n404), .A2(new_n405), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  OAI211_X1 g0575(.A(new_n775), .B(new_n210), .C1(G45), .C2(new_n226), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n772), .B1(G116), .B2(new_n210), .C1(new_n773), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(G13), .A2(G33), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT96), .Z(new_n779));
  NOR2_X1   g0579(.A1(new_n779), .A2(G20), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n222), .B1(G20), .B2(new_n310), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n769), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n207), .A2(new_n332), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  NOR3_X1   g0585(.A1(new_n785), .A2(G190), .A3(G200), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NOR3_X1   g0587(.A1(new_n785), .A2(new_n339), .A3(G200), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  OAI221_X1 g0589(.A(new_n253), .B1(new_n787), .B2(new_n255), .C1(new_n395), .C2(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n339), .A2(G179), .A3(G200), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n791), .A2(new_n207), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n207), .A2(G179), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n793), .A2(G190), .A3(G200), .ZN(new_n794));
  OAI22_X1  g0594(.A1(new_n792), .A2(new_n456), .B1(new_n794), .B2(new_n525), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n793), .A2(new_n339), .A3(new_n337), .ZN(new_n796));
  INV_X1    g0596(.A(G159), .ZN(new_n797));
  NOR3_X1   g0597(.A1(new_n796), .A2(KEYINPUT32), .A3(new_n797), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n793), .A2(new_n339), .A3(G200), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(new_n323), .ZN(new_n800));
  NOR4_X1   g0600(.A1(new_n790), .A2(new_n795), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n796), .A2(new_n797), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT32), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n784), .A2(G190), .A3(G200), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n802), .A2(new_n803), .B1(new_n202), .B2(new_n804), .ZN(new_n805));
  NAND3_X1  g0605(.A1(new_n784), .A2(new_n339), .A3(G200), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n805), .B1(G68), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n796), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n786), .A2(G311), .B1(G329), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  OAI211_X1 g0611(.A(new_n810), .B(new_n414), .C1(new_n811), .C2(new_n789), .ZN(new_n812));
  INV_X1    g0612(.A(G317), .ZN(new_n813));
  NAND2_X1  g0613(.A1(new_n813), .A2(KEYINPUT33), .ZN(new_n814));
  OR2_X1    g0614(.A1(new_n813), .A2(KEYINPUT33), .ZN(new_n815));
  NAND3_X1  g0615(.A1(new_n807), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n816), .B1(new_n817), .B2(new_n799), .C1(new_n568), .C2(new_n794), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n812), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n792), .ZN(new_n820));
  INV_X1    g0620(.A(new_n804), .ZN(new_n821));
  AOI22_X1  g0621(.A1(G294), .A2(new_n820), .B1(new_n821), .B2(G326), .ZN(new_n822));
  XOR2_X1   g0622(.A(new_n822), .B(KEYINPUT97), .Z(new_n823));
  AOI22_X1  g0623(.A1(new_n801), .A2(new_n808), .B1(new_n819), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n781), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n783), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g0626(.A(new_n826), .B(KEYINPUT98), .Z(new_n827));
  INV_X1    g0627(.A(new_n780), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n827), .B1(new_n702), .B2(new_n828), .ZN(new_n829));
  AND2_X1   g0629(.A1(new_n768), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G396));
  OAI22_X1  g0631(.A1(new_n804), .A2(new_n568), .B1(new_n794), .B2(new_n323), .ZN(new_n832));
  INV_X1    g0632(.A(new_n799), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(G87), .B2(new_n833), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n253), .B1(new_n788), .B2(G294), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n786), .A2(G116), .B1(G311), .B2(new_n809), .ZN(new_n836));
  AOI22_X1  g0636(.A1(G97), .A2(new_n820), .B1(new_n807), .B2(G283), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n834), .A2(new_n835), .A3(new_n836), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G143), .A2(new_n788), .B1(new_n786), .B2(G159), .ZN(new_n839));
  INV_X1    g0639(.A(G137), .ZN(new_n840));
  INV_X1    g0640(.A(G150), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n839), .B1(new_n840), .B2(new_n804), .C1(new_n841), .C2(new_n806), .ZN(new_n842));
  INV_X1    g0642(.A(KEYINPUT34), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n775), .B1(G132), .B2(new_n809), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n794), .A2(new_n202), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n799), .A2(new_n243), .ZN(new_n847));
  AOI211_X1 g0647(.A(new_n846), .B(new_n847), .C1(G58), .C2(new_n820), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n844), .A2(new_n845), .A3(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n842), .A2(new_n843), .ZN(new_n850));
  OAI21_X1  g0650(.A(new_n838), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(new_n781), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n781), .A2(new_n778), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n852), .B(new_n766), .C1(G77), .C2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n336), .A2(new_n697), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n321), .A2(new_n697), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n335), .B1(new_n341), .B2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n779), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n336), .A2(new_n341), .A3(new_n696), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n724), .A2(new_n862), .ZN(new_n863));
  AND2_X1   g0663(.A1(new_n856), .A2(new_n858), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n863), .B1(new_n720), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(new_n760), .ZN(new_n866));
  OR2_X1    g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n766), .B1(new_n865), .B2(new_n866), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n861), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(new_n869), .ZN(G384));
  NOR2_X1   g0670(.A1(new_n763), .A2(new_n206), .ZN(new_n871));
  INV_X1    g0671(.A(new_n694), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n422), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND4_X1  g0674(.A1(new_n439), .A2(new_n873), .A3(new_n874), .A4(new_n448), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n397), .B1(new_n407), .B2(new_n243), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(new_n409), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n877), .A2(new_n283), .A3(new_n408), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n878), .A2(new_n421), .B1(new_n437), .B2(new_n433), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n694), .B1(new_n878), .B2(new_n421), .ZN(new_n880));
  AND4_X1   g0680(.A1(new_n418), .A2(new_n444), .A3(new_n421), .A4(new_n445), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n875), .B1(new_n882), .B2(new_n874), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n880), .B1(new_n443), .B2(new_n451), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(KEYINPUT102), .B1(new_n755), .B2(new_n758), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT102), .ZN(new_n891));
  AOI211_X1 g0691(.A(new_n891), .B(KEYINPUT31), .C1(new_n754), .C2(new_n696), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n859), .B1(new_n757), .B2(new_n893), .ZN(new_n894));
  NAND4_X1  g0694(.A1(new_n394), .A2(new_n365), .A3(new_n363), .A4(new_n366), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n389), .A2(new_n697), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g0699(.A(new_n896), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n391), .A2(new_n394), .A3(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n895), .A2(KEYINPUT100), .A3(new_n896), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n899), .A2(new_n901), .A3(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n889), .A2(new_n894), .A3(new_n903), .ZN(new_n904));
  XNOR2_X1  g0704(.A(KEYINPUT101), .B(KEYINPUT40), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n743), .A2(new_n744), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n759), .A2(new_n891), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n756), .A2(KEYINPUT31), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n755), .A2(KEYINPUT102), .A3(new_n758), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n906), .A2(new_n907), .A3(new_n908), .A4(new_n909), .ZN(new_n910));
  AND3_X1   g0710(.A1(new_n910), .A2(new_n864), .A3(new_n903), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n422), .B(new_n872), .C1(new_n443), .C2(new_n451), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n439), .A2(new_n873), .A3(new_n448), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT37), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n915), .A2(new_n875), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n917), .A2(new_n886), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n912), .B1(new_n918), .B2(new_n888), .ZN(new_n919));
  AOI22_X1  g0719(.A1(new_n904), .A2(new_n905), .B1(new_n911), .B2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  INV_X1    g0721(.A(new_n910), .ZN(new_n922));
  OR2_X1    g0722(.A1(new_n453), .A2(new_n922), .ZN(new_n923));
  AND2_X1   g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n921), .A2(new_n923), .ZN(new_n925));
  NOR3_X1   g0725(.A1(new_n924), .A2(new_n925), .A3(new_n742), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n721), .A2(new_n728), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n453), .B1(new_n740), .B2(new_n737), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n930), .A2(new_n682), .ZN(new_n931));
  INV_X1    g0731(.A(new_n903), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(new_n863), .B2(new_n856), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n889), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n443), .A2(new_n694), .ZN(new_n935));
  INV_X1    g0735(.A(KEYINPUT39), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n883), .A2(new_n884), .A3(KEYINPUT38), .ZN(new_n937));
  AOI21_X1  g0737(.A(KEYINPUT38), .B1(new_n913), .B2(new_n916), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n936), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n391), .A2(new_n696), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n939), .B(new_n940), .C1(new_n889), .C2(new_n936), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n931), .B(new_n942), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n871), .B1(new_n927), .B2(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n944), .B1(new_n943), .B2(new_n927), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT35), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n459), .A2(new_n946), .ZN(new_n947));
  AOI211_X1 g0747(.A(new_n556), .B(new_n224), .C1(new_n459), .C2(new_n946), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n947), .B1(new_n949), .B2(KEYINPUT99), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT99), .B2(new_n949), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n951), .B(KEYINPUT36), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n716), .B(G77), .C1(new_n395), .C2(new_n213), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n242), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n954), .A2(G1), .A3(new_n385), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n945), .A2(new_n952), .A3(new_n955), .ZN(G367));
  AND2_X1   g0756(.A1(new_n494), .A2(new_n497), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n732), .B2(new_n697), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n733), .A2(new_n663), .A3(new_n696), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n960), .A2(new_n707), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT45), .Z(new_n962));
  NOR2_X1   g0762(.A1(new_n960), .A2(new_n707), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n962), .A2(new_n964), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(new_n705), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n690), .A2(new_n706), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n699), .B2(new_n706), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n704), .A2(KEYINPUT103), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n968), .B(new_n969), .Z(new_n970));
  NAND3_X1  g0770(.A1(new_n966), .A2(new_n761), .A3(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n971), .A2(new_n761), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n712), .B(KEYINPUT41), .Z(new_n974));
  OAI21_X1  g0774(.A(new_n764), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n960), .ZN(new_n976));
  NOR2_X1   g0776(.A1(new_n976), .A2(new_n967), .ZN(new_n977));
  XNOR2_X1  g0777(.A(new_n977), .B(KEYINPUT42), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n497), .B1(new_n976), .B2(new_n638), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n697), .ZN(new_n980));
  OR2_X1    g0780(.A1(new_n551), .A2(new_n697), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n659), .A2(new_n981), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n981), .A2(new_n651), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  AOI22_X1  g0784(.A1(new_n978), .A2(new_n980), .B1(KEYINPUT43), .B2(new_n984), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n984), .A2(KEYINPUT43), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n985), .B(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n705), .A2(new_n976), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n987), .B(new_n988), .Z(new_n989));
  NAND3_X1  g0789(.A1(new_n982), .A2(new_n780), .A3(new_n983), .ZN(new_n990));
  INV_X1    g0790(.A(G311), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n775), .B1(new_n991), .B2(new_n804), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n789), .A2(new_n568), .B1(new_n787), .B2(new_n817), .ZN(new_n993));
  AOI211_X1 g0793(.A(new_n992), .B(new_n993), .C1(G317), .C2(new_n809), .ZN(new_n994));
  INV_X1    g0794(.A(G294), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n792), .A2(new_n323), .B1(new_n806), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(G97), .B2(new_n833), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT46), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n998), .B1(new_n794), .B2(new_n556), .ZN(new_n999));
  INV_X1    g0799(.A(new_n794), .ZN(new_n1000));
  NAND3_X1  g0800(.A1(new_n1000), .A2(KEYINPUT46), .A3(G116), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n994), .A2(new_n997), .A3(new_n999), .A4(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n253), .B1(new_n789), .B2(new_n841), .ZN(new_n1003));
  AOI21_X1  g0803(.A(new_n1003), .B1(G137), .B2(new_n809), .ZN(new_n1004));
  INV_X1    g0804(.A(G143), .ZN(new_n1005));
  OAI22_X1  g0805(.A1(new_n804), .A2(new_n1005), .B1(new_n794), .B2(new_n395), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n792), .A2(new_n243), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n799), .A2(new_n255), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n786), .A2(G50), .B1(new_n807), .B2(G159), .ZN(new_n1010));
  OR2_X1    g0810(.A1(new_n1010), .A2(KEYINPUT105), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(KEYINPUT105), .ZN(new_n1012));
  NAND4_X1  g0812(.A1(new_n1004), .A2(new_n1009), .A3(new_n1011), .A4(new_n1012), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n1002), .A2(new_n1013), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1014), .A2(KEYINPUT47), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1014), .A2(KEYINPUT47), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1015), .A2(new_n781), .A3(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n775), .A2(new_n210), .ZN(new_n1018));
  OAI221_X1 g0818(.A(new_n782), .B1(new_n210), .B2(new_n319), .C1(new_n1018), .C2(new_n236), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(new_n766), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT104), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1017), .A2(new_n1021), .ZN(new_n1022));
  XOR2_X1   g0822(.A(new_n1022), .B(KEYINPUT106), .Z(new_n1023));
  AOI22_X1  g0823(.A1(new_n975), .A2(new_n989), .B1(new_n990), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(G387));
  INV_X1    g0825(.A(new_n712), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1026), .B1(new_n761), .B2(new_n970), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n761), .B2(new_n970), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n233), .A2(G45), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1029), .B(KEYINPUT107), .ZN(new_n1030));
  AOI211_X1 g0830(.A(G45), .B(new_n714), .C1(G68), .C2(G77), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n285), .A2(G50), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1018), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n1035), .B1(G107), .B2(new_n210), .C1(new_n713), .C2(new_n770), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n769), .B1(new_n1036), .B2(new_n782), .ZN(new_n1037));
  OAI21_X1  g0837(.A(new_n1037), .B1(new_n699), .B2(new_n828), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n789), .A2(new_n202), .B1(new_n787), .B2(new_n243), .ZN(new_n1039));
  AOI21_X1  g0839(.A(new_n1039), .B1(G150), .B2(new_n809), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n521), .A2(new_n820), .B1(new_n821), .B2(G159), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n286), .A2(new_n807), .B1(new_n1000), .B2(G77), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n775), .B1(G97), .B2(new_n833), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n774), .B1(G326), .B2(new_n809), .ZN(new_n1045));
  AOI22_X1  g0845(.A1(new_n820), .A2(G283), .B1(new_n1000), .B2(G294), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(G303), .A2(new_n786), .B1(new_n788), .B2(G317), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n1047), .B1(new_n991), .B2(new_n806), .C1(new_n811), .C2(new_n804), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT108), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1046), .B1(new_n1050), .B2(KEYINPUT48), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1051), .B1(KEYINPUT48), .B2(new_n1050), .ZN(new_n1052));
  XNOR2_X1  g0852(.A(new_n1052), .B(KEYINPUT49), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT109), .ZN(new_n1054));
  OAI221_X1 g0854(.A(new_n1045), .B1(new_n556), .B2(new_n799), .C1(new_n1053), .C2(new_n1054), .ZN(new_n1055));
  AND2_X1   g0855(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1044), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1038), .B1(new_n1057), .B2(new_n781), .ZN(new_n1058));
  AOI21_X1  g0858(.A(new_n1058), .B1(new_n765), .B2(new_n970), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1028), .A2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n971), .A2(new_n712), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n966), .B1(new_n761), .B2(new_n970), .ZN(new_n1062));
  OR2_X1    g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n976), .A2(new_n780), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n782), .B1(new_n456), .B2(new_n210), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n1018), .A2(new_n240), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n766), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n788), .A2(G311), .B1(new_n821), .B2(G317), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT52), .Z(new_n1069));
  OAI21_X1  g0869(.A(new_n414), .B1(new_n796), .B2(new_n811), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n800), .B(new_n1070), .C1(G283), .C2(new_n1000), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(G294), .A2(new_n786), .B1(new_n820), .B2(G116), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1073), .B1(new_n568), .B2(new_n806), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT110), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n788), .A2(G159), .B1(new_n821), .B2(G150), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT51), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n792), .A2(new_n255), .B1(new_n806), .B2(new_n202), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n525), .A2(new_n799), .B1(new_n794), .B2(new_n213), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  AOI22_X1  g0880(.A1(new_n786), .A2(new_n286), .B1(G143), .B2(new_n809), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1080), .A2(new_n774), .A3(new_n1081), .ZN(new_n1082));
  OAI22_X1  g0882(.A1(new_n1072), .A2(new_n1075), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1083));
  AOI21_X1  g0883(.A(new_n1067), .B1(new_n1083), .B2(new_n781), .ZN(new_n1084));
  AOI22_X1  g0884(.A1(new_n966), .A2(new_n765), .B1(new_n1064), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1063), .A2(new_n1085), .ZN(G390));
  NOR3_X1   g0886(.A1(new_n453), .A2(new_n922), .A3(new_n742), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n1087), .ZN(new_n1088));
  NAND3_X1  g0888(.A1(new_n930), .A2(new_n682), .A3(new_n1088), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n910), .A2(G330), .A3(new_n864), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1090), .A2(new_n932), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n760), .A2(new_n864), .A3(new_n903), .ZN(new_n1092));
  AND2_X1   g0892(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n697), .B(new_n858), .C1(new_n735), .C2(new_n657), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1094), .A2(new_n856), .ZN(new_n1095));
  INV_X1    g0895(.A(KEYINPUT111), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1094), .A2(KEYINPUT111), .A3(new_n856), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n724), .A2(new_n862), .B1(new_n336), .B2(new_n697), .ZN(new_n1100));
  INV_X1    g0900(.A(new_n1100), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n668), .A2(new_n957), .A3(new_n697), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1102), .A2(new_n643), .B1(new_n758), .B2(new_n755), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n759), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n864), .B(G330), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n932), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n894), .A2(G330), .A3(new_n903), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(new_n1093), .A2(new_n1099), .B1(new_n1101), .B2(new_n1108), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1089), .A2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n1110), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1097), .A2(new_n903), .A3(new_n1098), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n940), .B1(new_n918), .B2(new_n888), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n939), .B1(new_n889), .B2(new_n936), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n933), .B2(new_n940), .ZN(new_n1116));
  NAND3_X1  g0916(.A1(new_n1114), .A2(new_n1116), .A3(new_n1092), .ZN(new_n1117));
  OAI22_X1  g0917(.A1(new_n1100), .A2(new_n932), .B1(new_n391), .B2(new_n696), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n1112), .A2(new_n1113), .B1(new_n1118), .B2(new_n1115), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1117), .B1(new_n1119), .B2(new_n1107), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1026), .B1(new_n1111), .B2(new_n1120), .ZN(new_n1121));
  AND3_X1   g0921(.A1(new_n1114), .A2(new_n1116), .A3(new_n1092), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1107), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1124), .A2(new_n1110), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n765), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n766), .B1(new_n286), .B2(new_n854), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n794), .A2(new_n525), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n414), .B1(new_n796), .B2(new_n995), .C1(new_n789), .C2(new_n556), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n792), .A2(new_n255), .B1(new_n804), .B2(new_n817), .ZN(new_n1131));
  OR4_X1    g0931(.A1(new_n1129), .A2(new_n1130), .A3(new_n847), .A4(new_n1131), .ZN(new_n1132));
  AOI22_X1  g0932(.A1(new_n786), .A2(G97), .B1(new_n807), .B2(G107), .ZN(new_n1133));
  XNOR2_X1  g0933(.A(new_n1133), .B(KEYINPUT112), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(KEYINPUT54), .B(G143), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n253), .B1(new_n787), .B2(new_n1135), .ZN(new_n1136));
  INV_X1    g0936(.A(G132), .ZN(new_n1137));
  INV_X1    g0937(.A(G125), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n789), .A2(new_n1137), .B1(new_n796), .B2(new_n1138), .ZN(new_n1139));
  OAI22_X1  g0939(.A1(new_n792), .A2(new_n797), .B1(new_n806), .B2(new_n840), .ZN(new_n1140));
  INV_X1    g0940(.A(G128), .ZN(new_n1141));
  OAI22_X1  g0941(.A1(new_n804), .A2(new_n1141), .B1(new_n799), .B2(new_n202), .ZN(new_n1142));
  OR4_X1    g0942(.A1(new_n1136), .A2(new_n1139), .A3(new_n1140), .A4(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1000), .A2(G150), .ZN(new_n1144));
  XNOR2_X1  g0944(.A(new_n1144), .B(KEYINPUT53), .ZN(new_n1145));
  OAI22_X1  g0945(.A1(new_n1132), .A2(new_n1134), .B1(new_n1143), .B2(new_n1145), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1128), .B1(new_n1146), .B2(new_n781), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1115), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1147), .B1(new_n1148), .B2(new_n779), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1126), .A2(new_n1127), .A3(new_n1149), .ZN(G378));
  AND3_X1   g0950(.A1(new_n934), .A2(new_n935), .A3(new_n941), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n295), .A2(new_n694), .ZN(new_n1152));
  INV_X1    g0952(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1153), .B1(new_n307), .B2(new_n313), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1154), .ZN(new_n1155));
  AOI211_X1 g0955(.A(new_n1152), .B(new_n312), .C1(new_n302), .C2(new_n306), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1155), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1158), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1160), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1161));
  NAND3_X1  g0961(.A1(new_n1159), .A2(new_n1161), .A3(KEYINPUT116), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1163), .B1(new_n920), .B2(G330), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT115), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1158), .B1(new_n1155), .B2(new_n1157), .ZN(new_n1166));
  NOR3_X1   g0966(.A1(new_n1154), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1165), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1159), .A2(new_n1161), .A3(KEYINPUT115), .A4(KEYINPUT116), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n911), .A2(new_n919), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n910), .A2(new_n864), .A3(new_n903), .ZN(new_n1172));
  AOI21_X1  g0972(.A(KEYINPUT38), .B1(new_n883), .B2(new_n884), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n937), .A2(new_n1173), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n905), .B1(new_n1172), .B2(new_n1174), .ZN(new_n1175));
  AND4_X1   g0975(.A1(G330), .A2(new_n1170), .A3(new_n1171), .A4(new_n1175), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1151), .B1(new_n1164), .B2(new_n1176), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1171), .A2(new_n1175), .A3(G330), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1178), .A2(new_n1162), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n920), .A2(G330), .A3(new_n1170), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1179), .A2(new_n1180), .A3(new_n942), .ZN(new_n1181));
  AOI21_X1  g0981(.A(new_n764), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n250), .A2(new_n266), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT113), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n202), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(new_n266), .B2(new_n775), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n788), .A2(G107), .B1(G283), .B2(new_n809), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n319), .B2(new_n787), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n1007), .B(new_n1188), .C1(G77), .C2(new_n1000), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n804), .A2(new_n556), .B1(new_n799), .B2(new_n395), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G97), .B2(new_n807), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n266), .A3(new_n775), .A4(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT58), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1186), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1184), .B1(G124), .B2(new_n809), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n806), .A2(new_n1137), .B1(new_n804), .B2(new_n1138), .ZN(new_n1196));
  AOI22_X1  g0996(.A1(G128), .A2(new_n788), .B1(new_n786), .B2(G137), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1197), .B1(new_n794), .B2(new_n1135), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n1196), .B(new_n1198), .C1(G150), .C2(new_n820), .ZN(new_n1199));
  INV_X1    g0999(.A(KEYINPUT59), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1195), .B1(new_n797), .B2(new_n799), .C1(new_n1199), .C2(new_n1200), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1199), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n1202), .A2(KEYINPUT59), .ZN(new_n1203));
  OAI221_X1 g1003(.A(new_n1194), .B1(new_n1193), .B2(new_n1192), .C1(new_n1201), .C2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1204), .A2(new_n781), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT114), .ZN(new_n1206));
  AOI211_X1 g1006(.A(new_n769), .B(new_n1206), .C1(new_n202), .C2(new_n853), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1168), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1166), .A2(new_n1167), .A3(new_n1165), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n860), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1207), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(new_n1211), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1182), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1087), .B(new_n681), .C1(new_n928), .C2(new_n929), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n1120), .B2(new_n1109), .ZN(new_n1216));
  INV_X1    g1016(.A(KEYINPUT57), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1217), .B1(new_n1177), .B2(new_n1181), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1026), .B1(new_n1216), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1177), .A2(new_n1181), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1216), .A2(new_n1220), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n1219), .A2(KEYINPUT117), .B1(new_n1221), .B2(new_n1217), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1089), .B1(new_n1124), .B2(new_n1110), .ZN(new_n1223));
  AND3_X1   g1023(.A1(new_n1179), .A2(new_n1180), .A3(new_n942), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n942), .B1(new_n1179), .B2(new_n1180), .ZN(new_n1225));
  OAI21_X1  g1025(.A(KEYINPUT57), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n712), .B1(new_n1223), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT117), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1214), .B1(new_n1222), .B2(new_n1229), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(G375));
  INV_X1    g1031(.A(KEYINPUT118), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1108), .A2(new_n1101), .ZN(new_n1233));
  INV_X1    g1033(.A(new_n1099), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1233), .B1(new_n1234), .B2(new_n1235), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1232), .B1(new_n1215), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n974), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1089), .A2(KEYINPUT118), .A3(new_n1109), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1237), .A2(new_n1238), .A3(new_n1239), .A4(new_n1111), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n932), .A2(new_n778), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n766), .B1(G68), .B2(new_n854), .ZN(new_n1242));
  OAI22_X1  g1042(.A1(new_n806), .A2(new_n556), .B1(new_n804), .B2(new_n995), .ZN(new_n1243));
  AOI21_X1  g1043(.A(new_n1243), .B1(G97), .B2(new_n1000), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n253), .B1(new_n809), .B2(G303), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(G107), .A2(new_n786), .B1(new_n788), .B2(G283), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1008), .B1(new_n521), .B2(new_n820), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1244), .A2(new_n1245), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  OAI22_X1  g1048(.A1(new_n395), .A2(new_n799), .B1(new_n794), .B2(new_n797), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n774), .B1(new_n1141), .B2(new_n796), .C1(new_n787), .C2(new_n841), .ZN(new_n1250));
  AOI211_X1 g1050(.A(new_n1249), .B(new_n1250), .C1(G50), .C2(new_n820), .ZN(new_n1251));
  XNOR2_X1  g1051(.A(new_n1251), .B(KEYINPUT119), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n788), .A2(G137), .ZN(new_n1253));
  OAI221_X1 g1053(.A(new_n1253), .B1(new_n806), .B2(new_n1135), .C1(new_n1137), .C2(new_n804), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1248), .B1(new_n1252), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1242), .B1(new_n1255), .B2(new_n781), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(new_n1236), .A2(new_n765), .B1(new_n1241), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1240), .A2(new_n1257), .ZN(G381));
  XNOR2_X1  g1058(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1259));
  OR4_X1    g1059(.A1(G387), .A2(G381), .A3(G390), .A4(G378), .ZN(new_n1260));
  NOR2_X1   g1060(.A1(G393), .A2(G396), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1261), .A2(new_n869), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(new_n1262), .B(KEYINPUT120), .ZN(new_n1263));
  OR3_X1    g1063(.A1(new_n1259), .A2(new_n1260), .A3(new_n1263), .ZN(G407));
  NAND2_X1  g1064(.A1(new_n1127), .A2(new_n1149), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1125), .B2(new_n1121), .ZN(new_n1266));
  INV_X1    g1066(.A(G213), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(G343), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(new_n1259), .C2(new_n1269), .ZN(G409));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  OAI211_X1 g1071(.A(KEYINPUT117), .B(new_n712), .C1(new_n1223), .C2(new_n1226), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1221), .A2(new_n1217), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1219), .A2(KEYINPUT117), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1213), .C1(new_n1274), .C2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(KEYINPUT122), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n1277), .B1(new_n1182), .B2(new_n1212), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n765), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1279), .A2(new_n1211), .A3(KEYINPUT122), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1216), .A2(new_n1220), .A3(new_n1238), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1278), .A2(new_n1280), .A3(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1282), .A2(new_n1266), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1276), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1268), .ZN(new_n1285));
  OAI21_X1  g1085(.A(KEYINPUT60), .B1(new_n1089), .B2(new_n1109), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1237), .A2(new_n1286), .A3(new_n1239), .ZN(new_n1287));
  NOR2_X1   g1087(.A1(new_n1215), .A2(new_n1236), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1026), .B1(new_n1288), .B2(KEYINPUT60), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G384), .B1(new_n1290), .B2(new_n1257), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1257), .ZN(new_n1292));
  AOI211_X1 g1092(.A(new_n869), .B(new_n1292), .C1(new_n1287), .C2(new_n1289), .ZN(new_n1293));
  NOR2_X1   g1093(.A1(new_n1291), .A2(new_n1293), .ZN(new_n1294));
  NAND4_X1  g1094(.A1(new_n1284), .A2(KEYINPUT63), .A3(new_n1285), .A4(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT125), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1295), .A2(new_n1296), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1268), .B1(new_n1276), .B2(new_n1283), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1298), .A2(KEYINPUT125), .A3(KEYINPUT63), .A4(new_n1294), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(G393), .A2(G396), .ZN(new_n1301));
  INV_X1    g1101(.A(new_n1301), .ZN(new_n1302));
  OAI211_X1 g1102(.A(new_n1063), .B(new_n1085), .C1(new_n1302), .C2(new_n1261), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1261), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(G390), .A2(new_n1301), .A3(new_n1304), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(G387), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1303), .A2(new_n1305), .A3(new_n1024), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT61), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1307), .A2(new_n1308), .A3(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1290), .A2(new_n1257), .ZN(new_n1311));
  NAND2_X1  g1111(.A1(new_n1311), .A2(new_n869), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1290), .A2(G384), .A3(new_n1257), .ZN(new_n1313));
  INV_X1    g1113(.A(G2897), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1285), .A2(new_n1314), .ZN(new_n1315));
  NAND3_X1  g1115(.A1(new_n1312), .A2(new_n1313), .A3(new_n1315), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1315), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1317), .B1(new_n1291), .B2(new_n1293), .ZN(new_n1318));
  AND2_X1   g1118(.A1(new_n1316), .A2(new_n1318), .ZN(new_n1319));
  AOI21_X1  g1119(.A(new_n1319), .B1(new_n1298), .B2(KEYINPUT124), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT124), .ZN(new_n1321));
  AND2_X1   g1121(.A1(new_n1282), .A2(new_n1266), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1322), .B1(new_n1230), .B2(G378), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1321), .B1(new_n1323), .B2(new_n1268), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n1310), .B1(new_n1320), .B2(new_n1324), .ZN(new_n1325));
  NAND2_X1  g1125(.A1(new_n1300), .A2(new_n1325), .ZN(new_n1326));
  AOI211_X1 g1126(.A(KEYINPUT123), .B(KEYINPUT63), .C1(new_n1298), .C2(new_n1294), .ZN(new_n1327));
  INV_X1    g1127(.A(KEYINPUT123), .ZN(new_n1328));
  NAND3_X1  g1128(.A1(new_n1284), .A2(new_n1285), .A3(new_n1294), .ZN(new_n1329));
  INV_X1    g1129(.A(KEYINPUT63), .ZN(new_n1330));
  AOI21_X1  g1130(.A(new_n1328), .B1(new_n1329), .B2(new_n1330), .ZN(new_n1331));
  NOR2_X1   g1131(.A1(new_n1327), .A2(new_n1331), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1271), .B1(new_n1326), .B2(new_n1332), .ZN(new_n1333));
  NAND2_X1  g1133(.A1(new_n1329), .A2(new_n1330), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1334), .A2(KEYINPUT123), .ZN(new_n1335));
  NAND3_X1  g1135(.A1(new_n1329), .A2(new_n1328), .A3(new_n1330), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND4_X1  g1137(.A1(new_n1337), .A2(KEYINPUT126), .A3(new_n1300), .A4(new_n1325), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1333), .A2(new_n1338), .ZN(new_n1339));
  NAND2_X1  g1139(.A1(new_n1307), .A2(new_n1308), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1341));
  OAI211_X1 g1141(.A(new_n1341), .B(new_n1309), .C1(new_n1298), .C2(new_n1319), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1329), .A2(KEYINPUT62), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1340), .B1(new_n1342), .B2(new_n1343), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1339), .A2(new_n1344), .ZN(G405));
  NAND2_X1  g1145(.A1(G375), .A2(new_n1266), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(new_n1276), .ZN(new_n1347));
  OR2_X1    g1147(.A1(new_n1347), .A2(new_n1294), .ZN(new_n1348));
  OR2_X1    g1148(.A1(new_n1340), .A2(KEYINPUT127), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1347), .A2(new_n1294), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1348), .A2(new_n1349), .A3(new_n1350), .ZN(new_n1351));
  NAND2_X1  g1151(.A1(new_n1340), .A2(KEYINPUT127), .ZN(new_n1352));
  XOR2_X1   g1152(.A(new_n1351), .B(new_n1352), .Z(G402));
endmodule


