//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 1 0 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:21 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n959, new_n960, new_n961, new_n962, new_n963, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NOR2_X1   g003(.A1(new_n189), .A2(G104), .ZN(new_n190));
  INV_X1    g004(.A(G104), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G107), .ZN(new_n192));
  OAI21_X1  g006(.A(G101), .B1(new_n190), .B2(new_n192), .ZN(new_n193));
  OAI21_X1  g007(.A(KEYINPUT3), .B1(new_n191), .B2(G107), .ZN(new_n194));
  AOI21_X1  g008(.A(G101), .B1(new_n191), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(new_n189), .A3(G104), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n194), .A2(new_n195), .A3(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n193), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n203), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n202), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n200), .A2(G143), .ZN(new_n208));
  OAI211_X1 g022(.A(G128), .B(new_n206), .C1(new_n207), .C2(new_n208), .ZN(new_n209));
  NAND4_X1  g023(.A1(new_n199), .A2(KEYINPUT73), .A3(new_n205), .A4(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT10), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n209), .A2(new_n205), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n193), .A2(new_n198), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n210), .A2(new_n211), .A3(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n191), .A2(G107), .ZN(new_n217));
  NAND3_X1  g031(.A1(new_n194), .A2(new_n197), .A3(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n218), .A2(G101), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT72), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n218), .A2(KEYINPUT72), .A3(G101), .ZN(new_n222));
  AND2_X1   g036(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT4), .ZN(new_n225));
  AND3_X1   g039(.A1(new_n218), .A2(new_n225), .A3(G101), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n201), .A2(new_n203), .A3(KEYINPUT0), .A4(G128), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n207), .A2(new_n208), .ZN(new_n228));
  XNOR2_X1  g042(.A(KEYINPUT0), .B(G128), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n227), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n224), .A2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n209), .A2(new_n205), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(KEYINPUT10), .A3(new_n199), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT11), .ZN(new_n235));
  INV_X1    g049(.A(G134), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n235), .B1(new_n236), .B2(G137), .ZN(new_n237));
  INV_X1    g051(.A(G137), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n238), .A2(KEYINPUT11), .A3(G134), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n236), .A2(G137), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n237), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(G131), .ZN(new_n242));
  INV_X1    g056(.A(G131), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n237), .A2(new_n239), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n242), .A2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT74), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT74), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n242), .A2(new_n247), .A3(new_n244), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n216), .A2(new_n232), .A3(new_n234), .A4(new_n249), .ZN(new_n250));
  XNOR2_X1  g064(.A(G110), .B(G140), .ZN(new_n251));
  INV_X1    g065(.A(G953), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n252), .A2(G227), .ZN(new_n253));
  XOR2_X1   g067(.A(new_n251), .B(new_n253), .Z(new_n254));
  INV_X1    g068(.A(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(KEYINPUT76), .B1(new_n233), .B2(new_n199), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT76), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n213), .A2(new_n214), .A3(new_n258), .ZN(new_n259));
  NAND4_X1  g073(.A1(new_n257), .A2(new_n210), .A3(new_n215), .A4(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT12), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(KEYINPUT75), .ZN(new_n262));
  NOR2_X1   g076(.A1(new_n262), .A2(KEYINPUT12), .ZN(new_n263));
  INV_X1    g077(.A(new_n263), .ZN(new_n264));
  AND2_X1   g078(.A1(new_n245), .A2(KEYINPUT75), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n260), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n260), .A2(new_n265), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(new_n263), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n256), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND3_X1  g083(.A1(new_n216), .A2(new_n232), .A3(new_n234), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n245), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n255), .B1(new_n271), .B2(new_n250), .ZN(new_n272));
  OAI211_X1 g086(.A(new_n187), .B(new_n188), .C1(new_n269), .C2(new_n272), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n187), .A2(new_n188), .ZN(new_n274));
  INV_X1    g088(.A(new_n274), .ZN(new_n275));
  AND2_X1   g089(.A1(new_n250), .A2(new_n255), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(new_n271), .ZN(new_n277));
  INV_X1    g091(.A(new_n250), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n278), .B1(new_n268), .B2(new_n266), .ZN(new_n279));
  OAI211_X1 g093(.A(new_n277), .B(G469), .C1(new_n279), .C2(new_n255), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n273), .A2(new_n275), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT77), .ZN(new_n282));
  INV_X1    g096(.A(G221), .ZN(new_n283));
  XOR2_X1   g097(.A(KEYINPUT9), .B(G234), .Z(new_n284));
  AOI21_X1  g098(.A(new_n283), .B1(new_n284), .B2(new_n188), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AND3_X1   g100(.A1(new_n281), .A2(new_n282), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n282), .B1(new_n281), .B2(new_n286), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(G217), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n290), .B1(G234), .B2(new_n188), .ZN(new_n291));
  XNOR2_X1  g105(.A(KEYINPUT22), .B(G137), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n292), .B(new_n293), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n204), .A2(G119), .ZN(new_n296));
  NAND2_X1  g110(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G119), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G128), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n296), .B1(new_n303), .B2(new_n297), .ZN(new_n304));
  OAI21_X1  g118(.A(G110), .B1(new_n301), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n296), .A2(new_n300), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT24), .B(G110), .ZN(new_n307));
  OR2_X1    g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G140), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G125), .ZN(new_n310));
  INV_X1    g124(.A(G125), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(G140), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n310), .A2(new_n312), .A3(KEYINPUT16), .ZN(new_n313));
  OR3_X1    g127(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n314));
  AOI21_X1  g128(.A(G146), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n313), .A2(G146), .A3(new_n314), .ZN(new_n316));
  OAI211_X1 g130(.A(new_n305), .B(new_n308), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n299), .A2(G128), .ZN(new_n318));
  AND2_X1   g132(.A1(KEYINPUT67), .A2(KEYINPUT23), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n318), .B1(new_n319), .B2(new_n302), .ZN(new_n320));
  INV_X1    g134(.A(G110), .ZN(new_n321));
  NAND4_X1  g135(.A1(new_n320), .A2(new_n321), .A3(new_n300), .A4(new_n298), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT68), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n306), .A2(new_n307), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n322), .A2(new_n323), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n310), .A2(new_n312), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n326), .A2(G146), .ZN(new_n327));
  NOR3_X1   g141(.A1(new_n311), .A2(KEYINPUT16), .A3(G140), .ZN(new_n328));
  XNOR2_X1  g142(.A(G125), .B(G140), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n328), .B1(new_n329), .B2(KEYINPUT16), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n327), .B1(new_n330), .B2(G146), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n325), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g146(.A(new_n323), .B1(new_n322), .B2(new_n324), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n317), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT69), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  OAI211_X1 g150(.A(new_n317), .B(KEYINPUT69), .C1(new_n332), .C2(new_n333), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n295), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n295), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT25), .B1(new_n341), .B2(new_n188), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT25), .ZN(new_n343));
  NOR4_X1   g157(.A1(new_n338), .A2(new_n340), .A3(new_n343), .A4(G902), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n291), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT71), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n291), .A2(G902), .ZN(new_n347));
  XOR2_X1   g161(.A(new_n347), .B(KEYINPUT70), .Z(new_n348));
  AOI21_X1  g162(.A(new_n346), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n348), .ZN(new_n350));
  NOR4_X1   g164(.A1(new_n338), .A2(new_n340), .A3(KEYINPUT71), .A4(new_n350), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NOR2_X1   g167(.A1(G237), .A2(G953), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G210), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n355), .B(KEYINPUT27), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT26), .B(G101), .ZN(new_n357));
  XNOR2_X1  g171(.A(new_n356), .B(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(new_n230), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n245), .ZN(new_n360));
  INV_X1    g174(.A(G113), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT2), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT2), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n363), .A2(G113), .ZN(new_n364));
  AND2_X1   g178(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n299), .A2(G116), .ZN(new_n366));
  INV_X1    g180(.A(G116), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G119), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  OAI21_X1  g183(.A(KEYINPUT66), .B1(new_n365), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n362), .A2(new_n364), .ZN(new_n371));
  XNOR2_X1  g185(.A(G116), .B(G119), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT66), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n370), .A2(new_n374), .B1(new_n369), .B2(new_n365), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n236), .A2(G137), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n238), .A2(G134), .ZN(new_n377));
  OAI21_X1  g191(.A(G131), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n209), .A2(new_n244), .A3(new_n378), .A4(new_n205), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n360), .A2(new_n375), .A3(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n380), .B(KEYINPUT28), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n244), .A2(new_n378), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n233), .A2(new_n382), .A3(KEYINPUT65), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT65), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n379), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n383), .A2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT64), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n230), .A2(new_n387), .ZN(new_n388));
  XOR2_X1   g202(.A(KEYINPUT0), .B(G128), .Z(new_n389));
  OAI21_X1  g203(.A(new_n389), .B1(new_n207), .B2(new_n208), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n390), .A2(KEYINPUT64), .A3(new_n227), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n388), .A2(new_n391), .A3(new_n245), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n365), .A2(new_n369), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n371), .A2(new_n372), .A3(new_n373), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n373), .B1(new_n371), .B2(new_n372), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n394), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n393), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n358), .B1(new_n381), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT31), .ZN(new_n400));
  AOI21_X1  g214(.A(KEYINPUT30), .B1(new_n386), .B2(new_n392), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n230), .B1(new_n244), .B2(new_n242), .ZN(new_n402));
  INV_X1    g216(.A(new_n379), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT30), .ZN(new_n404));
  NOR3_X1   g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  NOR3_X1   g219(.A1(new_n401), .A2(new_n375), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n380), .A2(new_n358), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n400), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n405), .ZN(new_n409));
  AND2_X1   g223(.A1(new_n388), .A2(new_n391), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n410), .A2(new_n245), .B1(new_n383), .B2(new_n385), .ZN(new_n411));
  OAI211_X1 g225(.A(new_n397), .B(new_n409), .C1(new_n411), .C2(KEYINPUT30), .ZN(new_n412));
  INV_X1    g226(.A(new_n407), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n412), .A2(KEYINPUT31), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n399), .B1(new_n408), .B2(new_n414), .ZN(new_n415));
  NOR2_X1   g229(.A1(G472), .A2(G902), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g231(.A(KEYINPUT32), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(new_n399), .ZN(new_n419));
  NOR3_X1   g233(.A1(new_n406), .A2(new_n400), .A3(new_n407), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT31), .B1(new_n412), .B2(new_n413), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n419), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT32), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n422), .A2(new_n423), .A3(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n418), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n397), .B1(new_n402), .B2(new_n403), .ZN(new_n426));
  AND2_X1   g240(.A1(new_n381), .A2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n358), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT29), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(G902), .B1(new_n427), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n380), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n406), .A2(new_n432), .ZN(new_n433));
  NOR2_X1   g247(.A1(new_n433), .A2(new_n358), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n381), .A2(new_n398), .A3(new_n358), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(new_n429), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n431), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(G472), .ZN(new_n438));
  AOI21_X1  g252(.A(new_n353), .B1(new_n425), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n214), .B1(new_n370), .B2(new_n374), .ZN(new_n440));
  NAND2_X1  g254(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n441));
  INV_X1    g255(.A(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n443));
  OAI211_X1 g257(.A(new_n366), .B(new_n368), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  OR2_X1    g258(.A1(KEYINPUT79), .A2(KEYINPUT5), .ZN(new_n445));
  NAND4_X1  g259(.A1(new_n445), .A2(G116), .A3(new_n299), .A4(new_n441), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n446), .A3(G113), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n440), .A2(new_n447), .ZN(new_n448));
  INV_X1    g262(.A(new_n226), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n397), .A2(new_n449), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n218), .A2(KEYINPUT72), .A3(G101), .ZN(new_n451));
  AOI21_X1  g265(.A(KEYINPUT72), .B1(new_n218), .B2(G101), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n453));
  NOR3_X1   g267(.A1(new_n451), .A2(new_n452), .A3(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n448), .B1(new_n450), .B2(new_n454), .ZN(new_n455));
  XNOR2_X1  g269(.A(G110), .B(G122), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(new_n448), .B(new_n456), .C1(new_n450), .C2(new_n454), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n311), .B1(new_n390), .B2(new_n227), .ZN(new_n461));
  AOI21_X1  g275(.A(G125), .B1(new_n209), .B2(new_n205), .ZN(new_n462));
  NOR2_X1   g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(G224), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XOR2_X1   g279(.A(new_n463), .B(new_n465), .Z(new_n466));
  INV_X1    g280(.A(KEYINPUT6), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n455), .A2(new_n467), .A3(new_n457), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n460), .A2(new_n466), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n372), .A2(KEYINPUT5), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n470), .A2(G113), .A3(new_n446), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n447), .B1(new_n395), .B2(new_n396), .ZN(new_n472));
  AOI22_X1  g286(.A1(new_n440), .A2(new_n471), .B1(new_n472), .B2(new_n214), .ZN(new_n473));
  XOR2_X1   g287(.A(KEYINPUT80), .B(KEYINPUT8), .Z(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n456), .ZN(new_n475));
  INV_X1    g289(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g290(.A(KEYINPUT81), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT81), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n370), .A2(new_n374), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n479), .A2(new_n199), .A3(new_n471), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n199), .B1(new_n479), .B2(new_n447), .ZN(new_n481));
  OAI211_X1 g295(.A(new_n478), .B(new_n475), .C1(new_n480), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n477), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT7), .ZN(new_n484));
  OAI22_X1  g298(.A1(new_n461), .A2(new_n462), .B1(new_n484), .B2(new_n465), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n230), .A2(G125), .ZN(new_n486));
  NOR2_X1   g300(.A1(new_n465), .A2(new_n484), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n486), .B(new_n487), .C1(new_n233), .C2(G125), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n226), .B1(new_n479), .B2(new_n394), .ZN(new_n490));
  AOI22_X1  g304(.A1(new_n490), .A2(new_n224), .B1(new_n447), .B2(new_n440), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n491), .B2(new_n456), .ZN(new_n492));
  AOI21_X1  g306(.A(G902), .B1(new_n483), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n469), .A2(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(G210), .B1(G237), .B2(G902), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n494), .A2(new_n496), .ZN(new_n497));
  NAND3_X1  g311(.A1(new_n469), .A2(new_n493), .A3(new_n495), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  XNOR2_X1  g313(.A(G113), .B(G122), .ZN(new_n500));
  XNOR2_X1  g314(.A(new_n500), .B(new_n191), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n354), .A2(G214), .ZN(new_n503));
  NOR2_X1   g317(.A1(KEYINPUT82), .A2(G143), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n354), .B(G214), .C1(KEYINPUT82), .C2(G143), .ZN(new_n506));
  AND2_X1   g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(KEYINPUT18), .A2(G131), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n329), .A2(new_n200), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n326), .A2(G146), .ZN(new_n510));
  AOI22_X1  g324(.A1(new_n507), .A2(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n505), .A2(new_n506), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(KEYINPUT18), .A3(G131), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(KEYINPUT17), .A3(G131), .ZN(new_n514));
  INV_X1    g328(.A(new_n315), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n330), .A2(G146), .ZN(new_n516));
  AND3_X1   g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n505), .A2(new_n506), .A3(new_n243), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT83), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n512), .A2(G131), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT17), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n505), .A2(new_n506), .A3(KEYINPUT83), .A4(new_n243), .ZN(new_n523));
  NAND4_X1  g337(.A1(new_n520), .A2(new_n521), .A3(new_n522), .A4(new_n523), .ZN(new_n524));
  AOI221_X4 g338(.A(new_n502), .B1(new_n511), .B2(new_n513), .C1(new_n517), .C2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n517), .A2(new_n524), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n511), .A2(new_n513), .ZN(new_n527));
  AOI21_X1  g341(.A(new_n501), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n188), .B1(new_n525), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT87), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT87), .B(new_n188), .C1(new_n525), .C2(new_n528), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(G475), .A3(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(G475), .A2(G902), .ZN(new_n534));
  XOR2_X1   g348(.A(new_n534), .B(KEYINPUT86), .Z(new_n535));
  INV_X1    g349(.A(KEYINPUT84), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n310), .A2(new_n312), .A3(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT19), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT19), .B1(new_n329), .B2(new_n536), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n200), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI21_X1  g355(.A(new_n316), .B1(new_n541), .B2(KEYINPUT85), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n520), .A2(new_n523), .A3(new_n521), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n537), .B(new_n538), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT85), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n544), .A2(new_n545), .A3(new_n200), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n542), .A2(new_n543), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g361(.A(new_n501), .B1(new_n547), .B2(new_n527), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n535), .B1(new_n548), .B2(new_n525), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT20), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT20), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n551), .B(new_n535), .C1(new_n548), .C2(new_n525), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n533), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n202), .A2(G128), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n204), .A2(G143), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n555), .A2(new_n556), .A3(new_n236), .ZN(new_n557));
  INV_X1    g371(.A(G122), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(G116), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n367), .A2(G122), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n561), .A2(G107), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n559), .A2(new_n560), .A3(new_n189), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n557), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT13), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n555), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n556), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n555), .A2(new_n565), .ZN(new_n568));
  OAI21_X1  g382(.A(G134), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n564), .A2(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n367), .A2(KEYINPUT14), .A3(G122), .ZN(new_n571));
  OAI211_X1 g385(.A(G107), .B(new_n571), .C1(new_n561), .C2(KEYINPUT14), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n236), .B1(new_n555), .B2(new_n556), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n572), .B(new_n563), .C1(new_n557), .C2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n284), .A2(G217), .A3(new_n252), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n570), .A2(new_n574), .A3(new_n576), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(G902), .ZN(new_n581));
  INV_X1    g395(.A(G478), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n582), .A2(KEYINPUT15), .ZN(new_n583));
  XNOR2_X1  g397(.A(new_n581), .B(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(G234), .A2(G237), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n586), .A2(G902), .A3(G953), .ZN(new_n587));
  XOR2_X1   g401(.A(new_n587), .B(KEYINPUT88), .Z(new_n588));
  XNOR2_X1  g402(.A(KEYINPUT21), .B(G898), .ZN(new_n589));
  AND2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AND3_X1   g404(.A1(new_n586), .A2(G952), .A3(new_n252), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G214), .B1(G237), .B2(G902), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT78), .ZN(new_n594));
  OR2_X1    g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  NOR4_X1   g409(.A1(new_n499), .A2(new_n554), .A3(new_n585), .A4(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n289), .A2(new_n439), .A3(new_n596), .ZN(new_n597));
  XNOR2_X1  g411(.A(new_n597), .B(G101), .ZN(G3));
  INV_X1    g412(.A(new_n592), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n497), .A2(KEYINPUT89), .A3(new_n498), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n578), .A2(new_n601), .A3(new_n579), .ZN(new_n602));
  NOR2_X1   g416(.A1(new_n582), .A2(G902), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT91), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n604), .B1(new_n575), .B2(KEYINPUT90), .ZN(new_n605));
  INV_X1    g419(.A(KEYINPUT90), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n576), .B2(KEYINPUT91), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n605), .A2(new_n576), .B1(new_n575), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g422(.A(new_n602), .B(new_n603), .C1(new_n608), .C2(new_n601), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n582), .B1(new_n580), .B2(G902), .ZN(new_n610));
  AND2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n611), .B1(new_n553), .B2(new_n533), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT89), .ZN(new_n613));
  NAND4_X1  g427(.A1(new_n469), .A2(new_n493), .A3(new_n613), .A4(new_n495), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n614), .A2(new_n593), .ZN(new_n615));
  AND4_X1   g429(.A1(new_n599), .A2(new_n600), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  OAI21_X1  g430(.A(G472), .B1(new_n415), .B2(G902), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n422), .A2(new_n416), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n619), .A2(new_n353), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n289), .A2(new_n616), .A3(new_n620), .ZN(new_n621));
  XOR2_X1   g435(.A(KEYINPUT34), .B(G104), .Z(new_n622));
  XNOR2_X1  g436(.A(new_n621), .B(new_n622), .ZN(G6));
  NAND2_X1  g437(.A1(new_n600), .A2(new_n615), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT92), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n553), .A2(new_n625), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n550), .A2(KEYINPUT92), .A3(new_n552), .ZN(new_n627));
  NAND4_X1  g441(.A1(new_n626), .A2(new_n533), .A3(new_n585), .A4(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n624), .A2(new_n628), .ZN(new_n629));
  AND4_X1   g443(.A1(new_n289), .A2(new_n599), .A3(new_n620), .A4(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT35), .B(G107), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(KEYINPUT93), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n334), .B(new_n633), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n295), .A2(KEYINPUT36), .ZN(new_n635));
  OR2_X1    g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(new_n345), .B1(new_n350), .B2(new_n639), .ZN(new_n640));
  NAND4_X1  g454(.A1(new_n640), .A2(KEYINPUT94), .A3(new_n618), .A4(new_n617), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT94), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n350), .B1(new_n636), .B2(new_n637), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n336), .A2(new_n337), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n294), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n645), .A2(new_n188), .A3(new_n339), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(new_n343), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n341), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n643), .B1(new_n649), .B2(new_n291), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n642), .B1(new_n619), .B2(new_n650), .ZN(new_n651));
  NAND4_X1  g465(.A1(new_n289), .A2(new_n641), .A3(new_n596), .A4(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT37), .B(G110), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G12));
  INV_X1    g468(.A(G900), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n591), .B1(new_n588), .B2(new_n655), .ZN(new_n656));
  XOR2_X1   g470(.A(new_n656), .B(KEYINPUT95), .Z(new_n657));
  NOR3_X1   g471(.A1(new_n624), .A2(new_n628), .A3(new_n657), .ZN(new_n658));
  AOI21_X1  g472(.A(new_n650), .B1(new_n425), .B2(new_n438), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n289), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n657), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n289), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n663), .B(KEYINPUT40), .ZN(new_n664));
  OR2_X1    g478(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n664), .A2(KEYINPUT97), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n499), .B(KEYINPUT38), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n358), .B1(new_n426), .B2(new_n380), .ZN(new_n668));
  XOR2_X1   g482(.A(new_n668), .B(KEYINPUT96), .Z(new_n669));
  NOR2_X1   g483(.A1(new_n406), .A2(new_n407), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n188), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(G472), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n425), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n673), .A2(new_n650), .ZN(new_n674));
  INV_X1    g488(.A(new_n593), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n554), .A2(new_n585), .ZN(new_n676));
  NOR4_X1   g490(.A1(new_n667), .A2(new_n674), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n665), .A2(new_n666), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT98), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n665), .A2(new_n666), .A3(KEYINPUT98), .A4(new_n677), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(new_n202), .ZN(G45));
  INV_X1    g497(.A(new_n657), .ZN(new_n684));
  AND4_X1   g498(.A1(new_n600), .A2(new_n612), .A3(new_n615), .A4(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n288), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n260), .A2(new_n264), .A3(new_n265), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n264), .B1(new_n260), .B2(new_n265), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n250), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  AOI22_X1  g503(.A1(new_n689), .A2(new_n254), .B1(new_n271), .B2(new_n276), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n274), .B1(new_n690), .B2(G469), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n285), .B1(new_n691), .B2(new_n273), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n282), .ZN(new_n693));
  NAND4_X1  g507(.A1(new_n659), .A2(new_n685), .A3(new_n686), .A4(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  OAI21_X1  g509(.A(new_n188), .B1(new_n269), .B2(new_n272), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n286), .A3(new_n273), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n439), .A2(new_n616), .A3(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND4_X1  g516(.A1(new_n439), .A2(new_n629), .A3(new_n599), .A4(new_n699), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n425), .A2(new_n438), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n706), .A2(new_n640), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n533), .A2(new_n553), .A3(new_n584), .A4(new_n599), .ZN(new_n708));
  INV_X1    g522(.A(new_n708), .ZN(new_n709));
  NAND4_X1  g523(.A1(new_n699), .A2(new_n600), .A3(new_n615), .A4(new_n709), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n705), .B1(new_n707), .B2(new_n710), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n624), .A2(new_n698), .A3(new_n708), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(KEYINPUT99), .A3(new_n659), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G119), .ZN(G21));
  NOR2_X1   g529(.A1(new_n624), .A2(new_n676), .ZN(new_n716));
  OAI22_X1  g530(.A1(new_n420), .A2(new_n421), .B1(new_n427), .B2(new_n358), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n416), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n617), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n353), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n716), .A2(new_n720), .A3(new_n599), .A4(new_n699), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G122), .ZN(G24));
  NOR2_X1   g536(.A1(new_n624), .A2(new_n698), .ZN(new_n723));
  NOR2_X1   g537(.A1(new_n719), .A2(new_n650), .ZN(new_n724));
  INV_X1    g538(.A(new_n612), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n725), .A2(new_n657), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(KEYINPUT100), .B(G125), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n727), .B(new_n728), .ZN(G27));
  AND3_X1   g543(.A1(new_n612), .A2(KEYINPUT42), .A3(new_n684), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n439), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT101), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n281), .A2(new_n732), .A3(new_n286), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n732), .B1(new_n281), .B2(new_n286), .ZN(new_n734));
  INV_X1    g548(.A(KEYINPUT102), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n497), .A2(new_n498), .A3(new_n593), .ZN(new_n736));
  NOR4_X1   g550(.A1(new_n733), .A2(new_n734), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n281), .A2(new_n286), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n736), .B1(new_n738), .B2(KEYINPUT101), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n692), .A2(new_n732), .ZN(new_n740));
  AOI21_X1  g554(.A(KEYINPUT102), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(new_n731), .B1(new_n737), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(KEYINPUT104), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n731), .B(new_n744), .C1(new_n737), .C2(new_n741), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(new_n439), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n739), .A2(new_n740), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n750), .A2(new_n735), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n739), .A2(KEYINPUT102), .A3(new_n740), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n748), .B1(new_n753), .B2(new_n726), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT105), .B1(new_n746), .B2(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n439), .B1(new_n737), .B2(new_n741), .ZN(new_n756));
  INV_X1    g570(.A(new_n726), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n747), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g572(.A(KEYINPUT105), .ZN(new_n759));
  NAND4_X1  g573(.A1(new_n758), .A2(new_n743), .A3(new_n759), .A4(new_n745), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n243), .ZN(G33));
  NAND2_X1  g576(.A1(new_n626), .A2(new_n627), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n763), .A2(new_n657), .ZN(new_n764));
  AND3_X1   g578(.A1(new_n764), .A2(new_n533), .A3(new_n585), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n439), .B(new_n765), .C1(new_n737), .C2(new_n741), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G134), .ZN(G36));
  INV_X1    g581(.A(KEYINPUT43), .ZN(new_n768));
  OAI22_X1  g582(.A1(new_n554), .A2(new_n611), .B1(KEYINPUT106), .B2(new_n768), .ZN(new_n769));
  OR2_X1    g583(.A1(new_n554), .A2(new_n611), .ZN(new_n770));
  XNOR2_X1  g584(.A(KEYINPUT106), .B(KEYINPUT43), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n769), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n772), .A2(new_n619), .A3(new_n640), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  NOR2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(KEYINPUT107), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n690), .A2(KEYINPUT45), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n690), .B2(KEYINPUT45), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT46), .B1(new_n780), .B2(new_n275), .ZN(new_n781));
  INV_X1    g595(.A(new_n273), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n780), .A2(KEYINPUT46), .A3(new_n275), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n285), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n736), .B1(new_n773), .B2(new_n774), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n776), .A2(new_n662), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  XOR2_X1   g602(.A(new_n785), .B(KEYINPUT47), .Z(new_n789));
  INV_X1    g603(.A(new_n353), .ZN(new_n790));
  OR4_X1    g604(.A1(new_n706), .A2(new_n757), .A3(new_n790), .A4(new_n736), .ZN(new_n791));
  OR2_X1    g605(.A1(new_n789), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G140), .ZN(G42));
  NOR2_X1   g607(.A1(new_n738), .A2(new_n657), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n716), .A2(new_n673), .A3(new_n794), .A4(new_n650), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n660), .A2(new_n694), .A3(new_n727), .A4(new_n795), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT110), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n796), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n798), .B1(new_n796), .B2(new_n797), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT52), .ZN(new_n802));
  AND2_X1   g616(.A1(new_n796), .A2(new_n802), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n796), .A2(new_n802), .ZN(new_n804));
  OAI22_X1  g618(.A1(new_n800), .A2(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n796), .A2(new_n797), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n806), .A2(KEYINPUT111), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n796), .A2(new_n802), .ZN(new_n808));
  AND2_X1   g622(.A1(new_n660), .A2(new_n727), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n809), .A2(KEYINPUT52), .A3(new_n694), .A4(new_n795), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n807), .A2(new_n808), .A3(new_n810), .A4(new_n799), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n805), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n758), .A2(new_n743), .A3(new_n745), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n499), .A2(new_n595), .ZN(new_n814));
  INV_X1    g628(.A(new_n554), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n585), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n816), .A2(new_n725), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n289), .A2(new_n814), .A3(new_n620), .A4(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n652), .A2(new_n818), .A3(new_n597), .ZN(new_n819));
  OAI211_X1 g633(.A(new_n726), .B(new_n724), .C1(new_n737), .C2(new_n741), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n533), .A2(new_n584), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n736), .A2(new_n821), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n289), .A2(new_n659), .A3(new_n764), .A4(new_n822), .ZN(new_n823));
  NAND4_X1  g637(.A1(new_n819), .A2(new_n766), .A3(new_n820), .A4(new_n823), .ZN(new_n824));
  INV_X1    g638(.A(new_n824), .ZN(new_n825));
  AND3_X1   g639(.A1(new_n712), .A2(KEYINPUT99), .A3(new_n659), .ZN(new_n826));
  AOI21_X1  g640(.A(KEYINPUT99), .B1(new_n712), .B2(new_n659), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT53), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n703), .A2(new_n721), .A3(new_n700), .ZN(new_n830));
  NOR3_X1   g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n812), .A2(new_n813), .A3(new_n825), .A4(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT54), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT108), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n828), .A2(new_n834), .A3(new_n830), .ZN(new_n835));
  AND3_X1   g649(.A1(new_n703), .A2(new_n700), .A3(new_n721), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT108), .B1(new_n836), .B2(new_n714), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n835), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n755), .A2(new_n838), .A3(new_n760), .A4(new_n825), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n803), .A2(new_n804), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n829), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n832), .A2(new_n833), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT109), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n839), .A2(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n824), .A2(new_n835), .A3(new_n837), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(KEYINPUT109), .A3(new_n755), .A4(new_n760), .ZN(new_n846));
  NAND3_X1  g660(.A1(new_n844), .A2(new_n846), .A3(new_n812), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(new_n829), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n839), .A2(new_n829), .A3(new_n840), .ZN(new_n849));
  INV_X1    g663(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n848), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n842), .B1(new_n851), .B2(KEYINPUT54), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n667), .A2(new_n675), .A3(new_n699), .ZN(new_n853));
  XOR2_X1   g667(.A(new_n853), .B(KEYINPUT112), .Z(new_n854));
  NAND3_X1  g668(.A1(new_n772), .A2(new_n591), .A3(new_n720), .ZN(new_n855));
  NOR2_X1   g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT114), .ZN(new_n857));
  XNOR2_X1  g671(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n858));
  OR3_X1    g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  OAI21_X1  g673(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n856), .A2(KEYINPUT50), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n859), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(new_n673), .ZN(new_n863));
  INV_X1    g677(.A(new_n591), .ZN(new_n864));
  NOR3_X1   g678(.A1(new_n698), .A2(new_n736), .A3(new_n864), .ZN(new_n865));
  AND3_X1   g679(.A1(new_n863), .A2(new_n790), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n866), .A2(new_n815), .A3(new_n611), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n772), .A2(new_n724), .A3(new_n865), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n697), .A2(new_n273), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n789), .B1(new_n286), .B2(new_n870), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n855), .A2(new_n736), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n869), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n862), .A2(KEYINPUT51), .A3(new_n873), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT51), .B1(new_n862), .B2(new_n873), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n772), .A2(new_n439), .A3(new_n865), .ZN(new_n876));
  XOR2_X1   g690(.A(new_n876), .B(KEYINPUT48), .Z(new_n877));
  INV_X1    g691(.A(G952), .ZN(new_n878));
  AOI211_X1 g692(.A(new_n878), .B(G953), .C1(new_n866), .C2(new_n612), .ZN(new_n879));
  INV_X1    g693(.A(new_n723), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n879), .B1(new_n880), .B2(new_n855), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n875), .A2(new_n877), .A3(new_n881), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n852), .A2(new_n874), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n883), .B1(G952), .B2(G953), .ZN(new_n884));
  XOR2_X1   g698(.A(new_n870), .B(KEYINPUT49), .Z(new_n885));
  NOR4_X1   g699(.A1(new_n770), .A2(new_n353), .A3(new_n285), .A4(new_n594), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n885), .A2(new_n886), .A3(new_n863), .A4(new_n667), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n884), .A2(new_n887), .ZN(G75));
  INV_X1    g702(.A(KEYINPUT116), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n188), .B1(new_n832), .B2(new_n841), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT56), .B1(new_n890), .B2(G210), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n460), .A2(new_n468), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(KEYINPUT115), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n466), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n891), .A2(new_n895), .ZN(new_n896));
  INV_X1    g710(.A(new_n896), .ZN(new_n897));
  OAI22_X1  g711(.A1(new_n891), .A2(new_n895), .B1(G952), .B2(new_n252), .ZN(new_n898));
  OAI21_X1  g712(.A(new_n889), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n252), .A2(G952), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n890), .A2(G210), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT56), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(new_n895), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n900), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n905), .A2(KEYINPUT116), .A3(new_n896), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n899), .A2(new_n906), .ZN(G51));
  XNOR2_X1  g721(.A(new_n274), .B(KEYINPUT57), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n833), .B1(new_n832), .B2(new_n841), .ZN(new_n909));
  OAI21_X1  g723(.A(new_n908), .B1(new_n842), .B2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT117), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g726(.A(KEYINPUT117), .B(new_n908), .C1(new_n842), .C2(new_n909), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n912), .B(new_n913), .C1(new_n272), .C2(new_n269), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n890), .A2(new_n779), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n900), .B1(new_n914), .B2(new_n915), .ZN(G54));
  AND3_X1   g730(.A1(new_n890), .A2(KEYINPUT58), .A3(G475), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n548), .A2(new_n525), .ZN(new_n918));
  INV_X1    g732(.A(new_n918), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT118), .B1(new_n917), .B2(new_n919), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n900), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n917), .A2(KEYINPUT118), .A3(new_n919), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n922), .A2(new_n923), .ZN(G60));
  NAND2_X1  g738(.A1(G478), .A2(G902), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT121), .ZN(new_n926));
  XOR2_X1   g740(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n927));
  XNOR2_X1  g741(.A(new_n926), .B(new_n927), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n805), .A2(new_n811), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n839), .B2(new_n843), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT53), .B1(new_n930), .B2(new_n846), .ZN(new_n931));
  OAI21_X1  g745(.A(KEYINPUT54), .B1(new_n931), .B2(new_n849), .ZN(new_n932));
  NAND3_X1  g746(.A1(new_n832), .A2(new_n833), .A3(new_n841), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n928), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  OAI21_X1  g748(.A(new_n602), .B1(new_n608), .B2(new_n601), .ZN(new_n935));
  XOR2_X1   g749(.A(new_n935), .B(KEYINPUT119), .Z(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(KEYINPUT122), .B1(new_n934), .B2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT122), .ZN(new_n939));
  OAI211_X1 g753(.A(new_n939), .B(new_n936), .C1(new_n852), .C2(new_n928), .ZN(new_n940));
  OR2_X1    g754(.A1(new_n842), .A2(new_n909), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n936), .A2(new_n928), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n900), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  AND3_X1   g757(.A1(new_n938), .A2(new_n940), .A3(new_n943), .ZN(G63));
  NAND2_X1  g758(.A1(new_n832), .A2(new_n841), .ZN(new_n945));
  NAND2_X1  g759(.A1(G217), .A2(G902), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n946), .B(KEYINPUT60), .Z(new_n947));
  NAND2_X1  g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n341), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n900), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n945), .A2(new_n638), .A3(new_n947), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT61), .ZN(new_n953));
  OR2_X1    g767(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(KEYINPUT123), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n952), .A2(new_n954), .A3(new_n955), .ZN(new_n956));
  NAND4_X1  g770(.A1(new_n950), .A2(KEYINPUT123), .A3(new_n953), .A4(new_n951), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n956), .A2(new_n957), .ZN(G66));
  OAI21_X1  g772(.A(G953), .B1(new_n589), .B2(new_n464), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n838), .A2(new_n819), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n961), .B2(G953), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n893), .B1(G898), .B2(new_n252), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n962), .B(new_n963), .ZN(G69));
  NOR2_X1   g778(.A1(new_n401), .A2(new_n405), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n544), .B(KEYINPUT124), .Z(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n787), .A2(new_n766), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n809), .A2(new_n694), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT125), .Z(new_n971));
  NAND4_X1  g785(.A1(new_n785), .A2(new_n439), .A3(new_n662), .A4(new_n716), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n972), .B(KEYINPUT126), .ZN(new_n973));
  AND4_X1   g787(.A1(new_n792), .A2(new_n969), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n761), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n252), .A3(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(G900), .A2(G953), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n968), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n968), .A2(new_n252), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n680), .A2(new_n681), .A3(new_n971), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n980), .A2(KEYINPUT62), .ZN(new_n981));
  INV_X1    g795(.A(new_n817), .ZN(new_n982));
  OR4_X1    g796(.A1(new_n749), .A2(new_n663), .A3(new_n736), .A4(new_n982), .ZN(new_n983));
  AND3_X1   g797(.A1(new_n792), .A2(new_n787), .A3(new_n983), .ZN(new_n984));
  AND2_X1   g798(.A1(new_n981), .A2(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT62), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n680), .A2(new_n986), .A3(new_n681), .A4(new_n971), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n979), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n978), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n252), .B1(G227), .B2(G900), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n989), .B(new_n990), .ZN(G72));
  NOR2_X1   g805(.A1(new_n433), .A2(new_n428), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n981), .A2(new_n984), .A3(new_n961), .A4(new_n987), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  AND3_X1   g809(.A1(new_n993), .A2(KEYINPUT127), .A3(new_n995), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT127), .B1(new_n993), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n851), .B(new_n995), .C1(new_n670), .C2(new_n434), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n974), .A2(new_n975), .A3(new_n961), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n1000), .A2(new_n995), .ZN(new_n1001));
  NOR3_X1   g815(.A1(new_n406), .A2(new_n432), .A3(new_n358), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n900), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n998), .A2(new_n999), .A3(new_n1003), .ZN(G57));
endmodule


