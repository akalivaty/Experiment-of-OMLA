//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 0 1 1 0 1 0 1 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n601,
    new_n602, new_n603, new_n604, new_n606, new_n607, new_n608, new_n609,
    new_n610, new_n611, new_n612, new_n613, new_n614, new_n615, new_n616,
    new_n617, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n665, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n839, new_n840, new_n841,
    new_n842, new_n844, new_n845, new_n846, new_n847, new_n849, new_n850,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n859, new_n860, new_n861, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921;
  INV_X1    g000(.A(G119), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G116), .ZN(new_n188));
  INV_X1    g002(.A(G116), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G119), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT2), .B(G113), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n192), .A2(new_n194), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n191), .A2(new_n193), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n195), .A2(new_n196), .ZN(new_n197));
  INV_X1    g011(.A(KEYINPUT30), .ZN(new_n198));
  NAND2_X1  g012(.A1(KEYINPUT0), .A2(G128), .ZN(new_n199));
  INV_X1    g013(.A(G143), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n200), .A2(G146), .ZN(new_n201));
  XNOR2_X1  g015(.A(KEYINPUT64), .B(G143), .ZN(new_n202));
  AOI211_X1 g016(.A(new_n199), .B(new_n201), .C1(new_n202), .C2(G146), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(new_n199), .ZN(new_n205));
  NOR2_X1   g019(.A1(KEYINPUT0), .A2(G128), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n200), .A2(KEYINPUT64), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT64), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G143), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G146), .ZN(new_n212));
  NOR2_X1   g026(.A1(new_n212), .A2(G143), .ZN(new_n213));
  OAI211_X1 g027(.A(KEYINPUT65), .B(new_n207), .C1(new_n211), .C2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n213), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n216), .B1(new_n202), .B2(G146), .ZN(new_n217));
  AOI21_X1  g031(.A(KEYINPUT65), .B1(new_n217), .B2(new_n207), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n204), .B1(new_n215), .B2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT68), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT65), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n208), .A2(new_n210), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n213), .B1(new_n223), .B2(new_n212), .ZN(new_n224));
  INV_X1    g038(.A(new_n207), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n222), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n203), .B1(new_n226), .B2(new_n214), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(KEYINPUT68), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n231), .A2(new_n233), .A3(new_n237), .A4(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT66), .ZN(new_n239));
  AND2_X1   g053(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n238), .A2(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n236), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT69), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(new_n238), .B(new_n239), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .A3(new_n236), .ZN(new_n246));
  NAND4_X1  g060(.A1(new_n221), .A2(new_n228), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n201), .B1(new_n202), .B2(G146), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT1), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(new_n249), .A3(G128), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  INV_X1    g065(.A(new_n201), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n251), .B1(new_n252), .B2(KEYINPUT1), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n250), .B1(new_n224), .B2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n232), .A2(G134), .ZN(new_n255));
  AOI21_X1  g069(.A(new_n237), .B1(new_n255), .B2(new_n234), .ZN(new_n256));
  XNOR2_X1  g070(.A(new_n256), .B(KEYINPUT67), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n254), .A2(new_n245), .A3(new_n257), .ZN(new_n258));
  AOI21_X1  g072(.A(new_n198), .B1(new_n247), .B2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n242), .ZN(new_n260));
  OAI211_X1 g074(.A(new_n258), .B(new_n198), .C1(new_n260), .C2(new_n219), .ZN(new_n261));
  INV_X1    g075(.A(new_n261), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n197), .B1(new_n259), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n258), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n226), .A2(new_n214), .ZN(new_n265));
  AOI21_X1  g079(.A(KEYINPUT68), .B1(new_n265), .B2(new_n204), .ZN(new_n266));
  AOI211_X1 g080(.A(new_n220), .B(new_n203), .C1(new_n226), .C2(new_n214), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(new_n244), .A2(new_n246), .ZN(new_n269));
  AOI21_X1  g083(.A(new_n264), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(new_n197), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g086(.A(G210), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n273), .A2(G237), .A3(G953), .ZN(new_n274));
  XNOR2_X1  g088(.A(new_n274), .B(KEYINPUT27), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n275), .B(KEYINPUT70), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT26), .B(G101), .ZN(new_n277));
  XNOR2_X1  g091(.A(new_n276), .B(new_n277), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n263), .A2(new_n272), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(KEYINPUT31), .ZN(new_n280));
  OAI21_X1  g094(.A(new_n258), .B1(new_n260), .B2(new_n219), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(new_n197), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT28), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n283), .B1(new_n270), .B2(new_n271), .ZN(new_n284));
  AND4_X1   g098(.A1(new_n283), .A2(new_n247), .A3(new_n271), .A4(new_n258), .ZN(new_n285));
  OAI21_X1  g099(.A(new_n282), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  INV_X1    g100(.A(new_n278), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT31), .ZN(new_n289));
  NAND4_X1  g103(.A1(new_n263), .A2(new_n289), .A3(new_n272), .A4(new_n278), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n280), .A2(new_n288), .A3(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(G472), .A2(G902), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT71), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT32), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(KEYINPUT71), .A3(new_n292), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n295), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n292), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n284), .A2(new_n285), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n270), .A2(new_n271), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT29), .ZN(new_n303));
  NOR2_X1   g117(.A1(new_n287), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(G902), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n303), .B1(new_n286), .B2(new_n287), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n263), .A2(new_n272), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(new_n278), .ZN(new_n308));
  OAI21_X1  g122(.A(new_n305), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(G472), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n298), .A2(new_n299), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT72), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT72), .ZN(new_n313));
  NAND4_X1  g127(.A1(new_n298), .A2(new_n313), .A3(new_n310), .A4(new_n299), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(G902), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT79), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n317), .A2(KEYINPUT25), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n187), .A2(G128), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT75), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n319), .A2(new_n320), .A3(KEYINPUT23), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n187), .A2(G128), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n321), .B(new_n322), .C1(new_n320), .C2(KEYINPUT23), .ZN(new_n323));
  INV_X1    g137(.A(new_n322), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n324), .A2(new_n319), .A3(new_n320), .A4(KEYINPUT23), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT76), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(KEYINPUT76), .B1(new_n323), .B2(new_n325), .ZN(new_n329));
  OAI21_X1  g143(.A(G110), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  OR2_X1    g144(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(KEYINPUT77), .ZN(new_n332));
  XNOR2_X1  g146(.A(G125), .B(G140), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n333), .A2(KEYINPUT16), .ZN(new_n334));
  INV_X1    g148(.A(G125), .ZN(new_n335));
  OR3_X1    g149(.A1(new_n335), .A2(KEYINPUT16), .A3(G140), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(G146), .A3(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(new_n337), .ZN(new_n338));
  AOI21_X1  g152(.A(G146), .B1(new_n334), .B2(new_n336), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(KEYINPUT74), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n322), .B1(new_n341), .B2(new_n319), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n341), .B2(new_n319), .ZN(new_n343));
  XNOR2_X1  g157(.A(KEYINPUT24), .B(G110), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n340), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n331), .A2(new_n332), .A3(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n343), .A2(new_n344), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT78), .ZN(new_n349));
  AOI21_X1  g163(.A(G110), .B1(new_n323), .B2(new_n325), .ZN(new_n350));
  OR3_X1    g164(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n349), .B1(new_n348), .B2(new_n350), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n333), .A2(new_n212), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n351), .A2(new_n352), .A3(new_n353), .A4(new_n337), .ZN(new_n354));
  XNOR2_X1  g168(.A(KEYINPUT22), .B(G137), .ZN(new_n355));
  INV_X1    g169(.A(G221), .ZN(new_n356));
  INV_X1    g170(.A(G234), .ZN(new_n357));
  NOR3_X1   g171(.A1(new_n356), .A2(new_n357), .A3(G953), .ZN(new_n358));
  XOR2_X1   g172(.A(new_n355), .B(new_n358), .Z(new_n359));
  INV_X1    g173(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n347), .A2(new_n354), .A3(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(new_n360), .B1(new_n347), .B2(new_n354), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n316), .B(new_n318), .C1(new_n362), .C2(new_n363), .ZN(new_n364));
  OAI21_X1  g178(.A(G217), .B1(new_n357), .B2(G902), .ZN(new_n365));
  XNOR2_X1  g179(.A(new_n365), .B(KEYINPUT73), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n347), .A2(new_n354), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n369), .A2(new_n359), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n361), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n318), .B1(new_n371), .B2(new_n316), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n366), .A2(new_n316), .ZN(new_n373));
  XOR2_X1   g187(.A(new_n373), .B(KEYINPUT80), .Z(new_n374));
  INV_X1    g188(.A(new_n371), .ZN(new_n375));
  OAI22_X1  g189(.A1(new_n368), .A2(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT9), .B(G234), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n378), .B(KEYINPUT81), .ZN(new_n379));
  AOI21_X1  g193(.A(new_n356), .B1(new_n379), .B2(new_n316), .ZN(new_n380));
  XNOR2_X1  g194(.A(G110), .B(G140), .ZN(new_n381));
  INV_X1    g195(.A(G953), .ZN(new_n382));
  NAND2_X1  g196(.A1(new_n382), .A2(G227), .ZN(new_n383));
  XNOR2_X1  g197(.A(new_n381), .B(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(new_n384), .B(KEYINPUT82), .Z(new_n385));
  INV_X1    g199(.A(G104), .ZN(new_n386));
  NOR3_X1   g200(.A1(new_n386), .A2(KEYINPUT3), .A3(G107), .ZN(new_n387));
  XOR2_X1   g201(.A(KEYINPUT83), .B(G104), .Z(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(G107), .ZN(new_n389));
  XNOR2_X1  g203(.A(KEYINPUT83), .B(G104), .ZN(new_n390));
  INV_X1    g204(.A(G107), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(KEYINPUT3), .ZN(new_n393));
  INV_X1    g207(.A(G101), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n389), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(G104), .B2(new_n391), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G101), .ZN(new_n397));
  AND2_X1   g211(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g212(.A(new_n250), .ZN(new_n399));
  OAI21_X1  g213(.A(KEYINPUT1), .B1(new_n202), .B2(G146), .ZN(new_n400));
  AOI21_X1  g214(.A(new_n248), .B1(G128), .B2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n398), .B1(new_n399), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n402), .B1(new_n254), .B2(new_n398), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n269), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT12), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n260), .A2(new_n405), .ZN(new_n406));
  AOI22_X1  g220(.A1(new_n404), .A2(new_n405), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT10), .ZN(new_n408));
  AND2_X1   g222(.A1(new_n254), .A2(KEYINPUT10), .ZN(new_n409));
  AOI22_X1  g223(.A1(new_n402), .A2(new_n408), .B1(new_n398), .B2(new_n409), .ZN(new_n410));
  OR3_X1    g224(.A1(new_n386), .A2(KEYINPUT3), .A3(G107), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n390), .B2(new_n391), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n412), .B1(KEYINPUT3), .B2(new_n392), .ZN(new_n413));
  NOR2_X1   g227(.A1(new_n413), .A2(new_n394), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n389), .A2(new_n393), .ZN(new_n418));
  XNOR2_X1  g232(.A(KEYINPUT84), .B(KEYINPUT4), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND3_X1  g234(.A1(new_n418), .A2(G101), .A3(new_n420), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n417), .A2(new_n221), .A3(new_n228), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n269), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n410), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(new_n424), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n385), .B1(new_n407), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n410), .A2(new_n422), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n269), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n424), .A3(new_n384), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n430), .A2(new_n316), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(G469), .ZN(new_n432));
  INV_X1    g246(.A(G469), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n424), .A2(new_n384), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n407), .A2(new_n434), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n384), .B1(new_n428), .B2(new_n424), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n433), .B(new_n316), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n380), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(G214), .B1(G237), .B2(G902), .ZN(new_n439));
  INV_X1    g253(.A(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n395), .A2(KEYINPUT4), .ZN(new_n441));
  OAI211_X1 g255(.A(new_n197), .B(new_n421), .C1(new_n414), .C2(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n192), .A2(KEYINPUT5), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n188), .A2(KEYINPUT5), .ZN(new_n444));
  INV_X1    g258(.A(G113), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  AOI22_X1  g260(.A1(new_n443), .A2(new_n446), .B1(new_n192), .B2(new_n194), .ZN(new_n447));
  AND3_X1   g261(.A1(new_n447), .A2(new_n395), .A3(new_n397), .ZN(new_n448));
  INV_X1    g262(.A(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(G110), .B(G122), .ZN(new_n450));
  AND3_X1   g264(.A1(new_n442), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(new_n450), .B(KEYINPUT85), .Z(new_n452));
  AOI21_X1  g266(.A(new_n452), .B1(new_n442), .B2(new_n449), .ZN(new_n453));
  OAI21_X1  g267(.A(KEYINPUT6), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  OR2_X1    g268(.A1(new_n453), .A2(KEYINPUT6), .ZN(new_n455));
  XNOR2_X1  g269(.A(KEYINPUT86), .B(G224), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n382), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n227), .A2(G125), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT87), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n254), .A2(new_n335), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n459), .A2(new_n460), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(new_n462), .ZN(new_n463));
  AOI21_X1  g277(.A(new_n460), .B1(new_n459), .B2(new_n461), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n458), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n464), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n457), .A3(new_n462), .ZN(new_n467));
  AOI22_X1  g281(.A1(new_n454), .A2(new_n455), .B1(new_n465), .B2(new_n467), .ZN(new_n468));
  XNOR2_X1  g282(.A(new_n450), .B(KEYINPUT8), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n447), .B1(new_n395), .B2(new_n397), .ZN(new_n470));
  OAI21_X1  g284(.A(new_n469), .B1(new_n448), .B2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT88), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n459), .A2(new_n461), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT89), .ZN(new_n475));
  XNOR2_X1  g289(.A(new_n457), .B(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n474), .A2(KEYINPUT7), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n457), .A2(KEYINPUT7), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n459), .A2(new_n461), .A3(new_n478), .ZN(new_n479));
  OAI211_X1 g293(.A(KEYINPUT88), .B(new_n469), .C1(new_n448), .C2(new_n470), .ZN(new_n480));
  NAND4_X1  g294(.A1(new_n473), .A2(new_n477), .A3(new_n479), .A4(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(new_n316), .B1(new_n481), .B2(new_n451), .ZN(new_n482));
  OAI21_X1  g296(.A(G210), .B1(G237), .B2(G902), .ZN(new_n483));
  INV_X1    g297(.A(new_n483), .ZN(new_n484));
  NOR3_X1   g298(.A1(new_n468), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n484), .B1(new_n468), .B2(new_n482), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n440), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G237), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n489), .A2(new_n382), .A3(G214), .ZN(new_n490));
  OR2_X1    g304(.A1(new_n490), .A2(new_n200), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n202), .A2(new_n490), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT90), .ZN(new_n495));
  NOR2_X1   g309(.A1(KEYINPUT90), .A2(KEYINPUT91), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  OAI211_X1 g311(.A(KEYINPUT18), .B(G131), .C1(new_n495), .C2(new_n497), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n333), .A2(G146), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n333), .A2(G146), .ZN(new_n500));
  AOI21_X1  g314(.A(KEYINPUT91), .B1(KEYINPUT18), .B2(G131), .ZN(new_n501));
  AOI211_X1 g315(.A(new_n499), .B(new_n500), .C1(new_n494), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n493), .A2(KEYINPUT17), .A3(G131), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n493), .B(G131), .ZN(new_n505));
  OAI211_X1 g319(.A(new_n340), .B(new_n504), .C1(new_n505), .C2(KEYINPUT17), .ZN(new_n506));
  XNOR2_X1  g320(.A(G113), .B(G122), .ZN(new_n507));
  XNOR2_X1  g321(.A(new_n507), .B(new_n386), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n503), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n508), .B1(new_n503), .B2(new_n506), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n316), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(G475), .ZN(new_n513));
  AND2_X1   g327(.A1(new_n505), .A2(new_n337), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n333), .B(KEYINPUT19), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n212), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n516), .B(KEYINPUT92), .ZN(new_n517));
  AOI22_X1  g331(.A1(new_n514), .A2(new_n517), .B1(new_n498), .B2(new_n502), .ZN(new_n518));
  OAI21_X1  g332(.A(new_n509), .B1(new_n518), .B2(new_n508), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT20), .ZN(new_n520));
  NOR2_X1   g334(.A1(G475), .A2(G902), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n520), .B1(new_n519), .B2(new_n521), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(G952), .ZN(new_n526));
  AOI211_X1 g340(.A(G953), .B(new_n526), .C1(G234), .C2(G237), .ZN(new_n527));
  OAI211_X1 g341(.A(G902), .B(G953), .C1(new_n357), .C2(new_n489), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT96), .ZN(new_n529));
  XNOR2_X1  g343(.A(KEYINPUT21), .B(G898), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n200), .A2(G128), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n534), .B1(new_n202), .B2(G128), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n535), .A2(KEYINPUT13), .ZN(new_n536));
  OR3_X1    g350(.A1(new_n223), .A2(KEYINPUT13), .A3(new_n251), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(G134), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n535), .A2(new_n230), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT93), .ZN(new_n541));
  NAND4_X1  g355(.A1(new_n536), .A2(new_n537), .A3(new_n541), .A4(G134), .ZN(new_n542));
  INV_X1    g356(.A(G122), .ZN(new_n543));
  NOR2_X1   g357(.A1(new_n543), .A2(G116), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n189), .A2(G122), .ZN(new_n545));
  OR3_X1    g359(.A1(new_n544), .A2(new_n545), .A3(G107), .ZN(new_n546));
  OAI21_X1  g360(.A(G107), .B1(new_n544), .B2(new_n545), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n539), .A2(new_n540), .A3(new_n542), .A4(new_n548), .ZN(new_n549));
  XNOR2_X1  g363(.A(new_n535), .B(new_n230), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT14), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n544), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n545), .A2(KEYINPUT14), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n552), .B1(new_n553), .B2(new_n544), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT94), .ZN(new_n555));
  AND3_X1   g369(.A1(new_n554), .A2(new_n555), .A3(G107), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n555), .B1(new_n554), .B2(G107), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n550), .B(new_n546), .C1(new_n556), .C2(new_n557), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n379), .A2(G217), .A3(new_n382), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n549), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n559), .B1(new_n549), .B2(new_n558), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n560), .B1(new_n561), .B2(KEYINPUT95), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT95), .ZN(new_n563));
  AOI211_X1 g377(.A(new_n563), .B(new_n559), .C1(new_n549), .C2(new_n558), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n316), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(G478), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n566), .A2(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  OAI221_X1 g382(.A(new_n316), .B1(KEYINPUT15), .B2(new_n566), .C1(new_n562), .C2(new_n564), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NOR2_X1   g384(.A1(new_n533), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n438), .A2(new_n488), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n315), .A2(new_n377), .A3(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(KEYINPUT97), .B(G101), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n574), .B(new_n575), .ZN(G3));
  AND2_X1   g390(.A1(new_n295), .A2(new_n297), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n291), .A2(new_n316), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(G472), .ZN(new_n579));
  NAND4_X1  g393(.A1(new_n577), .A2(new_n438), .A3(new_n377), .A4(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n487), .B1(new_n485), .B2(new_n582), .ZN(new_n583));
  NOR4_X1   g397(.A1(new_n468), .A2(new_n482), .A3(KEYINPUT98), .A4(new_n484), .ZN(new_n584));
  OR2_X1    g398(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n439), .ZN(new_n586));
  AND2_X1   g400(.A1(new_n561), .A2(KEYINPUT99), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n560), .B1(new_n561), .B2(KEYINPUT99), .ZN(new_n588));
  OAI21_X1  g402(.A(KEYINPUT33), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OR2_X1    g403(.A1(new_n562), .A2(new_n564), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n589), .B1(new_n590), .B2(KEYINPUT33), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n591), .A2(G478), .A3(new_n316), .ZN(new_n592));
  INV_X1    g406(.A(new_n565), .ZN(new_n593));
  XOR2_X1   g407(.A(KEYINPUT100), .B(G478), .Z(new_n594));
  OAI21_X1  g408(.A(new_n592), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n524), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n586), .A2(new_n596), .A3(new_n531), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n581), .A2(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT34), .B(G104), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G6));
  INV_X1    g414(.A(new_n570), .ZN(new_n601));
  NOR3_X1   g415(.A1(new_n586), .A2(new_n601), .A3(new_n533), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n581), .A2(new_n602), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT35), .B(G107), .Z(new_n604));
  XNOR2_X1  g418(.A(new_n603), .B(new_n604), .ZN(G9));
  AND2_X1   g419(.A1(new_n577), .A2(new_n579), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n360), .A2(KEYINPUT36), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n369), .B(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n374), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n610), .B1(new_n368), .B2(new_n372), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT101), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT101), .ZN(new_n613));
  OAI211_X1 g427(.A(new_n613), .B(new_n610), .C1(new_n368), .C2(new_n372), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n606), .A2(new_n573), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT37), .B(G110), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G12));
  NOR2_X1   g432(.A1(new_n586), .A2(new_n601), .ZN(new_n619));
  INV_X1    g433(.A(G900), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n527), .B1(new_n529), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n524), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(new_n615), .ZN(new_n623));
  INV_X1    g437(.A(new_n438), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n315), .A2(new_n619), .A3(new_n622), .A4(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G128), .ZN(G30));
  INV_X1    g441(.A(new_n301), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n278), .B1(new_n628), .B2(new_n272), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n629), .B1(new_n307), .B2(new_n278), .ZN(new_n630));
  OAI21_X1  g444(.A(G472), .B1(new_n630), .B2(G902), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n298), .A2(new_n299), .A3(new_n631), .ZN(new_n632));
  XNOR2_X1  g446(.A(new_n632), .B(KEYINPUT102), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n621), .B(KEYINPUT39), .Z(new_n634));
  NAND2_X1  g448(.A1(new_n438), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT103), .B(KEYINPUT40), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n486), .A2(new_n487), .ZN(new_n639));
  XNOR2_X1  g453(.A(new_n639), .B(KEYINPUT38), .ZN(new_n640));
  AND3_X1   g454(.A1(new_n524), .A2(new_n570), .A3(new_n439), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n638), .A2(new_n623), .A3(new_n640), .A4(new_n641), .ZN(new_n642));
  OR3_X1    g456(.A1(new_n633), .A2(new_n637), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(new_n223), .ZN(G45));
  NAND3_X1  g458(.A1(new_n585), .A2(new_n439), .A3(new_n615), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n596), .ZN(new_n647));
  INV_X1    g461(.A(new_n621), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  NAND4_X1  g464(.A1(new_n315), .A2(new_n438), .A3(new_n646), .A4(new_n650), .ZN(new_n651));
  XNOR2_X1  g465(.A(KEYINPUT104), .B(G146), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n651), .B(new_n652), .ZN(G48));
  OAI21_X1  g467(.A(new_n316), .B1(new_n435), .B2(new_n436), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G469), .ZN(new_n655));
  INV_X1    g469(.A(new_n380), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n655), .A2(new_n656), .A3(new_n437), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT105), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND4_X1  g473(.A1(new_n655), .A2(KEYINPUT105), .A3(new_n656), .A4(new_n437), .ZN(new_n660));
  AND2_X1   g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n315), .A2(new_n377), .A3(new_n597), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT41), .B(G113), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G15));
  NAND4_X1  g478(.A1(new_n315), .A2(new_n377), .A3(new_n602), .A4(new_n661), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G116), .ZN(G18));
  NOR3_X1   g480(.A1(new_n657), .A2(new_n570), .A3(new_n533), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n315), .A2(new_n646), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  AND3_X1   g483(.A1(new_n659), .A2(new_n532), .A3(new_n660), .ZN(new_n670));
  OAI21_X1  g484(.A(new_n641), .B1(new_n583), .B2(new_n584), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(KEYINPUT106), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT106), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n641), .B(new_n673), .C1(new_n583), .C2(new_n584), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  OAI211_X1 g489(.A(new_n280), .B(new_n290), .C1(new_n302), .C2(new_n278), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(new_n292), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n579), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(new_n376), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(KEYINPUT107), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n670), .A2(new_n675), .A3(new_n679), .A4(KEYINPUT107), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(new_n684), .B(G122), .ZN(G24));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n686));
  OAI21_X1  g500(.A(new_n686), .B1(new_n623), .B2(new_n678), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n615), .A2(new_n579), .A3(KEYINPUT108), .A4(new_n677), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g503(.A1(new_n586), .A2(new_n657), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n689), .A2(new_n650), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(G125), .ZN(G27));
  NOR2_X1   g506(.A1(new_n639), .A2(new_n440), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g508(.A1(new_n624), .A2(new_n694), .ZN(new_n695));
  NAND4_X1  g509(.A1(new_n315), .A2(new_n377), .A3(new_n650), .A4(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT42), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n310), .A2(new_n299), .ZN(new_n698));
  AOI21_X1  g512(.A(KEYINPUT32), .B1(new_n291), .B2(new_n292), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n377), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n700), .B(KEYINPUT109), .ZN(new_n701));
  NOR4_X1   g515(.A1(new_n649), .A2(new_n624), .A3(new_n697), .A4(new_n694), .ZN(new_n702));
  AOI22_X1  g516(.A1(new_n696), .A2(new_n697), .B1(new_n701), .B2(new_n702), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(new_n237), .ZN(G33));
  INV_X1    g518(.A(new_n622), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n705), .A2(new_n601), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(KEYINPUT110), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n315), .A2(new_n377), .A3(new_n695), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  NAND2_X1  g523(.A1(new_n595), .A2(new_n525), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT43), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n606), .A2(new_n711), .A3(new_n623), .ZN(new_n712));
  OR2_X1    g526(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n430), .B(KEYINPUT45), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(G469), .ZN(new_n716));
  NAND2_X1  g530(.A1(G469), .A2(G902), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n716), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n718), .A2(new_n437), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT46), .B1(new_n716), .B2(new_n717), .ZN(new_n720));
  OAI21_X1  g534(.A(new_n656), .B1(new_n719), .B2(new_n720), .ZN(new_n721));
  INV_X1    g535(.A(new_n634), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND4_X1  g537(.A1(new_n713), .A2(new_n693), .A3(new_n714), .A4(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G137), .ZN(G39));
  XNOR2_X1  g539(.A(new_n721), .B(KEYINPUT47), .ZN(new_n726));
  NAND3_X1  g540(.A1(new_n650), .A2(new_n376), .A3(new_n693), .ZN(new_n727));
  OR3_X1    g541(.A1(new_n726), .A2(new_n315), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G140), .ZN(G42));
  INV_X1    g543(.A(new_n527), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n711), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n731), .A2(new_n679), .ZN(new_n732));
  AND2_X1   g546(.A1(new_n655), .A2(new_n437), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(new_n380), .ZN(new_n734));
  AOI211_X1 g548(.A(new_n694), .B(new_n732), .C1(new_n726), .C2(new_n734), .ZN(new_n735));
  NOR4_X1   g549(.A1(new_n732), .A2(new_n439), .A3(new_n640), .A4(new_n657), .ZN(new_n736));
  XOR2_X1   g550(.A(new_n736), .B(KEYINPUT50), .Z(new_n737));
  NOR2_X1   g551(.A1(new_n694), .A2(new_n657), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(KEYINPUT118), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n739), .A2(new_n731), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(KEYINPUT119), .ZN(new_n741));
  AOI211_X1 g555(.A(new_n735), .B(new_n737), .C1(new_n689), .C2(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n633), .A2(new_n739), .A3(new_n377), .A4(new_n527), .ZN(new_n743));
  XOR2_X1   g557(.A(new_n743), .B(KEYINPUT120), .Z(new_n744));
  NOR2_X1   g558(.A1(new_n595), .A2(new_n524), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n742), .A2(KEYINPUT51), .A3(new_n746), .ZN(new_n747));
  AOI21_X1  g561(.A(KEYINPUT51), .B1(new_n742), .B2(new_n746), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n741), .A2(new_n701), .ZN(new_n749));
  OR3_X1    g563(.A1(new_n749), .A2(KEYINPUT121), .A3(KEYINPUT48), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n749), .A2(KEYINPUT48), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT122), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n749), .A2(KEYINPUT122), .A3(KEYINPUT48), .ZN(new_n754));
  OAI21_X1  g568(.A(KEYINPUT121), .B1(new_n749), .B2(KEYINPUT48), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n750), .A2(new_n753), .A3(new_n754), .A4(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n744), .A2(new_n647), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n732), .A2(new_n586), .A3(new_n657), .ZN(new_n758));
  NOR3_X1   g572(.A1(new_n758), .A2(new_n526), .A3(G953), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(new_n757), .A3(new_n759), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n747), .A2(new_n748), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n662), .A2(new_n665), .A3(new_n668), .A4(new_n684), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT112), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n645), .B1(new_n312), .B2(new_n314), .ZN(new_n765));
  AOI22_X1  g579(.A1(new_n765), .A2(new_n667), .B1(new_n682), .B2(new_n683), .ZN(new_n766));
  NAND4_X1  g580(.A1(new_n766), .A2(KEYINPUT112), .A3(new_n662), .A4(new_n665), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  AOI211_X1 g582(.A(new_n376), .B(new_n572), .C1(new_n312), .C2(new_n314), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n488), .A2(new_n532), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n580), .A2(new_n596), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n769), .A2(KEYINPUT113), .A3(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT113), .ZN(new_n773));
  INV_X1    g587(.A(new_n771), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n773), .B1(new_n574), .B2(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n570), .B(KEYINPUT114), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n776), .A2(new_n525), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n580), .A2(new_n770), .A3(new_n777), .ZN(new_n778));
  OR2_X1    g592(.A1(new_n616), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g593(.A1(new_n772), .A2(new_n775), .A3(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n776), .A2(new_n705), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n693), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(KEYINPUT115), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT115), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(new_n784), .A3(new_n693), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n315), .A2(new_n625), .A3(new_n783), .A4(new_n785), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n689), .A2(new_n650), .A3(new_n695), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n708), .A2(new_n786), .A3(new_n787), .ZN(new_n788));
  NOR2_X1   g602(.A1(new_n703), .A2(new_n788), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n768), .A2(new_n780), .A3(new_n789), .ZN(new_n790));
  INV_X1    g604(.A(KEYINPUT116), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n768), .A2(new_n780), .A3(new_n789), .A4(KEYINPUT116), .ZN(new_n793));
  AND3_X1   g607(.A1(new_n626), .A2(new_n651), .A3(new_n691), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n624), .A2(new_n611), .A3(new_n621), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n795), .A2(new_n632), .A3(new_n675), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n794), .A2(KEYINPUT52), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n626), .A2(new_n651), .A3(new_n691), .A4(new_n796), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n797), .A2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n792), .A2(new_n793), .A3(new_n801), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(KEYINPUT53), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT117), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n801), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n797), .A2(KEYINPUT117), .A3(new_n800), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT53), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n807), .A2(new_n792), .A3(new_n808), .A4(new_n793), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n803), .A2(KEYINPUT54), .A3(new_n809), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n762), .A2(new_n808), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n780), .A2(new_n789), .A3(new_n811), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n812), .B1(new_n805), .B2(new_n806), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n813), .B1(new_n802), .B2(new_n808), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT54), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n761), .A2(new_n810), .A3(new_n816), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n817), .B1(G952), .B2(G953), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n640), .A2(new_n710), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n377), .A2(new_n656), .A3(new_n439), .ZN(new_n820));
  XNOR2_X1  g634(.A(new_n820), .B(KEYINPUT111), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n733), .B(KEYINPUT49), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n633), .A2(new_n819), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n818), .A2(new_n823), .ZN(G75));
  NOR2_X1   g638(.A1(new_n382), .A2(G952), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT56), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n802), .A2(new_n808), .ZN(new_n827));
  INV_X1    g641(.A(new_n813), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(G902), .ZN(new_n830));
  OAI21_X1  g644(.A(new_n826), .B1(new_n830), .B2(new_n273), .ZN(new_n831));
  AND4_X1   g645(.A1(new_n465), .A2(new_n454), .A3(new_n455), .A4(new_n467), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n832), .A2(new_n468), .ZN(new_n833));
  XNOR2_X1  g647(.A(new_n833), .B(KEYINPUT55), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n825), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  OAI211_X1 g650(.A(new_n826), .B(new_n834), .C1(new_n830), .C2(new_n273), .ZN(new_n837));
  AND2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(G51));
  XNOR2_X1  g652(.A(new_n814), .B(KEYINPUT54), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n717), .B(KEYINPUT57), .ZN(new_n840));
  OAI22_X1  g654(.A1(new_n839), .A2(new_n840), .B1(new_n436), .B2(new_n435), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n830), .A2(new_n716), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n825), .B1(new_n841), .B2(new_n842), .ZN(G54));
  INV_X1    g657(.A(new_n830), .ZN(new_n844));
  AND2_X1   g658(.A1(KEYINPUT58), .A2(G475), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n844), .A2(new_n519), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n519), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n846), .A2(new_n847), .A3(new_n825), .ZN(G60));
  INV_X1    g662(.A(new_n825), .ZN(new_n849));
  NAND2_X1  g663(.A1(G478), .A2(G902), .ZN(new_n850));
  XOR2_X1   g664(.A(new_n850), .B(KEYINPUT59), .Z(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n816), .B2(new_n810), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n849), .B1(new_n852), .B2(new_n591), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n829), .A2(KEYINPUT54), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n854), .A2(new_n816), .ZN(new_n855));
  INV_X1    g669(.A(new_n851), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n591), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(KEYINPUT123), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT123), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n855), .A2(new_n860), .A3(new_n857), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n853), .B1(new_n859), .B2(new_n861), .ZN(G63));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n863));
  INV_X1    g677(.A(KEYINPUT61), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n608), .ZN(new_n866));
  NAND2_X1  g680(.A1(G217), .A2(G902), .ZN(new_n867));
  XNOR2_X1  g681(.A(new_n867), .B(KEYINPUT60), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n814), .A2(new_n866), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n865), .B1(new_n869), .B2(new_n864), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n375), .B1(new_n814), .B2(new_n868), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n870), .A2(new_n849), .A3(new_n871), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n863), .B1(new_n871), .B2(new_n849), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n868), .B1(new_n827), .B2(new_n828), .ZN(new_n874));
  AOI21_X1  g688(.A(KEYINPUT124), .B1(new_n874), .B2(new_n608), .ZN(new_n875));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n876));
  NOR4_X1   g690(.A1(new_n814), .A2(new_n876), .A3(new_n866), .A4(new_n868), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n873), .A2(new_n875), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n872), .B1(new_n878), .B2(KEYINPUT61), .ZN(G66));
  INV_X1    g693(.A(new_n456), .ZN(new_n880));
  OAI21_X1  g694(.A(G953), .B1(new_n880), .B2(new_n530), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n768), .A2(new_n780), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n882), .B2(G953), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n454), .B(new_n455), .C1(G898), .C2(new_n382), .ZN(new_n884));
  XNOR2_X1  g698(.A(new_n883), .B(new_n884), .ZN(G69));
  AOI21_X1  g699(.A(new_n382), .B1(G227), .B2(G900), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n723), .A2(new_n701), .A3(new_n675), .ZN(new_n887));
  AND4_X1   g701(.A1(new_n708), .A2(new_n728), .A3(new_n724), .A4(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(new_n703), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n794), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n890), .A2(KEYINPUT127), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT127), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n888), .A2(new_n892), .A3(new_n889), .A4(new_n794), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n891), .A2(new_n382), .A3(new_n893), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n259), .A2(new_n262), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(new_n515), .ZN(new_n896));
  AOI21_X1  g710(.A(new_n896), .B1(G900), .B2(G953), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n894), .A2(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT126), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n886), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n728), .A2(new_n724), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n794), .A2(new_n643), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT62), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n315), .A2(new_n377), .ZN(new_n904));
  INV_X1    g718(.A(new_n904), .ZN(new_n905));
  AOI211_X1 g719(.A(new_n694), .B(new_n635), .C1(new_n596), .C2(new_n777), .ZN(new_n906));
  AOI211_X1 g720(.A(new_n901), .B(new_n903), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n896), .B1(new_n907), .B2(G953), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n898), .ZN(new_n909));
  XOR2_X1   g723(.A(new_n900), .B(new_n909), .Z(G72));
  AND3_X1   g724(.A1(new_n891), .A2(new_n882), .A3(new_n893), .ZN(new_n911));
  NAND2_X1  g725(.A1(G472), .A2(G902), .ZN(new_n912));
  XOR2_X1   g726(.A(new_n912), .B(KEYINPUT63), .Z(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n307), .B(new_n287), .C1(new_n911), .C2(new_n914), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n907), .B2(new_n882), .ZN(new_n916));
  OR2_X1    g730(.A1(new_n307), .A2(new_n287), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n915), .B(new_n849), .C1(new_n916), .C2(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n803), .A2(new_n809), .ZN(new_n919));
  INV_X1    g733(.A(new_n308), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n914), .B1(new_n920), .B2(new_n279), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n918), .B1(new_n919), .B2(new_n921), .ZN(G57));
endmodule


