//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 1 1 1 1 0 1 1 0 1 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 1 0 0 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:35:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1215, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1285, new_n1286;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G13), .ZN(new_n204));
  OAI211_X1 g0004(.A(new_n204), .B(G250), .C1(G257), .C2(G264), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT0), .Z(new_n206));
  AOI22_X1  g0006(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n207));
  INV_X1    g0007(.A(G50), .ZN(new_n208));
  INV_X1    g0008(.A(G226), .ZN(new_n209));
  INV_X1    g0009(.A(G77), .ZN(new_n210));
  INV_X1    g0010(.A(G244), .ZN(new_n211));
  OAI221_X1 g0011(.A(new_n207), .B1(new_n208), .B2(new_n209), .C1(new_n210), .C2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G97), .B2(G257), .ZN(new_n213));
  INV_X1    g0013(.A(G58), .ZN(new_n214));
  INV_X1    g0014(.A(G232), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  XNOR2_X1  g0016(.A(KEYINPUT65), .B(G68), .ZN(new_n217));
  OAI221_X1 g0017(.A(new_n213), .B1(new_n214), .B2(new_n215), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g0021(.A(new_n203), .B1(new_n218), .B2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT1), .ZN(new_n223));
  NAND2_X1  g0023(.A1(G1), .A2(G13), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G20), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT64), .ZN(new_n227));
  NOR2_X1   g0027(.A1(G58), .A2(G68), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  NAND2_X1  g0029(.A1(new_n229), .A2(G50), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  AOI211_X1 g0031(.A(new_n206), .B(new_n223), .C1(new_n227), .C2(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G250), .B(G257), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G264), .ZN(new_n234));
  XOR2_X1   g0034(.A(new_n234), .B(G270), .Z(new_n235));
  XOR2_X1   g0035(.A(G238), .B(G244), .Z(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G226), .B(G232), .Z(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n235), .B(new_n240), .Z(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G107), .B(G116), .Z(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  XNOR2_X1  g0048(.A(KEYINPUT3), .B(G33), .ZN(new_n249));
  INV_X1    g0049(.A(G1698), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n250), .A2(G222), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G223), .A2(G1698), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n249), .A2(new_n251), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(new_n224), .B1(G33), .B2(G41), .ZN(new_n254));
  OAI211_X1 g0054(.A(new_n253), .B(new_n254), .C1(G77), .C2(new_n249), .ZN(new_n255));
  INV_X1    g0055(.A(new_n254), .ZN(new_n256));
  INV_X1    g0056(.A(G41), .ZN(new_n257));
  INV_X1    g0057(.A(G45), .ZN(new_n258));
  AOI21_X1  g0058(.A(G1), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(KEYINPUT67), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(G41), .B2(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(KEYINPUT67), .ZN(new_n264));
  NAND4_X1  g0064(.A1(new_n256), .A2(new_n261), .A3(G274), .A4(new_n264), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n254), .A2(new_n259), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n255), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  OAI22_X1  g0070(.A1(new_n268), .A2(new_n269), .B1(KEYINPUT74), .B2(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n262), .A2(G13), .A3(G20), .ZN(new_n272));
  INV_X1    g0072(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(new_n208), .ZN(new_n274));
  NAND3_X1  g0074(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n224), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n276), .B1(new_n262), .B2(G20), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G50), .ZN(new_n278));
  INV_X1    g0078(.A(G20), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n279), .B1(new_n228), .B2(new_n208), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G20), .A2(G33), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n280), .B1(G150), .B2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT8), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n283), .A2(KEYINPUT68), .A3(G58), .ZN(new_n284));
  XOR2_X1   g0084(.A(KEYINPUT8), .B(G58), .Z(new_n285));
  OAI21_X1  g0085(.A(new_n284), .B1(new_n285), .B2(KEYINPUT68), .ZN(new_n286));
  INV_X1    g0086(.A(G33), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n287), .A2(G20), .ZN(new_n288));
  INV_X1    g0088(.A(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n282), .B1(new_n286), .B2(new_n289), .ZN(new_n290));
  AOI21_X1  g0090(.A(KEYINPUT69), .B1(new_n290), .B2(new_n276), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n276), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT69), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n274), .B(new_n278), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n270), .A2(KEYINPUT74), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n296), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n271), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n268), .A2(G200), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT75), .ZN(new_n302));
  OAI211_X1 g0102(.A(new_n300), .B(new_n301), .C1(new_n302), .C2(KEYINPUT10), .ZN(new_n303));
  INV_X1    g0103(.A(new_n271), .ZN(new_n304));
  INV_X1    g0104(.A(new_n299), .ZN(new_n305));
  OAI211_X1 g0105(.A(new_n301), .B(new_n304), .C1(new_n305), .C2(new_n297), .ZN(new_n306));
  OAI211_X1 g0106(.A(new_n302), .B(new_n304), .C1(new_n305), .C2(new_n297), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT10), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n306), .A2(new_n307), .A3(new_n308), .ZN(new_n309));
  AND2_X1   g0109(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n268), .A2(G179), .ZN(new_n311));
  INV_X1    g0111(.A(G169), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n311), .B1(new_n312), .B2(new_n268), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n295), .A2(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n249), .A2(G232), .A3(new_n250), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n315), .B(KEYINPUT70), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n249), .A2(G238), .A3(G1698), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n249), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n254), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n266), .A2(G244), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n320), .A2(new_n265), .A3(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n322), .A2(new_n312), .ZN(new_n323));
  XOR2_X1   g0123(.A(KEYINPUT15), .B(G87), .Z(new_n324));
  NAND2_X1  g0124(.A1(new_n324), .A2(new_n288), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT71), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n285), .A2(new_n281), .B1(G20), .B2(G77), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT71), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n324), .A2(new_n328), .A3(new_n288), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n326), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n276), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n273), .A2(new_n210), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n277), .A2(G77), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT72), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND4_X1  g0136(.A1(new_n331), .A2(KEYINPUT72), .A3(new_n332), .A4(new_n333), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n265), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n339), .B1(new_n319), .B2(new_n254), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(new_n341), .A3(new_n321), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n323), .A2(new_n338), .A3(new_n342), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n310), .A2(new_n314), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n266), .A2(G238), .ZN(new_n345));
  NOR2_X1   g0145(.A1(G226), .A2(G1698), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n346), .B1(new_n215), .B2(G1698), .ZN(new_n347));
  AOI22_X1  g0147(.A1(new_n347), .A2(new_n249), .B1(G33), .B2(G97), .ZN(new_n348));
  OAI211_X1 g0148(.A(new_n345), .B(new_n265), .C1(new_n348), .C2(new_n256), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(KEYINPUT76), .ZN(new_n351));
  OR3_X1    g0151(.A1(new_n349), .A2(KEYINPUT77), .A3(new_n351), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n351), .B1(new_n349), .B2(KEYINPUT77), .ZN(new_n353));
  OAI21_X1  g0153(.A(KEYINPUT77), .B1(new_n349), .B2(KEYINPUT13), .ZN(new_n354));
  NAND4_X1  g0154(.A1(new_n352), .A2(G190), .A3(new_n353), .A4(new_n354), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n349), .B(KEYINPUT13), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(G200), .ZN(new_n357));
  AND2_X1   g0157(.A1(KEYINPUT65), .A2(G68), .ZN(new_n358));
  NOR2_X1   g0158(.A1(KEYINPUT65), .A2(G68), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(KEYINPUT12), .B1(new_n360), .B2(new_n272), .ZN(new_n361));
  XNOR2_X1  g0161(.A(new_n361), .B(KEYINPUT78), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n272), .A2(KEYINPUT12), .A3(G68), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n277), .A2(G68), .ZN(new_n365));
  AOI22_X1  g0165(.A1(new_n217), .A2(G20), .B1(G50), .B2(new_n281), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n210), .B2(new_n289), .ZN(new_n367));
  INV_X1    g0167(.A(KEYINPUT11), .ZN(new_n368));
  AND3_X1   g0168(.A1(new_n367), .A2(new_n368), .A3(new_n276), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n368), .B1(new_n367), .B2(new_n276), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n364), .B(new_n365), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT79), .ZN(new_n372));
  AND2_X1   g0172(.A1(new_n371), .A2(new_n372), .ZN(new_n373));
  NOR2_X1   g0173(.A1(new_n371), .A2(new_n372), .ZN(new_n374));
  OAI211_X1 g0174(.A(new_n355), .B(new_n357), .C1(new_n373), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(KEYINPUT80), .ZN(new_n376));
  XNOR2_X1  g0176(.A(new_n371), .B(new_n372), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT80), .ZN(new_n378));
  NAND4_X1  g0178(.A1(new_n377), .A2(new_n378), .A3(new_n355), .A4(new_n357), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n376), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n356), .A2(G169), .ZN(new_n381));
  OR2_X1    g0181(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n352), .A2(G179), .A3(new_n353), .A4(new_n354), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n382), .A2(new_n383), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n377), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n380), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT3), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(KEYINPUT81), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT81), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT3), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(new_n392), .A3(G33), .ZN(new_n393));
  NOR2_X1   g0193(.A1(KEYINPUT3), .A2(G33), .ZN(new_n394));
  INV_X1    g0194(.A(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n279), .A3(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(KEYINPUT7), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT7), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n393), .A2(new_n398), .A3(new_n279), .A4(new_n395), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n397), .A2(G68), .A3(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n229), .B1(new_n217), .B2(new_n214), .ZN(new_n401));
  AOI22_X1  g0201(.A1(new_n401), .A2(G20), .B1(G159), .B2(new_n281), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n400), .A2(KEYINPUT16), .A3(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT16), .ZN(new_n404));
  AND2_X1   g0204(.A1(KEYINPUT3), .A2(G33), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n405), .A2(G20), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT81), .B(KEYINPUT3), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n406), .B(KEYINPUT7), .C1(new_n407), .C2(G33), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n398), .B1(new_n249), .B2(G20), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n217), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n228), .B1(new_n360), .B2(G58), .ZN(new_n411));
  INV_X1    g0211(.A(G159), .ZN(new_n412));
  INV_X1    g0212(.A(new_n281), .ZN(new_n413));
  OAI22_X1  g0213(.A1(new_n411), .A2(new_n279), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n404), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n403), .A2(new_n276), .A3(new_n415), .ZN(new_n416));
  INV_X1    g0216(.A(new_n277), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n417), .A2(new_n286), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n418), .B1(new_n273), .B2(new_n286), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n266), .A2(G232), .ZN(new_n421));
  NAND2_X1  g0221(.A1(G33), .A2(G87), .ZN(new_n422));
  XOR2_X1   g0222(.A(new_n422), .B(KEYINPUT82), .Z(new_n423));
  NOR2_X1   g0223(.A1(new_n250), .A2(G226), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n424), .B1(new_n393), .B2(new_n395), .ZN(new_n425));
  NOR2_X1   g0225(.A1(G223), .A2(G1698), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n423), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n265), .B(new_n421), .C1(new_n428), .C2(new_n256), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n429), .A2(G169), .ZN(new_n430));
  AOI211_X1 g0230(.A(new_n426), .B(new_n424), .C1(new_n393), .C2(new_n395), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n254), .B1(new_n431), .B2(new_n423), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n432), .A2(G179), .A3(new_n265), .A4(new_n421), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n420), .A2(new_n434), .ZN(new_n435));
  XOR2_X1   g0235(.A(KEYINPUT83), .B(KEYINPUT18), .Z(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  INV_X1    g0238(.A(new_n419), .ZN(new_n439));
  INV_X1    g0239(.A(new_n276), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n408), .A2(new_n409), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n360), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n402), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n440), .B1(new_n443), .B2(new_n404), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n439), .B1(new_n444), .B2(new_n403), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n429), .A2(G200), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n432), .A2(G190), .A3(new_n265), .A4(new_n421), .ZN(new_n447));
  NAND4_X1  g0247(.A1(new_n445), .A2(KEYINPUT17), .A3(new_n446), .A4(new_n447), .ZN(new_n448));
  NAND4_X1  g0248(.A1(new_n416), .A2(new_n446), .A3(new_n447), .A4(new_n419), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT17), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n420), .A2(new_n434), .A3(new_n436), .ZN(new_n452));
  NAND4_X1  g0252(.A1(new_n438), .A2(new_n448), .A3(new_n451), .A4(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n388), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n338), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n322), .A2(G200), .ZN(new_n456));
  INV_X1    g0256(.A(KEYINPUT73), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(G200), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n459), .B1(new_n340), .B2(new_n321), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT73), .B1(new_n460), .B2(new_n338), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n340), .A2(G190), .A3(new_n321), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n458), .A2(new_n461), .A3(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n454), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n272), .A2(G97), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n262), .A2(G33), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n440), .A2(new_n272), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT84), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n440), .A2(KEYINPUT84), .A3(new_n272), .A4(new_n467), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n470), .A2(G97), .A3(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n413), .A2(new_n210), .ZN(new_n473));
  INV_X1    g0273(.A(KEYINPUT6), .ZN(new_n474));
  INV_X1    g0274(.A(G97), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n318), .ZN(new_n476));
  NOR2_X1   g0276(.A1(G97), .A2(G107), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n474), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n318), .A2(KEYINPUT6), .A3(G97), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n279), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  AOI211_X1 g0280(.A(new_n473), .B(new_n480), .C1(G107), .C2(new_n441), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n466), .B(new_n472), .C1(new_n481), .C2(new_n440), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n258), .A2(G1), .ZN(new_n483));
  NOR2_X1   g0283(.A1(KEYINPUT5), .A2(G41), .ZN(new_n484));
  AND2_X1   g0284(.A1(KEYINPUT5), .A2(G41), .ZN(new_n485));
  OAI211_X1 g0285(.A(new_n483), .B(G274), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g0286(.A(new_n486), .B(KEYINPUT85), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT4), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n394), .B1(new_n407), .B2(G33), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n489), .B1(new_n490), .B2(new_n211), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n249), .A2(KEYINPUT4), .A3(G244), .A4(new_n250), .ZN(new_n492));
  NOR2_X1   g0292(.A1(new_n405), .A2(new_n394), .ZN(new_n493));
  OAI21_X1  g0293(.A(KEYINPUT4), .B1(new_n493), .B2(new_n220), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(G1698), .ZN(new_n495));
  NAND2_X1  g0295(.A1(G33), .A2(G283), .ZN(new_n496));
  NAND4_X1  g0296(.A1(new_n491), .A2(new_n492), .A3(new_n495), .A4(new_n496), .ZN(new_n497));
  AOI21_X1  g0297(.A(new_n488), .B1(new_n497), .B2(new_n254), .ZN(new_n498));
  OR2_X1    g0298(.A1(new_n485), .A2(new_n484), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n254), .B1(new_n499), .B2(new_n483), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G257), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n312), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n211), .B1(new_n393), .B2(new_n395), .ZN(new_n503));
  OAI21_X1  g0303(.A(new_n492), .B1(new_n503), .B2(KEYINPUT4), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n489), .B1(new_n249), .B2(G250), .ZN(new_n505));
  OAI21_X1  g0305(.A(new_n496), .B1(new_n505), .B2(new_n250), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n254), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n507), .A2(G179), .A3(new_n501), .A4(new_n487), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n482), .B1(new_n502), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT86), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT86), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n512), .B(new_n482), .C1(new_n502), .C2(new_n509), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(new_n482), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n507), .A2(new_n501), .A3(new_n487), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n516), .A2(G200), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n515), .B(new_n517), .C1(new_n269), .C2(new_n516), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT94), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n393), .A2(new_n395), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n220), .A2(new_n250), .ZN(new_n521));
  OR2_X1    g0321(.A1(new_n250), .A2(G257), .ZN(new_n522));
  AND3_X1   g0322(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(G294), .ZN(new_n524));
  NOR2_X1   g0324(.A1(new_n287), .A2(new_n524), .ZN(new_n525));
  OAI21_X1  g0325(.A(new_n519), .B1(new_n523), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n527));
  OAI211_X1 g0327(.A(new_n527), .B(KEYINPUT94), .C1(new_n287), .C2(new_n524), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n526), .A2(new_n254), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n500), .A2(G264), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n487), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G200), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(G190), .A3(new_n487), .A4(new_n530), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n470), .A2(G107), .A3(new_n471), .ZN(new_n534));
  OAI211_X1 g0334(.A(KEYINPUT92), .B(KEYINPUT25), .C1(new_n272), .C2(G107), .ZN(new_n535));
  XOR2_X1   g0335(.A(KEYINPUT92), .B(KEYINPUT25), .Z(new_n536));
  NAND3_X1  g0336(.A1(new_n536), .A2(new_n318), .A3(new_n273), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT93), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n534), .A2(KEYINPUT93), .A3(new_n535), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT91), .B1(new_n318), .B2(G20), .ZN(new_n543));
  XOR2_X1   g0343(.A(new_n543), .B(KEYINPUT23), .Z(new_n544));
  NAND2_X1  g0344(.A1(new_n288), .A2(G116), .ZN(new_n545));
  NOR2_X1   g0345(.A1(KEYINPUT22), .A2(G20), .ZN(new_n546));
  OAI211_X1 g0346(.A(G87), .B(new_n546), .C1(new_n405), .C2(new_n394), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT90), .ZN(new_n548));
  OR2_X1    g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n547), .A2(new_n548), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(new_n393), .B2(new_n395), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G87), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n544), .B(new_n545), .C1(new_n551), .C2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(KEYINPUT24), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI211_X1 g0357(.A(G20), .B(new_n219), .C1(new_n393), .C2(new_n395), .ZN(new_n558));
  OAI211_X1 g0358(.A(new_n550), .B(new_n549), .C1(new_n558), .C2(new_n552), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n559), .A2(KEYINPUT24), .A3(new_n544), .A4(new_n545), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n557), .A2(new_n276), .A3(new_n560), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n532), .A2(new_n533), .A3(new_n542), .A4(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n542), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n531), .A2(new_n312), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n529), .A2(new_n341), .A3(new_n487), .A4(new_n530), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(new_n566));
  NAND4_X1  g0366(.A1(new_n514), .A2(new_n518), .A3(new_n562), .A4(new_n566), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n500), .A2(G270), .ZN(new_n568));
  INV_X1    g0368(.A(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n520), .A2(G264), .A3(G1698), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n571));
  AOI21_X1  g0371(.A(G1698), .B1(new_n393), .B2(new_n395), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n572), .A2(G257), .B1(G303), .B2(new_n493), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT89), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n520), .A2(new_n574), .A3(G264), .A4(G1698), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n571), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  AOI211_X1 g0376(.A(new_n488), .B(new_n569), .C1(new_n576), .C2(new_n254), .ZN(new_n577));
  INV_X1    g0377(.A(G116), .ZN(new_n578));
  OR2_X1    g0378(.A1(new_n468), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n273), .A2(new_n578), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n496), .B(new_n279), .C1(G33), .C2(new_n475), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n581), .B(new_n276), .C1(new_n279), .C2(G116), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT20), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n582), .A2(new_n583), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n579), .B(new_n580), .C1(new_n584), .C2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(G169), .ZN(new_n587));
  OAI21_X1  g0387(.A(KEYINPUT21), .B1(new_n577), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n488), .B1(new_n576), .B2(new_n254), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n568), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT21), .ZN(new_n591));
  INV_X1    g0391(.A(new_n587), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n590), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(new_n586), .ZN(new_n594));
  NOR2_X1   g0394(.A1(new_n590), .A2(new_n594), .ZN(new_n595));
  AOI22_X1  g0395(.A1(new_n588), .A2(new_n593), .B1(new_n595), .B2(G179), .ZN(new_n596));
  NAND3_X1  g0396(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n279), .A2(new_n597), .B1(new_n477), .B2(new_n219), .ZN(new_n598));
  XNOR2_X1  g0398(.A(new_n598), .B(KEYINPUT87), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n553), .A2(G68), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT19), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n289), .B2(new_n475), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n599), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n324), .ZN(new_n604));
  AOI22_X1  g0404(.A1(new_n603), .A2(new_n276), .B1(new_n273), .B2(new_n604), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n470), .A2(new_n324), .A3(new_n471), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR3_X1    g0407(.A1(new_n258), .A2(G1), .A3(G274), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n256), .B(new_n608), .C1(G250), .C2(new_n483), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n393), .A2(new_n395), .B1(new_n211), .B2(G1698), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n216), .A2(new_n250), .ZN(new_n611));
  AOI22_X1  g0411(.A1(new_n610), .A2(new_n611), .B1(G33), .B2(G116), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n609), .B1(new_n612), .B2(new_n256), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n613), .A2(new_n312), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n607), .B(new_n614), .C1(G179), .C2(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n470), .A2(G87), .A3(new_n471), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n605), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(G200), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(KEYINPUT88), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  OR2_X1    g0420(.A1(new_n613), .A2(new_n269), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT88), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n605), .A2(new_n618), .A3(new_n622), .A4(new_n616), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n620), .A2(new_n621), .A3(new_n623), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n589), .A2(G190), .A3(new_n568), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n625), .B(new_n594), .C1(new_n459), .C2(new_n577), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n596), .A2(new_n615), .A3(new_n624), .A4(new_n626), .ZN(new_n627));
  NOR4_X1   g0427(.A1(new_n344), .A2(new_n464), .A3(new_n567), .A4(new_n627), .ZN(G372));
  NOR2_X1   g0428(.A1(new_n344), .A2(new_n464), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n517), .B1(new_n269), .B2(new_n516), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n630), .A2(new_n482), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n511), .B2(new_n513), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n588), .A2(new_n593), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n595), .A2(G179), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n566), .A2(new_n633), .A3(new_n634), .ZN(new_n635));
  NAND4_X1  g0435(.A1(new_n621), .A2(new_n605), .A3(new_n618), .A4(new_n616), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n615), .A2(new_n636), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n632), .A2(new_n635), .A3(new_n562), .A4(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n624), .A2(new_n615), .ZN(new_n639));
  OAI21_X1  g0439(.A(KEYINPUT26), .B1(new_n514), .B2(new_n639), .ZN(new_n640));
  AND3_X1   g0440(.A1(new_n507), .A2(new_n501), .A3(new_n487), .ZN(new_n641));
  OAI21_X1  g0441(.A(new_n508), .B1(new_n641), .B2(new_n312), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT95), .ZN(new_n643));
  XNOR2_X1  g0443(.A(new_n642), .B(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(KEYINPUT26), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n644), .A2(new_n637), .A3(new_n645), .A4(new_n482), .ZN(new_n646));
  NAND4_X1  g0446(.A1(new_n638), .A2(new_n615), .A3(new_n640), .A4(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n629), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g0448(.A(new_n449), .B(KEYINPUT17), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n343), .B1(new_n376), .B2(new_n379), .ZN(new_n650));
  INV_X1    g0450(.A(new_n387), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT18), .ZN(new_n653));
  AND3_X1   g0453(.A1(new_n420), .A2(new_n434), .A3(KEYINPUT96), .ZN(new_n654));
  AOI21_X1  g0454(.A(KEYINPUT96), .B1(new_n420), .B2(new_n434), .ZN(new_n655));
  OAI21_X1  g0455(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT96), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n435), .A2(new_n657), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n420), .A2(new_n434), .A3(KEYINPUT96), .ZN(new_n659));
  NAND3_X1  g0459(.A1(new_n658), .A2(KEYINPUT18), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n652), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n663), .A2(new_n310), .B1(new_n295), .B2(new_n313), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n648), .A2(new_n664), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT97), .Z(G369));
  NAND3_X1  g0466(.A1(new_n633), .A2(new_n634), .A3(new_n626), .ZN(new_n667));
  INV_X1    g0467(.A(G13), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n668), .A2(G20), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n669), .A2(new_n224), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  OR2_X1    g0471(.A1(new_n671), .A2(KEYINPUT98), .ZN(new_n672));
  INV_X1    g0472(.A(G213), .ZN(new_n673));
  AOI21_X1  g0473(.A(new_n673), .B1(new_n670), .B2(KEYINPUT27), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(KEYINPUT98), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n672), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(G343), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n679), .A2(new_n594), .ZN(new_n680));
  MUX2_X1   g0480(.A(new_n667), .B(new_n596), .S(new_n680), .Z(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT99), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n563), .A2(new_n678), .ZN(new_n683));
  AND2_X1   g0483(.A1(new_n562), .A2(new_n683), .ZN(new_n684));
  MUX2_X1   g0484(.A(new_n678), .B(new_n684), .S(new_n566), .Z(new_n685));
  NAND3_X1  g0485(.A1(new_n682), .A2(G330), .A3(new_n685), .ZN(new_n686));
  INV_X1    g0486(.A(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n596), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n688), .A2(new_n684), .A3(new_n566), .A4(new_n679), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n566), .B2(new_n678), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n687), .A2(new_n690), .ZN(G399));
  INV_X1    g0491(.A(new_n204), .ZN(new_n692));
  NOR2_X1   g0492(.A1(new_n692), .A2(G41), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NOR4_X1   g0494(.A1(G87), .A2(G97), .A3(G107), .A4(G116), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n694), .A2(G1), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n696), .B1(new_n230), .B2(new_n694), .ZN(new_n697));
  XNOR2_X1  g0497(.A(new_n697), .B(KEYINPUT28), .ZN(new_n698));
  AND2_X1   g0498(.A1(new_n644), .A2(new_n482), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n637), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(KEYINPUT26), .ZN(new_n701));
  OR3_X1    g0501(.A1(new_n514), .A2(new_n639), .A3(KEYINPUT26), .ZN(new_n702));
  NAND4_X1  g0502(.A1(new_n701), .A2(new_n615), .A3(new_n638), .A4(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(new_n679), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(KEYINPUT29), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n647), .A2(new_n679), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n705), .B1(KEYINPUT29), .B2(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  AND4_X1   g0508(.A1(new_n341), .A2(new_n590), .A3(new_n516), .A4(new_n531), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n529), .A2(new_n530), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n710), .A2(new_n613), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n711), .A2(new_n509), .A3(new_n577), .ZN(new_n712));
  INV_X1    g0512(.A(KEYINPUT30), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n613), .A2(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  INV_X1    g0514(.A(new_n714), .ZN(new_n715));
  AND2_X1   g0515(.A1(new_n715), .A2(KEYINPUT100), .ZN(new_n716));
  OR2_X1    g0516(.A1(new_n712), .A2(new_n713), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n717), .B1(new_n715), .B2(KEYINPUT100), .ZN(new_n718));
  OAI211_X1 g0518(.A(KEYINPUT31), .B(new_n678), .C1(new_n716), .C2(new_n718), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n679), .B1(new_n714), .B2(new_n717), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR3_X1   g0521(.A1(new_n567), .A2(new_n627), .A3(new_n678), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT31), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  AOI21_X1  g0524(.A(new_n708), .B1(new_n719), .B2(new_n724), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n707), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n698), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(G13), .A2(G33), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n682), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n249), .A2(G355), .A3(new_n204), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n244), .A2(new_n258), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n520), .A2(new_n692), .ZN(new_n735));
  OAI21_X1  g0535(.A(new_n735), .B1(G45), .B2(new_n230), .ZN(new_n736));
  OAI221_X1 g0536(.A(new_n733), .B1(G116), .B2(new_n204), .C1(new_n734), .C2(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n224), .B1(G20), .B2(new_n312), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n730), .A2(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n669), .A2(G45), .ZN(new_n741));
  NAND3_X1  g0541(.A1(new_n694), .A2(G1), .A3(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n279), .A2(new_n341), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n744), .A2(G190), .A3(new_n459), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n214), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n341), .A2(G200), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT101), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(G20), .A3(G190), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n750), .A2(G87), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n744), .A2(G200), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n752), .A2(new_n269), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(KEYINPUT102), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n755), .B1(new_n752), .B2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR3_X1   g0557(.A1(new_n752), .A2(new_n755), .A3(G190), .ZN(new_n758));
  OR2_X1    g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(G68), .ZN(new_n761));
  OAI221_X1 g0561(.A(new_n751), .B1(new_n208), .B2(new_n754), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n748), .A2(G20), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(G190), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NOR2_X1   g0565(.A1(G190), .A2(G200), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n766), .A2(G20), .A3(G179), .ZN(new_n767));
  OAI22_X1  g0567(.A1(new_n765), .A2(new_n318), .B1(new_n210), .B2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n269), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n279), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n766), .A2(G20), .A3(new_n341), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n412), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  OAI221_X1 g0573(.A(new_n249), .B1(new_n770), .B2(new_n475), .C1(new_n773), .C2(KEYINPUT32), .ZN(new_n774));
  OR4_X1    g0574(.A1(new_n746), .A2(new_n762), .A3(new_n768), .A4(new_n774), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(KEYINPUT32), .B2(new_n773), .ZN(new_n776));
  INV_X1    g0576(.A(G303), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n749), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(G322), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n493), .B1(new_n745), .B2(new_n779), .ZN(new_n780));
  XNOR2_X1  g0580(.A(KEYINPUT33), .B(G317), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n780), .B1(new_n759), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n764), .A2(G283), .ZN(new_n783));
  INV_X1    g0583(.A(new_n770), .ZN(new_n784));
  INV_X1    g0584(.A(new_n767), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n784), .A2(G294), .B1(G311), .B2(new_n785), .ZN(new_n786));
  XOR2_X1   g0586(.A(new_n771), .B(KEYINPUT103), .Z(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n788), .A2(G329), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n782), .A2(new_n783), .A3(new_n786), .A4(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n778), .B(new_n790), .C1(G326), .C2(new_n753), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n738), .B1(new_n776), .B2(new_n791), .ZN(new_n792));
  NAND4_X1  g0592(.A1(new_n732), .A2(new_n740), .A3(new_n743), .A4(new_n792), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n682), .A2(G330), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n682), .A2(G330), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n795), .A3(new_n742), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n793), .A2(new_n796), .ZN(G396));
  NOR2_X1   g0597(.A1(new_n725), .A2(KEYINPUT106), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n343), .A2(new_n678), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n463), .B1(new_n455), .B2(new_n679), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n799), .B1(new_n800), .B2(new_n343), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n706), .A2(new_n802), .ZN(new_n803));
  NAND3_X1  g0603(.A1(new_n647), .A2(new_n801), .A3(new_n679), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n798), .A2(new_n805), .ZN(new_n806));
  AOI22_X1  g0606(.A1(new_n725), .A2(KEYINPUT106), .B1(new_n803), .B2(new_n804), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n806), .B(new_n742), .C1(new_n807), .C2(new_n798), .ZN(new_n808));
  INV_X1    g0608(.A(new_n745), .ZN(new_n809));
  AOI22_X1  g0609(.A1(G137), .A2(new_n753), .B1(new_n809), .B2(G143), .ZN(new_n810));
  INV_X1    g0610(.A(G150), .ZN(new_n811));
  OAI221_X1 g0611(.A(new_n810), .B1(new_n412), .B2(new_n767), .C1(new_n760), .C2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  OAI22_X1  g0613(.A1(new_n813), .A2(KEYINPUT34), .B1(new_n761), .B2(new_n765), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n490), .B(new_n814), .C1(KEYINPUT34), .C2(new_n813), .ZN(new_n815));
  INV_X1    g0615(.A(G132), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n214), .B2(new_n770), .C1(new_n816), .C2(new_n787), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n749), .A2(new_n208), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n754), .A2(new_n777), .B1(new_n578), .B2(new_n767), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n819), .B1(new_n759), .B2(G283), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT104), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n764), .A2(G87), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n249), .B1(new_n750), .B2(G107), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT105), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n770), .A2(new_n475), .B1(new_n745), .B2(new_n524), .ZN(new_n825));
  AOI22_X1  g0625(.A1(new_n788), .A2(G311), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND4_X1  g0626(.A1(new_n821), .A2(new_n822), .A3(new_n823), .A4(new_n826), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n825), .A2(new_n824), .ZN(new_n828));
  OAI22_X1  g0628(.A1(new_n817), .A2(new_n818), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n738), .ZN(new_n830));
  NOR2_X1   g0630(.A1(new_n738), .A2(new_n728), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n831), .A2(new_n210), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n802), .A2(new_n728), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n830), .A2(new_n743), .A3(new_n832), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n808), .A2(new_n834), .ZN(G384));
  NOR2_X1   g0635(.A1(new_n387), .A2(new_n678), .ZN(new_n836));
  INV_X1    g0636(.A(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n676), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n403), .A2(new_n276), .ZN(new_n839));
  AOI21_X1  g0639(.A(KEYINPUT16), .B1(new_n400), .B2(new_n402), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n419), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g0641(.A1(new_n453), .A2(new_n838), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n420), .A2(new_n838), .ZN(new_n843));
  INV_X1    g0643(.A(KEYINPUT37), .ZN(new_n844));
  NAND4_X1  g0644(.A1(new_n435), .A2(new_n843), .A3(new_n844), .A4(new_n449), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n841), .B1(new_n434), .B2(new_n838), .ZN(new_n846));
  AND2_X1   g0646(.A1(new_n846), .A2(new_n449), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n845), .B1(new_n847), .B2(new_n844), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n842), .A2(new_n848), .A3(KEYINPUT38), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n656), .A2(new_n660), .A3(new_n649), .ZN(new_n851));
  INV_X1    g0651(.A(new_n843), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n658), .A2(new_n449), .A3(new_n659), .ZN(new_n854));
  INV_X1    g0654(.A(KEYINPUT109), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n852), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g0656(.A1(new_n658), .A2(KEYINPUT109), .A3(new_n449), .A4(new_n659), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n844), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n845), .B(KEYINPUT110), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n853), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT38), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n850), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT111), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT39), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n842), .A2(new_n848), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(new_n862), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n868), .A2(KEYINPUT108), .A3(new_n849), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT108), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n867), .A2(new_n870), .A3(new_n862), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n869), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n872), .A2(KEYINPUT111), .ZN(new_n873));
  AOI211_X1 g0673(.A(KEYINPUT39), .B(new_n850), .C1(new_n861), .C2(new_n862), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n866), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n875), .A2(KEYINPUT112), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n851), .A2(new_n852), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n854), .A2(new_n855), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n878), .A2(new_n843), .A3(new_n857), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n880), .B2(new_n859), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n865), .B(new_n849), .C1(new_n881), .C2(KEYINPUT38), .ZN(new_n882));
  NAND3_X1  g0682(.A1(new_n882), .A2(KEYINPUT111), .A3(new_n872), .ZN(new_n883));
  INV_X1    g0683(.A(KEYINPUT112), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n883), .A2(new_n884), .A3(new_n866), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n837), .B1(new_n876), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n799), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n804), .A2(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n386), .A2(new_n678), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n889), .B1(new_n380), .B2(new_n387), .ZN(new_n890));
  INV_X1    g0690(.A(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n380), .A2(new_n387), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n888), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n869), .A2(new_n871), .ZN(new_n895));
  OAI22_X1  g0695(.A1(new_n894), .A2(new_n895), .B1(new_n662), .B2(new_n838), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n886), .A2(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n707), .A2(new_n629), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n664), .ZN(new_n899));
  XNOR2_X1  g0699(.A(new_n897), .B(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n513), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n512), .B1(new_n642), .B2(new_n482), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n518), .B(new_n562), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n667), .A2(new_n639), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n904), .A2(new_n905), .A3(new_n566), .A4(new_n679), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n720), .B1(new_n906), .B2(KEYINPUT31), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n720), .A2(KEYINPUT31), .ZN(new_n908));
  INV_X1    g0708(.A(new_n908), .ZN(new_n909));
  OAI211_X1 g0709(.A(new_n801), .B(new_n893), .C1(new_n907), .C2(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(KEYINPUT40), .B1(new_n910), .B2(new_n863), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT40), .ZN(new_n912));
  AND3_X1   g0712(.A1(new_n869), .A2(new_n912), .A3(new_n871), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n802), .B1(new_n724), .B2(new_n908), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n913), .A2(new_n914), .A3(new_n893), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n911), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n724), .A2(new_n908), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n629), .A2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n916), .B(new_n918), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n919), .A2(G330), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n900), .B(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(new_n262), .B2(new_n669), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n231), .B1(new_n217), .B2(new_n214), .ZN(new_n923));
  OAI22_X1  g0723(.A1(new_n923), .A2(new_n210), .B1(G50), .B2(new_n761), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n924), .A2(G1), .A3(new_n668), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n478), .A2(new_n479), .ZN(new_n926));
  INV_X1    g0726(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g0727(.A(new_n578), .B1(new_n927), .B2(KEYINPUT35), .ZN(new_n928));
  OAI211_X1 g0728(.A(new_n928), .B(new_n227), .C1(KEYINPUT35), .C2(new_n927), .ZN(new_n929));
  XOR2_X1   g0729(.A(KEYINPUT107), .B(KEYINPUT36), .Z(new_n930));
  XNOR2_X1  g0730(.A(new_n929), .B(new_n930), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n922), .A2(new_n925), .A3(new_n931), .ZN(G367));
  NAND2_X1  g0732(.A1(new_n699), .A2(new_n678), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n632), .B1(new_n515), .B2(new_n679), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n514), .B1(new_n935), .B2(new_n566), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n679), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n689), .A2(new_n934), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT42), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n937), .A2(KEYINPUT43), .A3(new_n939), .ZN(new_n940));
  INV_X1    g0740(.A(new_n637), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n617), .A2(new_n678), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT113), .ZN(new_n943));
  MUX2_X1   g0743(.A(new_n941), .B(new_n615), .S(new_n943), .Z(new_n944));
  AND2_X1   g0744(.A1(new_n940), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n937), .A2(new_n939), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT43), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OR2_X1    g0748(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n945), .A2(new_n948), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n686), .A2(KEYINPUT114), .A3(new_n935), .ZN(new_n952));
  OAI21_X1  g0752(.A(KEYINPUT114), .B1(new_n686), .B2(new_n935), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT115), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g0756(.A1(new_n952), .A2(KEYINPUT115), .A3(new_n953), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n949), .B(new_n950), .C1(new_n957), .C2(new_n954), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n693), .B(KEYINPUT41), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n935), .A2(new_n690), .ZN(new_n961));
  XNOR2_X1  g0761(.A(new_n961), .B(KEYINPUT45), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n935), .A2(new_n690), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n962), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n966), .A2(KEYINPUT116), .A3(new_n687), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n685), .B1(new_n688), .B2(new_n679), .ZN(new_n968));
  INV_X1    g0768(.A(new_n689), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n795), .B(new_n970), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n687), .A2(KEYINPUT116), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n972), .A2(new_n962), .A3(new_n965), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n967), .A2(new_n726), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n960), .B1(new_n974), .B2(new_n726), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n741), .A2(G1), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n956), .B(new_n958), .C1(new_n975), .C2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n764), .A2(G77), .ZN(new_n978));
  OAI221_X1 g0778(.A(new_n978), .B1(new_n208), .B2(new_n767), .C1(new_n214), .C2(new_n749), .ZN(new_n979));
  INV_X1    g0779(.A(G137), .ZN(new_n980));
  OAI221_X1 g0780(.A(new_n249), .B1(new_n980), .B2(new_n771), .C1(new_n760), .C2(new_n412), .ZN(new_n981));
  AOI211_X1 g0781(.A(new_n979), .B(new_n981), .C1(G143), .C2(new_n753), .ZN(new_n982));
  OAI221_X1 g0782(.A(new_n982), .B1(new_n761), .B2(new_n770), .C1(new_n811), .C2(new_n745), .ZN(new_n983));
  XOR2_X1   g0783(.A(KEYINPUT117), .B(G317), .Z(new_n984));
  OAI22_X1  g0784(.A1(new_n765), .A2(new_n475), .B1(new_n771), .B2(new_n984), .ZN(new_n985));
  INV_X1    g0785(.A(G311), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n490), .B1(new_n754), .B2(new_n986), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n770), .A2(new_n318), .B1(new_n745), .B2(new_n777), .ZN(new_n988));
  NOR3_X1   g0788(.A1(new_n985), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(G283), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n989), .B1(new_n990), .B2(new_n767), .C1(new_n524), .C2(new_n760), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n749), .A2(new_n578), .ZN(new_n992));
  XNOR2_X1  g0792(.A(new_n992), .B(KEYINPUT46), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n983), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  XNOR2_X1  g0794(.A(new_n994), .B(KEYINPUT47), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n738), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n944), .A2(new_n730), .ZN(new_n997));
  INV_X1    g0797(.A(new_n735), .ZN(new_n998));
  OAI221_X1 g0798(.A(new_n739), .B1(new_n204), .B2(new_n604), .C1(new_n235), .C2(new_n998), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n996), .A2(new_n743), .A3(new_n997), .A4(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n977), .A2(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n971), .A2(new_n976), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n1002), .B(KEYINPUT118), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n760), .A2(new_n286), .B1(new_n761), .B2(new_n767), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT119), .B(G150), .Z(new_n1005));
  OAI22_X1  g0805(.A1(new_n765), .A2(new_n475), .B1(new_n771), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n749), .A2(new_n210), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1006), .A2(new_n490), .A3(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g0808(.A(new_n1008), .B(KEYINPUT120), .ZN(new_n1009));
  AOI211_X1 g0809(.A(new_n1004), .B(new_n1009), .C1(new_n324), .C2(new_n784), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n208), .B2(new_n745), .C1(new_n412), .C2(new_n754), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n759), .A2(G311), .B1(G303), .B2(new_n785), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n779), .B2(new_n754), .C1(new_n745), .C2(new_n984), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n1014), .B1(new_n990), .B2(new_n770), .C1(new_n524), .C2(new_n749), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT49), .ZN(new_n1016));
  OR2_X1    g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n764), .A2(G116), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n771), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1019), .A2(G326), .ZN(new_n1020));
  NAND4_X1  g0820(.A1(new_n1017), .A2(new_n490), .A3(new_n1018), .A4(new_n1020), .ZN(new_n1021));
  AND2_X1   g0821(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1011), .B1(new_n1021), .B2(new_n1022), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n240), .A2(G45), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n249), .A2(new_n204), .ZN(new_n1025));
  OAI22_X1  g0825(.A1(new_n1024), .A2(new_n998), .B1(new_n695), .B2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n285), .A2(new_n208), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT50), .Z(new_n1028));
  NAND2_X1  g0828(.A1(G68), .A2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1028), .A2(new_n258), .A3(new_n1029), .A4(new_n695), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1026), .A2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n692), .A2(new_n318), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n1023), .A2(new_n738), .B1(new_n739), .B2(new_n1033), .ZN(new_n1034));
  OAI211_X1 g0834(.A(new_n1034), .B(new_n743), .C1(new_n685), .C2(new_n731), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n726), .A2(new_n971), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n726), .A2(new_n971), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1037), .A2(new_n693), .ZN(new_n1038));
  OAI211_X1 g0838(.A(new_n1003), .B(new_n1035), .C1(new_n1036), .C2(new_n1038), .ZN(G393));
  AOI21_X1  g0839(.A(new_n742), .B1(new_n935), .B2(new_n730), .ZN(new_n1040));
  OAI221_X1 g0840(.A(new_n739), .B1(new_n475), .B2(new_n204), .C1(new_n998), .C2(new_n247), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G150), .A2(new_n753), .B1(new_n809), .B2(G159), .ZN(new_n1042));
  NOR2_X1   g0842(.A1(new_n1042), .A2(KEYINPUT51), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(G77), .B2(new_n784), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n750), .A2(new_n360), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n490), .B1(G143), .B2(new_n1019), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1044), .A2(new_n822), .A3(new_n1045), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n759), .A2(G50), .B1(new_n285), .B2(new_n785), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT121), .Z(new_n1049));
  AOI211_X1 g0849(.A(new_n1047), .B(new_n1049), .C1(KEYINPUT51), .C2(new_n1042), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G107), .A2(new_n764), .B1(new_n750), .B2(G283), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n249), .B1(new_n785), .B2(G294), .ZN(new_n1052));
  OAI211_X1 g0852(.A(new_n1051), .B(new_n1052), .C1(new_n779), .C2(new_n771), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT52), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n753), .A2(G317), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1055), .B1(new_n986), .B2(new_n745), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n760), .A2(new_n777), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AND2_X1   g0857(.A1(new_n1056), .A2(new_n1054), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n770), .A2(new_n578), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1053), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n738), .B1(new_n1050), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1040), .A2(new_n1041), .A3(new_n1061), .ZN(new_n1062));
  XNOR2_X1  g0862(.A(new_n966), .B(new_n687), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n976), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n1062), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  AND3_X1   g0865(.A1(new_n726), .A2(new_n973), .A3(new_n971), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1037), .A2(new_n1063), .B1(new_n1066), .B2(new_n967), .ZN(new_n1067));
  AOI21_X1  g0867(.A(new_n1065), .B1(new_n1067), .B2(new_n693), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1068), .ZN(G390));
  AOI21_X1  g0869(.A(KEYINPUT122), .B1(new_n894), .B2(new_n837), .ZN(new_n1070));
  AND3_X1   g0870(.A1(new_n380), .A2(new_n387), .A3(new_n889), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n890), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1072), .B1(new_n804), .B2(new_n887), .ZN(new_n1073));
  INV_X1    g0873(.A(KEYINPUT122), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1073), .A2(new_n1074), .A3(new_n836), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1070), .A2(new_n1075), .ZN(new_n1076));
  NAND3_X1  g0876(.A1(new_n1076), .A2(new_n876), .A3(new_n885), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n800), .A2(new_n343), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n703), .A2(new_n679), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n887), .ZN(new_n1080));
  AOI211_X1 g0880(.A(new_n863), .B(new_n836), .C1(new_n1080), .C2(new_n893), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n725), .A2(new_n801), .A3(new_n893), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  AND3_X1   g0884(.A1(new_n1077), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n910), .A2(new_n708), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n1077), .B2(new_n1082), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n976), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n883), .A2(new_n884), .A3(new_n866), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n884), .B1(new_n883), .B2(new_n866), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1091), .A2(new_n728), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n286), .A2(new_n831), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n249), .B1(new_n767), .B2(new_n1094), .C1(new_n760), .C2(new_n980), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1095), .B1(G125), .B2(new_n788), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n784), .A2(G159), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n749), .A2(new_n1005), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT53), .ZN(new_n1099));
  AOI22_X1  g0899(.A1(new_n764), .A2(G50), .B1(G128), .B2(new_n753), .ZN(new_n1100));
  NAND4_X1  g0900(.A1(new_n1096), .A2(new_n1097), .A3(new_n1099), .A4(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1101), .B1(G132), .B2(new_n809), .ZN(new_n1102));
  AOI22_X1  g0902(.A1(new_n788), .A2(G294), .B1(new_n750), .B2(G87), .ZN(new_n1103));
  OAI221_X1 g0903(.A(new_n1103), .B1(new_n761), .B2(new_n765), .C1(new_n210), .C2(new_n770), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n493), .B1(new_n475), .B2(new_n767), .C1(new_n760), .C2(new_n318), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n754), .A2(new_n990), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n745), .A2(new_n578), .ZN(new_n1107));
  NOR4_X1   g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1106), .A4(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n738), .B1(new_n1102), .B2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1092), .A2(new_n743), .A3(new_n1093), .A4(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1088), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1086), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n894), .A2(KEYINPUT122), .A3(new_n837), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n1074), .B1(new_n1073), .B2(new_n836), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  NOR3_X1   g0915(.A1(new_n1089), .A2(new_n1115), .A3(new_n1090), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1112), .B1(new_n1116), .B2(new_n1081), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1077), .A2(new_n1082), .A3(new_n1084), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n629), .A2(new_n917), .A3(G330), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n898), .A2(new_n664), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1080), .ZN(new_n1122));
  AND2_X1   g0922(.A1(new_n914), .A2(G330), .ZN(new_n1123));
  OAI211_X1 g0923(.A(new_n1122), .B(new_n1083), .C1(new_n1123), .C2(new_n893), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n893), .B1(new_n725), .B2(new_n801), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n888), .B1(new_n1125), .B2(new_n1086), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1121), .A2(new_n1127), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1117), .A2(new_n1118), .A3(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n1081), .B1(new_n1091), .B2(new_n1076), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1130), .B2(new_n1086), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1127), .ZN(new_n1132));
  NOR2_X1   g0932(.A1(new_n1132), .A2(new_n1120), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n694), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1111), .B1(new_n1129), .B2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1135), .ZN(G378));
  NAND3_X1  g0936(.A1(new_n303), .A2(new_n309), .A3(new_n314), .ZN(new_n1137));
  XOR2_X1   g0937(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1138));
  XNOR2_X1  g0938(.A(new_n1137), .B(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n295), .A2(new_n838), .ZN(new_n1140));
  XNOR2_X1  g0940(.A(new_n1139), .B(new_n1140), .ZN(new_n1141));
  AND3_X1   g0941(.A1(new_n916), .A2(G330), .A3(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1141), .B1(new_n916), .B2(G330), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n886), .A2(new_n896), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n836), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1141), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n849), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n914), .A2(new_n1147), .A3(new_n893), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n910), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1148), .A2(KEYINPUT40), .B1(new_n1149), .B2(new_n913), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1146), .B1(new_n1150), .B2(new_n708), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n896), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n916), .A2(new_n1141), .A3(G330), .ZN(new_n1153));
  NAND4_X1  g0953(.A1(new_n1145), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n831), .A2(new_n208), .ZN(new_n1157));
  NOR2_X1   g0957(.A1(new_n1146), .A2(new_n729), .ZN(new_n1158));
  INV_X1    g0958(.A(G124), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n287), .B1(new_n771), .B2(new_n1159), .ZN(new_n1160));
  OAI22_X1  g0960(.A1(new_n749), .A2(new_n1094), .B1(new_n811), .B2(new_n770), .ZN(new_n1161));
  NOR2_X1   g0961(.A1(new_n760), .A2(new_n816), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(G125), .C2(new_n753), .ZN(new_n1163));
  INV_X1    g0963(.A(G128), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1163), .B1(new_n1164), .B2(new_n745), .C1(new_n980), .C2(new_n767), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G41), .B(new_n1160), .C1(new_n1165), .C2(KEYINPUT59), .ZN(new_n1166));
  OAI221_X1 g0966(.A(new_n1166), .B1(KEYINPUT59), .B2(new_n1165), .C1(new_n412), .C2(new_n765), .ZN(new_n1167));
  OAI22_X1  g0967(.A1(new_n770), .A2(new_n761), .B1(new_n745), .B2(new_n318), .ZN(new_n1168));
  AOI211_X1 g0968(.A(new_n394), .B(new_n1007), .C1(G283), .C2(new_n788), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n604), .B2(new_n767), .ZN(new_n1170));
  AOI211_X1 g0970(.A(new_n1168), .B(new_n1170), .C1(G116), .C2(new_n753), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n393), .A2(new_n257), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n764), .B2(G58), .ZN(new_n1173));
  OAI211_X1 g0973(.A(new_n1171), .B(new_n1173), .C1(new_n475), .C2(new_n760), .ZN(new_n1174));
  XNOR2_X1  g0974(.A(new_n1174), .B(KEYINPUT58), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1172), .A2(new_n208), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1167), .A2(new_n1175), .A3(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g0977(.A(new_n1177), .B(KEYINPUT123), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n742), .B(new_n1158), .C1(new_n738), .C2(new_n1178), .ZN(new_n1179));
  AOI22_X1  g0979(.A1(new_n1156), .A2(new_n976), .B1(new_n1157), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g0980(.A(new_n1133), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(new_n1121), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1182), .B2(new_n1156), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1120), .B1(new_n1131), .B2(new_n1133), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n1144), .A2(new_n1154), .A3(KEYINPUT57), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n693), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1180), .B1(new_n1183), .B2(new_n1186), .ZN(G375));
  NAND2_X1  g0987(.A1(new_n1132), .A2(new_n1120), .ZN(new_n1188));
  NAND3_X1  g0988(.A1(new_n1188), .A2(new_n1128), .A3(new_n959), .ZN(new_n1189));
  AOI22_X1  g0989(.A1(new_n759), .A2(G116), .B1(G107), .B2(new_n785), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1190), .A2(KEYINPUT124), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n524), .B2(new_n754), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n749), .A2(new_n475), .ZN(new_n1193));
  NOR2_X1   g0993(.A1(new_n1190), .A2(KEYINPUT124), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n788), .A2(G303), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n324), .A2(new_n784), .B1(new_n809), .B2(G283), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1195), .A2(new_n978), .A3(new_n493), .A4(new_n1196), .ZN(new_n1197));
  NOR4_X1   g0997(.A1(new_n1192), .A2(new_n1193), .A3(new_n1194), .A4(new_n1197), .ZN(new_n1198));
  AOI22_X1  g0998(.A1(new_n764), .A2(G58), .B1(G137), .B2(new_n809), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(new_n208), .B2(new_n770), .C1(new_n412), .C2(new_n749), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n520), .B1(new_n816), .B2(new_n754), .C1(new_n760), .C2(new_n1094), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n787), .A2(new_n1164), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n767), .A2(new_n811), .ZN(new_n1203));
  NOR4_X1   g1003(.A1(new_n1200), .A2(new_n1201), .A3(new_n1202), .A4(new_n1203), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n738), .B1(new_n1198), .B2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n743), .B(new_n1205), .C1(new_n893), .C2(new_n729), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1206), .B1(new_n761), .B2(new_n831), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n1207), .B1(new_n1127), .B2(new_n976), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1189), .A2(new_n1208), .ZN(G381));
  NOR2_X1   g1009(.A1(G375), .A2(G378), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(G381), .A2(G384), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1068), .A2(new_n977), .A3(new_n1000), .ZN(new_n1212));
  NOR3_X1   g1012(.A1(new_n1212), .A2(G396), .A3(G393), .ZN(new_n1213));
  NAND3_X1  g1013(.A1(new_n1210), .A2(new_n1211), .A3(new_n1213), .ZN(G407));
  AOI21_X1  g1014(.A(new_n673), .B1(new_n1210), .B2(new_n677), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(G407), .ZN(G409));
  NOR2_X1   g1016(.A1(new_n673), .A2(G343), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(G2897), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  INV_X1    g1019(.A(KEYINPUT60), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1188), .A2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1132), .A2(KEYINPUT60), .A3(new_n1120), .ZN(new_n1222));
  NAND4_X1  g1022(.A1(new_n1221), .A2(new_n693), .A3(new_n1128), .A4(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(KEYINPUT125), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n808), .A2(new_n1224), .A3(new_n834), .ZN(new_n1225));
  INV_X1    g1025(.A(new_n1225), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1223), .A2(new_n1208), .A3(new_n1226), .ZN(new_n1227));
  AND2_X1   g1027(.A1(new_n1223), .A2(new_n1208), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(G384), .A2(KEYINPUT125), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1225), .ZN(new_n1230));
  OAI211_X1 g1030(.A(new_n1219), .B(new_n1227), .C1(new_n1228), .C2(new_n1230), .ZN(new_n1231));
  AND3_X1   g1031(.A1(new_n1223), .A2(new_n1208), .A3(new_n1226), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1230), .B1(new_n1223), .B2(new_n1208), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1218), .B1(new_n1232), .B2(new_n1233), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1217), .B1(G375), .B2(G378), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1128), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1237));
  OAI211_X1 g1037(.A(new_n1156), .B(new_n959), .C1(new_n1237), .C2(new_n1120), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1135), .A2(new_n1180), .A3(new_n1238), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1235), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  AND3_X1   g1040(.A1(new_n1144), .A2(new_n1154), .A3(KEYINPUT57), .ZN(new_n1241));
  OAI21_X1  g1041(.A(new_n1241), .B1(new_n1237), .B2(new_n1120), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1155), .B1(new_n1181), .B2(new_n1121), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1242), .B(new_n693), .C1(new_n1243), .C2(KEYINPUT57), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1135), .B1(new_n1244), .B2(new_n1180), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n1111), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1134), .A2(new_n1129), .ZN(new_n1247));
  AND4_X1   g1047(.A1(new_n1246), .A2(new_n1247), .A3(new_n1238), .A4(new_n1180), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n1232), .A2(new_n1233), .ZN(new_n1249));
  NOR4_X1   g1049(.A1(new_n1245), .A2(new_n1248), .A3(new_n1217), .A4(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT63), .B1(new_n1240), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1217), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1179), .A2(new_n1157), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1254), .B1(new_n1155), .B2(new_n1064), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n694), .B1(new_n1182), .B2(new_n1241), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT57), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1257), .B1(new_n1184), .B2(new_n1155), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1255), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1253), .B(new_n1239), .C1(new_n1259), .C2(new_n1135), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n1252), .B1(new_n1260), .B2(new_n1249), .ZN(new_n1261));
  XNOR2_X1  g1061(.A(G393), .B(G396), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1212), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1068), .B1(new_n977), .B2(new_n1000), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1263), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT61), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(G390), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1268), .A2(new_n1212), .A3(new_n1262), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1266), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT126), .ZN(new_n1271));
  XNOR2_X1  g1071(.A(new_n1270), .B(new_n1271), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1251), .A2(new_n1261), .A3(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(KEYINPUT62), .B1(new_n1260), .B2(new_n1249), .ZN(new_n1274));
  XOR2_X1   g1074(.A(KEYINPUT127), .B(KEYINPUT61), .Z(new_n1275));
  AND2_X1   g1075(.A1(new_n1231), .A2(new_n1234), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1260), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT62), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1249), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1236), .A2(new_n1278), .A3(new_n1239), .A4(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1274), .A2(new_n1277), .A3(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1266), .A2(new_n1269), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1273), .A2(new_n1283), .ZN(G405));
  XNOR2_X1  g1084(.A(new_n1282), .B(new_n1279), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1210), .A2(new_n1245), .ZN(new_n1286));
  XNOR2_X1  g1086(.A(new_n1285), .B(new_n1286), .ZN(G402));
endmodule


