//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n223, new_n224,
    new_n225, new_n226, new_n227, new_n228, new_n229, new_n230, new_n232,
    new_n233, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1245, new_n1246, new_n1247, new_n1248,
    new_n1250, new_n1251, new_n1252, new_n1253, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  AOI22_X1  g0003(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n204));
  AOI22_X1  g0004(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n207));
  AOI22_X1  g0007(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g0009(.A(new_n203), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT1), .ZN(new_n211));
  OR3_X1    g0011(.A1(new_n203), .A2(KEYINPUT64), .A3(G13), .ZN(new_n212));
  OAI21_X1  g0012(.A(KEYINPUT64), .B1(new_n203), .B2(G13), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  OAI211_X1 g0014(.A(new_n214), .B(G250), .C1(G257), .C2(G264), .ZN(new_n215));
  XOR2_X1   g0015(.A(new_n215), .B(KEYINPUT0), .Z(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(G50), .B1(G58), .B2(G68), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  AOI211_X1 g0021(.A(new_n211), .B(new_n216), .C1(new_n219), .C2(new_n221), .ZN(G361));
  XNOR2_X1  g0022(.A(G238), .B(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G232), .ZN(new_n224));
  XNOR2_X1  g0024(.A(new_n223), .B(new_n224), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT2), .B(G226), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n225), .B(new_n226), .ZN(new_n227));
  XNOR2_X1  g0027(.A(G250), .B(G257), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G264), .B(G270), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n227), .B(new_n230), .ZN(G358));
  XOR2_X1   g0031(.A(G87), .B(G97), .Z(new_n232));
  XOR2_X1   g0032(.A(G107), .B(G116), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(G50), .ZN(new_n235));
  NAND2_X1  g0035(.A1(new_n235), .A2(G68), .ZN(new_n236));
  INV_X1    g0036(.A(G68), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n237), .A2(G50), .ZN(new_n238));
  NAND2_X1  g0038(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n234), .B(new_n241), .Z(G351));
  INV_X1    g0042(.A(G13), .ZN(new_n243));
  NOR3_X1   g0043(.A1(new_n243), .A2(new_n218), .A3(G1), .ZN(new_n244));
  NAND3_X1  g0044(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(new_n217), .ZN(new_n246));
  NOR2_X1   g0046(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  INV_X1    g0048(.A(G58), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n249), .A2(KEYINPUT8), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT8), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(new_n244), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n248), .A2(new_n256), .B1(new_n257), .B2(new_n253), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT73), .ZN(new_n259));
  INV_X1    g0059(.A(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n260), .A2(KEYINPUT72), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT72), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n262), .A2(G33), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n265));
  NOR2_X1   g0065(.A1(KEYINPUT3), .A2(G33), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n259), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT3), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n269), .B1(new_n261), .B2(new_n263), .ZN(new_n270));
  NOR3_X1   g0070(.A1(new_n270), .A2(KEYINPUT73), .A3(new_n266), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n218), .B1(new_n268), .B2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT74), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT7), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  OAI21_X1  g0075(.A(KEYINPUT73), .B1(new_n270), .B2(new_n266), .ZN(new_n276));
  XNOR2_X1  g0076(.A(KEYINPUT72), .B(G33), .ZN(new_n277));
  OAI211_X1 g0077(.A(new_n259), .B(new_n267), .C1(new_n277), .C2(new_n269), .ZN(new_n278));
  AOI21_X1  g0078(.A(G20), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(KEYINPUT74), .B1(new_n279), .B2(KEYINPUT7), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n267), .B1(new_n277), .B2(new_n269), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(KEYINPUT7), .A3(new_n218), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n275), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n284), .A2(G68), .ZN(new_n285));
  XNOR2_X1  g0085(.A(G58), .B(G68), .ZN(new_n286));
  NOR2_X1   g0086(.A1(G20), .A2(G33), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n286), .A2(G20), .B1(G159), .B2(new_n287), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n285), .A2(KEYINPUT16), .A3(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n246), .ZN(new_n290));
  AND2_X1   g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NOR3_X1   g0091(.A1(new_n291), .A2(new_n274), .A3(G20), .ZN(new_n292));
  OAI21_X1  g0092(.A(new_n292), .B1(new_n264), .B2(KEYINPUT3), .ZN(new_n293));
  XNOR2_X1  g0093(.A(KEYINPUT3), .B(G33), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n274), .B1(new_n294), .B2(G20), .ZN(new_n295));
  AND2_X1   g0095(.A1(new_n293), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n288), .B1(new_n296), .B2(new_n237), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT16), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n290), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n258), .B1(new_n289), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(KEYINPUT78), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(KEYINPUT17), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(G41), .ZN(new_n304));
  OAI211_X1 g0104(.A(G1), .B(G13), .C1(new_n260), .C2(new_n304), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n254), .B1(G41), .B2(G45), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n308), .A2(KEYINPUT75), .A3(G232), .ZN(new_n309));
  INV_X1    g0109(.A(KEYINPUT75), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n310), .B1(new_n307), .B2(new_n224), .ZN(new_n311));
  INV_X1    g0111(.A(G45), .ZN(new_n312));
  AOI21_X1  g0112(.A(G1), .B1(new_n304), .B2(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n305), .A2(G274), .A3(new_n313), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n309), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT76), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT76), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n309), .A2(new_n311), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  INV_X1    g0118(.A(G226), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(G1698), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n320), .B1(G223), .B2(G1698), .ZN(new_n321));
  INV_X1    g0121(.A(G87), .ZN(new_n322));
  OAI22_X1  g0122(.A1(new_n282), .A2(new_n321), .B1(new_n260), .B2(new_n322), .ZN(new_n323));
  AOI21_X1  g0123(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g0125(.A1(new_n316), .A2(new_n318), .A3(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(G200), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n328), .B1(G190), .B2(new_n326), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n301), .A2(KEYINPUT17), .ZN(new_n330));
  NAND4_X1  g0130(.A1(new_n300), .A2(new_n303), .A3(new_n329), .A4(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n258), .ZN(new_n332));
  INV_X1    g0132(.A(new_n288), .ZN(new_n333));
  AOI211_X1 g0133(.A(new_n298), .B(new_n333), .C1(new_n284), .C2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(new_n299), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n329), .B(new_n332), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n336), .A2(new_n302), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n331), .A2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(G244), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n314), .B1(new_n307), .B2(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G1698), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n294), .A2(G232), .A3(new_n341), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n294), .A2(G238), .A3(G1698), .ZN(new_n343));
  INV_X1    g0143(.A(G107), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n342), .B(new_n343), .C1(new_n344), .C2(new_n294), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n340), .B1(new_n345), .B2(new_n324), .ZN(new_n346));
  INV_X1    g0146(.A(G179), .ZN(new_n347));
  AOI21_X1  g0147(.A(KEYINPUT67), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(KEYINPUT67), .A3(new_n347), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n247), .A2(G77), .A3(new_n255), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n352), .B1(G77), .B2(new_n257), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n253), .A2(new_n287), .B1(G20), .B2(G77), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n218), .A2(G33), .ZN(new_n355));
  XNOR2_X1  g0155(.A(KEYINPUT15), .B(G87), .ZN(new_n356));
  OAI21_X1  g0156(.A(new_n354), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n353), .B1(new_n357), .B2(new_n246), .ZN(new_n358));
  INV_X1    g0158(.A(new_n346), .ZN(new_n359));
  INV_X1    g0159(.A(G169), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n358), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n351), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n346), .A2(G190), .ZN(new_n363));
  XOR2_X1   g0163(.A(KEYINPUT66), .B(G200), .Z(new_n364));
  OAI211_X1 g0164(.A(new_n358), .B(new_n363), .C1(new_n364), .C2(new_n346), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n362), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n294), .A2(G232), .A3(G1698), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n294), .A2(G226), .A3(new_n341), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G33), .A2(G97), .ZN(new_n369));
  NAND3_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n370), .A2(new_n324), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n305), .A2(G238), .A3(new_n306), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT70), .ZN(new_n373));
  AND3_X1   g0173(.A1(new_n314), .A2(new_n372), .A3(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n373), .B1(new_n314), .B2(new_n372), .ZN(new_n375));
  OAI21_X1  g0175(.A(new_n371), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(KEYINPUT13), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT13), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n371), .B(new_n378), .C1(new_n374), .C2(new_n375), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n377), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(G169), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n381), .A2(KEYINPUT14), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n377), .A2(G179), .A3(new_n379), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n380), .A2(new_n384), .A3(G169), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n287), .A2(G50), .B1(G20), .B2(new_n237), .ZN(new_n387));
  INV_X1    g0187(.A(G77), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n355), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n389), .A2(new_n246), .ZN(new_n390));
  OR2_X1    g0190(.A1(new_n390), .A2(KEYINPUT11), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n244), .A2(new_n237), .ZN(new_n392));
  XNOR2_X1  g0192(.A(new_n392), .B(KEYINPUT12), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(KEYINPUT11), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n247), .A2(G68), .A3(new_n255), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n391), .A2(new_n393), .A3(new_n394), .A4(new_n395), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n366), .B1(new_n386), .B2(new_n396), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n294), .A2(G222), .A3(new_n341), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n294), .A2(G223), .A3(G1698), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n398), .B(new_n399), .C1(new_n388), .C2(new_n294), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n400), .A2(new_n324), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n314), .B1(new_n307), .B2(new_n319), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(G190), .A3(new_n403), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n402), .B1(new_n400), .B2(new_n324), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n404), .B1(new_n364), .B2(new_n405), .ZN(new_n406));
  XNOR2_X1  g0206(.A(KEYINPUT8), .B(G58), .ZN(new_n407));
  INV_X1    g0207(.A(G150), .ZN(new_n408));
  INV_X1    g0208(.A(new_n287), .ZN(new_n409));
  OAI22_X1  g0209(.A1(new_n407), .A2(new_n355), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(G58), .A2(G68), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n218), .B1(new_n411), .B2(new_n235), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n246), .B1(new_n410), .B2(new_n412), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n235), .B1(new_n254), .B2(G20), .ZN(new_n414));
  AOI22_X1  g0214(.A1(new_n247), .A2(new_n414), .B1(new_n235), .B2(new_n244), .ZN(new_n415));
  AND3_X1   g0215(.A1(new_n413), .A2(KEYINPUT68), .A3(new_n415), .ZN(new_n416));
  AOI21_X1  g0216(.A(KEYINPUT68), .B1(new_n413), .B2(new_n415), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n406), .B1(KEYINPUT9), .B2(new_n418), .ZN(new_n419));
  OR2_X1    g0219(.A1(new_n416), .A2(new_n417), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT9), .ZN(new_n421));
  AOI21_X1  g0221(.A(KEYINPUT69), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT69), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n418), .A2(new_n423), .A3(KEYINPUT9), .ZN(new_n424));
  OAI21_X1  g0224(.A(new_n419), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT10), .ZN(new_n426));
  INV_X1    g0226(.A(KEYINPUT10), .ZN(new_n427));
  OAI211_X1 g0227(.A(new_n419), .B(new_n427), .C1(new_n422), .C2(new_n424), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n413), .A2(new_n415), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n430), .B1(new_n405), .B2(G169), .ZN(new_n431));
  AOI21_X1  g0231(.A(new_n431), .B1(new_n347), .B2(new_n405), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n380), .A2(G200), .ZN(new_n434));
  INV_X1    g0234(.A(new_n396), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n377), .A2(G190), .A3(new_n379), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT71), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(KEYINPUT71), .A3(new_n435), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n397), .A2(new_n429), .A3(new_n433), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n326), .A2(G169), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(new_n347), .B2(new_n326), .ZN(new_n444));
  INV_X1    g0244(.A(new_n444), .ZN(new_n445));
  NOR3_X1   g0245(.A1(new_n300), .A2(new_n445), .A3(KEYINPUT18), .ZN(new_n446));
  INV_X1    g0246(.A(KEYINPUT18), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n447), .B1(new_n448), .B2(new_n444), .ZN(new_n449));
  OAI21_X1  g0249(.A(KEYINPUT77), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n333), .B1(new_n284), .B2(G68), .ZN(new_n451));
  AOI21_X1  g0251(.A(new_n335), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n452));
  OAI21_X1  g0252(.A(new_n444), .B1(new_n452), .B2(new_n258), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(KEYINPUT18), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT77), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n448), .A2(new_n447), .A3(new_n444), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n338), .B(new_n442), .C1(new_n450), .C2(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(G33), .A2(G283), .ZN(new_n459));
  INV_X1    g0259(.A(G97), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n459), .B(new_n218), .C1(G33), .C2(new_n460), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(new_n246), .C1(new_n218), .C2(G116), .ZN(new_n462));
  XNOR2_X1  g0262(.A(new_n462), .B(KEYINPUT20), .ZN(new_n463));
  INV_X1    g0263(.A(G116), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n244), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n247), .B1(G1), .B2(new_n260), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(new_n464), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n463), .A2(new_n467), .ZN(new_n468));
  XNOR2_X1  g0268(.A(KEYINPUT5), .B(G41), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n312), .A2(G1), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n471), .A2(G270), .A3(new_n305), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n469), .A2(new_n305), .A3(G274), .A4(new_n470), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(G264), .B(G1698), .C1(new_n270), .C2(new_n266), .ZN(new_n475));
  OAI211_X1 g0275(.A(G257), .B(new_n341), .C1(new_n270), .C2(new_n266), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n291), .A2(new_n266), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G303), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n479), .B2(new_n324), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n468), .A2(new_n480), .A3(new_n360), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(KEYINPUT21), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n480), .A2(G190), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n468), .B1(new_n480), .B2(new_n327), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT85), .ZN(new_n487));
  AOI211_X1 g0287(.A(new_n347), .B(new_n474), .C1(new_n479), .C2(new_n324), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n480), .A2(new_n360), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n488), .B1(new_n489), .B2(KEYINPUT21), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n487), .B1(new_n490), .B2(new_n468), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n479), .A2(new_n324), .ZN(new_n492));
  OAI211_X1 g0292(.A(KEYINPUT21), .B(G169), .C1(new_n492), .C2(new_n474), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n480), .A2(G179), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  INV_X1    g0295(.A(new_n468), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n495), .A2(KEYINPUT85), .A3(new_n496), .ZN(new_n497));
  AOI211_X1 g0297(.A(new_n482), .B(new_n486), .C1(new_n491), .C2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT6), .ZN(new_n499));
  NOR3_X1   g0299(.A1(new_n499), .A2(new_n460), .A3(G107), .ZN(new_n500));
  XNOR2_X1  g0300(.A(G97), .B(G107), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n500), .B1(new_n499), .B2(new_n501), .ZN(new_n502));
  OAI22_X1  g0302(.A1(new_n502), .A2(new_n218), .B1(new_n388), .B2(new_n409), .ZN(new_n503));
  AOI21_X1  g0303(.A(new_n344), .B1(new_n293), .B2(new_n295), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n246), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NOR2_X1   g0305(.A1(new_n257), .A2(G97), .ZN(new_n506));
  INV_X1    g0306(.A(new_n466), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n506), .B1(new_n507), .B2(G97), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n324), .B1(new_n470), .B2(new_n469), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(G257), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(new_n473), .ZN(new_n512));
  OAI211_X1 g0312(.A(G250), .B(G1698), .C1(new_n291), .C2(new_n266), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n459), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT4), .ZN(new_n515));
  NOR2_X1   g0315(.A1(new_n515), .A2(new_n339), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n294), .A2(new_n341), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT79), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT79), .ZN(new_n519));
  NAND4_X1  g0319(.A1(new_n294), .A2(new_n519), .A3(new_n341), .A4(new_n516), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n514), .B1(new_n518), .B2(new_n520), .ZN(new_n521));
  OAI211_X1 g0321(.A(G244), .B(new_n341), .C1(new_n270), .C2(new_n266), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n515), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n512), .B1(new_n524), .B2(new_n324), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n509), .B1(new_n525), .B2(G190), .ZN(new_n526));
  OAI21_X1  g0326(.A(KEYINPUT80), .B1(new_n525), .B2(new_n327), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT80), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n305), .B1(new_n521), .B2(new_n523), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n528), .B(G200), .C1(new_n529), .C2(new_n512), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n526), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n524), .A2(new_n324), .ZN(new_n532));
  INV_X1    g0332(.A(new_n512), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n360), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n525), .A2(new_n347), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n536), .A3(new_n509), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n531), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n538), .A2(KEYINPUT81), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT81), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n531), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(G250), .B(new_n341), .C1(new_n270), .C2(new_n266), .ZN(new_n543));
  OAI211_X1 g0343(.A(G257), .B(G1698), .C1(new_n270), .C2(new_n266), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n264), .A2(G294), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n543), .A2(new_n544), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n324), .ZN(new_n547));
  INV_X1    g0347(.A(G190), .ZN(new_n548));
  AND3_X1   g0348(.A1(new_n471), .A2(G264), .A3(new_n305), .ZN(new_n549));
  INV_X1    g0349(.A(new_n549), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n547), .A2(new_n548), .A3(new_n473), .A4(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(new_n473), .ZN(new_n552));
  AOI211_X1 g0352(.A(new_n552), .B(new_n549), .C1(new_n546), .C2(new_n324), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n551), .B(KEYINPUT88), .C1(new_n553), .C2(G200), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n549), .B1(new_n546), .B2(new_n324), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n473), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT88), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n327), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT25), .ZN(new_n559));
  NOR3_X1   g0359(.A1(new_n257), .A2(new_n559), .A3(G107), .ZN(new_n560));
  AOI21_X1  g0360(.A(KEYINPUT25), .B1(new_n244), .B2(new_n344), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n466), .A2(new_n344), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT22), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(new_n322), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n564), .B1(new_n270), .B2(new_n266), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n277), .A2(new_n464), .ZN(new_n566));
  INV_X1    g0366(.A(new_n566), .ZN(new_n567));
  AOI21_X1  g0367(.A(G20), .B1(new_n565), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n218), .A2(G87), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n563), .B1(new_n477), .B2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(KEYINPUT23), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(new_n344), .A3(G20), .ZN(new_n572));
  INV_X1    g0372(.A(KEYINPUT87), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n571), .A2(new_n344), .A3(KEYINPUT87), .A4(G20), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT86), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(KEYINPUT23), .B1(new_n344), .B2(G20), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n578), .B1(new_n577), .B2(KEYINPUT23), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n570), .A2(new_n576), .A3(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(KEYINPUT24), .B1(new_n568), .B2(new_n580), .ZN(new_n581));
  AND3_X1   g0381(.A1(new_n570), .A2(new_n576), .A3(new_n579), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT24), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n566), .B1(new_n281), .B2(new_n564), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n582), .B(new_n583), .C1(G20), .C2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g0386(.A(new_n562), .B1(new_n586), .B2(new_n246), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n554), .A2(new_n558), .A3(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(new_n470), .ZN(new_n589));
  AND2_X1   g0389(.A1(new_n589), .A2(G250), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n305), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n305), .A2(G274), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n592), .B2(new_n589), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n281), .A2(G244), .A3(G1698), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n281), .A2(G238), .A3(new_n341), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n594), .A2(new_n595), .A3(new_n567), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n593), .B1(new_n596), .B2(new_n324), .ZN(new_n597));
  OAI21_X1  g0397(.A(KEYINPUT84), .B1(new_n597), .B2(new_n364), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(G190), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n356), .ZN(new_n601));
  NOR2_X1   g0401(.A1(new_n601), .A2(new_n257), .ZN(new_n602));
  INV_X1    g0402(.A(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n237), .A2(G20), .ZN(new_n604));
  NOR3_X1   g0404(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n605));
  AOI21_X1  g0405(.A(G20), .B1(G33), .B2(G97), .ZN(new_n606));
  OAI21_X1  g0406(.A(KEYINPUT19), .B1(new_n605), .B2(new_n606), .ZN(new_n607));
  INV_X1    g0407(.A(KEYINPUT19), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(new_n218), .A3(G33), .A4(G97), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n281), .A2(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT82), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n246), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n604), .B1(new_n270), .B2(new_n266), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n607), .A2(new_n609), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n613), .A2(new_n611), .A3(new_n614), .ZN(new_n615));
  INV_X1    g0415(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n603), .B1(new_n612), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(KEYINPUT83), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n613), .A2(new_n614), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT82), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n246), .A3(new_n615), .ZN(new_n621));
  INV_X1    g0421(.A(KEYINPUT83), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n621), .A2(new_n622), .A3(new_n603), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n618), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n507), .A2(G87), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n597), .A2(KEYINPUT84), .A3(G190), .ZN(new_n626));
  NAND4_X1  g0426(.A1(new_n600), .A2(new_n624), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n556), .A2(new_n360), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n553), .A2(new_n347), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n290), .B1(new_n581), .B2(new_n585), .ZN(new_n630));
  OAI211_X1 g0430(.A(new_n628), .B(new_n629), .C1(new_n630), .C2(new_n562), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n507), .A2(new_n601), .ZN(new_n632));
  AOI21_X1  g0432(.A(new_n290), .B1(new_n619), .B2(KEYINPUT82), .ZN(new_n633));
  AOI211_X1 g0433(.A(KEYINPUT83), .B(new_n602), .C1(new_n633), .C2(new_n615), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n622), .B1(new_n621), .B2(new_n603), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n632), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n597), .A2(new_n347), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n597), .A2(G169), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  AND4_X1   g0440(.A1(new_n588), .A2(new_n627), .A3(new_n631), .A4(new_n640), .ZN(new_n641));
  AND4_X1   g0441(.A1(new_n458), .A2(new_n498), .A3(new_n542), .A4(new_n641), .ZN(G372));
  NAND2_X1  g0442(.A1(new_n596), .A2(new_n324), .ZN(new_n643));
  INV_X1    g0443(.A(new_n593), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n364), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  OAI211_X1 g0447(.A(new_n647), .B(new_n625), .C1(new_n634), .C2(new_n635), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT89), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n624), .A2(KEYINPUT89), .A3(new_n647), .A4(new_n625), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n650), .A2(new_n651), .A3(new_n599), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n588), .A2(new_n531), .A3(new_n537), .ZN(new_n653));
  INV_X1    g0453(.A(new_n482), .ZN(new_n654));
  OAI211_X1 g0454(.A(new_n631), .B(new_n654), .C1(new_n468), .C2(new_n490), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n652), .A2(new_n653), .A3(new_n655), .A4(new_n640), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT26), .ZN(new_n657));
  AND3_X1   g0457(.A1(new_n535), .A2(new_n536), .A3(new_n509), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n652), .A2(new_n657), .A3(new_n658), .A4(new_n640), .ZN(new_n659));
  INV_X1    g0459(.A(new_n640), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n627), .A2(new_n640), .A3(new_n658), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(KEYINPUT26), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n656), .A2(new_n659), .A3(new_n662), .ZN(new_n663));
  AND2_X1   g0463(.A1(new_n458), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n454), .A2(new_n456), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n386), .A2(new_n396), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n437), .A2(new_n351), .A3(new_n361), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(KEYINPUT90), .ZN(new_n669));
  XNOR2_X1  g0469(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n338), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n665), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(new_n429), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n433), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  OR2_X1    g0474(.A1(new_n664), .A2(new_n674), .ZN(G369));
  NAND2_X1  g0475(.A1(new_n491), .A2(new_n497), .ZN(new_n676));
  INV_X1    g0476(.A(new_n486), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n254), .A2(new_n218), .A3(G13), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n678), .A2(KEYINPUT27), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G213), .A3(new_n680), .ZN(new_n681));
  OR2_X1    g0481(.A1(new_n681), .A2(KEYINPUT91), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n681), .A2(KEYINPUT91), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(G343), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n686), .A2(new_n496), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n676), .A2(new_n654), .A3(new_n677), .A4(new_n687), .ZN(new_n688));
  OAI211_X1 g0488(.A(new_n496), .B(new_n686), .C1(new_n482), .C2(new_n495), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  INV_X1    g0491(.A(new_n691), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n686), .B1(new_n630), .B2(new_n562), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n588), .A2(new_n631), .A3(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(KEYINPUT92), .ZN(new_n695));
  INV_X1    g0495(.A(KEYINPUT92), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n588), .A2(new_n631), .A3(new_n696), .A4(new_n693), .ZN(new_n697));
  NAND2_X1  g0497(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g0498(.A(new_n631), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n692), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n686), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(KEYINPUT85), .B1(new_n495), .B2(new_n496), .ZN(new_n705));
  AOI211_X1 g0505(.A(new_n487), .B(new_n468), .C1(new_n493), .C2(new_n494), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n654), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND4_X1  g0507(.A1(new_n695), .A2(new_n707), .A3(new_n703), .A4(new_n697), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n702), .A2(new_n704), .A3(new_n708), .ZN(G399));
  NAND2_X1  g0509(.A1(new_n214), .A2(new_n304), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT93), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n605), .A2(new_n464), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n254), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n713), .B1(new_n221), .B2(new_n711), .ZN(new_n714));
  XOR2_X1   g0514(.A(new_n714), .B(KEYINPUT28), .Z(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n542), .A2(new_n641), .A3(new_n498), .A4(new_n703), .ZN(new_n717));
  AND2_X1   g0517(.A1(new_n525), .A2(new_n555), .ZN(new_n718));
  NAND4_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .A3(new_n488), .A4(new_n597), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n597), .A2(new_n480), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n720), .A2(new_n534), .A3(new_n347), .A4(new_n556), .ZN(new_n721));
  INV_X1    g0521(.A(KEYINPUT30), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n525), .A2(new_n555), .A3(new_n597), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n722), .B1(new_n723), .B2(new_n494), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  AND3_X1   g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n686), .ZN(new_n726));
  AOI21_X1  g0526(.A(KEYINPUT31), .B1(new_n725), .B2(new_n686), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n716), .B1(new_n717), .B2(new_n728), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n663), .A2(new_n703), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT29), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND4_X1  g0532(.A1(new_n652), .A2(KEYINPUT26), .A3(new_n658), .A4(new_n640), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n661), .A2(new_n657), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n654), .B(new_n631), .C1(new_n705), .C2(new_n706), .ZN(new_n736));
  NAND4_X1  g0536(.A1(new_n736), .A2(new_n652), .A3(new_n653), .A4(new_n640), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n640), .ZN(new_n738));
  OAI211_X1 g0538(.A(KEYINPUT29), .B(new_n703), .C1(new_n735), .C2(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n729), .B1(new_n732), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n715), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n218), .A2(new_n548), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n347), .A2(G200), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(G322), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n477), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n218), .A2(new_n347), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n548), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  INV_X1    g0550(.A(G326), .ZN(new_n751));
  INV_X1    g0551(.A(G294), .ZN(new_n752));
  NOR3_X1   g0552(.A1(new_n548), .A2(G179), .A3(G200), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n218), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n218), .A2(G190), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(new_n743), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI211_X1 g0558(.A(new_n746), .B(new_n755), .C1(G311), .C2(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n756), .A2(new_n347), .A3(new_n327), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT98), .ZN(new_n761));
  OR2_X1    g0561(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n761), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g0564(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n765), .A2(G329), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n646), .A2(new_n347), .A3(new_n742), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n646), .A2(new_n347), .A3(new_n756), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G303), .A2(new_n768), .B1(new_n770), .B2(G283), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n747), .A2(new_n548), .A3(G200), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n772), .A2(KEYINPUT99), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n772), .A2(KEYINPUT99), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  XNOR2_X1  g0576(.A(KEYINPUT33), .B(G317), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n759), .A2(new_n766), .A3(new_n771), .A4(new_n778), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n754), .A2(new_n460), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n294), .B1(new_n757), .B2(new_n388), .C1(new_n249), .C2(new_n744), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n780), .B(new_n781), .C1(G50), .C2(new_n749), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G87), .A2(new_n768), .B1(new_n770), .B2(G107), .ZN(new_n783));
  OAI211_X1 g0583(.A(new_n782), .B(new_n783), .C1(new_n237), .C2(new_n775), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n765), .A2(G159), .ZN(new_n785));
  XNOR2_X1  g0585(.A(new_n785), .B(KEYINPUT32), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n779), .B1(new_n784), .B2(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n217), .B1(G20), .B2(new_n360), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n243), .A2(G20), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n254), .B1(new_n790), .B2(G45), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n711), .A2(new_n792), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n214), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n477), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n796), .A2(G355), .B1(new_n464), .B2(new_n795), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n268), .A2(new_n271), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n798), .A2(new_n795), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n800), .B1(new_n312), .B2(new_n221), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n802), .B1(new_n312), .B2(new_n241), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n801), .A2(KEYINPUT95), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n797), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g0605(.A1(G13), .A2(G33), .ZN(new_n806));
  INV_X1    g0606(.A(new_n806), .ZN(new_n807));
  NOR2_X1   g0607(.A1(new_n807), .A2(G20), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n808), .A2(new_n788), .ZN(new_n809));
  XOR2_X1   g0609(.A(new_n809), .B(KEYINPUT96), .Z(new_n810));
  AOI21_X1  g0610(.A(new_n794), .B1(new_n805), .B2(new_n810), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n789), .B1(new_n811), .B2(KEYINPUT97), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n812), .B1(KEYINPUT97), .B2(new_n811), .ZN(new_n813));
  INV_X1    g0613(.A(new_n808), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n813), .B1(new_n690), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(KEYINPUT94), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(new_n690), .B2(G330), .ZN(new_n817));
  AOI211_X1 g0617(.A(KEYINPUT94), .B(new_n716), .C1(new_n688), .C2(new_n689), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n819), .B(new_n794), .C1(G330), .C2(new_n690), .ZN(new_n820));
  AND2_X1   g0620(.A1(new_n815), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(G396));
  NOR2_X1   g0622(.A1(new_n703), .A2(new_n358), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n362), .A2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n366), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n824), .B1(new_n825), .B2(new_n823), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT100), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT100), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n828), .B(new_n824), .C1(new_n825), .C2(new_n823), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n730), .A2(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n663), .A2(new_n830), .A3(new_n703), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n729), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n793), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n835), .B2(new_n834), .ZN(new_n837));
  INV_X1    g0637(.A(new_n788), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n838), .A2(new_n807), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n793), .B1(G77), .B2(new_n839), .ZN(new_n840));
  OAI221_X1 g0640(.A(new_n477), .B1(new_n757), .B2(new_n464), .C1(new_n752), .C2(new_n744), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n780), .B(new_n841), .C1(G303), .C2(new_n749), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n765), .A2(G311), .ZN(new_n843));
  AOI22_X1  g0643(.A1(G107), .A2(new_n768), .B1(new_n770), .B2(G87), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n776), .A2(G283), .ZN(new_n845));
  NAND4_X1  g0645(.A1(new_n842), .A2(new_n843), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  INV_X1    g0646(.A(new_n744), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G143), .A2(new_n847), .B1(new_n758), .B2(G159), .ZN(new_n848));
  INV_X1    g0648(.A(G137), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n848), .B1(new_n849), .B2(new_n750), .C1(new_n775), .C2(new_n408), .ZN(new_n850));
  XOR2_X1   g0650(.A(new_n850), .B(KEYINPUT34), .Z(new_n851));
  AOI22_X1  g0651(.A1(new_n765), .A2(G132), .B1(G50), .B2(new_n768), .ZN(new_n852));
  INV_X1    g0652(.A(new_n754), .ZN(new_n853));
  AOI22_X1  g0653(.A1(new_n770), .A2(G68), .B1(G58), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n852), .A2(new_n798), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n846), .B1(new_n851), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n840), .B1(new_n856), .B2(new_n788), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n857), .B1(new_n830), .B2(new_n807), .ZN(new_n858));
  AND2_X1   g0658(.A1(new_n837), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n859), .ZN(G384));
  INV_X1    g0660(.A(new_n502), .ZN(new_n861));
  OR2_X1    g0661(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(KEYINPUT35), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n862), .A2(G116), .A3(new_n219), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g0664(.A(new_n864), .B(KEYINPUT36), .Z(new_n865));
  OAI211_X1 g0665(.A(new_n221), .B(G77), .C1(new_n249), .C2(new_n237), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n254), .B(G13), .C1(new_n866), .C2(new_n236), .ZN(new_n867));
  NOR2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g0668(.A1(new_n351), .A2(new_n361), .A3(new_n703), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n833), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n435), .A2(new_n703), .ZN(new_n871));
  INV_X1    g0671(.A(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n666), .A2(new_n437), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n386), .B1(new_n439), .B2(new_n440), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n873), .B1(new_n874), .B2(new_n872), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n870), .A2(new_n875), .ZN(new_n876));
  OR2_X1    g0676(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n285), .A2(new_n288), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n298), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n290), .B1(new_n451), .B2(KEYINPUT16), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n258), .B1(new_n879), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n336), .B1(new_n881), .B2(new_n684), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n445), .ZN(new_n883));
  OAI21_X1  g0683(.A(KEYINPUT37), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  XOR2_X1   g0684(.A(new_n684), .B(KEYINPUT102), .Z(new_n885));
  OAI21_X1  g0685(.A(new_n885), .B1(new_n452), .B2(new_n258), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT37), .ZN(new_n887));
  NAND4_X1  g0687(.A1(new_n453), .A2(new_n886), .A3(new_n887), .A4(new_n336), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g0689(.A(new_n338), .B1(new_n450), .B2(new_n457), .ZN(new_n890));
  OR2_X1    g0690(.A1(new_n881), .A2(new_n684), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n889), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT38), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n889), .B(KEYINPUT38), .C1(new_n890), .C2(new_n891), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n876), .A2(KEYINPUT101), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n877), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n453), .A2(new_n886), .A3(new_n336), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n899), .A2(KEYINPUT37), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n900), .A2(KEYINPUT103), .A3(new_n888), .ZN(new_n901));
  INV_X1    g0701(.A(new_n886), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n902), .B1(new_n665), .B2(new_n338), .ZN(new_n903));
  INV_X1    g0703(.A(KEYINPUT103), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n899), .A2(new_n904), .A3(KEYINPUT37), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n901), .A2(new_n903), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n893), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n895), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT39), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g0710(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n911));
  INV_X1    g0711(.A(new_n666), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n912), .A2(new_n703), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n910), .A2(new_n911), .A3(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n885), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n665), .A2(new_n916), .ZN(new_n917));
  AND3_X1   g0717(.A1(new_n898), .A2(new_n915), .A3(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n458), .A2(new_n732), .A3(new_n739), .ZN(new_n919));
  INV_X1    g0719(.A(KEYINPUT104), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n458), .A2(new_n732), .A3(new_n739), .A4(KEYINPUT104), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n674), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n918), .B(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  INV_X1    g0725(.A(new_n875), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n831), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n717), .A2(new_n728), .ZN(new_n928));
  AND2_X1   g0728(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n925), .B1(new_n908), .B2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n927), .A2(new_n925), .A3(new_n928), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n931), .B1(new_n894), .B2(new_n895), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n458), .A2(new_n928), .ZN(new_n935));
  AOI21_X1  g0735(.A(new_n716), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n935), .B2(new_n934), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n924), .A2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n254), .B2(new_n790), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n924), .A2(new_n937), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n868), .B1(new_n939), .B2(new_n940), .ZN(G367));
  OAI21_X1  g0741(.A(new_n809), .B1(new_n214), .B2(new_n356), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n942), .B1(new_n799), .B2(new_n230), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n768), .A2(G116), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT46), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n754), .A2(new_n344), .ZN(new_n946));
  INV_X1    g0746(.A(G303), .ZN(new_n947));
  INV_X1    g0747(.A(G283), .ZN(new_n948));
  OAI22_X1  g0748(.A1(new_n744), .A2(new_n947), .B1(new_n757), .B2(new_n948), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n946), .B(new_n949), .C1(G311), .C2(new_n749), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n765), .A2(G317), .B1(G97), .B2(new_n770), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n798), .B1(new_n776), .B2(G294), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n945), .A2(new_n950), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n769), .A2(new_n388), .ZN(new_n954));
  OAI221_X1 g0754(.A(new_n294), .B1(new_n235), .B2(new_n757), .C1(new_n767), .C2(new_n249), .ZN(new_n955));
  XNOR2_X1  g0755(.A(KEYINPUT111), .B(G137), .ZN(new_n956));
  AOI211_X1 g0756(.A(new_n954), .B(new_n955), .C1(new_n765), .C2(new_n956), .ZN(new_n957));
  INV_X1    g0757(.A(G159), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n957), .B1(new_n958), .B2(new_n775), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n749), .A2(G143), .B1(new_n847), .B2(G150), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n960), .B1(new_n237), .B2(new_n754), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n961), .B(KEYINPUT110), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n953), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  XNOR2_X1  g0763(.A(new_n963), .B(KEYINPUT47), .ZN(new_n964));
  AOI211_X1 g0764(.A(new_n794), .B(new_n943), .C1(new_n964), .C2(new_n788), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n703), .B1(new_n624), .B2(new_n625), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n966), .A2(new_n640), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n652), .A2(new_n640), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n967), .B1(new_n968), .B2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT105), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n965), .B1(new_n970), .B2(new_n814), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n708), .A2(new_n704), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n686), .A2(new_n509), .ZN(new_n973));
  OAI22_X1  g0773(.A1(new_n538), .A2(new_n973), .B1(new_n537), .B2(new_n703), .ZN(new_n974));
  INV_X1    g0774(.A(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n972), .A2(KEYINPUT44), .A3(new_n975), .ZN(new_n979));
  NAND4_X1  g0779(.A1(new_n708), .A2(KEYINPUT45), .A3(new_n704), .A4(new_n974), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n708), .A2(new_n704), .A3(new_n974), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n978), .A2(new_n979), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(KEYINPUT107), .B1(new_n984), .B2(new_n702), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(new_n980), .ZN(new_n986));
  AOI21_X1  g0786(.A(KEYINPUT44), .B1(new_n972), .B2(new_n975), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n977), .B(new_n974), .C1(new_n708), .C2(new_n704), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n986), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT107), .ZN(new_n990));
  INV_X1    g0790(.A(new_n702), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n989), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n691), .A2(KEYINPUT94), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n707), .A2(new_n703), .ZN(new_n994));
  NAND3_X1  g0794(.A1(new_n698), .A2(new_n700), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n995), .A2(new_n708), .ZN(new_n996));
  INV_X1    g0796(.A(KEYINPUT108), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n690), .A2(new_n816), .A3(G330), .ZN(new_n998));
  NAND4_X1  g0798(.A1(new_n993), .A2(new_n996), .A3(new_n997), .A4(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n692), .A2(new_n708), .A3(new_n995), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n997), .B1(new_n819), .B2(new_n996), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n1001), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g0803(.A1(new_n985), .A2(new_n992), .A3(new_n740), .A4(new_n1003), .ZN(new_n1004));
  OAI211_X1 g0804(.A(new_n986), .B(new_n702), .C1(new_n987), .C2(new_n988), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT109), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n978), .A2(new_n979), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1008), .A2(KEYINPUT109), .A3(new_n702), .A4(new_n986), .ZN(new_n1009));
  AND2_X1   g0809(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n740), .B1(new_n1004), .B2(new_n1010), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n711), .B(KEYINPUT41), .Z(new_n1012));
  INV_X1    g0812(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n792), .B1(new_n1011), .B2(new_n1013), .ZN(new_n1014));
  NAND2_X1  g0814(.A1(new_n970), .A2(KEYINPUT43), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n969), .A2(KEYINPUT105), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT43), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n969), .A2(KEYINPUT105), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1016), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(KEYINPUT42), .B1(new_n708), .B2(new_n975), .ZN(new_n1020));
  NOR3_X1   g0820(.A1(new_n538), .A2(new_n631), .A3(new_n973), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n703), .B1(new_n1021), .B2(new_n658), .ZN(new_n1022));
  AND2_X1   g0822(.A1(new_n1020), .A2(new_n1022), .ZN(new_n1023));
  OR3_X1    g0823(.A1(new_n708), .A2(new_n975), .A3(KEYINPUT42), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g0825(.A1(new_n1015), .A2(new_n1019), .A3(new_n1025), .ZN(new_n1026));
  XOR2_X1   g0826(.A(new_n969), .B(KEYINPUT105), .Z(new_n1027));
  NAND4_X1  g0827(.A1(new_n1027), .A2(new_n1023), .A3(new_n1017), .A4(new_n1024), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n702), .A2(new_n975), .ZN(new_n1029));
  NAND3_X1  g0829(.A1(new_n1026), .A2(new_n1028), .A3(new_n1029), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(KEYINPUT106), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT106), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1026), .A2(new_n1028), .A3(new_n1032), .A4(new_n1029), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1029), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1034), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n971), .B1(new_n1014), .B2(new_n1038), .ZN(G387));
  NAND2_X1  g0839(.A1(new_n1003), .A2(new_n740), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n732), .A2(new_n739), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n1041), .A2(new_n729), .B1(new_n1001), .B2(new_n1002), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n711), .B(KEYINPUT112), .ZN(new_n1043));
  NAND3_X1  g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n800), .B1(G45), .B2(new_n227), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1045), .B1(new_n712), .B2(new_n796), .ZN(new_n1046));
  NOR3_X1   g0846(.A1(new_n407), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT50), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n253), .B2(new_n235), .ZN(new_n1049));
  OAI21_X1  g0849(.A(new_n312), .B1(new_n237), .B2(new_n388), .ZN(new_n1050));
  NOR4_X1   g0850(.A1(new_n1047), .A2(new_n1049), .A3(new_n712), .A4(new_n1050), .ZN(new_n1051));
  OAI22_X1  g0851(.A1(new_n1046), .A2(new_n1051), .B1(G107), .B2(new_n214), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n794), .B1(new_n1052), .B2(new_n810), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n744), .A2(new_n235), .B1(new_n757), .B2(new_n237), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G159), .B2(new_n749), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n1055), .B(new_n798), .C1(new_n356), .C2(new_n754), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n764), .A2(new_n408), .B1(new_n460), .B2(new_n769), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n775), .A2(new_n407), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n767), .A2(new_n388), .ZN(new_n1059));
  NOR4_X1   g0859(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  OAI22_X1  g0860(.A1(new_n764), .A2(new_n751), .B1(new_n464), .B2(new_n769), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G317), .A2(new_n847), .B1(new_n758), .B2(G303), .ZN(new_n1062));
  INV_X1    g0862(.A(G311), .ZN(new_n1063));
  OAI221_X1 g0863(.A(new_n1062), .B1(new_n745), .B2(new_n750), .C1(new_n775), .C2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT48), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n768), .A2(G294), .B1(G283), .B2(new_n853), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1066), .A2(new_n1067), .A3(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(new_n1069), .ZN(new_n1070));
  AOI211_X1 g0870(.A(new_n798), .B(new_n1061), .C1(new_n1070), .C2(KEYINPUT49), .ZN(new_n1071));
  OR2_X1    g0871(.A1(new_n1070), .A2(KEYINPUT49), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n1060), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1053), .B1(new_n1073), .B2(new_n838), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n701), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1074), .B1(new_n1075), .B2(new_n808), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1076), .B1(new_n1003), .B2(new_n792), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1044), .A2(new_n1077), .ZN(G393));
  AOI22_X1  g0878(.A1(new_n1007), .A2(new_n1009), .B1(new_n991), .B2(new_n989), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(new_n792), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n809), .B1(new_n214), .B2(new_n460), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1081), .B1(new_n799), .B2(new_n234), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n767), .A2(new_n237), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n754), .A2(new_n388), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1084), .B1(new_n253), .B2(new_n758), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1085), .B1(new_n322), .B2(new_n769), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n1083), .B(new_n1086), .C1(G143), .C2(new_n765), .ZN(new_n1087));
  AOI22_X1  g0887(.A1(new_n749), .A2(G150), .B1(new_n847), .B2(G159), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1088), .B(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n776), .A2(G50), .ZN(new_n1091));
  NAND4_X1  g0891(.A1(new_n1087), .A2(new_n798), .A3(new_n1090), .A4(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n294), .B1(new_n770), .B2(G107), .ZN(new_n1093));
  OAI221_X1 g0893(.A(new_n1093), .B1(new_n948), .B2(new_n767), .C1(new_n745), .C2(new_n764), .ZN(new_n1094));
  XOR2_X1   g0894(.A(new_n1094), .B(KEYINPUT114), .Z(new_n1095));
  AOI22_X1  g0895(.A1(new_n749), .A2(G317), .B1(new_n847), .B2(G311), .ZN(new_n1096));
  XOR2_X1   g0896(.A(new_n1096), .B(KEYINPUT52), .Z(new_n1097));
  AOI22_X1  g0897(.A1(new_n853), .A2(G116), .B1(new_n758), .B2(G294), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(new_n947), .C2(new_n775), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1092), .B1(new_n1095), .B2(new_n1099), .ZN(new_n1100));
  AOI211_X1 g0900(.A(new_n794), .B(new_n1082), .C1(new_n1100), .C2(new_n788), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n814), .B2(new_n974), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1007), .A2(new_n1009), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n993), .A2(new_n996), .A3(new_n998), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1104), .A2(KEYINPUT108), .ZN(new_n1105));
  AND4_X1   g0905(.A1(new_n740), .A2(new_n1105), .A3(new_n1000), .A4(new_n999), .ZN(new_n1106));
  NAND4_X1  g0906(.A1(new_n1103), .A2(new_n1106), .A3(new_n992), .A4(new_n985), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n1043), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n1079), .A2(new_n1106), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1080), .B(new_n1102), .C1(new_n1108), .C2(new_n1109), .ZN(G390));
  AOI21_X1  g0910(.A(new_n914), .B1(new_n870), .B2(new_n875), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n1111), .ZN(new_n1112));
  AND3_X1   g0912(.A1(new_n894), .A2(KEYINPUT39), .A3(new_n895), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT39), .B1(new_n907), .B2(new_n895), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n1112), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n928), .A2(G330), .A3(new_n875), .A4(new_n830), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n830), .B(new_n703), .C1(new_n735), .C2(new_n738), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n869), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n875), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n908), .A2(new_n1119), .A3(new_n913), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1115), .A2(new_n1116), .A3(new_n1120), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1116), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1111), .B1(new_n910), .B2(new_n911), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1120), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1122), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n729), .A2(new_n830), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n926), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1127), .A2(new_n869), .A3(new_n1116), .A4(new_n1117), .ZN(new_n1128));
  INV_X1    g0928(.A(KEYINPUT115), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1116), .A2(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n875), .B1(new_n729), .B2(new_n830), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n870), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1129), .B(new_n875), .C1(new_n729), .C2(new_n830), .ZN(new_n1133));
  OAI21_X1  g0933(.A(new_n1128), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n458), .A2(new_n729), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1134), .A2(new_n923), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n1121), .A2(new_n1125), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(KEYINPUT116), .ZN(new_n1138));
  INV_X1    g0938(.A(KEYINPUT116), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1121), .A2(new_n1125), .A3(new_n1136), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1043), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1121), .A2(new_n1125), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1136), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1142), .B1(new_n1143), .B2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1141), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1143), .A2(new_n791), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n806), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n793), .B1(new_n253), .B2(new_n839), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n477), .B1(new_n757), .B2(new_n460), .C1(new_n464), .C2(new_n744), .ZN(new_n1150));
  AOI211_X1 g0950(.A(new_n1084), .B(new_n1150), .C1(G283), .C2(new_n749), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n765), .A2(G294), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G87), .A2(new_n768), .B1(new_n770), .B2(G68), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n776), .A2(G107), .ZN(new_n1154));
  NAND4_X1  g0954(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .A4(new_n1154), .ZN(new_n1155));
  AOI22_X1  g0955(.A1(new_n765), .A2(G125), .B1(G50), .B2(new_n770), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n776), .A2(new_n956), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT54), .B(G143), .ZN(new_n1158));
  OAI21_X1  g0958(.A(new_n294), .B1(new_n757), .B2(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1159), .B1(G132), .B2(new_n847), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G159), .A2(new_n853), .B1(new_n749), .B2(G128), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .A4(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n768), .A2(G150), .ZN(new_n1163));
  XNOR2_X1  g0963(.A(new_n1163), .B(KEYINPUT53), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1155), .B1(new_n1162), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1149), .B1(new_n1165), .B2(new_n788), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1147), .B1(new_n1148), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1146), .A2(new_n1167), .ZN(G378));
  NAND2_X1  g0968(.A1(new_n429), .A2(new_n433), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n418), .A2(new_n684), .ZN(new_n1170));
  XNOR2_X1  g0970(.A(new_n1169), .B(new_n1170), .ZN(new_n1171));
  XNOR2_X1  g0971(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(new_n1171), .B(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n806), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n793), .B1(G50), .B2(new_n839), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n847), .A2(G107), .B1(new_n758), .B2(new_n601), .ZN(new_n1176));
  OAI221_X1 g0976(.A(new_n1176), .B1(new_n237), .B2(new_n754), .C1(new_n464), .C2(new_n750), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(G97), .B2(new_n776), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n798), .A2(G41), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n769), .A2(new_n249), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1059), .B(new_n1180), .C1(new_n765), .C2(G283), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1178), .A2(new_n1179), .A3(new_n1181), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(new_n1182), .B(KEYINPUT58), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n767), .A2(new_n1158), .ZN(new_n1184));
  INV_X1    g0984(.A(KEYINPUT117), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(new_n776), .A2(G132), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  NOR2_X1   g0986(.A1(new_n754), .A2(new_n408), .ZN(new_n1187));
  INV_X1    g0987(.A(G128), .ZN(new_n1188));
  OAI22_X1  g0988(.A1(new_n744), .A2(new_n1188), .B1(new_n757), .B2(new_n849), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1187), .B(new_n1189), .C1(G125), .C2(new_n749), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n1186), .B(new_n1190), .C1(new_n1185), .C2(new_n1184), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(KEYINPUT59), .ZN(new_n1193));
  OAI211_X1 g0993(.A(new_n260), .B(new_n304), .C1(new_n769), .C2(new_n958), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G124), .B2(new_n765), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1196));
  OAI21_X1  g0996(.A(new_n235), .B1(G33), .B2(G41), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1183), .B1(new_n1192), .B2(new_n1196), .C1(new_n1179), .C2(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT118), .ZN(new_n1199));
  OR2_X1    g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(new_n838), .B1(new_n1198), .B2(new_n1199), .ZN(new_n1201));
  AOI21_X1  g1001(.A(new_n1175), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1174), .A2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1173), .B1(new_n933), .B2(new_n716), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1173), .ZN(new_n1205));
  OAI211_X1 g1005(.A(G330), .B(new_n1205), .C1(new_n930), .C2(new_n932), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n918), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n918), .B1(new_n1206), .B2(new_n1204), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1203), .B1(new_n1209), .B2(new_n791), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n1210), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n923), .A2(new_n1135), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1141), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1209), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT57), .B1(new_n1214), .B2(new_n1215), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1212), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1217));
  OAI21_X1  g1017(.A(KEYINPUT57), .B1(new_n1207), .B2(new_n1208), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n1043), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  OAI21_X1  g1019(.A(new_n1211), .B1(new_n1216), .B2(new_n1219), .ZN(G375));
  OAI22_X1  g1020(.A1(new_n750), .A2(new_n752), .B1(new_n356), .B2(new_n754), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n477), .B1(new_n757), .B2(new_n344), .C1(new_n948), .C2(new_n744), .ZN(new_n1222));
  OR3_X1    g1022(.A1(new_n1221), .A2(new_n954), .A3(new_n1222), .ZN(new_n1223));
  OAI22_X1  g1023(.A1(new_n764), .A2(new_n947), .B1(new_n460), .B2(new_n767), .ZN(new_n1224));
  XOR2_X1   g1024(.A(new_n1224), .B(KEYINPUT120), .Z(new_n1225));
  AOI211_X1 g1025(.A(new_n1223), .B(new_n1225), .C1(G116), .C2(new_n776), .ZN(new_n1226));
  AOI22_X1  g1026(.A1(new_n765), .A2(G128), .B1(G159), .B2(new_n768), .ZN(new_n1227));
  AOI22_X1  g1027(.A1(new_n749), .A2(G132), .B1(new_n847), .B2(new_n956), .ZN(new_n1228));
  OAI211_X1 g1028(.A(new_n1227), .B(new_n1228), .C1(new_n249), .C2(new_n769), .ZN(new_n1229));
  OAI22_X1  g1029(.A1(new_n754), .A2(new_n235), .B1(new_n408), .B2(new_n757), .ZN(new_n1230));
  XNOR2_X1  g1030(.A(new_n1230), .B(KEYINPUT121), .ZN(new_n1231));
  OAI21_X1  g1031(.A(new_n798), .B1(new_n775), .B2(new_n1158), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1229), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n788), .B1(new_n1226), .B2(new_n1233), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n793), .B1(G68), .B2(new_n839), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1234), .B(new_n1236), .C1(new_n875), .C2(new_n807), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1134), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1238), .A2(new_n791), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1237), .B1(new_n1239), .B2(KEYINPUT119), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n1240), .B1(KEYINPUT119), .B2(new_n1239), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1212), .A2(new_n1238), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1144), .A2(new_n1013), .A3(new_n1242), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1241), .A2(new_n1243), .ZN(G381));
  INV_X1    g1044(.A(G390), .ZN(new_n1245));
  AND3_X1   g1045(.A1(new_n1044), .A2(new_n821), .A3(new_n1077), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1245), .A2(new_n859), .A3(new_n1246), .ZN(new_n1247));
  OR3_X1    g1047(.A1(G381), .A2(new_n1247), .A3(G387), .ZN(new_n1248));
  OR3_X1    g1048(.A1(G375), .A2(G378), .A3(new_n1248), .ZN(G407));
  INV_X1    g1049(.A(G378), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n685), .A2(G213), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1251), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G407), .B(G213), .C1(G375), .C2(new_n1253), .ZN(G409));
  AOI21_X1  g1054(.A(new_n821), .B1(new_n1044), .B2(new_n1077), .ZN(new_n1255));
  OAI21_X1  g1055(.A(KEYINPUT122), .B1(new_n1246), .B2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(G393), .A2(G396), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT122), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1044), .A2(new_n821), .A3(new_n1077), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1257), .A2(new_n1258), .A3(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1261));
  AOI22_X1  g1061(.A1(new_n1031), .A2(new_n1033), .B1(new_n1036), .B2(new_n1035), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1012), .B1(new_n1107), .B2(new_n740), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1262), .B1(new_n1263), .B2(new_n792), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1264), .A2(new_n971), .A3(G390), .ZN(new_n1265));
  AOI21_X1  g1065(.A(G390), .B1(new_n1264), .B2(new_n971), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1261), .B1(new_n1265), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(G387), .A2(new_n1245), .ZN(new_n1268));
  AND2_X1   g1068(.A1(new_n1256), .A2(new_n1260), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1264), .A2(new_n971), .A3(G390), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1268), .A2(new_n1269), .A3(new_n1270), .ZN(new_n1271));
  AND2_X1   g1071(.A1(new_n1267), .A2(new_n1271), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT125), .ZN(new_n1273));
  OAI211_X1 g1073(.A(G378), .B(new_n1211), .C1(new_n1216), .C2(new_n1219), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1217), .A2(new_n1209), .A3(new_n1012), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1250), .B1(new_n1275), .B2(new_n1210), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1274), .A2(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n1251), .ZN(new_n1278));
  INV_X1    g1078(.A(KEYINPUT60), .ZN(new_n1279));
  AOI211_X1 g1079(.A(new_n1142), .B(new_n1136), .C1(new_n1279), .C2(new_n1242), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1280), .B1(new_n1279), .B2(new_n1242), .ZN(new_n1281));
  AND3_X1   g1081(.A1(new_n1281), .A2(G384), .A3(new_n1241), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G384), .B1(new_n1281), .B2(new_n1241), .ZN(new_n1283));
  OAI211_X1 g1083(.A(G2897), .B(new_n1252), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1281), .A2(new_n1241), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1285), .A2(new_n859), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1281), .A2(G384), .A3(new_n1241), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1252), .A2(G2897), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1286), .A2(new_n1287), .A3(new_n1288), .ZN(new_n1289));
  AND2_X1   g1089(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1278), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1282), .A2(new_n1283), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1277), .A2(new_n1251), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(new_n1293), .A2(KEYINPUT62), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1273), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT61), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1267), .A2(new_n1298), .A3(new_n1271), .ZN(new_n1299));
  INV_X1    g1099(.A(KEYINPUT123), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1299), .A2(new_n1300), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1267), .A2(new_n1271), .A3(KEYINPUT123), .A4(new_n1298), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1252), .B1(new_n1274), .B2(new_n1276), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1284), .A2(new_n1289), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1303), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  AOI21_X1  g1106(.A(KEYINPUT63), .B1(new_n1304), .B2(new_n1292), .ZN(new_n1307));
  NOR2_X1   g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  NAND3_X1  g1108(.A1(new_n1304), .A2(KEYINPUT63), .A3(new_n1292), .ZN(new_n1309));
  AOI21_X1  g1109(.A(KEYINPUT124), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1310));
  AND2_X1   g1110(.A1(new_n1301), .A2(new_n1302), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1311), .B1(new_n1278), .B2(new_n1290), .ZN(new_n1312));
  INV_X1    g1112(.A(KEYINPUT63), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1293), .A2(new_n1313), .ZN(new_n1314));
  AND4_X1   g1114(.A1(KEYINPUT124), .A2(new_n1312), .A3(new_n1309), .A4(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1297), .B1(new_n1310), .B2(new_n1315), .ZN(G405));
  NAND3_X1  g1116(.A1(new_n1286), .A2(KEYINPUT126), .A3(new_n1287), .ZN(new_n1317));
  XNOR2_X1  g1117(.A(new_n1317), .B(KEYINPUT127), .ZN(new_n1318));
  XNOR2_X1  g1118(.A(G375), .B(G378), .ZN(new_n1319));
  OR2_X1    g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1321));
  AND3_X1   g1121(.A1(new_n1320), .A2(new_n1272), .A3(new_n1321), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n1272), .B1(new_n1320), .B2(new_n1321), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1322), .A2(new_n1323), .ZN(G402));
endmodule


