//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 1 1 1 1 0 0 1 0 0 0 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n718, new_n719, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n783, new_n784,
    new_n785, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n795, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n813, new_n814, new_n815, new_n817,
    new_n818, new_n819, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1004, new_n1005, new_n1006, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1016, new_n1017,
    new_n1018, new_n1019, new_n1020, new_n1021, new_n1022, new_n1023,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1051, new_n1052;
  INV_X1    g000(.A(G228gat), .ZN(new_n202));
  INV_X1    g001(.A(G233gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT2), .B1(new_n205), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G141gat), .ZN(new_n208));
  NOR2_X1   g007(.A1(new_n208), .A2(G148gat), .ZN(new_n209));
  INV_X1    g008(.A(G148gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G141gat), .ZN(new_n211));
  OAI211_X1 g010(.A(new_n207), .B(KEYINPUT79), .C1(new_n209), .C2(new_n211), .ZN(new_n212));
  XNOR2_X1  g011(.A(G155gat), .B(G162gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XOR2_X1   g014(.A(G141gat), .B(G148gat), .Z(new_n216));
  NAND4_X1  g015(.A1(new_n216), .A2(KEYINPUT79), .A3(new_n213), .A4(new_n207), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT29), .ZN(new_n220));
  XNOR2_X1  g019(.A(KEYINPUT71), .B(G197gat), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(G204gat), .ZN(new_n222));
  INV_X1    g021(.A(G211gat), .ZN(new_n223));
  INV_X1    g022(.A(G218gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND2_X1  g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT73), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT72), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n225), .A2(KEYINPUT73), .A3(new_n226), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT22), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n222), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g035(.A(new_n232), .B1(new_n222), .B2(new_n234), .ZN(new_n237));
  OAI21_X1  g036(.A(new_n220), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT3), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n219), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n222), .A2(new_n234), .ZN(new_n241));
  INV_X1    g040(.A(new_n232), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n243), .A2(new_n235), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n215), .A2(new_n239), .A3(new_n217), .ZN(new_n245));
  XNOR2_X1  g044(.A(KEYINPUT74), .B(KEYINPUT29), .ZN(new_n246));
  AND2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NOR2_X1   g046(.A1(new_n244), .A2(new_n247), .ZN(new_n248));
  OAI21_X1  g047(.A(new_n204), .B1(new_n240), .B2(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(G78gat), .B(G106gat), .Z(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT84), .ZN(new_n251));
  XNOR2_X1  g050(.A(new_n251), .B(G50gat), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  AND3_X1   g052(.A1(new_n215), .A2(KEYINPUT81), .A3(new_n217), .ZN(new_n254));
  AOI21_X1  g053(.A(KEYINPUT81), .B1(new_n215), .B2(new_n217), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n229), .A2(new_n231), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n241), .A2(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n222), .A2(new_n229), .A3(new_n231), .A4(new_n234), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(new_n246), .A3(new_n259), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n256), .B1(new_n260), .B2(new_n239), .ZN(new_n261));
  INV_X1    g060(.A(new_n204), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(new_n244), .B2(new_n247), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n249), .B(new_n253), .C1(new_n261), .C2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(KEYINPUT29), .B1(new_n243), .B2(new_n235), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n218), .B1(new_n265), .B2(KEYINPUT3), .ZN(new_n266));
  INV_X1    g065(.A(new_n248), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n262), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n261), .A2(new_n263), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n252), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n271));
  INV_X1    g070(.A(G22gat), .ZN(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  AND3_X1   g072(.A1(new_n264), .A2(new_n270), .A3(new_n273), .ZN(new_n274));
  AOI21_X1  g073(.A(new_n273), .B1(new_n264), .B2(new_n270), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT67), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT67), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G120gat), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n278), .A2(new_n280), .A3(G113gat), .ZN(new_n281));
  INV_X1    g080(.A(G113gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n282), .A2(KEYINPUT68), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT68), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(G113gat), .ZN(new_n285));
  NAND3_X1  g084(.A1(new_n283), .A2(new_n285), .A3(G120gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT1), .ZN(new_n288));
  INV_X1    g087(.A(G127gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(G134gat), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n290), .B1(new_n289), .B2(G134gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  AOI21_X1  g091(.A(KEYINPUT1), .B1(new_n282), .B2(new_n277), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(new_n282), .B2(new_n277), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n289), .A2(KEYINPUT66), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT66), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(G127gat), .ZN(new_n297));
  AND3_X1   g096(.A1(new_n295), .A2(new_n297), .A3(G134gat), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT65), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n299), .B1(new_n289), .B2(G134gat), .ZN(new_n300));
  INV_X1    g099(.A(G134gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n301), .A2(KEYINPUT65), .A3(G127gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n300), .A2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n294), .B1(new_n298), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT69), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n292), .A2(new_n304), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n305), .B1(new_n292), .B2(new_n304), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G190gat), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n309), .A2(G183gat), .ZN(new_n310));
  INV_X1    g109(.A(G183gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n311), .A2(G190gat), .ZN(new_n312));
  OAI21_X1  g111(.A(KEYINPUT24), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(G169gat), .A2(G176gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n319), .B1(new_n320), .B2(KEYINPUT24), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n313), .A2(new_n318), .A3(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT25), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n311), .A2(G190gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n309), .A2(G183gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n321), .B1(new_n328), .B2(KEYINPUT24), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT25), .A3(new_n318), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n314), .A2(KEYINPUT26), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT26), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n319), .A2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n331), .B(new_n320), .C1(new_n333), .C2(new_n314), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT28), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n311), .A2(KEYINPUT27), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT27), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(G183gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n338), .A3(new_n309), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT64), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n334), .B1(new_n335), .B2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT28), .ZN(new_n343));
  AOI22_X1  g142(.A1(new_n325), .A2(new_n330), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n308), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n341), .A2(new_n335), .ZN(new_n346));
  INV_X1    g145(.A(new_n334), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n343), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g147(.A(KEYINPUT25), .B1(new_n329), .B2(new_n318), .ZN(new_n349));
  AND4_X1   g148(.A1(KEYINPUT25), .A2(new_n313), .A3(new_n318), .A4(new_n322), .ZN(new_n350));
  OAI21_X1  g149(.A(new_n348), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n307), .B2(new_n306), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n345), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G227gat), .A2(G233gat), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(KEYINPUT33), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g155(.A(G15gat), .B(G43gat), .ZN(new_n357));
  XNOR2_X1  g156(.A(G71gat), .B(G99gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n356), .A2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT34), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(new_n354), .B2(KEYINPUT70), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n362), .B1(new_n353), .B2(new_n355), .ZN(new_n363));
  INV_X1    g162(.A(new_n362), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n345), .A2(new_n352), .A3(new_n354), .A4(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n360), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n365), .B(new_n363), .C1(new_n356), .C2(new_n359), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n353), .A2(new_n355), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT32), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n371), .B1(new_n367), .B2(new_n368), .ZN(new_n374));
  NOR3_X1   g173(.A1(new_n276), .A2(new_n373), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(G226gat), .A2(G233gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n246), .ZN(new_n377));
  OAI211_X1 g176(.A(KEYINPUT75), .B(new_n376), .C1(new_n344), .C2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(new_n376), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n351), .B2(new_n246), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n381), .B1(new_n351), .B2(new_n379), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n244), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(KEYINPUT76), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT76), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(G64gat), .B(G92gat), .ZN(new_n391));
  XOR2_X1   g190(.A(new_n390), .B(new_n391), .Z(new_n392));
  OAI21_X1  g191(.A(new_n376), .B1(new_n344), .B2(KEYINPUT29), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n325), .A2(new_n330), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n376), .B1(new_n394), .B2(new_n348), .ZN(new_n395));
  INV_X1    g194(.A(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n393), .A2(new_n396), .A3(new_n244), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT77), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  NAND4_X1  g198(.A1(new_n393), .A2(new_n396), .A3(KEYINPUT77), .A4(new_n244), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND4_X1  g200(.A1(new_n389), .A2(KEYINPUT30), .A3(new_n392), .A4(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n383), .A2(new_n387), .A3(new_n384), .ZN(new_n403));
  AOI21_X1  g202(.A(new_n387), .B1(new_n383), .B2(new_n384), .ZN(new_n404));
  OAI21_X1  g203(.A(new_n401), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(new_n392), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n402), .A2(new_n407), .A3(KEYINPUT78), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT78), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n392), .B(new_n401), .C1(new_n403), .C2(new_n404), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT30), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n392), .B1(new_n389), .B2(new_n401), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n409), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(G1gat), .B(G29gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT0), .ZN(new_n416));
  XNOR2_X1  g215(.A(G57gat), .B(G85gat), .ZN(new_n417));
  XOR2_X1   g216(.A(new_n416), .B(new_n417), .Z(new_n418));
  NAND2_X1  g217(.A1(new_n218), .A2(KEYINPUT3), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n292), .A2(new_n304), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n419), .A2(new_n420), .A3(new_n245), .ZN(new_n421));
  NAND2_X1  g220(.A1(G225gat), .A2(G233gat), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(KEYINPUT5), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  AND2_X1   g224(.A1(new_n421), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n427), .B1(new_n308), .B2(new_n256), .ZN(new_n428));
  INV_X1    g227(.A(new_n420), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT82), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT4), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n429), .A2(new_n219), .A3(new_n430), .A4(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n292), .A2(new_n304), .A3(new_n215), .A4(new_n217), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT82), .B1(new_n433), .B2(KEYINPUT4), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  OAI21_X1  g234(.A(new_n426), .B1(new_n428), .B2(new_n435), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n218), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n433), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n423), .B1(new_n438), .B2(new_n424), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n433), .A2(KEYINPUT4), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT81), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n218), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n215), .A2(KEYINPUT81), .A3(new_n217), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n292), .A2(new_n304), .A3(new_n305), .ZN(new_n446));
  NAND4_X1  g245(.A1(new_n442), .A2(new_n444), .A3(new_n445), .A4(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n427), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n441), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(KEYINPUT5), .B1(new_n449), .B2(new_n421), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n418), .B1(new_n440), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n449), .A2(new_n421), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n452), .A2(new_n424), .ZN(new_n453));
  INV_X1    g252(.A(new_n418), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n453), .A2(new_n454), .A3(new_n439), .A4(new_n436), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT6), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n451), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n440), .A2(new_n450), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n458), .A2(KEYINPUT6), .A3(new_n454), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n457), .A2(new_n459), .B1(new_n411), .B2(new_n410), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n375), .A2(new_n408), .A3(new_n414), .A4(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n374), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(new_n372), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n410), .A2(new_n411), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(new_n402), .A3(new_n407), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n457), .A2(new_n459), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n468), .A2(new_n276), .A3(KEYINPUT35), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n461), .A2(KEYINPUT35), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n379), .B1(new_n351), .B2(new_n220), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n384), .B1(new_n471), .B2(new_n395), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT85), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(KEYINPUT85), .B(new_n384), .C1(new_n471), .C2(new_n395), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n378), .B(new_n244), .C1(new_n380), .C2(new_n382), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n474), .A2(new_n475), .A3(new_n476), .ZN(new_n477));
  AOI21_X1  g276(.A(KEYINPUT38), .B1(new_n477), .B2(KEYINPUT37), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT37), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n392), .A2(new_n479), .ZN(new_n480));
  OAI211_X1 g279(.A(KEYINPUT86), .B(new_n478), .C1(new_n413), .C2(new_n480), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n478), .B(new_n406), .C1(new_n405), .C2(KEYINPUT37), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n457), .A2(new_n459), .A3(new_n410), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n481), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT87), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n481), .A2(new_n484), .A3(new_n485), .A4(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT38), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n407), .B1(new_n479), .B2(new_n392), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n405), .A2(KEYINPUT37), .ZN(new_n492));
  AOI21_X1  g291(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n487), .A2(new_n489), .A3(new_n494), .ZN(new_n495));
  AOI21_X1  g294(.A(new_n422), .B1(new_n449), .B2(new_n421), .ZN(new_n496));
  OAI21_X1  g295(.A(KEYINPUT39), .B1(new_n438), .B2(new_n423), .ZN(new_n497));
  OR2_X1    g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT39), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n454), .B1(new_n496), .B2(new_n499), .ZN(new_n500));
  AND2_X1   g299(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n501), .A2(KEYINPUT40), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(KEYINPUT40), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n465), .A2(new_n502), .A3(new_n455), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n276), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g305(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n495), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n414), .A2(new_n408), .A3(new_n460), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n509), .A2(new_n276), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT36), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n463), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n462), .A2(KEYINPUT36), .A3(new_n372), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n510), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n470), .B1(new_n508), .B2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G43gat), .B(G50gat), .ZN(new_n518));
  AOI22_X1  g317(.A1(new_n518), .A2(KEYINPUT15), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT14), .ZN(new_n520));
  INV_X1    g319(.A(G29gat), .ZN(new_n521));
  INV_X1    g320(.A(G36gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g322(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT15), .ZN(new_n526));
  INV_X1    g325(.A(G43gat), .ZN(new_n527));
  AND2_X1   g326(.A1(new_n527), .A2(G50gat), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n527), .A2(G50gat), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n526), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n519), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n524), .A2(KEYINPUT88), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT88), .ZN(new_n533));
  OAI211_X1 g332(.A(new_n533), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n532), .A2(new_n534), .A3(new_n523), .ZN(new_n535));
  NAND2_X1  g334(.A1(G29gat), .A2(G36gat), .ZN(new_n536));
  AND2_X1   g335(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n518), .A2(KEYINPUT15), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n531), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(G1gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT16), .ZN(new_n541));
  OR2_X1    g340(.A1(G15gat), .A2(G22gat), .ZN(new_n542));
  NAND2_X1  g341(.A1(G15gat), .A2(G22gat), .ZN(new_n543));
  AOI21_X1  g342(.A(new_n541), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n546));
  OR2_X1    g345(.A1(KEYINPUT90), .A2(G8gat), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n542), .A2(G1gat), .A3(new_n543), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .A4(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n548), .ZN(new_n550));
  OAI211_X1 g349(.A(KEYINPUT90), .B(G8gat), .C1(new_n550), .C2(new_n544), .ZN(new_n551));
  NAND4_X1  g350(.A1(new_n539), .A2(KEYINPUT91), .A3(new_n549), .A4(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n535), .A2(new_n536), .ZN(new_n554));
  INV_X1    g353(.A(new_n538), .ZN(new_n555));
  XOR2_X1   g354(.A(G43gat), .B(G50gat), .Z(new_n556));
  AOI22_X1  g355(.A1(new_n556), .A2(new_n526), .B1(new_n524), .B2(new_n523), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n554), .A2(new_n555), .B1(new_n557), .B2(new_n519), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n549), .A2(new_n551), .ZN(new_n559));
  OAI21_X1  g358(.A(new_n553), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n552), .A2(new_n560), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n561), .A2(KEYINPUT92), .B1(new_n558), .B2(new_n559), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n552), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  XOR2_X1   g365(.A(new_n566), .B(KEYINPUT13), .Z(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(G113gat), .B(G141gat), .ZN(new_n569));
  XNOR2_X1  g368(.A(new_n569), .B(G197gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT11), .B(G169gat), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n570), .B(new_n571), .Z(new_n572));
  XOR2_X1   g371(.A(new_n572), .B(KEYINPUT12), .Z(new_n573));
  INV_X1    g372(.A(new_n573), .ZN(new_n574));
  XNOR2_X1  g373(.A(KEYINPUT89), .B(KEYINPUT17), .ZN(new_n575));
  AND4_X1   g374(.A1(new_n538), .A2(new_n530), .A3(new_n536), .A4(new_n525), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n538), .B1(new_n535), .B2(new_n536), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n575), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n531), .B(KEYINPUT17), .C1(new_n537), .C2(new_n538), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(new_n579), .A3(new_n559), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n566), .A3(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT18), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n561), .A2(KEYINPUT18), .A3(new_n566), .A4(new_n580), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n568), .A2(new_n574), .A3(new_n583), .A4(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n583), .A2(new_n584), .ZN(new_n586));
  INV_X1    g385(.A(new_n567), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n587), .B1(new_n562), .B2(new_n564), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n573), .B1(new_n586), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n585), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n517), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n593), .B(new_n205), .ZN(new_n594));
  XNOR2_X1  g393(.A(G183gat), .B(G211gat), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n594), .B(new_n595), .Z(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(G71gat), .ZN(new_n598));
  INV_X1    g397(.A(G78gat), .ZN(new_n599));
  OAI21_X1  g398(.A(KEYINPUT93), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OR2_X1    g399(.A1(G57gat), .A2(G64gat), .ZN(new_n601));
  NAND2_X1  g400(.A1(G57gat), .A2(G64gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n600), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(G71gat), .B(G78gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n598), .A2(new_n599), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n601), .B(new_n602), .C1(new_n609), .C2(KEYINPUT9), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n610), .B2(new_n600), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT21), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n559), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n617), .A2(new_n289), .ZN(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(new_n617), .A2(new_n289), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n614), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  INV_X1    g421(.A(new_n614), .ZN(new_n623));
  NOR3_X1   g422(.A1(new_n622), .A2(new_n623), .A3(new_n618), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n597), .B1(new_n621), .B2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n622), .B2(new_n618), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n619), .A2(new_n614), .A3(new_n620), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n627), .A3(new_n596), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n625), .A2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n629), .ZN(new_n630));
  XOR2_X1   g429(.A(G134gat), .B(G162gat), .Z(new_n631));
  AND2_X1   g430(.A1(G232gat), .A2(G233gat), .ZN(new_n632));
  NOR2_X1   g431(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT96), .ZN(new_n635));
  INV_X1    g434(.A(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT95), .ZN(new_n637));
  NAND2_X1  g436(.A1(G85gat), .A2(G92gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT7), .ZN(new_n639));
  XNOR2_X1  g438(.A(G99gat), .B(G106gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(G99gat), .A2(G106gat), .ZN(new_n641));
  INV_X1    g440(.A(G85gat), .ZN(new_n642));
  INV_X1    g441(.A(G92gat), .ZN(new_n643));
  AOI22_X1  g442(.A1(KEYINPUT8), .A2(new_n641), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  AND3_X1   g443(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n640), .B1(new_n639), .B2(new_n644), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n539), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n632), .A2(KEYINPUT41), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n637), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n649), .ZN(new_n651));
  AOI211_X1 g450(.A(KEYINPUT95), .B(new_n651), .C1(new_n539), .C2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n639), .A2(new_n644), .ZN(new_n653));
  INV_X1    g452(.A(new_n640), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n644), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n578), .A2(new_n579), .A3(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT94), .ZN(new_n659));
  OAI22_X1  g458(.A1(new_n650), .A2(new_n652), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n658), .A2(new_n659), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(G190gat), .B(G218gat), .Z(new_n663));
  NOR3_X1   g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n663), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n637), .A3(new_n649), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n649), .B1(new_n558), .B2(new_n657), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(KEYINPUT95), .ZN(new_n668));
  AND3_X1   g467(.A1(new_n578), .A2(new_n579), .A3(new_n657), .ZN(new_n669));
  AOI22_X1  g468(.A1(new_n666), .A2(new_n668), .B1(new_n669), .B2(KEYINPUT94), .ZN(new_n670));
  AOI21_X1  g469(.A(new_n665), .B1(new_n670), .B2(new_n661), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n636), .B1(new_n664), .B2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n663), .B1(new_n660), .B2(new_n662), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n670), .A2(new_n661), .A3(new_n665), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n634), .A2(KEYINPUT96), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n630), .A2(new_n678), .ZN(new_n679));
  OAI211_X1 g478(.A(new_n655), .B(new_n656), .C1(new_n608), .C2(new_n611), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n605), .A2(new_n607), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n610), .A2(new_n606), .A3(new_n600), .ZN(new_n682));
  OAI211_X1 g481(.A(new_n681), .B(new_n682), .C1(new_n645), .C2(new_n646), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT10), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n680), .A2(new_n683), .A3(new_n684), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n647), .B(KEYINPUT10), .C1(new_n611), .C2(new_n608), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(G230gat), .A2(G233gat), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n680), .A2(new_n683), .ZN(new_n690));
  INV_X1    g489(.A(new_n688), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(G120gat), .B(G148gat), .ZN(new_n694));
  XNOR2_X1  g493(.A(G176gat), .B(G204gat), .ZN(new_n695));
  XOR2_X1   g494(.A(new_n694), .B(new_n695), .Z(new_n696));
  INV_X1    g495(.A(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n693), .A2(new_n697), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n689), .A2(new_n692), .A3(new_n696), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n592), .A2(new_n679), .A3(new_n701), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n467), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(new_n540), .ZN(G1324gat));
  INV_X1    g503(.A(new_n702), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n705), .A2(new_n465), .ZN(new_n706));
  AND2_X1   g505(.A1(new_n706), .A2(G8gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(KEYINPUT16), .B(G8gat), .ZN(new_n708));
  NOR2_X1   g507(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(KEYINPUT42), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n710), .B1(KEYINPUT42), .B2(new_n709), .ZN(G1325gat));
  INV_X1    g510(.A(new_n463), .ZN(new_n712));
  AOI21_X1  g511(.A(G15gat), .B1(new_n705), .B2(new_n712), .ZN(new_n713));
  INV_X1    g512(.A(new_n514), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n714), .A2(G15gat), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT97), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n713), .B1(new_n705), .B2(new_n716), .ZN(G1326gat));
  NOR2_X1   g516(.A1(new_n702), .A2(new_n505), .ZN(new_n718));
  XOR2_X1   g517(.A(KEYINPUT43), .B(G22gat), .Z(new_n719));
  XNOR2_X1  g518(.A(new_n718), .B(new_n719), .ZN(G1327gat));
  NAND2_X1  g519(.A1(new_n461), .A2(KEYINPUT35), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n469), .A2(new_n466), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n493), .B1(new_n486), .B2(KEYINPUT87), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n506), .B1(new_n724), .B2(new_n489), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n723), .B1(new_n725), .B2(new_n515), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n630), .A2(new_n701), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n677), .ZN(new_n728));
  XNOR2_X1  g527(.A(new_n728), .B(KEYINPUT98), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n726), .A2(new_n590), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n731), .A2(new_n521), .A3(new_n468), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT45), .ZN(new_n733));
  OAI21_X1  g532(.A(KEYINPUT44), .B1(new_n517), .B2(new_n677), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT44), .ZN(new_n735));
  AND3_X1   g534(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n736));
  AOI21_X1  g535(.A(new_n635), .B1(new_n673), .B2(new_n674), .ZN(new_n737));
  OAI21_X1  g536(.A(KEYINPUT99), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT99), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n672), .A2(new_n739), .A3(new_n676), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n738), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n726), .A2(new_n735), .A3(new_n741), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n734), .A2(new_n742), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n591), .ZN(new_n744));
  AND2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n745), .A2(new_n468), .ZN(new_n746));
  INV_X1    g545(.A(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n733), .B1(new_n747), .B2(new_n521), .ZN(G1328gat));
  INV_X1    g547(.A(new_n465), .ZN(new_n749));
  NOR3_X1   g548(.A1(new_n730), .A2(G36gat), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT46), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n745), .A2(new_n465), .ZN(new_n752));
  INV_X1    g551(.A(KEYINPUT100), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(G36gat), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n752), .A2(new_n753), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n751), .B1(new_n755), .B2(new_n756), .ZN(G1329gat));
  NAND3_X1  g556(.A1(new_n745), .A2(G43gat), .A3(new_n714), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n527), .B1(new_n730), .B2(new_n463), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT47), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT47), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n762), .A3(new_n759), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1330gat));
  NAND3_X1  g563(.A1(new_n743), .A2(new_n276), .A3(new_n744), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT101), .ZN(new_n766));
  AOI211_X1 g565(.A(G50gat), .B(new_n505), .C1(new_n730), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n731), .A2(KEYINPUT101), .ZN(new_n768));
  AOI22_X1  g567(.A1(new_n765), .A2(G50gat), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT102), .B1(new_n765), .B2(G50gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT48), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n765), .A2(G50gat), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n767), .A2(new_n768), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT102), .ZN(new_n775));
  OAI211_X1 g574(.A(new_n773), .B(new_n774), .C1(new_n775), .C2(new_n771), .ZN(new_n776));
  INV_X1    g575(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n772), .A2(new_n777), .ZN(G1331gat));
  NAND3_X1  g577(.A1(new_n679), .A2(new_n591), .A3(new_n700), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n517), .A2(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(new_n468), .ZN(new_n781));
  XNOR2_X1  g580(.A(new_n781), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n465), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n783), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT49), .B(G64gat), .Z(new_n785));
  OAI21_X1  g584(.A(new_n784), .B1(new_n783), .B2(new_n785), .ZN(G1333gat));
  XNOR2_X1  g585(.A(new_n463), .B(KEYINPUT103), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n780), .A2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT104), .ZN(new_n789));
  AOI21_X1  g588(.A(G71gat), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n789), .B2(new_n788), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n780), .A2(G71gat), .A3(new_n714), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  XNOR2_X1  g592(.A(new_n793), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n276), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g595(.A1(new_n629), .A2(new_n590), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n515), .B1(new_n495), .B2(new_n507), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n678), .B(new_n797), .C1(new_n798), .C2(new_n470), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT51), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND4_X1  g600(.A1(new_n726), .A2(KEYINPUT51), .A3(new_n678), .A4(new_n797), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XOR2_X1   g602(.A(new_n803), .B(KEYINPUT105), .Z(new_n804));
  NOR3_X1   g603(.A1(new_n467), .A2(G85gat), .A3(new_n701), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT106), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n797), .A2(new_n700), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n743), .A2(new_n809), .ZN(new_n810));
  OAI21_X1  g609(.A(G85gat), .B1(new_n810), .B2(new_n467), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n807), .A2(new_n811), .ZN(G1336gat));
  OAI21_X1  g611(.A(G92gat), .B1(new_n810), .B2(new_n749), .ZN(new_n813));
  NAND4_X1  g612(.A1(new_n803), .A2(new_n643), .A3(new_n465), .A4(new_n700), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g614(.A(new_n815), .B(KEYINPUT52), .ZN(G1337gat));
  NOR3_X1   g615(.A1(new_n463), .A2(G99gat), .A3(new_n701), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n804), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G99gat), .B1(new_n810), .B2(new_n514), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(G1338gat));
  INV_X1    g619(.A(KEYINPUT108), .ZN(new_n821));
  AOI21_X1  g620(.A(new_n735), .B1(new_n726), .B2(new_n678), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n741), .A2(new_n735), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n508), .A2(new_n516), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n723), .ZN(new_n825));
  OAI211_X1 g624(.A(new_n276), .B(new_n809), .C1(new_n822), .C2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n505), .A2(G106gat), .A3(new_n701), .ZN(new_n827));
  XNOR2_X1  g626(.A(new_n827), .B(KEYINPUT107), .ZN(new_n828));
  AOI22_X1  g627(.A1(new_n826), .A2(G106gat), .B1(new_n803), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n821), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  INV_X1    g630(.A(G106gat), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n808), .B1(new_n734), .B2(new_n742), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n832), .B1(new_n833), .B2(new_n276), .ZN(new_n834));
  INV_X1    g633(.A(new_n828), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n835), .B1(new_n801), .B2(new_n802), .ZN(new_n836));
  OAI211_X1 g635(.A(KEYINPUT108), .B(KEYINPUT53), .C1(new_n834), .C2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n831), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n826), .A2(KEYINPUT110), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT110), .ZN(new_n840));
  NAND4_X1  g639(.A1(new_n743), .A2(new_n840), .A3(new_n276), .A4(new_n809), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n841), .A3(G106gat), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT111), .ZN(new_n843));
  XNOR2_X1  g642(.A(KEYINPUT109), .B(KEYINPUT53), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n844), .B1(new_n803), .B2(new_n827), .ZN(new_n845));
  AND3_X1   g644(.A1(new_n842), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n843), .B1(new_n842), .B2(new_n845), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n838), .B1(new_n846), .B2(new_n847), .ZN(G1339gat));
  NAND2_X1  g647(.A1(new_n561), .A2(KEYINPUT92), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n558), .A2(new_n559), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n849), .A2(new_n587), .A3(new_n564), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n561), .A2(new_n580), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(G229gat), .A3(G233gat), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n572), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT113), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  INV_X1    g656(.A(new_n572), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n858), .B1(new_n851), .B2(new_n853), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n859), .A2(KEYINPUT113), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n857), .A2(new_n585), .A3(new_n700), .A4(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n685), .A2(new_n686), .A3(new_n691), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n689), .A2(KEYINPUT54), .A3(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n691), .B1(new_n685), .B2(new_n686), .ZN(new_n864));
  INV_X1    g663(.A(KEYINPUT54), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n696), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n863), .A2(KEYINPUT55), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n699), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(KEYINPUT55), .B1(new_n863), .B2(new_n866), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT112), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  AOI211_X1 g671(.A(KEYINPUT112), .B(KEYINPUT55), .C1(new_n863), .C2(new_n866), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n869), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n861), .B1(new_n591), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n875), .A2(KEYINPUT115), .ZN(new_n876));
  NOR3_X1   g675(.A1(new_n736), .A2(new_n737), .A3(KEYINPUT99), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n739), .B1(new_n672), .B2(new_n676), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n861), .B(new_n880), .C1(new_n591), .C2(new_n874), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(KEYINPUT114), .ZN(new_n883));
  NOR2_X1   g682(.A1(new_n586), .A2(new_n588), .ZN(new_n884));
  AOI22_X1  g683(.A1(new_n884), .A2(new_n574), .B1(new_n859), .B2(KEYINPUT113), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT55), .ZN(new_n886));
  AND3_X1   g685(.A1(new_n685), .A2(new_n686), .A3(new_n691), .ZN(new_n887));
  NOR3_X1   g686(.A1(new_n887), .A2(new_n864), .A3(new_n865), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n687), .A2(new_n865), .A3(new_n688), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n889), .A2(new_n697), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n886), .B1(new_n888), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n870), .A2(new_n871), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n885), .A2(new_n894), .A3(new_n857), .A4(new_n869), .ZN(new_n895));
  OAI21_X1  g694(.A(new_n883), .B1(new_n879), .B2(new_n895), .ZN(new_n896));
  INV_X1    g695(.A(new_n874), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n857), .A2(new_n585), .A3(new_n860), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n741), .A2(new_n897), .A3(new_n898), .A4(KEYINPUT114), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n896), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n629), .B1(new_n882), .B2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n629), .A2(new_n677), .A3(new_n701), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n902), .A2(new_n590), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT116), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  INV_X1    g703(.A(new_n903), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT116), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n741), .B1(new_n875), .B2(KEYINPUT115), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n907), .A2(new_n881), .B1(new_n896), .B2(new_n899), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n905), .B(new_n906), .C1(new_n908), .C2(new_n629), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n904), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n910), .A2(new_n276), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(new_n468), .A3(new_n466), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n912), .A2(new_n590), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(G113gat), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT117), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT117), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n913), .A2(new_n916), .A3(G113gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n283), .A2(new_n285), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n915), .B(new_n917), .C1(new_n918), .C2(new_n913), .ZN(G1340gat));
  NAND2_X1  g718(.A1(new_n912), .A2(new_n700), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n920), .B1(new_n278), .B2(new_n280), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n277), .B2(new_n920), .ZN(G1341gat));
  NAND2_X1  g721(.A1(new_n912), .A2(new_n629), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n295), .A2(new_n297), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g724(.A(KEYINPUT118), .B1(new_n923), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n923), .A2(new_n925), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT118), .ZN(new_n928));
  NAND4_X1  g727(.A1(new_n912), .A2(new_n928), .A3(new_n924), .A4(new_n629), .ZN(new_n929));
  AND3_X1   g728(.A1(new_n926), .A2(new_n927), .A3(new_n929), .ZN(G1342gat));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n465), .A2(new_n677), .ZN(new_n932));
  NOR2_X1   g731(.A1(new_n463), .A2(G134gat), .ZN(new_n933));
  NAND4_X1  g732(.A1(new_n911), .A2(new_n468), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(new_n931), .B1(new_n934), .B2(KEYINPUT56), .ZN(new_n935));
  INV_X1    g734(.A(new_n932), .ZN(new_n936));
  NOR4_X1   g735(.A1(new_n910), .A2(new_n467), .A3(new_n276), .A4(new_n936), .ZN(new_n937));
  INV_X1    g736(.A(KEYINPUT56), .ZN(new_n938));
  NAND4_X1  g737(.A1(new_n937), .A2(KEYINPUT119), .A3(new_n938), .A4(new_n933), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n934), .A2(KEYINPUT56), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n911), .A2(new_n468), .A3(new_n712), .A4(new_n932), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G134gat), .ZN(new_n942));
  NAND4_X1  g741(.A1(new_n935), .A2(new_n939), .A3(new_n940), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n943), .A2(KEYINPUT120), .ZN(new_n944));
  AOI22_X1  g743(.A1(KEYINPUT56), .A2(new_n934), .B1(new_n941), .B2(G134gat), .ZN(new_n945));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n945), .A2(new_n946), .A3(new_n939), .A4(new_n935), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n944), .A2(new_n947), .ZN(G1343gat));
  NAND4_X1  g747(.A1(new_n514), .A2(new_n468), .A3(new_n276), .A4(new_n749), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n910), .A2(new_n949), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n950), .A2(new_n208), .A3(new_n590), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n904), .A2(new_n276), .A3(new_n909), .ZN(new_n952));
  INV_X1    g751(.A(KEYINPUT57), .ZN(new_n953));
  NAND2_X1  g752(.A1(new_n869), .A2(new_n891), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n861), .B1(new_n591), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n955), .A2(new_n677), .ZN(new_n956));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n900), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g758(.A1(new_n956), .A2(new_n957), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n630), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n961), .A2(new_n905), .ZN(new_n962));
  NOR2_X1   g761(.A1(new_n505), .A2(new_n953), .ZN(new_n963));
  AOI22_X1  g762(.A1(new_n952), .A2(new_n953), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n514), .A2(new_n468), .A3(new_n749), .ZN(new_n965));
  NOR3_X1   g764(.A1(new_n964), .A2(new_n591), .A3(new_n965), .ZN(new_n966));
  OAI21_X1  g765(.A(new_n951), .B1(new_n966), .B2(new_n208), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(KEYINPUT58), .ZN(G1344gat));
  NAND3_X1  g767(.A1(new_n950), .A2(new_n210), .A3(new_n700), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n964), .A2(new_n701), .A3(new_n965), .ZN(new_n970));
  NOR3_X1   g769(.A1(new_n970), .A2(KEYINPUT59), .A3(new_n210), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT59), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n904), .A2(new_n909), .A3(new_n963), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n903), .A2(KEYINPUT122), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT122), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n902), .B2(new_n590), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n956), .B1(new_n677), .B2(new_n895), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n977), .B1(new_n630), .B2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n953), .B1(new_n979), .B2(new_n505), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n973), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n701), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  AOI21_X1  g782(.A(new_n972), .B1(new_n983), .B2(G148gat), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n969), .B1(new_n971), .B2(new_n984), .ZN(G1345gat));
  NAND3_X1  g784(.A1(new_n950), .A2(new_n205), .A3(new_n629), .ZN(new_n986));
  NOR3_X1   g785(.A1(new_n964), .A2(new_n630), .A3(new_n965), .ZN(new_n987));
  OAI21_X1  g786(.A(new_n986), .B1(new_n987), .B2(new_n205), .ZN(G1346gat));
  NAND3_X1  g787(.A1(new_n950), .A2(new_n206), .A3(new_n678), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n964), .A2(new_n879), .A3(new_n965), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n989), .B1(new_n990), .B2(new_n206), .ZN(G1347gat));
  NOR2_X1   g790(.A1(new_n749), .A2(new_n468), .ZN(new_n992));
  NAND3_X1  g791(.A1(new_n911), .A2(new_n787), .A3(new_n992), .ZN(new_n993));
  INV_X1    g792(.A(G169gat), .ZN(new_n994));
  NOR3_X1   g793(.A1(new_n993), .A2(new_n994), .A3(new_n591), .ZN(new_n995));
  INV_X1    g794(.A(new_n992), .ZN(new_n996));
  NOR4_X1   g795(.A1(new_n910), .A2(new_n276), .A3(new_n463), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g796(.A(G169gat), .B1(new_n997), .B2(new_n590), .ZN(new_n998));
  NOR2_X1   g797(.A1(new_n995), .A2(new_n998), .ZN(G1348gat));
  OAI21_X1  g798(.A(G176gat), .B1(new_n993), .B2(new_n701), .ZN(new_n1000));
  INV_X1    g799(.A(G176gat), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n997), .A2(new_n1001), .A3(new_n700), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n1000), .A2(new_n1002), .ZN(G1349gat));
  OAI21_X1  g802(.A(G183gat), .B1(new_n993), .B2(new_n630), .ZN(new_n1004));
  NAND4_X1  g803(.A1(new_n997), .A2(new_n336), .A3(new_n338), .A4(new_n629), .ZN(new_n1005));
  NAND2_X1  g804(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  XNOR2_X1  g805(.A(new_n1006), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g806(.A1(new_n997), .A2(new_n309), .A3(new_n741), .ZN(new_n1008));
  INV_X1    g807(.A(KEYINPUT123), .ZN(new_n1009));
  XNOR2_X1  g808(.A(new_n1008), .B(new_n1009), .ZN(new_n1010));
  OAI21_X1  g809(.A(G190gat), .B1(new_n993), .B2(new_n677), .ZN(new_n1011));
  INV_X1    g810(.A(KEYINPUT61), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  OR2_X1    g812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  NAND3_X1  g813(.A1(new_n1010), .A2(new_n1013), .A3(new_n1014), .ZN(G1351gat));
  INV_X1    g814(.A(new_n952), .ZN(new_n1016));
  NOR2_X1   g815(.A1(new_n714), .A2(new_n996), .ZN(new_n1017));
  NAND2_X1  g816(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g817(.A(new_n1018), .ZN(new_n1019));
  AOI21_X1  g818(.A(G197gat), .B1(new_n1019), .B2(new_n590), .ZN(new_n1020));
  INV_X1    g819(.A(new_n1017), .ZN(new_n1021));
  AOI21_X1  g820(.A(new_n1021), .B1(new_n973), .B2(new_n980), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(G197gat), .A3(new_n590), .ZN(new_n1023));
  NOR2_X1   g822(.A1(new_n1020), .A2(new_n1023), .ZN(G1352gat));
  XOR2_X1   g823(.A(KEYINPUT124), .B(G204gat), .Z(new_n1025));
  NAND2_X1  g824(.A1(new_n700), .A2(new_n1025), .ZN(new_n1026));
  OR3_X1    g825(.A1(new_n1018), .A2(KEYINPUT62), .A3(new_n1026), .ZN(new_n1027));
  INV_X1    g826(.A(new_n1025), .ZN(new_n1028));
  INV_X1    g827(.A(new_n1022), .ZN(new_n1029));
  OAI21_X1  g828(.A(new_n1028), .B1(new_n1029), .B2(new_n701), .ZN(new_n1030));
  OAI21_X1  g829(.A(KEYINPUT62), .B1(new_n1018), .B2(new_n1026), .ZN(new_n1031));
  NAND3_X1  g830(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .ZN(new_n1032));
  NAND2_X1  g831(.A1(new_n1032), .A2(KEYINPUT125), .ZN(new_n1033));
  INV_X1    g832(.A(KEYINPUT125), .ZN(new_n1034));
  NAND4_X1  g833(.A1(new_n1027), .A2(new_n1030), .A3(new_n1034), .A4(new_n1031), .ZN(new_n1035));
  NAND2_X1  g834(.A1(new_n1033), .A2(new_n1035), .ZN(G1353gat));
  NAND3_X1  g835(.A1(new_n1019), .A2(new_n223), .A3(new_n629), .ZN(new_n1037));
  INV_X1    g836(.A(KEYINPUT63), .ZN(new_n1038));
  AOI21_X1  g837(.A(new_n223), .B1(KEYINPUT126), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g838(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g839(.A1(new_n1038), .A2(KEYINPUT126), .ZN(new_n1041));
  INV_X1    g840(.A(new_n1041), .ZN(new_n1042));
  AOI211_X1 g841(.A(new_n1040), .B(new_n1042), .C1(new_n1022), .C2(new_n629), .ZN(new_n1043));
  NAND3_X1  g842(.A1(new_n981), .A2(new_n629), .A3(new_n1017), .ZN(new_n1044));
  AOI21_X1  g843(.A(new_n1041), .B1(new_n1044), .B2(new_n1039), .ZN(new_n1045));
  OAI21_X1  g844(.A(new_n1037), .B1(new_n1043), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g845(.A(KEYINPUT127), .ZN(new_n1047));
  NAND2_X1  g846(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  OAI211_X1 g847(.A(KEYINPUT127), .B(new_n1037), .C1(new_n1043), .C2(new_n1045), .ZN(new_n1049));
  NAND2_X1  g848(.A1(new_n1048), .A2(new_n1049), .ZN(G1354gat));
  NAND3_X1  g849(.A1(new_n1019), .A2(new_n224), .A3(new_n741), .ZN(new_n1051));
  OAI21_X1  g850(.A(G218gat), .B1(new_n1029), .B2(new_n677), .ZN(new_n1052));
  NAND2_X1  g851(.A1(new_n1051), .A2(new_n1052), .ZN(G1355gat));
endmodule


