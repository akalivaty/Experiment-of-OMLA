//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 0 0 0 1 1 1 1 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:59 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n207, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1265, new_n1266,
    new_n1267, new_n1268, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1336, new_n1337, new_n1338, new_n1339, new_n1340, new_n1341,
    new_n1342, new_n1343, new_n1344;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(new_n205));
  XOR2_X1   g0005(.A(new_n205), .B(KEYINPUT64), .Z(G353));
  NOR2_X1   g0006(.A1(G97), .A2(G107), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n208), .A2(G87), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  INV_X1    g0012(.A(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n202), .A2(new_n203), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  INV_X1    g0015(.A(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(new_n212), .A2(new_n213), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G77), .A2(G244), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G50), .A2(G226), .B1(G107), .B2(G264), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G58), .A2(G232), .B1(G68), .B2(G238), .ZN(new_n225));
  NAND3_X1  g0025(.A1(new_n223), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI221_X1 g0027(.A(new_n220), .B1(new_n213), .B2(new_n212), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G226), .ZN(new_n232));
  XOR2_X1   g0032(.A(new_n232), .B(G232), .Z(new_n233));
  XOR2_X1   g0033(.A(new_n233), .B(KEYINPUT66), .Z(new_n234));
  XOR2_X1   g0034(.A(G250), .B(G257), .Z(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G68), .B(G77), .Z(new_n239));
  XNOR2_X1  g0039(.A(G50), .B(G58), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NOR2_X1   g0045(.A1(G20), .A2(G33), .ZN(new_n246));
  AOI22_X1  g0046(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n218), .A2(G33), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT8), .B(G58), .ZN(new_n249));
  OAI21_X1  g0049(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n217), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G1), .ZN(new_n254));
  NAND3_X1  g0054(.A1(new_n254), .A2(G13), .A3(G20), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(new_n201), .ZN(new_n256));
  AOI21_X1  g0056(.A(new_n252), .B1(new_n254), .B2(G20), .ZN(new_n257));
  OAI21_X1  g0057(.A(new_n256), .B1(new_n257), .B2(new_n201), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n253), .A2(new_n258), .ZN(new_n259));
  OR2_X1    g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NAND2_X1  g0060(.A1(KEYINPUT3), .A2(G33), .ZN(new_n261));
  AOI21_X1  g0061(.A(G1698), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AND2_X1   g0062(.A1(KEYINPUT3), .A2(G33), .ZN(new_n263));
  NOR2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n262), .A2(G222), .B1(new_n265), .B2(G77), .ZN(new_n266));
  INV_X1    g0066(.A(G223), .ZN(new_n267));
  INV_X1    g0067(.A(G1698), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n260), .B2(new_n261), .ZN(new_n269));
  INV_X1    g0069(.A(new_n269), .ZN(new_n270));
  OAI21_X1  g0070(.A(new_n266), .B1(new_n267), .B2(new_n270), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OAI211_X1 g0073(.A(new_n254), .B(G274), .C1(G41), .C2(G45), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT67), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g0076(.A(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G45), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g0079(.A1(new_n279), .A2(KEYINPUT67), .A3(new_n254), .A4(G274), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n276), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n217), .ZN(new_n282));
  NAND2_X1  g0082(.A1(G33), .A2(G41), .ZN(new_n283));
  AOI22_X1  g0083(.A1(new_n254), .A2(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT68), .B(G226), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n281), .B1(new_n284), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n273), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(G179), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G169), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n290), .B1(new_n273), .B2(new_n286), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n259), .B1(new_n289), .B2(new_n291), .ZN(new_n292));
  XNOR2_X1  g0092(.A(new_n292), .B(KEYINPUT69), .ZN(new_n293));
  INV_X1    g0093(.A(new_n293), .ZN(new_n294));
  XOR2_X1   g0094(.A(KEYINPUT8), .B(G58), .Z(new_n295));
  AND2_X1   g0095(.A1(new_n246), .A2(KEYINPUT70), .ZN(new_n296));
  NOR2_X1   g0096(.A1(new_n246), .A2(KEYINPUT70), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n295), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G77), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT15), .B(G87), .ZN(new_n300));
  OAI221_X1 g0100(.A(new_n298), .B1(new_n218), .B2(new_n299), .C1(new_n248), .C2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n252), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n255), .A2(G77), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(new_n257), .B2(G77), .ZN(new_n304));
  AND2_X1   g0104(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n262), .A2(G232), .B1(new_n265), .B2(G107), .ZN(new_n306));
  INV_X1    g0106(.A(G238), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n270), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(new_n272), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n281), .B1(G244), .B2(new_n284), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(new_n288), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(G169), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n305), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  XNOR2_X1  g0115(.A(new_n259), .B(KEYINPUT9), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n287), .A2(G200), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n273), .A2(G190), .A3(new_n286), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  OR2_X1    g0119(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(KEYINPUT10), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n315), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n311), .ZN(new_n323));
  INV_X1    g0123(.A(G200), .ZN(new_n324));
  OAI211_X1 g0124(.A(new_n305), .B(KEYINPUT71), .C1(new_n323), .C2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT71), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n324), .B1(new_n309), .B2(new_n310), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n302), .A2(new_n304), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n323), .A2(G190), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n325), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND3_X1   g0131(.A1(new_n294), .A2(new_n322), .A3(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(G33), .A2(G97), .ZN(new_n333));
  OAI211_X1 g0133(.A(G232), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n334));
  OAI211_X1 g0134(.A(G226), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n335));
  OAI211_X1 g0135(.A(new_n333), .B(new_n334), .C1(new_n335), .C2(KEYINPUT72), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT72), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n337), .B1(new_n262), .B2(G226), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n272), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT13), .ZN(new_n340));
  AOI22_X1  g0140(.A1(new_n284), .A2(G238), .B1(new_n276), .B2(new_n280), .ZN(new_n341));
  AND3_X1   g0141(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n340), .B1(new_n339), .B2(new_n341), .ZN(new_n343));
  OAI21_X1  g0143(.A(G169), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(KEYINPUT14), .ZN(new_n345));
  INV_X1    g0145(.A(KEYINPUT14), .ZN(new_n346));
  OAI211_X1 g0146(.A(new_n346), .B(G169), .C1(new_n342), .C2(new_n343), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n339), .A2(new_n341), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(KEYINPUT13), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n339), .A2(new_n340), .A3(new_n341), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n349), .A2(G179), .A3(new_n350), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n345), .A2(new_n347), .A3(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(G13), .ZN(new_n353));
  NOR2_X1   g0153(.A1(new_n353), .A2(G1), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n354), .A2(G20), .A3(new_n203), .ZN(new_n355));
  XNOR2_X1  g0155(.A(new_n355), .B(KEYINPUT12), .ZN(new_n356));
  INV_X1    g0156(.A(new_n257), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n248), .A2(new_n299), .B1(new_n218), .B2(G68), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT73), .ZN(new_n359));
  AND2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n246), .A2(G50), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n361), .B1(new_n358), .B2(new_n359), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n252), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT11), .ZN(new_n364));
  OAI221_X1 g0164(.A(new_n356), .B1(new_n203), .B2(new_n357), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n363), .A2(new_n364), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n352), .A2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n349), .A2(new_n350), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n370), .A2(G190), .ZN(new_n371));
  AOI21_X1  g0171(.A(G200), .B1(new_n349), .B2(new_n350), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n367), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AND2_X1   g0173(.A1(new_n369), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g0174(.A(G223), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n375));
  OAI211_X1 g0175(.A(G226), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n376));
  NAND2_X1  g0176(.A1(G33), .A2(G87), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n378), .A2(new_n272), .ZN(new_n379));
  AOI22_X1  g0179(.A1(new_n284), .A2(G232), .B1(new_n276), .B2(new_n280), .ZN(new_n380));
  AOI21_X1  g0180(.A(G200), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n379), .A2(new_n380), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(G190), .ZN(new_n384));
  INV_X1    g0184(.A(new_n383), .ZN(new_n385));
  INV_X1    g0185(.A(G190), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n385), .A2(KEYINPUT76), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n255), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n295), .A2(new_n389), .ZN(new_n390));
  AOI21_X1  g0190(.A(new_n390), .B1(new_n357), .B2(new_n295), .ZN(new_n391));
  NAND2_X1  g0191(.A1(G58), .A2(G68), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT75), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND3_X1  g0194(.A1(KEYINPUT75), .A2(G58), .A3(G68), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n394), .A2(new_n214), .A3(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(G20), .B1(G159), .B2(new_n246), .ZN(new_n397));
  NOR3_X1   g0197(.A1(new_n263), .A2(new_n264), .A3(G20), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(G68), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT74), .B(KEYINPUT7), .ZN(new_n401));
  AND3_X1   g0201(.A1(new_n265), .A2(new_n401), .A3(new_n218), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT16), .B(new_n397), .C1(new_n400), .C2(new_n402), .ZN(new_n403));
  AND2_X1   g0203(.A1(new_n403), .A2(new_n252), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n260), .A2(new_n399), .A3(new_n218), .A4(new_n261), .ZN(new_n405));
  OAI211_X1 g0205(.A(G68), .B(new_n405), .C1(new_n398), .C2(new_n401), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT16), .B1(new_n406), .B2(new_n397), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n391), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT17), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n410), .A2(KEYINPUT77), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n388), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  INV_X1    g0212(.A(new_n391), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n403), .A2(new_n252), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n407), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n415), .B1(new_n387), .B2(new_n384), .ZN(new_n416));
  XOR2_X1   g0216(.A(KEYINPUT77), .B(KEYINPUT17), .Z(new_n417));
  OAI21_X1  g0217(.A(new_n412), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(G169), .B1(new_n379), .B2(new_n380), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n385), .B2(new_n288), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n415), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n421), .A2(KEYINPUT18), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT18), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n415), .A2(new_n420), .A3(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n418), .A2(new_n425), .ZN(new_n426));
  AND3_X1   g0226(.A1(new_n332), .A2(new_n374), .A3(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n218), .B(G87), .C1(new_n263), .C2(new_n264), .ZN(new_n429));
  OR2_X1    g0229(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(KEYINPUT84), .A2(KEYINPUT22), .ZN(new_n432));
  XOR2_X1   g0232(.A(new_n432), .B(KEYINPUT85), .Z(new_n433));
  NAND2_X1  g0233(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT24), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n432), .B(KEYINPUT85), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n436), .A2(new_n429), .A3(new_n430), .ZN(new_n437));
  OR3_X1    g0237(.A1(new_n218), .A2(KEYINPUT23), .A3(G107), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n218), .A2(G33), .A3(G116), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT23), .B1(new_n218), .B2(G107), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  INV_X1    g0241(.A(new_n441), .ZN(new_n442));
  NAND4_X1  g0242(.A1(new_n434), .A2(new_n435), .A3(new_n437), .A4(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n443), .A2(KEYINPUT86), .ZN(new_n444));
  AOI21_X1  g0244(.A(new_n441), .B1(new_n431), .B2(new_n433), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT86), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n435), .A4(new_n437), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n434), .A2(new_n437), .A3(new_n442), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT24), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n252), .ZN(new_n451));
  INV_X1    g0251(.A(G107), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n354), .A2(G20), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT25), .ZN(new_n454));
  OR3_X1    g0254(.A1(new_n453), .A2(KEYINPUT87), .A3(new_n454), .ZN(new_n455));
  OAI21_X1  g0255(.A(KEYINPUT87), .B1(new_n453), .B2(new_n454), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n453), .A2(new_n454), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n455), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n254), .A2(G33), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n255), .A2(new_n459), .A3(new_n217), .A4(new_n251), .ZN(new_n460));
  INV_X1    g0260(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G107), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n458), .A2(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(G257), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G294), .ZN(new_n467));
  OAI21_X1  g0267(.A(G250), .B1(new_n263), .B2(new_n264), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n272), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n254), .A2(G45), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT5), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n472), .A2(new_n277), .ZN(new_n473));
  NAND2_X1  g0273(.A1(KEYINPUT5), .A2(G41), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n471), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n475), .A2(new_n272), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(G264), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n475), .A2(G274), .ZN(new_n478));
  NAND3_X1  g0278(.A1(new_n470), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(KEYINPUT88), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n469), .A2(new_n272), .B1(new_n476), .B2(G264), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT88), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n481), .A2(new_n482), .A3(new_n478), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n480), .A2(G169), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n481), .A2(G179), .A3(new_n478), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n465), .A2(new_n486), .ZN(new_n487));
  AND4_X1   g0287(.A1(new_n482), .A2(new_n470), .A3(new_n477), .A4(new_n478), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n482), .B1(new_n481), .B2(new_n478), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n386), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n479), .A2(new_n324), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n463), .B1(new_n450), .B2(new_n252), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n487), .A2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n255), .A2(new_n459), .ZN(new_n496));
  INV_X1    g0296(.A(new_n252), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n496), .A2(KEYINPUT83), .A3(new_n497), .A4(G116), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  INV_X1    g0299(.A(G116), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n460), .B2(new_n500), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n498), .A2(new_n501), .B1(new_n500), .B2(new_n389), .ZN(new_n502));
  INV_X1    g0302(.A(G33), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n503), .A2(G97), .ZN(new_n504));
  NAND2_X1  g0304(.A1(G33), .A2(G283), .ZN(new_n505));
  AOI21_X1  g0305(.A(G20), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(new_n218), .A2(new_n500), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n252), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT20), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  OAI211_X1 g0310(.A(KEYINPUT20), .B(new_n252), .C1(new_n506), .C2(new_n507), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n502), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  OAI211_X1 g0314(.A(G257), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n260), .A2(G303), .A3(new_n261), .ZN(new_n516));
  OAI211_X1 g0316(.A(G264), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT82), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n515), .B(new_n516), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  AOI21_X1  g0319(.A(KEYINPUT82), .B1(new_n269), .B2(G264), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n272), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NOR2_X1   g0321(.A1(new_n278), .A2(G1), .ZN(new_n522));
  INV_X1    g0322(.A(new_n474), .ZN(new_n523));
  NOR2_X1   g0323(.A1(KEYINPUT5), .A2(G41), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n282), .A2(new_n283), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n525), .A2(G270), .A3(new_n526), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(new_n478), .ZN(new_n528));
  INV_X1    g0328(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n521), .A2(new_n529), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n530), .A2(KEYINPUT21), .A3(G169), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n269), .A2(KEYINPUT82), .A3(G264), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n517), .A2(new_n518), .ZN(new_n533));
  NAND4_X1  g0333(.A1(new_n532), .A2(new_n533), .A3(new_n515), .A4(new_n516), .ZN(new_n534));
  AOI21_X1  g0334(.A(new_n528), .B1(new_n534), .B2(new_n272), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n535), .A2(G179), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n514), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n530), .A2(new_n324), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n386), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n513), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n290), .B1(new_n521), .B2(new_n529), .ZN(new_n541));
  AOI21_X1  g0341(.A(KEYINPUT21), .B1(new_n541), .B2(new_n513), .ZN(new_n542));
  NOR3_X1   g0342(.A1(new_n537), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G238), .B(new_n268), .C1(new_n263), .C2(new_n264), .ZN(new_n544));
  OAI211_X1 g0344(.A(G244), .B(G1698), .C1(new_n263), .C2(new_n264), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n272), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n471), .A2(G250), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n254), .A2(G45), .A3(G274), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n549), .A2(new_n550), .B1(new_n282), .B2(new_n283), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT80), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n548), .A2(KEYINPUT80), .A3(new_n552), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n555), .A2(new_n288), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(KEYINPUT80), .B1(new_n548), .B2(new_n552), .ZN(new_n558));
  AOI211_X1 g0358(.A(new_n554), .B(new_n551), .C1(new_n547), .C2(new_n272), .ZN(new_n559));
  OAI21_X1  g0359(.A(new_n290), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n260), .A2(new_n261), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n561), .A2(new_n218), .A3(G68), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n218), .B1(new_n333), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(G87), .ZN(new_n565));
  INV_X1    g0365(.A(G97), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n564), .B1(G107), .B2(new_n567), .ZN(new_n568));
  OAI21_X1  g0368(.A(new_n563), .B1(new_n333), .B2(G20), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n562), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n252), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n300), .A2(new_n389), .ZN(new_n572));
  OAI211_X1 g0372(.A(new_n571), .B(new_n572), .C1(new_n300), .C2(new_n460), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n557), .A2(new_n560), .A3(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n555), .A2(G190), .A3(new_n556), .ZN(new_n575));
  OAI21_X1  g0375(.A(G200), .B1(new_n558), .B2(new_n559), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n460), .A2(new_n565), .ZN(new_n577));
  OR2_X1    g0377(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n577), .A2(KEYINPUT81), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n571), .A2(new_n578), .A3(new_n572), .A4(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n575), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g0381(.A1(new_n574), .A2(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT79), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT4), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n584), .A2(G1698), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n585), .B(G244), .C1(new_n264), .C2(new_n263), .ZN(new_n586));
  INV_X1    g0386(.A(G244), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n260), .B2(new_n261), .ZN(new_n588));
  OAI211_X1 g0388(.A(new_n586), .B(new_n505), .C1(new_n588), .C2(KEYINPUT4), .ZN(new_n589));
  AOI21_X1  g0389(.A(new_n268), .B1(new_n468), .B2(KEYINPUT4), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n272), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n525), .A2(G257), .A3(new_n526), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n478), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n583), .B1(new_n595), .B2(G179), .ZN(new_n596));
  INV_X1    g0396(.A(G250), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n260), .B2(new_n261), .ZN(new_n598));
  OAI21_X1  g0398(.A(G1698), .B1(new_n598), .B2(new_n584), .ZN(new_n599));
  OAI21_X1  g0399(.A(G244), .B1(new_n263), .B2(new_n264), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n600), .A2(new_n584), .B1(G33), .B2(G283), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n599), .A2(new_n601), .A3(new_n586), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n593), .B1(new_n602), .B2(new_n272), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(KEYINPUT79), .A3(new_n288), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n596), .A2(new_n604), .ZN(new_n605));
  OAI211_X1 g0405(.A(G107), .B(new_n405), .C1(new_n398), .C2(new_n401), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G97), .A2(G107), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  OAI22_X1  g0408(.A1(new_n608), .A2(new_n207), .B1(KEYINPUT78), .B2(KEYINPUT6), .ZN(new_n609));
  NOR2_X1   g0409(.A1(KEYINPUT78), .A2(KEYINPUT6), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n208), .A2(new_n607), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n566), .A2(KEYINPUT6), .ZN(new_n612));
  NAND4_X1  g0412(.A1(new_n609), .A2(new_n611), .A3(G20), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n246), .A2(G77), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n606), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n252), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n255), .A2(new_n566), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(new_n461), .B2(new_n566), .ZN(new_n618));
  AOI22_X1  g0418(.A1(new_n595), .A2(new_n290), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n615), .A2(new_n252), .ZN(new_n620));
  INV_X1    g0420(.A(new_n618), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n591), .A2(new_n386), .A3(new_n594), .ZN(new_n623));
  OAI21_X1  g0423(.A(new_n623), .B1(new_n603), .B2(G200), .ZN(new_n624));
  AOI22_X1  g0424(.A1(new_n605), .A2(new_n619), .B1(new_n622), .B2(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n543), .A2(new_n582), .A3(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n428), .A2(new_n495), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n627), .B(KEYINPUT89), .ZN(G372));
  AND2_X1   g0428(.A1(new_n422), .A2(new_n424), .ZN(new_n629));
  AND3_X1   g0429(.A1(new_n388), .A2(new_n409), .A3(new_n411), .ZN(new_n630));
  AOI21_X1  g0430(.A(new_n417), .B1(new_n388), .B2(new_n409), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n632), .A2(new_n373), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n315), .B1(new_n352), .B2(new_n368), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n320), .A2(new_n321), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI21_X1  g0437(.A(KEYINPUT91), .B1(new_n637), .B2(new_n294), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT91), .ZN(new_n639));
  AOI211_X1 g0439(.A(new_n639), .B(new_n293), .C1(new_n635), .C2(new_n636), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  AOI22_X1  g0441(.A1(new_n451), .A2(new_n464), .B1(new_n484), .B2(new_n485), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n537), .B2(new_n542), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n541), .A2(new_n513), .ZN(new_n645));
  INV_X1    g0445(.A(KEYINPUT21), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  AOI22_X1  g0447(.A1(new_n541), .A2(KEYINPUT21), .B1(new_n535), .B2(G179), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n647), .B(KEYINPUT90), .C1(new_n514), .C2(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n642), .B1(new_n644), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n553), .A2(new_n290), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n557), .A2(new_n573), .A3(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n553), .A2(G200), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n575), .A2(new_n580), .A3(new_n653), .ZN(new_n654));
  AND2_X1   g0454(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n494), .A3(new_n625), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n574), .A2(new_n581), .ZN(new_n658));
  AOI21_X1  g0458(.A(KEYINPUT79), .B1(new_n603), .B2(new_n288), .ZN(new_n659));
  AND4_X1   g0459(.A1(KEYINPUT79), .A2(new_n591), .A3(new_n288), .A4(new_n594), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n619), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  OAI21_X1  g0461(.A(KEYINPUT26), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  OAI22_X1  g0462(.A1(new_n620), .A2(new_n621), .B1(new_n603), .B2(G169), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n596), .B2(new_n604), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT26), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n664), .A2(new_n665), .A3(new_n652), .A4(new_n654), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n662), .A2(new_n666), .A3(new_n652), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n427), .B1(new_n657), .B2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n641), .A2(new_n668), .ZN(G369));
  NAND2_X1  g0469(.A1(new_n354), .A2(new_n218), .ZN(new_n670));
  OR2_X1    g0470(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(KEYINPUT27), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n671), .A2(G213), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(G343), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n514), .A2(new_n676), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n543), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n644), .A2(new_n649), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n677), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n678), .A2(new_n680), .A3(G330), .ZN(new_n681));
  INV_X1    g0481(.A(new_n681), .ZN(new_n682));
  AOI21_X1  g0482(.A(new_n642), .B1(new_n493), .B2(new_n492), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n465), .A2(new_n675), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n685), .B1(new_n487), .B2(new_n676), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n682), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n531), .A2(new_n536), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n542), .B1(new_n688), .B2(new_n513), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n689), .A2(new_n675), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n690), .A2(new_n487), .A3(new_n494), .A4(new_n684), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT92), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n642), .A2(new_n676), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n696));
  OAI21_X1  g0496(.A(new_n687), .B1(new_n695), .B2(new_n696), .ZN(G399));
  INV_X1    g0497(.A(new_n211), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n698), .A2(G41), .ZN(new_n699));
  INV_X1    g0499(.A(new_n699), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n567), .A2(G107), .A3(G116), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n700), .A2(G1), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g0502(.A(new_n702), .B1(new_n215), .B2(new_n700), .ZN(new_n703));
  XNOR2_X1  g0503(.A(new_n703), .B(KEYINPUT28), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n652), .A2(new_n654), .ZN(new_n705));
  OAI21_X1  g0505(.A(KEYINPUT26), .B1(new_n705), .B2(new_n661), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n664), .A2(new_n665), .A3(new_n574), .A4(new_n581), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n706), .A2(new_n707), .A3(new_n652), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n647), .B1(new_n648), .B2(new_n514), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT93), .B1(new_n642), .B2(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT93), .ZN(new_n711));
  INV_X1    g0511(.A(new_n486), .ZN(new_n712));
  OAI211_X1 g0512(.A(new_n689), .B(new_n711), .C1(new_n712), .C2(new_n493), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n624), .A2(new_n622), .ZN(new_n714));
  AND4_X1   g0514(.A1(new_n661), .A2(new_n714), .A3(new_n652), .A4(new_n654), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n710), .A2(new_n713), .A3(new_n715), .A4(new_n494), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n708), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n717), .A2(KEYINPUT29), .A3(new_n676), .ZN(new_n718));
  INV_X1    g0518(.A(KEYINPUT94), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n675), .B1(new_n708), .B2(new_n716), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n722));
  INV_X1    g0522(.A(KEYINPUT29), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n679), .A2(new_n487), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n655), .A2(new_n494), .A3(new_n625), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  AND3_X1   g0526(.A1(new_n662), .A2(new_n666), .A3(new_n652), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n675), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n720), .A2(new_n722), .B1(new_n723), .B2(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n536), .ZN(new_n732));
  INV_X1    g0532(.A(new_n481), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n595), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g0534(.A1(new_n558), .A2(new_n559), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n732), .A2(KEYINPUT30), .A3(new_n734), .A4(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n603), .A2(new_n535), .ZN(new_n737));
  NAND4_X1  g0537(.A1(new_n737), .A2(new_n288), .A3(new_n479), .A4(new_n553), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR3_X1   g0539(.A1(new_n536), .A2(new_n733), .A3(new_n595), .ZN(new_n740));
  AOI21_X1  g0540(.A(KEYINPUT30), .B1(new_n740), .B2(new_n735), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n675), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NOR3_X1   g0542(.A1(new_n626), .A2(new_n495), .A3(new_n675), .ZN(new_n743));
  INV_X1    g0543(.A(KEYINPUT31), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n742), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  OAI211_X1 g0545(.A(KEYINPUT31), .B(new_n675), .C1(new_n739), .C2(new_n741), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n731), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n730), .A2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n704), .B1(new_n748), .B2(G1), .ZN(G364));
  AND2_X1   g0549(.A1(new_n678), .A2(new_n680), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n750), .A2(G330), .ZN(new_n751));
  NAND2_X1  g0551(.A1(new_n682), .A2(KEYINPUT95), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n353), .A2(G20), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G45), .ZN(new_n754));
  NAND3_X1  g0554(.A1(new_n700), .A2(G1), .A3(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(KEYINPUT95), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n681), .A2(new_n756), .ZN(new_n757));
  NAND4_X1  g0557(.A1(new_n751), .A2(new_n752), .A3(new_n755), .A4(new_n757), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n698), .A2(new_n561), .ZN(new_n759));
  AND2_X1   g0559(.A1(new_n241), .A2(G45), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n216), .A2(G45), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n759), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(G355), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n561), .A2(new_n211), .ZN(new_n764));
  OAI22_X1  g0564(.A1(new_n763), .A2(new_n764), .B1(G116), .B2(new_n211), .ZN(new_n765));
  XOR2_X1   g0565(.A(new_n765), .B(KEYINPUT96), .Z(new_n766));
  NAND2_X1  g0566(.A1(new_n762), .A2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(G13), .A2(G33), .ZN(new_n768));
  INV_X1    g0568(.A(new_n768), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(G20), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n217), .B1(G20), .B2(new_n290), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n755), .B1(new_n767), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n771), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n288), .A2(new_n324), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n218), .A2(new_n386), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n265), .B1(new_n778), .B2(G50), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT97), .B(G159), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n218), .A2(G190), .ZN(new_n781));
  NOR2_X1   g0581(.A1(G179), .A2(G200), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  OR3_X1    g0583(.A1(new_n780), .A2(new_n783), .A3(KEYINPUT32), .ZN(new_n784));
  OAI21_X1  g0584(.A(KEYINPUT32), .B1(new_n780), .B2(new_n783), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n779), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n288), .A2(G200), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n776), .A2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n781), .A2(new_n787), .ZN(new_n789));
  OAI22_X1  g0589(.A1(new_n788), .A2(new_n202), .B1(new_n789), .B2(new_n299), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n324), .A2(G179), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n776), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n565), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n781), .A2(new_n791), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n794), .A2(new_n452), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n786), .A2(new_n790), .A3(new_n793), .A4(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n775), .A2(new_n781), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n218), .B1(new_n782), .B2(G190), .ZN(new_n798));
  OAI22_X1  g0598(.A1(new_n797), .A2(new_n203), .B1(new_n798), .B2(new_n566), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT98), .Z(new_n800));
  INV_X1    g0600(.A(new_n789), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n778), .A2(G326), .B1(new_n801), .B2(G311), .ZN(new_n802));
  INV_X1    g0602(.A(G303), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n802), .B1(new_n803), .B2(new_n792), .ZN(new_n804));
  XNOR2_X1  g0604(.A(KEYINPUT33), .B(G317), .ZN(new_n805));
  OR2_X1    g0605(.A1(new_n805), .A2(KEYINPUT99), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n797), .B1(new_n805), .B2(KEYINPUT99), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n804), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n265), .B1(new_n794), .B2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(G322), .ZN(new_n811));
  INV_X1    g0611(.A(G329), .ZN(new_n812));
  OAI22_X1  g0612(.A1(new_n788), .A2(new_n811), .B1(new_n783), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n798), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n810), .B(new_n813), .C1(G294), .C2(new_n814), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n796), .A2(new_n800), .B1(new_n808), .B2(new_n815), .ZN(new_n816));
  INV_X1    g0616(.A(new_n770), .ZN(new_n817));
  OAI221_X1 g0617(.A(new_n773), .B1(new_n774), .B2(new_n816), .C1(new_n750), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n758), .A2(new_n818), .ZN(G396));
  NOR2_X1   g0619(.A1(new_n771), .A2(new_n768), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT100), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n755), .B1(new_n822), .B2(new_n299), .ZN(new_n823));
  INV_X1    g0623(.A(new_n780), .ZN(new_n824));
  AOI22_X1  g0624(.A1(G137), .A2(new_n778), .B1(new_n824), .B2(new_n801), .ZN(new_n825));
  INV_X1    g0625(.A(G150), .ZN(new_n826));
  XNOR2_X1  g0626(.A(KEYINPUT102), .B(G143), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n825), .B1(new_n826), .B2(new_n797), .C1(new_n788), .C2(new_n827), .ZN(new_n828));
  XNOR2_X1  g0628(.A(new_n828), .B(KEYINPUT34), .ZN(new_n829));
  INV_X1    g0629(.A(new_n792), .ZN(new_n830));
  INV_X1    g0630(.A(new_n794), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G50), .A2(new_n830), .B1(new_n831), .B2(G68), .ZN(new_n832));
  OAI21_X1  g0632(.A(new_n832), .B1(new_n202), .B2(new_n798), .ZN(new_n833));
  INV_X1    g0633(.A(new_n783), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n265), .B1(new_n834), .B2(G132), .ZN(new_n835));
  AND2_X1   g0635(.A1(new_n835), .A2(KEYINPUT103), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n835), .A2(KEYINPUT103), .ZN(new_n837));
  NOR3_X1   g0637(.A1(new_n833), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n777), .A2(new_n803), .B1(new_n789), .B2(new_n500), .ZN(new_n839));
  INV_X1    g0639(.A(new_n797), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n839), .B1(G283), .B2(new_n840), .ZN(new_n841));
  XNOR2_X1  g0641(.A(new_n841), .B(KEYINPUT101), .ZN(new_n842));
  OAI22_X1  g0642(.A1(new_n792), .A2(new_n452), .B1(new_n794), .B2(new_n565), .ZN(new_n843));
  INV_X1    g0643(.A(G294), .ZN(new_n844));
  OAI221_X1 g0644(.A(new_n265), .B1(new_n798), .B2(new_n566), .C1(new_n844), .C2(new_n788), .ZN(new_n845));
  AOI211_X1 g0645(.A(new_n843), .B(new_n845), .C1(G311), .C2(new_n834), .ZN(new_n846));
  AOI22_X1  g0646(.A1(new_n829), .A2(new_n838), .B1(new_n842), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n314), .ZN(new_n848));
  OAI211_X1 g0648(.A(new_n328), .B(new_n676), .C1(new_n848), .C2(new_n312), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n328), .A2(new_n675), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n331), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n315), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n850), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n823), .B1(new_n774), .B2(new_n847), .C1(new_n854), .C2(new_n769), .ZN(new_n855));
  INV_X1    g0655(.A(new_n755), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n729), .B(new_n854), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n856), .B1(new_n857), .B2(new_n747), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n857), .A2(new_n747), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n855), .B1(new_n859), .B2(new_n860), .ZN(G384));
  NOR2_X1   g0661(.A1(new_n753), .A2(new_n254), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  OR2_X1    g0663(.A1(new_n400), .A2(new_n402), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT16), .B1(new_n864), .B2(new_n397), .ZN(new_n865));
  OAI21_X1  g0665(.A(new_n413), .B1(new_n865), .B2(new_n414), .ZN(new_n866));
  INV_X1    g0666(.A(new_n673), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n868), .B1(new_n418), .B2(new_n425), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n388), .A2(new_n409), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT37), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n383), .A2(G179), .ZN(new_n872));
  OAI21_X1  g0672(.A(new_n673), .B1(new_n872), .B2(new_n419), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(new_n415), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n875));
  AOI22_X1  g0675(.A1(new_n409), .A2(new_n388), .B1(new_n866), .B2(new_n873), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n875), .B1(new_n871), .B2(new_n876), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n869), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(new_n878), .ZN(new_n879));
  AOI21_X1  g0679(.A(KEYINPUT38), .B1(new_n869), .B2(new_n877), .ZN(new_n880));
  OR2_X1    g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n746), .B(KEYINPUT106), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n745), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n368), .A2(new_n675), .ZN(new_n884));
  NAND3_X1  g0684(.A1(new_n369), .A2(new_n373), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n290), .B1(new_n349), .B2(new_n350), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n351), .B1(new_n886), .B2(new_n346), .ZN(new_n887));
  INV_X1    g0687(.A(new_n347), .ZN(new_n888));
  OAI211_X1 g0688(.A(new_n368), .B(new_n675), .C1(new_n887), .C2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT104), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT104), .ZN(new_n891));
  NAND4_X1  g0691(.A1(new_n352), .A2(new_n891), .A3(new_n368), .A4(new_n675), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n885), .A2(new_n890), .A3(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n854), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n881), .A2(new_n883), .A3(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT105), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n878), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n869), .A2(KEYINPUT105), .A3(KEYINPUT38), .A4(new_n877), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT38), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n415), .A2(new_n867), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n632), .B2(new_n629), .ZN(new_n904));
  INV_X1    g0704(.A(new_n875), .ZN(new_n905));
  AOI21_X1  g0705(.A(new_n871), .B1(new_n870), .B2(new_n874), .ZN(new_n906));
  NOR2_X1   g0706(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n902), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n900), .A2(new_n901), .A3(new_n908), .ZN(new_n909));
  NAND4_X1  g0709(.A1(new_n883), .A2(new_n909), .A3(new_n895), .A4(KEYINPUT40), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n898), .A2(new_n910), .ZN(new_n911));
  AND2_X1   g0711(.A1(new_n427), .A2(new_n883), .ZN(new_n912));
  OAI211_X1 g0712(.A(new_n863), .B(G330), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  NAND3_X1  g0713(.A1(new_n898), .A2(G330), .A3(new_n910), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n427), .A2(new_n883), .A3(G330), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n914), .A2(KEYINPUT107), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n911), .A2(new_n912), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n913), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n638), .A2(new_n640), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n919), .B1(new_n730), .B2(new_n427), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT39), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n900), .A2(new_n921), .A3(new_n908), .A4(new_n901), .ZN(new_n922));
  OAI21_X1  g0722(.A(KEYINPUT39), .B1(new_n879), .B2(new_n880), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n369), .A2(new_n675), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n885), .A2(new_n890), .A3(new_n892), .ZN(new_n927));
  OAI211_X1 g0727(.A(new_n676), .B(new_n854), .C1(new_n657), .C2(new_n667), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n927), .B1(new_n928), .B2(new_n849), .ZN(new_n929));
  AOI22_X1  g0729(.A1(new_n929), .A2(new_n881), .B1(new_n425), .B2(new_n673), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n926), .A2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n920), .B(new_n931), .Z(new_n932));
  AOI21_X1  g0732(.A(new_n862), .B1(new_n918), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n918), .B2(new_n932), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n216), .A2(G77), .A3(new_n394), .A4(new_n395), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n935), .B1(G50), .B2(new_n203), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n936), .A2(G1), .A3(new_n353), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n609), .A2(new_n611), .A3(new_n612), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT35), .ZN(new_n939));
  OR2_X1    g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n939), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n940), .A2(G116), .A3(new_n219), .A4(new_n941), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT36), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n934), .A2(new_n937), .A3(new_n943), .ZN(G367));
  INV_X1    g0744(.A(new_n759), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n237), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n772), .B1(new_n211), .B2(new_n300), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n856), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n798), .A2(new_n452), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n792), .A2(new_n500), .ZN(new_n950));
  OAI221_X1 g0750(.A(new_n265), .B1(new_n566), .B2(new_n794), .C1(new_n950), .C2(KEYINPUT46), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n949), .B(new_n951), .C1(KEYINPUT46), .C2(new_n950), .ZN(new_n952));
  AOI22_X1  g0752(.A1(G294), .A2(new_n840), .B1(new_n801), .B2(G283), .ZN(new_n953));
  INV_X1    g0753(.A(G317), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n953), .B1(new_n954), .B2(new_n783), .ZN(new_n955));
  INV_X1    g0755(.A(G311), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n777), .A2(new_n956), .B1(new_n788), .B2(new_n803), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT115), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n957), .A2(new_n958), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n955), .A2(new_n959), .A3(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n780), .A2(new_n797), .B1(new_n788), .B2(new_n826), .ZN(new_n962));
  OAI22_X1  g0762(.A1(new_n777), .A2(new_n827), .B1(new_n792), .B2(new_n202), .ZN(new_n963));
  NOR2_X1   g0763(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n831), .A2(G77), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n201), .B2(new_n789), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n798), .A2(new_n203), .ZN(new_n967));
  INV_X1    g0767(.A(G137), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n561), .B1(new_n783), .B2(new_n968), .ZN(new_n969));
  NOR3_X1   g0769(.A1(new_n966), .A2(new_n967), .A3(new_n969), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n952), .A2(new_n961), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  OR2_X1    g0771(.A1(new_n971), .A2(KEYINPUT47), .ZN(new_n972));
  AOI21_X1  g0772(.A(new_n774), .B1(new_n971), .B2(KEYINPUT47), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n948), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n580), .A2(new_n676), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n975), .B(KEYINPUT108), .Z(new_n976));
  INV_X1    g0776(.A(new_n652), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT109), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n976), .A2(KEYINPUT109), .A3(new_n977), .ZN(new_n981));
  OAI211_X1 g0781(.A(new_n980), .B(new_n981), .C1(new_n705), .C2(new_n976), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n974), .B1(new_n982), .B2(new_n817), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n754), .A2(G1), .ZN(new_n984));
  INV_X1    g0784(.A(new_n687), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n691), .A2(new_n693), .ZN(new_n986));
  NAND2_X1  g0786(.A1(new_n986), .A2(KEYINPUT92), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n625), .B1(new_n622), .B2(new_n676), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT110), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n661), .B2(new_n676), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n664), .A2(KEYINPUT110), .A3(new_n675), .ZN(new_n991));
  AND3_X1   g0791(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n987), .A2(new_n694), .A3(new_n992), .ZN(new_n993));
  NOR2_X1   g0793(.A1(KEYINPUT113), .A2(KEYINPUT44), .ZN(new_n994));
  INV_X1    g0794(.A(new_n994), .ZN(new_n995));
  OR2_X1    g0795(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n995), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n996), .A2(new_n997), .B1(KEYINPUT113), .B2(KEYINPUT44), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n988), .A2(new_n990), .A3(new_n991), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n999), .B1(new_n695), .B2(new_n696), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT45), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n985), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(KEYINPUT113), .A2(KEYINPUT44), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n997), .ZN(new_n1004));
  NOR2_X1   g0804(.A1(new_n993), .A2(new_n995), .ZN(new_n1005));
  OAI21_X1  g0805(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT45), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1000), .B(new_n1007), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1008), .A3(new_n687), .ZN(new_n1009));
  OAI21_X1  g0809(.A(new_n691), .B1(new_n686), .B2(new_n690), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n1010), .A2(new_n752), .A3(new_n757), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT114), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  NAND4_X1  g0813(.A1(new_n1010), .A2(new_n752), .A3(KEYINPUT114), .A4(new_n757), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1010), .A2(new_n681), .ZN(new_n1015));
  AND3_X1   g0815(.A1(new_n1013), .A2(new_n1014), .A3(new_n1015), .ZN(new_n1016));
  NAND4_X1  g0816(.A1(new_n1002), .A2(new_n1009), .A3(new_n748), .A4(new_n1016), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1017), .A2(new_n748), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n699), .B(KEYINPUT41), .Z(new_n1019));
  INV_X1    g0819(.A(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n984), .B1(new_n1018), .B2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n982), .B(KEYINPUT43), .Z(new_n1022));
  OAI21_X1  g0822(.A(new_n661), .B1(new_n992), .B2(new_n487), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n676), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT42), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n1025), .B1(new_n992), .B2(new_n691), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n495), .B1(new_n465), .B2(new_n675), .ZN(new_n1027));
  NAND4_X1  g0827(.A1(new_n1027), .A2(KEYINPUT42), .A3(new_n690), .A4(new_n999), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1026), .A2(new_n1028), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1024), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g0830(.A(KEYINPUT111), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n1024), .A2(new_n1029), .A3(KEYINPUT111), .ZN(new_n1033));
  AND3_X1   g0833(.A1(new_n1022), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n982), .A2(KEYINPUT43), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1035), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1037));
  NOR3_X1   g0837(.A1(new_n1034), .A2(new_n1037), .A3(KEYINPUT112), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT112), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1022), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1042));
  AOI21_X1  g0842(.A(new_n1039), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  OAI22_X1  g0843(.A1(new_n1038), .A2(new_n1043), .B1(new_n687), .B2(new_n992), .ZN(new_n1044));
  OAI21_X1  g0844(.A(KEYINPUT112), .B1(new_n1034), .B2(new_n1037), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1041), .A2(new_n1042), .A3(new_n1039), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n985), .A4(new_n999), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g0848(.A(new_n983), .B1(new_n1021), .B2(new_n1048), .ZN(G387));
  OR2_X1    g0849(.A1(new_n686), .A2(new_n817), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n764), .A2(new_n701), .B1(G107), .B2(new_n211), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n233), .A2(G45), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n701), .ZN(new_n1053));
  AOI211_X1 g0853(.A(G45), .B(new_n1053), .C1(G68), .C2(G77), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n249), .A2(G50), .ZN(new_n1055));
  XNOR2_X1  g0855(.A(new_n1055), .B(KEYINPUT50), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n945), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1051), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n772), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n856), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g0860(.A(new_n1060), .B(KEYINPUT116), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n792), .A2(new_n299), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n797), .A2(new_n249), .B1(new_n789), .B2(new_n203), .ZN(new_n1063));
  AOI211_X1 g0863(.A(new_n1062), .B(new_n1063), .C1(G159), .C2(new_n778), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n788), .A2(new_n201), .B1(new_n783), .B2(new_n826), .ZN(new_n1065));
  AOI211_X1 g0865(.A(new_n265), .B(new_n1065), .C1(G97), .C2(new_n831), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n300), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n814), .A2(new_n1067), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1064), .A2(new_n1066), .A3(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n834), .A2(G326), .ZN(new_n1070));
  AOI21_X1  g0870(.A(new_n561), .B1(new_n831), .B2(G116), .ZN(new_n1071));
  OAI22_X1  g0871(.A1(new_n792), .A2(new_n844), .B1(new_n798), .B2(new_n809), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n778), .A2(G322), .B1(new_n801), .B2(G303), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n1073), .B1(new_n956), .B2(new_n797), .C1(new_n954), .C2(new_n788), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT117), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1072), .B1(new_n1075), .B2(KEYINPUT48), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1076), .B1(KEYINPUT48), .B2(new_n1075), .ZN(new_n1077));
  INV_X1    g0877(.A(KEYINPUT49), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1070), .B(new_n1071), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1079));
  AND2_X1   g0879(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1069), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1061), .B1(new_n771), .B2(new_n1081), .ZN(new_n1082));
  AOI22_X1  g0882(.A1(new_n1016), .A2(new_n984), .B1(new_n1050), .B2(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1016), .A2(new_n748), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(new_n699), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n1016), .A2(new_n748), .ZN(new_n1086));
  OAI21_X1  g0886(.A(new_n1083), .B1(new_n1085), .B2(new_n1086), .ZN(G393));
  NOR3_X1   g0887(.A1(new_n998), .A2(new_n1001), .A3(new_n985), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n687), .B1(new_n1006), .B2(new_n1008), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n1084), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n1017), .A3(new_n699), .ZN(new_n1091));
  NAND3_X1  g0891(.A1(new_n1002), .A2(new_n1009), .A3(new_n984), .ZN(new_n1092));
  OAI221_X1 g0892(.A(new_n772), .B1(new_n566), .B2(new_n211), .C1(new_n244), .C2(new_n945), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n856), .ZN(new_n1094));
  OAI221_X1 g0894(.A(new_n265), .B1(new_n789), .B2(new_n844), .C1(new_n452), .C2(new_n794), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n792), .A2(new_n809), .B1(new_n783), .B2(new_n811), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1095), .B1(KEYINPUT118), .B2(new_n1096), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n777), .A2(new_n954), .B1(new_n788), .B2(new_n956), .ZN(new_n1098));
  XNOR2_X1  g0898(.A(new_n1098), .B(KEYINPUT52), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1097), .B(new_n1099), .C1(KEYINPUT118), .C2(new_n1096), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n797), .A2(new_n803), .B1(new_n798), .B2(new_n500), .ZN(new_n1101));
  XOR2_X1   g0901(.A(new_n1101), .B(KEYINPUT119), .Z(new_n1102));
  INV_X1    g0902(.A(G159), .ZN(new_n1103));
  OAI22_X1  g0903(.A1(new_n777), .A2(new_n826), .B1(new_n788), .B2(new_n1103), .ZN(new_n1104));
  XOR2_X1   g0904(.A(new_n1104), .B(KEYINPUT51), .Z(new_n1105));
  NAND2_X1  g0905(.A1(new_n814), .A2(G77), .ZN(new_n1106));
  OAI211_X1 g0906(.A(new_n1106), .B(new_n561), .C1(new_n565), .C2(new_n794), .ZN(new_n1107));
  OAI22_X1  g0907(.A1(new_n797), .A2(new_n201), .B1(new_n783), .B2(new_n827), .ZN(new_n1108));
  OAI22_X1  g0908(.A1(new_n792), .A2(new_n203), .B1(new_n789), .B2(new_n249), .ZN(new_n1109));
  OR3_X1    g0909(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1100), .A2(new_n1102), .B1(new_n1105), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1094), .B1(new_n1111), .B2(new_n771), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n1112), .B1(new_n999), .B2(new_n817), .ZN(new_n1113));
  AND2_X1   g0913(.A1(new_n1092), .A2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1091), .A2(new_n1114), .ZN(G390));
  AOI21_X1  g0915(.A(new_n850), .B1(new_n728), .B2(new_n854), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n742), .ZN(new_n1117));
  AND4_X1   g0917(.A1(new_n661), .A2(new_n714), .A3(new_n574), .A4(new_n581), .ZN(new_n1118));
  NAND4_X1  g0918(.A1(new_n683), .A2(new_n543), .A3(new_n1118), .A4(new_n676), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1117), .B1(new_n1119), .B2(KEYINPUT31), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n746), .ZN(new_n1121));
  OAI21_X1  g0921(.A(G330), .B1(new_n1120), .B2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n854), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n927), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n731), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT106), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n746), .B(new_n1126), .ZN(new_n1127));
  OAI211_X1 g0927(.A(new_n1125), .B(new_n893), .C1(new_n1120), .C2(new_n1127), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1116), .B1(new_n1124), .B2(new_n1128), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n315), .B1(new_n331), .B2(new_n851), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n850), .B1(new_n721), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n1122), .B2(new_n894), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n893), .B1(new_n883), .B2(new_n1125), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n920), .B(new_n915), .C1(new_n1129), .C2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n923), .B(new_n922), .C1(new_n929), .C2(new_n925), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n925), .ZN(new_n1138));
  OAI211_X1 g0938(.A(new_n909), .B(new_n1138), .C1(new_n1132), .C2(new_n927), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n747), .A2(new_n895), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1138), .B1(new_n1116), .B2(new_n927), .ZN(new_n1142));
  AND2_X1   g0942(.A1(new_n922), .A2(new_n923), .ZN(new_n1143));
  AND2_X1   g0943(.A1(new_n909), .A2(new_n1138), .ZN(new_n1144));
  AOI211_X1 g0944(.A(new_n675), .B(new_n1130), .C1(new_n708), .C2(new_n716), .ZN(new_n1145));
  OAI21_X1  g0945(.A(new_n893), .B1(new_n1145), .B2(new_n850), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n1142), .A2(new_n1143), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1141), .B1(new_n1147), .B2(new_n1128), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n700), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT120), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1136), .A2(new_n1148), .A3(new_n1150), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n729), .A2(new_n723), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n721), .A2(KEYINPUT94), .A3(KEYINPUT29), .ZN(new_n1153));
  AOI21_X1  g0953(.A(KEYINPUT94), .B1(new_n721), .B2(KEYINPUT29), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n427), .C1(new_n1153), .C2(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1155), .A2(new_n641), .A3(new_n915), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1135), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1116), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n893), .B1(new_n747), .B2(new_n854), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1128), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1158), .B1(new_n1159), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1156), .B1(new_n1157), .B2(new_n1161), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1128), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n1163), .A2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(KEYINPUT120), .B1(new_n1162), .B2(new_n1165), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n1149), .B1(new_n1151), .B2(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1165), .A2(new_n984), .ZN(new_n1168));
  INV_X1    g0968(.A(G132), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(new_n792), .A2(new_n826), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT53), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n561), .B1(new_n1169), .B2(new_n788), .C1(new_n1170), .C2(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n778), .A2(G128), .B1(new_n831), .B2(G50), .ZN(new_n1173));
  INV_X1    g0973(.A(G125), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1173), .B1(new_n1174), .B2(new_n783), .ZN(new_n1175));
  AOI211_X1 g0975(.A(new_n1172), .B(new_n1175), .C1(new_n1171), .C2(new_n1170), .ZN(new_n1176));
  XNOR2_X1  g0976(.A(KEYINPUT54), .B(G143), .ZN(new_n1177));
  OAI22_X1  g0977(.A1(new_n797), .A2(new_n968), .B1(new_n789), .B2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G159), .B2(new_n814), .ZN(new_n1179));
  XOR2_X1   g0979(.A(new_n1179), .B(KEYINPUT121), .Z(new_n1180));
  NAND2_X1  g0980(.A1(new_n1176), .A2(new_n1180), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n203), .A2(new_n794), .B1(new_n789), .B2(new_n566), .ZN(new_n1182));
  NOR3_X1   g0982(.A1(new_n1182), .A2(new_n561), .A3(new_n793), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n778), .A2(G283), .B1(new_n840), .B2(G107), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n788), .ZN(new_n1185));
  AOI22_X1  g0985(.A1(G116), .A2(new_n1185), .B1(new_n834), .B2(G294), .ZN(new_n1186));
  NAND4_X1  g0986(.A1(new_n1183), .A2(new_n1106), .A3(new_n1184), .A4(new_n1186), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n774), .B1(new_n1181), .B2(new_n1187), .ZN(new_n1188));
  AOI211_X1 g0988(.A(new_n755), .B(new_n1188), .C1(new_n249), .C2(new_n822), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1189), .B1(new_n924), .B2(new_n769), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1167), .A2(new_n1168), .A3(new_n1190), .ZN(G378));
  NAND2_X1  g0991(.A1(new_n259), .A2(new_n867), .ZN(new_n1192));
  NAND3_X1  g0992(.A1(new_n636), .A2(new_n292), .A3(new_n1192), .ZN(new_n1193));
  INV_X1    g0993(.A(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1192), .B1(new_n636), .B2(new_n292), .ZN(new_n1195));
  XOR2_X1   g0995(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1196));
  OR3_X1    g0996(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n1196), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n931), .A2(new_n1199), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n926), .A2(new_n930), .A3(new_n1197), .A4(new_n1198), .ZN(new_n1201));
  AND3_X1   g1001(.A1(new_n1200), .A2(new_n914), .A3(new_n1201), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n914), .B1(new_n1200), .B2(new_n1201), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1202), .A2(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n984), .ZN(new_n1205));
  NOR2_X1   g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n755), .B1(new_n822), .B2(new_n201), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n503), .B(new_n277), .C1(new_n780), .C2(new_n794), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n777), .A2(new_n1174), .B1(new_n797), .B2(new_n1169), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1185), .A2(G128), .ZN(new_n1210));
  OAI221_X1 g1010(.A(new_n1210), .B1(new_n968), .B2(new_n789), .C1(new_n792), .C2(new_n1177), .ZN(new_n1211));
  AOI211_X1 g1011(.A(new_n1209), .B(new_n1211), .C1(G150), .C2(new_n814), .ZN(new_n1212));
  INV_X1    g1012(.A(new_n1212), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1213), .A2(KEYINPUT59), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1208), .B(new_n1214), .C1(G124), .C2(new_n834), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(KEYINPUT59), .B2(new_n1213), .ZN(new_n1216));
  NOR2_X1   g1016(.A1(new_n788), .A2(new_n452), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT122), .ZN(new_n1218));
  AOI22_X1  g1018(.A1(new_n778), .A2(G116), .B1(new_n801), .B2(new_n1067), .ZN(new_n1219));
  OAI211_X1 g1019(.A(new_n1218), .B(new_n1219), .C1(new_n809), .C2(new_n783), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n265), .A2(new_n277), .ZN(new_n1221));
  OR2_X1    g1021(.A1(new_n1062), .A2(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n797), .A2(new_n566), .B1(new_n794), .B2(new_n202), .ZN(new_n1223));
  NOR4_X1   g1023(.A1(new_n1220), .A2(new_n967), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  OR2_X1    g1024(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT58), .ZN(new_n1226));
  OAI211_X1 g1026(.A(new_n1221), .B(new_n201), .C1(G33), .C2(G41), .ZN(new_n1227));
  AND4_X1   g1027(.A1(new_n1216), .A2(new_n1225), .A3(new_n1226), .A4(new_n1227), .ZN(new_n1228));
  OAI221_X1 g1028(.A(new_n1207), .B1(new_n1228), .B2(new_n774), .C1(new_n769), .C2(new_n1199), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT123), .Z(new_n1230));
  NOR2_X1   g1030(.A1(new_n1206), .A2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1231), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1156), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1151), .B2(new_n1166), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT57), .ZN(new_n1235));
  INV_X1    g1035(.A(new_n1204), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1234), .A2(new_n1235), .A3(new_n1236), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n1150), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1238));
  NAND3_X1  g1038(.A1(new_n1162), .A2(new_n1165), .A3(KEYINPUT120), .ZN(new_n1239));
  AOI21_X1  g1039(.A(new_n1156), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1240));
  OAI21_X1  g1040(.A(KEYINPUT57), .B1(new_n1240), .B2(new_n1204), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1232), .B1(new_n1242), .B2(new_n699), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1243), .ZN(G375));
  NOR2_X1   g1044(.A1(new_n1129), .A2(new_n1135), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(new_n1156), .ZN(new_n1246));
  NAND3_X1  g1046(.A1(new_n1246), .A2(new_n1020), .A3(new_n1136), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n927), .A2(new_n768), .ZN(new_n1248));
  OAI21_X1  g1048(.A(new_n856), .B1(new_n821), .B2(G68), .ZN(new_n1249));
  AOI22_X1  g1049(.A1(G150), .A2(new_n801), .B1(new_n834), .B2(G128), .ZN(new_n1250));
  OAI221_X1 g1050(.A(new_n1250), .B1(new_n1103), .B2(new_n792), .C1(new_n797), .C2(new_n1177), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(G132), .A2(new_n778), .B1(new_n1185), .B2(G137), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n265), .B1(new_n831), .B2(G58), .ZN(new_n1253));
  OAI211_X1 g1053(.A(new_n1252), .B(new_n1253), .C1(new_n201), .C2(new_n798), .ZN(new_n1254));
  AOI22_X1  g1054(.A1(G97), .A2(new_n830), .B1(new_n834), .B2(G303), .ZN(new_n1255));
  OAI221_X1 g1055(.A(new_n1255), .B1(new_n452), .B2(new_n789), .C1(new_n844), .C2(new_n777), .ZN(new_n1256));
  AOI22_X1  g1056(.A1(G116), .A2(new_n840), .B1(new_n1185), .B2(G283), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(new_n265), .A3(new_n965), .A4(new_n1068), .ZN(new_n1258));
  OAI22_X1  g1058(.A1(new_n1251), .A2(new_n1254), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1249), .B1(new_n1259), .B2(new_n771), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1248), .A2(new_n1260), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1261), .B1(new_n1245), .B2(new_n1205), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1262), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1247), .A2(new_n1263), .ZN(G381));
  INV_X1    g1064(.A(G378), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1243), .A2(new_n1265), .ZN(new_n1266));
  OR2_X1    g1066(.A1(G393), .A2(G396), .ZN(new_n1267));
  OR4_X1    g1067(.A1(G384), .A2(new_n1267), .A3(G381), .A4(G390), .ZN(new_n1268));
  OR3_X1    g1068(.A1(new_n1266), .A2(G387), .A3(new_n1268), .ZN(G407));
  OAI211_X1 g1069(.A(G407), .B(G213), .C1(G343), .C2(new_n1266), .ZN(G409));
  OAI211_X1 g1070(.A(new_n983), .B(G390), .C1(new_n1021), .C2(new_n1048), .ZN(new_n1271));
  INV_X1    g1071(.A(KEYINPUT124), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  XNOR2_X1  g1073(.A(G393), .B(G396), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1271), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1019), .B1(new_n1017), .B2(new_n748), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1047), .B(new_n1044), .C1(new_n1277), .C2(new_n984), .ZN(new_n1278));
  AOI21_X1  g1078(.A(G390), .B1(new_n1278), .B2(new_n983), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1273), .B(new_n1275), .C1(new_n1276), .C2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(G390), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(G387), .A2(new_n1281), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1282), .B(new_n1271), .C1(new_n1272), .C2(new_n1274), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(G384), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1246), .A2(KEYINPUT60), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT60), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1245), .A2(new_n1288), .A3(new_n1156), .ZN(new_n1289));
  AOI211_X1 g1089(.A(new_n700), .B(new_n1162), .C1(new_n1287), .C2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n1286), .B1(new_n1290), .B2(new_n1262), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(new_n699), .A3(new_n1136), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(G384), .A3(new_n1263), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1291), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n674), .A2(G213), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(G2897), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1295), .B(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1234), .A2(new_n1020), .A3(new_n1236), .ZN(new_n1300));
  AOI21_X1  g1100(.A(G378), .B1(new_n1300), .B2(new_n1231), .ZN(new_n1301));
  AOI21_X1  g1101(.A(new_n1301), .B1(new_n1243), .B2(G378), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1299), .B1(new_n1302), .B2(new_n1297), .ZN(new_n1303));
  INV_X1    g1103(.A(KEYINPUT61), .ZN(new_n1304));
  AOI21_X1  g1104(.A(new_n1235), .B1(new_n1234), .B2(new_n1236), .ZN(new_n1305));
  NOR3_X1   g1105(.A1(new_n1240), .A2(KEYINPUT57), .A3(new_n1204), .ZN(new_n1306));
  OAI21_X1  g1106(.A(new_n699), .B1(new_n1305), .B2(new_n1306), .ZN(new_n1307));
  NAND3_X1  g1107(.A1(new_n1307), .A2(G378), .A3(new_n1231), .ZN(new_n1308));
  INV_X1    g1108(.A(new_n1301), .ZN(new_n1309));
  AOI211_X1 g1109(.A(new_n1297), .B(new_n1295), .C1(new_n1308), .C2(new_n1309), .ZN(new_n1310));
  INV_X1    g1110(.A(KEYINPUT62), .ZN(new_n1311));
  OAI211_X1 g1111(.A(new_n1303), .B(new_n1304), .C1(new_n1310), .C2(new_n1311), .ZN(new_n1312));
  INV_X1    g1112(.A(new_n1295), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n700), .B1(new_n1237), .B2(new_n1241), .ZN(new_n1314));
  NOR3_X1   g1114(.A1(new_n1314), .A2(new_n1265), .A3(new_n1232), .ZN(new_n1315));
  OAI211_X1 g1115(.A(new_n1296), .B(new_n1313), .C1(new_n1315), .C2(new_n1301), .ZN(new_n1316));
  NOR2_X1   g1116(.A1(new_n1316), .A2(KEYINPUT62), .ZN(new_n1317));
  OAI21_X1  g1117(.A(new_n1285), .B1(new_n1312), .B2(new_n1317), .ZN(new_n1318));
  AOI21_X1  g1118(.A(new_n1297), .B1(new_n1308), .B2(new_n1309), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(new_n1303), .A2(KEYINPUT63), .B1(new_n1313), .B2(new_n1319), .ZN(new_n1320));
  INV_X1    g1120(.A(KEYINPUT125), .ZN(new_n1321));
  AOI21_X1  g1121(.A(KEYINPUT61), .B1(new_n1280), .B2(new_n1283), .ZN(new_n1322));
  INV_X1    g1122(.A(KEYINPUT63), .ZN(new_n1323));
  OAI21_X1  g1123(.A(new_n1322), .B1(new_n1316), .B2(new_n1323), .ZN(new_n1324));
  NOR3_X1   g1124(.A1(new_n1320), .A2(new_n1321), .A3(new_n1324), .ZN(new_n1325));
  NAND3_X1  g1125(.A1(new_n1295), .A2(G2897), .A3(new_n1297), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1291), .A2(new_n1294), .A3(new_n1298), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1326), .A2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1308), .A2(new_n1309), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1328), .B1(new_n1329), .B2(new_n1296), .ZN(new_n1330));
  OAI21_X1  g1130(.A(new_n1316), .B1(new_n1330), .B2(new_n1323), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1284), .A2(new_n1304), .ZN(new_n1332));
  AOI21_X1  g1132(.A(new_n1332), .B1(new_n1310), .B2(KEYINPUT63), .ZN(new_n1333));
  AOI21_X1  g1133(.A(KEYINPUT125), .B1(new_n1331), .B2(new_n1333), .ZN(new_n1334));
  OAI21_X1  g1134(.A(new_n1318), .B1(new_n1325), .B2(new_n1334), .ZN(G405));
  NAND2_X1  g1135(.A1(G375), .A2(new_n1265), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1313), .A2(KEYINPUT127), .ZN(new_n1337));
  NAND3_X1  g1137(.A1(new_n1336), .A2(new_n1308), .A3(new_n1337), .ZN(new_n1338));
  AND2_X1   g1138(.A1(new_n1338), .A2(new_n1285), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1338), .A2(new_n1285), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT127), .ZN(new_n1341));
  OAI21_X1  g1141(.A(new_n1341), .B1(new_n1295), .B2(KEYINPUT126), .ZN(new_n1342));
  OR3_X1    g1142(.A1(new_n1339), .A2(new_n1340), .A3(new_n1342), .ZN(new_n1343));
  OAI21_X1  g1143(.A(new_n1342), .B1(new_n1339), .B2(new_n1340), .ZN(new_n1344));
  NAND2_X1  g1144(.A1(new_n1343), .A2(new_n1344), .ZN(G402));
endmodule


