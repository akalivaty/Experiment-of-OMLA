//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 1 0 1 1 1 0 1 1 0 0 0 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:13 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n449, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n507, new_n508, new_n509, new_n510, new_n511, new_n512,
    new_n513, new_n514, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n541, new_n542, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1194, new_n1195, new_n1196,
    new_n1198;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT64), .Z(G217));
  NOR4_X1   g025(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT65), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n452), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(new_n452), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n457), .A2(G2106), .ZN(new_n458));
  INV_X1    g033(.A(new_n454), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n459), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n458), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  AND2_X1   g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  NOR2_X1   g039(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n465));
  OAI21_X1  g040(.A(G125), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n463), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  OAI211_X1 g043(.A(G137), .B(new_n463), .C1(new_n464), .C2(new_n465), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n463), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n468), .A2(new_n471), .ZN(G160));
  OR2_X1    g047(.A1(G100), .A2(G2105), .ZN(new_n473));
  OAI211_X1 g048(.A(new_n473), .B(G2104), .C1(G112), .C2(new_n463), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT67), .ZN(new_n475));
  XNOR2_X1  g050(.A(KEYINPUT3), .B(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G2105), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT66), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n476), .A2(new_n479), .A3(G2105), .ZN(new_n480));
  AND3_X1   g055(.A1(new_n478), .A2(G124), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n476), .A2(new_n463), .ZN(new_n482));
  INV_X1    g057(.A(new_n482), .ZN(new_n483));
  AOI211_X1 g058(.A(new_n475), .B(new_n481), .C1(G136), .C2(new_n483), .ZN(G162));
  OAI211_X1 g059(.A(G126), .B(G2105), .C1(new_n464), .C2(new_n465), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G114), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G2105), .ZN(new_n488));
  NAND3_X1  g063(.A1(new_n486), .A2(new_n488), .A3(G2104), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(G138), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n491), .A2(G2105), .ZN(new_n492));
  OAI21_X1  g067(.A(new_n492), .B1(new_n464), .B2(new_n465), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(KEYINPUT4), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT4), .ZN(new_n495));
  OAI211_X1 g070(.A(new_n492), .B(new_n495), .C1(new_n465), .C2(new_n464), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(G164));
  XNOR2_X1  g072(.A(KEYINPUT6), .B(G651), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(G50), .A3(G543), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT5), .B(G543), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(new_n498), .ZN(new_n501));
  INV_X1    g076(.A(G88), .ZN(new_n502));
  AOI22_X1  g077(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n503));
  INV_X1    g078(.A(G651), .ZN(new_n504));
  OAI221_X1 g079(.A(new_n499), .B1(new_n501), .B2(new_n502), .C1(new_n503), .C2(new_n504), .ZN(G303));
  INV_X1    g080(.A(G303), .ZN(G166));
  NAND3_X1  g081(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n507));
  XNOR2_X1  g082(.A(new_n507), .B(KEYINPUT7), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n498), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(G51), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AND2_X1   g086(.A1(KEYINPUT5), .A2(G543), .ZN(new_n512));
  NOR2_X1   g087(.A1(KEYINPUT5), .A2(G543), .ZN(new_n513));
  NOR2_X1   g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n498), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n514), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT68), .ZN(new_n518));
  OR3_X1    g093(.A1(new_n511), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n511), .B2(new_n517), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n519), .A2(new_n520), .ZN(G168));
  INV_X1    g096(.A(KEYINPUT69), .ZN(new_n522));
  INV_X1    g097(.A(G90), .ZN(new_n523));
  INV_X1    g098(.A(G52), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n501), .A2(new_n523), .B1(new_n509), .B2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n526), .A2(new_n504), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  NOR3_X1   g104(.A1(new_n525), .A2(new_n527), .A3(new_n522), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n529), .A2(new_n530), .ZN(G301));
  INV_X1    g106(.A(G301), .ZN(G171));
  INV_X1    g107(.A(G81), .ZN(new_n533));
  INV_X1    g108(.A(G43), .ZN(new_n534));
  OAI22_X1  g109(.A1(new_n501), .A2(new_n533), .B1(new_n509), .B2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n504), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n538), .A2(G860), .ZN(G153));
  NAND4_X1  g114(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g115(.A1(G1), .A2(G3), .ZN(new_n541));
  XNOR2_X1  g116(.A(new_n541), .B(KEYINPUT8), .ZN(new_n542));
  NAND4_X1  g117(.A1(G319), .A2(G483), .A3(G661), .A4(new_n542), .ZN(G188));
  NAND2_X1  g118(.A1(G78), .A2(G543), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n544), .B(KEYINPUT72), .ZN(new_n545));
  INV_X1    g120(.A(G65), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n545), .B1(new_n546), .B2(new_n514), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n549));
  INV_X1    g124(.A(KEYINPUT9), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n498), .A2(G53), .A3(G543), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT71), .ZN(new_n552));
  OAI211_X1 g127(.A(new_n549), .B(new_n550), .C1(new_n551), .C2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n501), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G91), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n548), .A2(new_n553), .A3(new_n555), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  OR2_X1    g132(.A1(new_n551), .A2(new_n549), .ZN(new_n558));
  OAI21_X1  g133(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(KEYINPUT9), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G299));
  INV_X1    g136(.A(G168), .ZN(G286));
  NAND2_X1  g137(.A1(new_n554), .A2(G87), .ZN(new_n563));
  INV_X1    g138(.A(new_n509), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G49), .ZN(new_n565));
  OAI21_X1  g140(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n566));
  AND3_X1   g141(.A1(new_n563), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G288));
  INV_X1    g143(.A(G86), .ZN(new_n569));
  INV_X1    g144(.A(G48), .ZN(new_n570));
  OAI22_X1  g145(.A1(new_n501), .A2(new_n569), .B1(new_n509), .B2(new_n570), .ZN(new_n571));
  INV_X1    g146(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(G73), .A2(G543), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT74), .ZN(new_n574));
  XNOR2_X1  g149(.A(new_n573), .B(new_n574), .ZN(new_n575));
  OAI211_X1 g150(.A(KEYINPUT73), .B(G61), .C1(new_n512), .C2(new_n513), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g152(.A(KEYINPUT73), .B1(new_n500), .B2(G61), .ZN(new_n578));
  OAI211_X1 g153(.A(KEYINPUT75), .B(G651), .C1(new_n577), .C2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT73), .ZN(new_n581));
  INV_X1    g156(.A(G61), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n514), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g158(.A1(new_n583), .A2(new_n576), .A3(new_n575), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT75), .B1(new_n584), .B2(G651), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n572), .B1(new_n580), .B2(new_n585), .ZN(G305));
  AND2_X1   g161(.A1(new_n500), .A2(G60), .ZN(new_n587));
  AND2_X1   g162(.A1(G72), .A2(G543), .ZN(new_n588));
  OAI21_X1  g163(.A(G651), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  AOI22_X1  g166(.A1(G85), .A2(new_n554), .B1(new_n564), .B2(G47), .ZN(new_n592));
  OAI211_X1 g167(.A(KEYINPUT76), .B(G651), .C1(new_n587), .C2(new_n588), .ZN(new_n593));
  NAND3_X1  g168(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT77), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND4_X1  g171(.A1(new_n591), .A2(new_n592), .A3(KEYINPUT77), .A4(new_n593), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n596), .A2(new_n597), .ZN(G290));
  AND3_X1   g173(.A1(new_n500), .A2(new_n498), .A3(G92), .ZN(new_n599));
  XNOR2_X1  g174(.A(new_n599), .B(KEYINPUT10), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n514), .B2(new_n602), .ZN(new_n603));
  AOI22_X1  g178(.A1(G54), .A2(new_n564), .B1(new_n603), .B2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n605), .A2(G868), .ZN(new_n606));
  AOI21_X1  g181(.A(new_n606), .B1(G171), .B2(G868), .ZN(G284));
  AOI21_X1  g182(.A(new_n606), .B1(G171), .B2(G868), .ZN(G321));
  MUX2_X1   g183(.A(G299), .B(G286), .S(G868), .Z(G280));
  XNOR2_X1  g184(.A(G280), .B(KEYINPUT78), .ZN(G297));
  INV_X1    g185(.A(new_n605), .ZN(new_n611));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(G860), .ZN(G148));
  OAI21_X1  g188(.A(KEYINPUT79), .B1(new_n538), .B2(G868), .ZN(new_n614));
  NAND2_X1  g189(.A1(new_n611), .A2(new_n612), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(G868), .ZN(new_n616));
  MUX2_X1   g191(.A(KEYINPUT79), .B(new_n614), .S(new_n616), .Z(G323));
  XNOR2_X1  g192(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND3_X1  g193(.A1(new_n478), .A2(G123), .A3(new_n480), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n483), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n463), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n623), .A2(G2096), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  XNOR2_X1  g200(.A(KEYINPUT80), .B(KEYINPUT12), .ZN(new_n626));
  NAND3_X1  g201(.A1(new_n463), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n626), .B(new_n627), .ZN(new_n628));
  XOR2_X1   g203(.A(new_n628), .B(KEYINPUT13), .Z(new_n629));
  AOI21_X1  g204(.A(new_n624), .B1(new_n625), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n623), .A2(G2096), .ZN(new_n631));
  OAI211_X1 g206(.A(new_n630), .B(new_n631), .C1(new_n625), .C2(new_n629), .ZN(G156));
  INV_X1    g207(.A(G14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2443), .B(G2446), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(KEYINPUT15), .B(G2435), .Z(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT81), .B(G2438), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2427), .B(G2430), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  OR2_X1    g216(.A1(new_n636), .A2(new_n637), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n636), .A2(new_n637), .ZN(new_n643));
  NAND3_X1  g218(.A1(new_n642), .A2(new_n639), .A3(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(KEYINPUT14), .A3(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT82), .ZN(new_n646));
  XNOR2_X1  g221(.A(G2451), .B(G2454), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n647), .B(KEYINPUT16), .Z(new_n648));
  NOR2_X1   g223(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  INV_X1    g224(.A(KEYINPUT82), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n645), .B(new_n650), .ZN(new_n651));
  INV_X1    g226(.A(new_n648), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n635), .B1(new_n649), .B2(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(G1341), .B(G1348), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n646), .A2(new_n648), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n651), .A2(new_n652), .ZN(new_n658));
  NAND3_X1  g233(.A1(new_n657), .A2(new_n658), .A3(new_n634), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n654), .A2(new_n656), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n660), .A2(KEYINPUT83), .ZN(new_n661));
  INV_X1    g236(.A(KEYINPUT83), .ZN(new_n662));
  NAND4_X1  g237(.A1(new_n654), .A2(new_n662), .A3(new_n659), .A4(new_n656), .ZN(new_n663));
  AOI21_X1  g238(.A(new_n633), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AND3_X1   g239(.A1(new_n657), .A2(new_n658), .A3(new_n634), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n634), .B1(new_n657), .B2(new_n658), .ZN(new_n666));
  OAI21_X1  g241(.A(new_n655), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT84), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  OAI211_X1 g244(.A(KEYINPUT84), .B(new_n655), .C1(new_n665), .C2(new_n666), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  AND2_X1   g246(.A1(new_n664), .A2(new_n671), .ZN(G401));
  INV_X1    g247(.A(KEYINPUT18), .ZN(new_n673));
  XOR2_X1   g248(.A(G2084), .B(G2090), .Z(new_n674));
  XNOR2_X1  g249(.A(G2067), .B(G2678), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(KEYINPUT17), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  OAI21_X1  g253(.A(new_n673), .B1(new_n677), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(new_n625), .ZN(new_n680));
  XOR2_X1   g255(.A(G2072), .B(G2078), .Z(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(new_n676), .B2(KEYINPUT18), .ZN(new_n682));
  XOR2_X1   g257(.A(new_n682), .B(G2096), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n680), .B(new_n683), .ZN(G227));
  XNOR2_X1  g259(.A(G1956), .B(G2474), .ZN(new_n685));
  INV_X1    g260(.A(KEYINPUT85), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  XOR2_X1   g262(.A(G1961), .B(G1966), .Z(new_n688));
  OR2_X1    g263(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(G1971), .B(G1976), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT19), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n687), .A2(new_n688), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n689), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n692), .A2(new_n691), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT20), .ZN(new_n695));
  NOR2_X1   g270(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NOR3_X1   g271(.A1(new_n692), .A2(KEYINPUT20), .A3(new_n691), .ZN(new_n697));
  OAI221_X1 g272(.A(new_n693), .B1(new_n691), .B2(new_n689), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1981), .B(G1986), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT87), .ZN(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  XNOR2_X1  g276(.A(new_n698), .B(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(KEYINPUT86), .ZN(new_n704));
  XNOR2_X1  g279(.A(G1991), .B(G1996), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT88), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n704), .B(new_n706), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n702), .A2(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n702), .A2(new_n707), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(G229));
  INV_X1    g285(.A(G16), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G24), .ZN(new_n712));
  INV_X1    g287(.A(G290), .ZN(new_n713));
  OAI21_X1  g288(.A(new_n712), .B1(new_n713), .B2(new_n711), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(G1986), .ZN(new_n715));
  INV_X1    g290(.A(KEYINPUT93), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(G1986), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n714), .B(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(KEYINPUT93), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n476), .A2(G131), .A3(new_n463), .ZN(new_n721));
  INV_X1    g296(.A(KEYINPUT90), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n721), .B(new_n722), .ZN(new_n723));
  NAND3_X1  g298(.A1(new_n478), .A2(G119), .A3(new_n480), .ZN(new_n724));
  OR2_X1    g299(.A1(G95), .A2(G2105), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n725), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n726));
  NAND3_X1  g301(.A1(new_n723), .A2(new_n724), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n727), .A2(G29), .ZN(new_n728));
  INV_X1    g303(.A(G29), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n729), .A2(G25), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n730), .B(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT35), .B(G1991), .Z(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT91), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(KEYINPUT92), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n732), .B(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n717), .A2(new_n720), .A3(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(G651), .B1(new_n577), .B2(new_n578), .ZN(new_n738));
  INV_X1    g313(.A(KEYINPUT75), .ZN(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI21_X1  g315(.A(new_n571), .B1(new_n740), .B2(new_n579), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n741), .A2(G16), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n742), .B1(G6), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT32), .B(G1981), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT94), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n745), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n711), .A2(G22), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G166), .B2(new_n711), .ZN(new_n749));
  INV_X1    g324(.A(G1971), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n711), .A2(G23), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n752), .B1(new_n567), .B2(new_n711), .ZN(new_n753));
  XNOR2_X1  g328(.A(KEYINPUT33), .B(G1976), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(KEYINPUT95), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n753), .B(new_n755), .Z(new_n756));
  NAND4_X1  g331(.A1(new_n746), .A2(new_n747), .A3(new_n751), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT34), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n737), .A2(new_n758), .ZN(new_n759));
  AND2_X1   g334(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G162), .A2(new_n729), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n729), .A2(G35), .ZN(new_n763));
  XOR2_X1   g338(.A(new_n763), .B(KEYINPUT102), .Z(new_n764));
  NOR2_X1   g339(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT29), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n766), .A2(G2090), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(KEYINPUT103), .ZN(new_n768));
  XNOR2_X1  g343(.A(KEYINPUT31), .B(G11), .ZN(new_n769));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n729), .B1(new_n770), .B2(G28), .ZN(new_n771));
  AND2_X1   g346(.A1(new_n771), .A2(KEYINPUT101), .ZN(new_n772));
  NAND2_X1  g347(.A1(new_n770), .A2(G28), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n773), .B1(new_n771), .B2(KEYINPUT101), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n769), .B1(new_n772), .B2(new_n774), .C1(new_n623), .C2(new_n729), .ZN(new_n775));
  NAND2_X1  g350(.A1(new_n483), .A2(G139), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n476), .A2(G127), .ZN(new_n778));
  NAND2_X1  g353(.A1(G115), .A2(G2104), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n463), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT25), .ZN(new_n782));
  NOR3_X1   g357(.A1(new_n777), .A2(new_n780), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n783), .A2(new_n729), .ZN(new_n784));
  AOI21_X1  g359(.A(new_n784), .B1(new_n729), .B2(G33), .ZN(new_n785));
  INV_X1    g360(.A(G2072), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n775), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(KEYINPUT24), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n729), .B1(new_n788), .B2(G34), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(new_n788), .B2(G34), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G160), .B2(G29), .ZN(new_n791));
  NOR2_X1   g366(.A1(new_n791), .A2(G2084), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G2084), .ZN(new_n793));
  NAND2_X1  g368(.A1(G164), .A2(G29), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n794), .B1(G27), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2078), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n793), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  NOR2_X1   g372(.A1(G16), .A2(G19), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n538), .B2(G16), .ZN(new_n799));
  AOI211_X1 g374(.A(new_n792), .B(new_n797), .C1(G1341), .C2(new_n799), .ZN(new_n800));
  OAI211_X1 g375(.A(new_n787), .B(new_n800), .C1(new_n766), .C2(G2090), .ZN(new_n801));
  NOR2_X1   g376(.A1(G171), .A2(new_n711), .ZN(new_n802));
  AOI21_X1  g377(.A(new_n802), .B1(G5), .B2(new_n711), .ZN(new_n803));
  INV_X1    g378(.A(G1961), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n799), .A2(G1341), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n796), .B2(new_n795), .ZN(new_n807));
  OAI211_X1 g382(.A(new_n805), .B(new_n807), .C1(new_n786), .C2(new_n785), .ZN(new_n808));
  NOR2_X1   g383(.A1(G4), .A2(G16), .ZN(new_n809));
  XNOR2_X1  g384(.A(new_n809), .B(KEYINPUT97), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n605), .B2(new_n711), .ZN(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT98), .B(G1348), .ZN(new_n812));
  INV_X1    g387(.A(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n811), .B(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n814), .B1(new_n803), .B2(new_n804), .ZN(new_n815));
  NOR3_X1   g390(.A1(new_n801), .A2(new_n808), .A3(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n729), .A2(G26), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT28), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n478), .A2(G128), .A3(new_n480), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n819), .A2(KEYINPUT99), .ZN(new_n820));
  INV_X1    g395(.A(KEYINPUT99), .ZN(new_n821));
  NAND4_X1  g396(.A1(new_n478), .A2(new_n821), .A3(G128), .A4(new_n480), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  OR2_X1    g398(.A1(G104), .A2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n824), .B(G2104), .C1(G116), .C2(new_n463), .ZN(new_n825));
  INV_X1    g400(.A(G140), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n825), .B1(new_n482), .B2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n823), .A2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n818), .B1(new_n830), .B2(new_n729), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(G2067), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n711), .A2(G20), .ZN(new_n833));
  XOR2_X1   g408(.A(new_n833), .B(KEYINPUT23), .Z(new_n834));
  AOI21_X1  g409(.A(new_n834), .B1(G299), .B2(G16), .ZN(new_n835));
  INV_X1    g410(.A(G1956), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NOR2_X1   g412(.A1(new_n832), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n478), .A2(G129), .A3(new_n480), .ZN(new_n839));
  NAND3_X1  g414(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n840));
  INV_X1    g415(.A(KEYINPUT26), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND3_X1  g417(.A1(new_n476), .A2(G141), .A3(new_n463), .ZN(new_n843));
  NAND3_X1  g418(.A1(new_n463), .A2(G105), .A3(G2104), .ZN(new_n844));
  AND3_X1   g419(.A1(new_n842), .A2(new_n843), .A3(new_n844), .ZN(new_n845));
  AND3_X1   g420(.A1(new_n839), .A2(new_n845), .A3(KEYINPUT100), .ZN(new_n846));
  AOI21_X1  g421(.A(KEYINPUT100), .B1(new_n839), .B2(new_n845), .ZN(new_n847));
  OR2_X1    g422(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  MUX2_X1   g423(.A(G32), .B(new_n848), .S(G29), .Z(new_n849));
  XNOR2_X1  g424(.A(KEYINPUT27), .B(G1996), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n849), .B(new_n850), .Z(new_n851));
  NOR2_X1   g426(.A1(G16), .A2(G21), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n852), .B1(G168), .B2(G16), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(G1966), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g430(.A1(new_n768), .A2(new_n816), .A3(new_n838), .A4(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n761), .A2(new_n856), .ZN(G311));
  OR2_X1    g432(.A1(new_n761), .A2(new_n856), .ZN(G150));
  NAND2_X1  g433(.A1(new_n611), .A2(G559), .ZN(new_n859));
  XNOR2_X1  g434(.A(new_n859), .B(KEYINPUT38), .ZN(new_n860));
  INV_X1    g435(.A(G93), .ZN(new_n861));
  INV_X1    g436(.A(G55), .ZN(new_n862));
  OAI22_X1  g437(.A1(new_n501), .A2(new_n861), .B1(new_n509), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g438(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n504), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(new_n538), .ZN(new_n867));
  INV_X1    g442(.A(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n860), .B(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT39), .ZN(new_n870));
  AOI21_X1  g445(.A(G860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n870), .B2(new_n869), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT104), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n866), .A2(G860), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT37), .Z(new_n875));
  NAND2_X1  g450(.A1(new_n873), .A2(new_n875), .ZN(G145));
  INV_X1    g451(.A(new_n496), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n495), .B1(new_n476), .B2(new_n492), .ZN(new_n878));
  OAI211_X1 g453(.A(new_n485), .B(new_n489), .C1(new_n877), .C2(new_n878), .ZN(new_n879));
  AOI21_X1  g454(.A(new_n879), .B1(new_n823), .B2(new_n828), .ZN(new_n880));
  AOI211_X1 g455(.A(G164), .B(new_n827), .C1(new_n820), .C2(new_n822), .ZN(new_n881));
  NOR2_X1   g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n839), .A2(new_n845), .ZN(new_n883));
  OR2_X1    g458(.A1(new_n783), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n783), .B1(new_n846), .B2(new_n847), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g461(.A1(new_n882), .A2(new_n886), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n884), .B(new_n885), .C1(new_n880), .C2(new_n881), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n727), .A2(new_n628), .ZN(new_n890));
  INV_X1    g465(.A(G142), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n463), .A2(G118), .ZN(new_n892));
  OAI21_X1  g467(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n893));
  OAI22_X1  g468(.A1(new_n482), .A2(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n478), .A2(G130), .A3(new_n480), .ZN(new_n895));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n478), .A2(KEYINPUT105), .A3(G130), .A4(new_n480), .ZN(new_n898));
  AOI21_X1  g473(.A(new_n894), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n628), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n723), .A2(new_n900), .A3(new_n724), .A4(new_n726), .ZN(new_n901));
  AND3_X1   g476(.A1(new_n890), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n899), .B1(new_n890), .B2(new_n901), .ZN(new_n903));
  OAI21_X1  g478(.A(new_n889), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n623), .B(G160), .ZN(new_n906));
  XNOR2_X1  g481(.A(new_n906), .B(G162), .ZN(new_n907));
  NOR2_X1   g482(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n902), .A2(new_n903), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n909), .A2(new_n887), .A3(new_n888), .ZN(new_n910));
  AOI21_X1  g485(.A(G37), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(KEYINPUT106), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT106), .ZN(new_n913));
  NAND4_X1  g488(.A1(new_n909), .A2(new_n887), .A3(new_n913), .A4(new_n888), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n912), .A2(new_n904), .A3(new_n914), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n915), .A2(KEYINPUT107), .A3(new_n907), .ZN(new_n916));
  AOI21_X1  g491(.A(KEYINPUT107), .B1(new_n915), .B2(new_n907), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g494(.A(KEYINPUT108), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n596), .A2(new_n567), .A3(new_n597), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n567), .B1(new_n596), .B2(new_n597), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n920), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(G290), .A2(G288), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n925), .A2(KEYINPUT108), .A3(new_n921), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n741), .B(G166), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n924), .A2(new_n926), .A3(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(new_n927), .ZN(new_n929));
  OAI211_X1 g504(.A(new_n929), .B(new_n920), .C1(new_n923), .C2(new_n922), .ZN(new_n930));
  AOI21_X1  g505(.A(KEYINPUT110), .B1(new_n928), .B2(new_n930), .ZN(new_n931));
  OR3_X1    g506(.A1(new_n931), .A2(KEYINPUT109), .A3(KEYINPUT42), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n928), .A2(new_n930), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT109), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n934), .B(KEYINPUT42), .C1(KEYINPUT109), .C2(new_n931), .ZN(new_n935));
  NOR2_X1   g510(.A1(G299), .A2(new_n605), .ZN(new_n936));
  AOI22_X1  g511(.A1(new_n557), .A2(new_n560), .B1(new_n600), .B2(new_n604), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  OAI21_X1  g515(.A(new_n940), .B1(new_n936), .B2(new_n937), .ZN(new_n941));
  INV_X1    g516(.A(new_n937), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n611), .A2(new_n560), .A3(new_n557), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(new_n943), .A3(KEYINPUT41), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n941), .A2(new_n944), .ZN(new_n945));
  XNOR2_X1  g520(.A(new_n867), .B(new_n615), .ZN(new_n946));
  MUX2_X1   g521(.A(new_n939), .B(new_n945), .S(new_n946), .Z(new_n947));
  AND3_X1   g522(.A1(new_n932), .A2(new_n935), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n947), .B1(new_n932), .B2(new_n935), .ZN(new_n949));
  OAI21_X1  g524(.A(G868), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(new_n866), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n950), .B1(G868), .B2(new_n951), .ZN(G295));
  OAI21_X1  g527(.A(new_n950), .B1(G868), .B2(new_n951), .ZN(G331));
  INV_X1    g528(.A(new_n530), .ZN(new_n954));
  NAND3_X1  g529(.A1(G168), .A2(new_n528), .A3(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n519), .B(new_n520), .C1(new_n529), .C2(new_n530), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n867), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  AOI21_X1  g532(.A(new_n867), .B1(new_n956), .B2(new_n955), .ZN(new_n958));
  OAI21_X1  g533(.A(new_n938), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n955), .A2(new_n956), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n868), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n867), .A2(new_n955), .A3(new_n956), .ZN(new_n962));
  NAND4_X1  g537(.A1(new_n961), .A2(new_n941), .A3(new_n944), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n959), .A2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n933), .A2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(G37), .ZN(new_n966));
  NAND4_X1  g541(.A1(new_n928), .A2(new_n930), .A3(new_n959), .A4(new_n963), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n965), .A2(new_n966), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT43), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT43), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n965), .A2(new_n970), .A3(new_n966), .A4(new_n967), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n969), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(KEYINPUT44), .B1(new_n970), .B2(KEYINPUT111), .ZN(new_n973));
  XNOR2_X1  g548(.A(new_n972), .B(new_n973), .ZN(G397));
  INV_X1    g549(.A(KEYINPUT124), .ZN(new_n975));
  INV_X1    g550(.A(G2084), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n494), .A2(new_n496), .ZN(new_n977));
  AND2_X1   g552(.A1(new_n485), .A2(new_n489), .ZN(new_n978));
  AOI21_X1  g553(.A(G1384), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT50), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  OAI21_X1  g556(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n982));
  INV_X1    g557(.A(G40), .ZN(new_n983));
  NOR3_X1   g558(.A1(new_n468), .A2(new_n471), .A3(new_n983), .ZN(new_n984));
  AND4_X1   g559(.A1(new_n976), .A2(new_n981), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  INV_X1    g560(.A(G1384), .ZN(new_n986));
  AOI21_X1  g561(.A(KEYINPUT45), .B1(new_n879), .B2(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(G160), .A2(G40), .ZN(new_n988));
  OAI21_X1  g563(.A(KEYINPUT118), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT118), .ZN(new_n990));
  OAI211_X1 g565(.A(new_n990), .B(new_n984), .C1(new_n979), .C2(KEYINPUT45), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n879), .A2(KEYINPUT45), .A3(new_n986), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G1966), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n985), .B1(new_n993), .B2(new_n994), .ZN(new_n995));
  INV_X1    g570(.A(G8), .ZN(new_n996));
  OAI21_X1  g571(.A(new_n975), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n991), .A2(new_n992), .ZN(new_n998));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n999), .B1(G164), .B2(G1384), .ZN(new_n1000));
  AOI21_X1  g575(.A(new_n990), .B1(new_n1000), .B2(new_n984), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n994), .B1(new_n998), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(new_n985), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1004), .A2(KEYINPUT124), .A3(G8), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G168), .A2(new_n996), .ZN(new_n1006));
  NOR2_X1   g581(.A1(new_n1006), .A2(KEYINPUT51), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n997), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g583(.A(KEYINPUT125), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n997), .A2(new_n1005), .A3(KEYINPUT125), .A4(new_n1007), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT51), .ZN(new_n1012));
  AOI211_X1 g587(.A(new_n1012), .B(new_n996), .C1(new_n995), .C2(G168), .ZN(new_n1013));
  INV_X1    g588(.A(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n1010), .A2(new_n1011), .A3(new_n1014), .ZN(new_n1015));
  AND2_X1   g590(.A1(new_n1004), .A2(new_n1006), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1015), .A2(new_n1017), .ZN(new_n1018));
  NAND4_X1  g593(.A1(new_n1000), .A2(new_n992), .A3(new_n796), .A4(new_n984), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1020), .A2(G2078), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1000), .A2(new_n992), .A3(new_n984), .A4(new_n1022), .ZN(new_n1023));
  AND3_X1   g598(.A1(new_n981), .A2(new_n982), .A3(new_n984), .ZN(new_n1024));
  OAI211_X1 g599(.A(new_n1021), .B(new_n1023), .C1(G1961), .C2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(G171), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n879), .A2(new_n986), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n988), .B1(new_n1027), .B2(KEYINPUT50), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n1028), .A2(new_n981), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1029), .A2(new_n804), .B1(new_n1019), .B2(new_n1020), .ZN(new_n1030));
  NAND4_X1  g605(.A1(new_n989), .A2(new_n991), .A3(new_n992), .A4(new_n1022), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n1030), .A2(G301), .A3(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1026), .A2(new_n1032), .A3(KEYINPUT54), .ZN(new_n1033));
  NAND2_X1  g608(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1034));
  OR2_X1    g609(.A1(KEYINPUT114), .A2(KEYINPUT55), .ZN(new_n1035));
  AOI22_X1  g610(.A1(G303), .A2(G8), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n503), .A2(new_n504), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n499), .B1(new_n501), .B2(new_n502), .ZN(new_n1038));
  OAI211_X1 g613(.A(G8), .B(new_n1035), .C1(new_n1037), .C2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1036), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1000), .A2(new_n984), .ZN(new_n1042));
  INV_X1    g617(.A(new_n992), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n750), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(G2090), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1028), .A2(new_n1045), .A3(new_n981), .ZN(new_n1046));
  AOI211_X1 g621(.A(new_n996), .B(new_n1041), .C1(new_n1044), .C2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT116), .B(new_n984), .C1(new_n979), .C2(new_n980), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(new_n981), .ZN(new_n1049));
  AOI21_X1  g624(.A(KEYINPUT116), .B1(new_n982), .B2(new_n984), .ZN(new_n1050));
  NOR3_X1   g625(.A1(new_n1049), .A2(new_n1050), .A3(G2090), .ZN(new_n1051));
  INV_X1    g626(.A(new_n1044), .ZN(new_n1052));
  OAI21_X1  g627(.A(G8), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1047), .B1(new_n1053), .B2(new_n1041), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT49), .ZN(new_n1055));
  INV_X1    g630(.A(G1981), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n740), .A2(new_n579), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1057), .B2(new_n572), .ZN(new_n1058));
  AOI211_X1 g633(.A(G1981), .B(new_n571), .C1(new_n740), .C2(new_n579), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1055), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(G305), .A2(G1981), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n741), .A2(new_n1056), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1061), .A2(new_n1062), .A3(KEYINPUT49), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n996), .B1(new_n979), .B2(new_n984), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1060), .A2(new_n1063), .A3(new_n1064), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n567), .A2(G1976), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1066), .A2(new_n1064), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT52), .ZN(new_n1068));
  OAI21_X1  g643(.A(new_n1068), .B1(new_n567), .B2(G1976), .ZN(new_n1069));
  NOR2_X1   g644(.A1(new_n1067), .A2(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1070), .B1(KEYINPUT52), .B2(new_n1067), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT117), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1065), .A2(new_n1071), .A3(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1072), .B1(new_n1065), .B2(new_n1071), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1033), .B(new_n1054), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT54), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1025), .A2(G171), .ZN(new_n1077));
  AOI21_X1  g652(.A(G301), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT126), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT126), .B(new_n1076), .C1(new_n1077), .C2(new_n1078), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1075), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  XOR2_X1   g658(.A(KEYINPUT122), .B(KEYINPUT61), .Z(new_n1084));
  OAI21_X1  g659(.A(new_n836), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1085));
  XNOR2_X1  g660(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1086));
  XNOR2_X1  g661(.A(new_n1086), .B(new_n786), .ZN(new_n1087));
  NAND4_X1  g662(.A1(new_n1000), .A2(new_n992), .A3(new_n984), .A4(new_n1087), .ZN(new_n1088));
  INV_X1    g663(.A(new_n560), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT57), .B1(new_n1089), .B2(new_n556), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT57), .ZN(new_n1091));
  AOI22_X1  g666(.A1(new_n547), .A2(G651), .B1(new_n554), .B2(G91), .ZN(new_n1092));
  NAND4_X1  g667(.A1(new_n560), .A2(new_n1091), .A3(new_n1092), .A4(new_n553), .ZN(new_n1093));
  AND2_X1   g668(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1085), .A2(new_n1088), .A3(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1094), .B1(new_n1085), .B2(new_n1088), .ZN(new_n1096));
  OAI21_X1  g671(.A(new_n1084), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT123), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT123), .B(new_n1084), .C1(new_n1095), .C2(new_n1096), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT60), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n813), .B1(new_n1028), .B2(new_n981), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n979), .A2(new_n984), .ZN(new_n1103));
  NOR2_X1   g678(.A1(new_n1103), .A2(G2067), .ZN(new_n1104));
  OAI21_X1  g679(.A(new_n611), .B1(new_n1102), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n1104), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1106), .B(new_n605), .C1(new_n1024), .C2(new_n813), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1101), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT59), .ZN(new_n1109));
  INV_X1    g684(.A(G1996), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1000), .A2(new_n992), .A3(new_n1110), .A4(new_n984), .ZN(new_n1111));
  XOR2_X1   g686(.A(KEYINPUT58), .B(G1341), .Z(new_n1112));
  NAND2_X1  g687(.A1(new_n1103), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1109), .B1(new_n1114), .B2(new_n538), .ZN(new_n1115));
  INV_X1    g690(.A(new_n538), .ZN(new_n1116));
  AOI211_X1 g691(.A(KEYINPUT59), .B(new_n1116), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1117));
  NOR2_X1   g692(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  NOR4_X1   g693(.A1(new_n1102), .A2(KEYINPUT60), .A3(new_n605), .A4(new_n1104), .ZN(new_n1119));
  NOR3_X1   g694(.A1(new_n1108), .A2(new_n1118), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(new_n1096), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1085), .A2(new_n1094), .A3(new_n1088), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1121), .A2(KEYINPUT61), .A3(new_n1122), .ZN(new_n1123));
  NAND4_X1  g698(.A1(new_n1099), .A2(new_n1100), .A3(new_n1120), .A4(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(new_n1105), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1122), .B1(new_n1096), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  OAI211_X1 g703(.A(KEYINPUT121), .B(new_n1122), .C1(new_n1096), .C2(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1124), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1018), .A2(new_n1083), .A3(new_n1131), .ZN(new_n1132));
  NOR3_X1   g707(.A1(new_n995), .A2(new_n996), .A3(G286), .ZN(new_n1133));
  OAI211_X1 g708(.A(new_n1054), .B(new_n1133), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1134));
  XOR2_X1   g709(.A(KEYINPUT119), .B(KEYINPUT63), .Z(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  AND2_X1   g711(.A1(new_n1065), .A2(new_n1071), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NOR2_X1   g713(.A1(new_n1047), .A2(new_n1138), .ZN(new_n1139));
  AND2_X1   g714(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n1041), .B1(new_n1140), .B2(new_n996), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1137), .A2(new_n1139), .A3(new_n1133), .A4(new_n1141), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1047), .A2(new_n1065), .A3(new_n1071), .ZN(new_n1143));
  NOR2_X1   g718(.A1(G288), .A2(G1976), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1059), .B1(new_n1065), .B2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(new_n1064), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1143), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT115), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT115), .ZN(new_n1149));
  OAI211_X1 g724(.A(new_n1149), .B(new_n1143), .C1(new_n1145), .C2(new_n1146), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1136), .A2(new_n1142), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  OAI211_X1 g726(.A(new_n1054), .B(new_n1078), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1152));
  INV_X1    g727(.A(new_n1152), .ZN(new_n1153));
  AOI21_X1  g728(.A(new_n1013), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1154));
  AOI21_X1  g729(.A(new_n1016), .B1(new_n1154), .B2(new_n1011), .ZN(new_n1155));
  INV_X1    g730(.A(KEYINPUT62), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1153), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AOI211_X1 g732(.A(KEYINPUT62), .B(new_n1016), .C1(new_n1154), .C2(new_n1011), .ZN(new_n1158));
  OAI211_X1 g733(.A(new_n1132), .B(new_n1151), .C1(new_n1157), .C2(new_n1158), .ZN(new_n1159));
  NOR2_X1   g734(.A1(new_n1000), .A2(new_n988), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1160), .A2(new_n1110), .ZN(new_n1161));
  NOR2_X1   g736(.A1(new_n1161), .A2(new_n848), .ZN(new_n1162));
  XNOR2_X1  g737(.A(new_n1162), .B(KEYINPUT113), .ZN(new_n1163));
  INV_X1    g738(.A(G2067), .ZN(new_n1164));
  XNOR2_X1  g739(.A(new_n829), .B(new_n1164), .ZN(new_n1165));
  INV_X1    g740(.A(new_n883), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n1165), .B1(new_n1110), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1163), .B1(new_n1160), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1160), .ZN(new_n1169));
  XOR2_X1   g744(.A(new_n727), .B(new_n734), .Z(new_n1170));
  OAI21_X1  g745(.A(new_n1168), .B1(new_n1169), .B2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n713), .A2(new_n718), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT112), .ZN(new_n1173));
  NOR2_X1   g748(.A1(G290), .A2(G1986), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1172), .A2(new_n1173), .A3(new_n1174), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1169), .B(new_n1175), .C1(new_n1173), .C2(new_n1172), .ZN(new_n1176));
  NOR2_X1   g751(.A1(new_n1171), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g752(.A1(new_n1159), .A2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1174), .A2(new_n1160), .ZN(new_n1179));
  XOR2_X1   g754(.A(new_n1179), .B(KEYINPUT48), .Z(new_n1180));
  NOR2_X1   g755(.A1(new_n1171), .A2(new_n1180), .ZN(new_n1181));
  NOR2_X1   g756(.A1(new_n727), .A2(new_n734), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1168), .A2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n830), .A2(new_n1164), .ZN(new_n1184));
  AOI21_X1  g759(.A(new_n1169), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1169), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1187));
  OR2_X1    g762(.A1(new_n1161), .A2(KEYINPUT46), .ZN(new_n1188));
  AOI21_X1  g763(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT47), .ZN(new_n1190));
  NOR3_X1   g765(.A1(new_n1181), .A2(new_n1185), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g766(.A1(new_n1178), .A2(new_n1191), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g767(.A1(G227), .A2(new_n461), .ZN(new_n1194));
  OAI21_X1  g768(.A(new_n1194), .B1(new_n708), .B2(new_n709), .ZN(new_n1195));
  AOI21_X1  g769(.A(new_n1195), .B1(new_n664), .B2(new_n671), .ZN(new_n1196));
  NAND3_X1  g770(.A1(new_n972), .A2(new_n918), .A3(new_n1196), .ZN(G225));
  INV_X1    g771(.A(KEYINPUT127), .ZN(new_n1198));
  XNOR2_X1  g772(.A(G225), .B(new_n1198), .ZN(G308));
endmodule


