//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n209, new_n210, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1223, new_n1224,
    new_n1226, new_n1227, new_n1228, new_n1229, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1290, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  NOR2_X1   g0007(.A1(G97), .A2(G107), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g0009(.A1(new_n209), .A2(G87), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0011(.A1(G1), .A2(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n203), .A2(new_n205), .ZN(new_n216));
  INV_X1    g0016(.A(G50), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G13), .ZN(new_n219));
  INV_X1    g0019(.A(G20), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g0022(.A(KEYINPUT66), .B(G238), .ZN(new_n223));
  NOR2_X1   g0023(.A1(new_n223), .A2(new_n202), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n212), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n215), .B(new_n222), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XOR2_X1   g0034(.A(KEYINPUT2), .B(G226), .Z(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n236), .B(new_n239), .Z(G358));
  XOR2_X1   g0040(.A(G87), .B(G97), .Z(new_n241));
  XNOR2_X1  g0041(.A(G107), .B(G116), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n217), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n202), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n243), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(KEYINPUT77), .ZN(new_n250));
  INV_X1    g0050(.A(KEYINPUT69), .ZN(new_n251));
  NOR2_X1   g0051(.A1(new_n251), .A2(G58), .ZN(new_n252));
  NOR2_X1   g0052(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n253));
  OAI21_X1  g0053(.A(G68), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n220), .B1(new_n206), .B2(new_n254), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  INV_X1    g0057(.A(G159), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n265), .A2(KEYINPUT7), .A3(new_n220), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  AOI21_X1  g0067(.A(KEYINPUT7), .B1(new_n265), .B2(new_n220), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(new_n260), .B1(new_n202), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT16), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n219), .B1(new_n212), .B2(new_n261), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  AND3_X1   g0074(.A1(new_n262), .A2(new_n264), .A3(KEYINPUT73), .ZN(new_n275));
  AOI21_X1  g0075(.A(KEYINPUT73), .B1(new_n262), .B2(new_n264), .ZN(new_n276));
  NOR2_X1   g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  AOI21_X1  g0077(.A(KEYINPUT7), .B1(new_n277), .B2(new_n220), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n266), .A2(KEYINPUT74), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT74), .ZN(new_n280));
  NAND4_X1  g0080(.A1(new_n265), .A2(new_n280), .A3(KEYINPUT7), .A4(new_n220), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n279), .A2(new_n281), .ZN(new_n282));
  OAI21_X1  g0082(.A(G68), .B1(new_n278), .B2(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(KEYINPUT75), .B1(new_n255), .B2(new_n259), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n251), .A2(G58), .ZN(new_n286));
  AOI21_X1  g0086(.A(new_n202), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  OAI21_X1  g0087(.A(G20), .B1(new_n287), .B2(new_n216), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT75), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n289), .C1(new_n258), .C2(new_n257), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g0091(.A1(new_n283), .A2(new_n291), .A3(KEYINPUT16), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT76), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  NOR3_X1   g0094(.A1(new_n275), .A2(new_n276), .A3(G20), .ZN(new_n295));
  OAI211_X1 g0095(.A(new_n279), .B(new_n281), .C1(new_n295), .C2(KEYINPUT7), .ZN(new_n296));
  AOI22_X1  g0096(.A1(new_n296), .A2(G68), .B1(new_n284), .B2(new_n290), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT76), .A3(KEYINPUT16), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n274), .B1(new_n294), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G1), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(KEYINPUT67), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT67), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G1), .ZN(new_n303));
  AND2_X1   g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g0104(.A(new_n273), .B1(new_n304), .B2(G20), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(KEYINPUT8), .A2(G58), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n285), .A2(new_n286), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n307), .B1(new_n308), .B2(KEYINPUT8), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g0110(.A1(new_n304), .A2(G13), .A3(G20), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n310), .B1(new_n309), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n250), .B1(new_n299), .B2(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(new_n273), .ZN(new_n316));
  AOI21_X1  g0116(.A(new_n316), .B1(new_n270), .B2(new_n271), .ZN(new_n317));
  AOI21_X1  g0117(.A(KEYINPUT76), .B1(new_n297), .B2(KEYINPUT16), .ZN(new_n318));
  AND4_X1   g0118(.A1(KEYINPUT76), .A2(new_n283), .A3(new_n291), .A4(KEYINPUT16), .ZN(new_n319));
  OAI21_X1  g0119(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n320), .A2(KEYINPUT77), .A3(new_n313), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n265), .A2(G1698), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n322), .A2(G223), .B1(G33), .B2(G87), .ZN(new_n323));
  INV_X1    g0123(.A(G226), .ZN(new_n324));
  INV_X1    g0124(.A(G1698), .ZN(new_n325));
  NOR2_X1   g0125(.A1(new_n265), .A2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI21_X1  g0127(.A(new_n323), .B1(new_n324), .B2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(G41), .ZN(new_n329));
  OAI211_X1 g0129(.A(G1), .B(G13), .C1(new_n261), .C2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g0132(.A(G45), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n329), .A2(new_n333), .ZN(new_n334));
  NAND3_X1  g0134(.A1(new_n334), .A2(new_n300), .A3(G274), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n331), .B1(new_n304), .B2(new_n334), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n336), .B1(new_n337), .B2(G232), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n332), .A2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(G169), .ZN(new_n340));
  INV_X1    g0140(.A(G179), .ZN(new_n341));
  OAI21_X1  g0141(.A(new_n340), .B1(new_n341), .B2(new_n339), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n315), .A2(new_n321), .A3(new_n342), .ZN(new_n343));
  OR2_X1    g0143(.A1(new_n343), .A2(KEYINPUT18), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n339), .A2(G200), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n332), .A2(G190), .A3(new_n338), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n320), .A2(new_n313), .A3(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT17), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  NAND4_X1  g0150(.A1(new_n320), .A2(new_n347), .A3(KEYINPUT17), .A4(new_n313), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(new_n352), .ZN(new_n353));
  NAND2_X1  g0153(.A1(new_n343), .A2(KEYINPUT18), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n344), .A2(new_n353), .A3(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n355), .B(KEYINPUT78), .Z(new_n356));
  NAND2_X1  g0156(.A1(new_n312), .A2(new_n202), .ZN(new_n357));
  XNOR2_X1  g0157(.A(new_n357), .B(KEYINPUT12), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n261), .A2(G20), .ZN(new_n359));
  INV_X1    g0159(.A(new_n359), .ZN(new_n360));
  INV_X1    g0160(.A(G77), .ZN(new_n361));
  OAI22_X1  g0161(.A1(new_n360), .A2(new_n361), .B1(new_n220), .B2(G68), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n257), .A2(new_n217), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n273), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  XNOR2_X1  g0164(.A(new_n364), .B(KEYINPUT11), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n305), .A2(G68), .ZN(new_n366));
  AND3_X1   g0166(.A1(new_n358), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g0167(.A(new_n367), .B(KEYINPUT71), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT13), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n262), .A2(new_n264), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(G232), .A3(G1698), .ZN(new_n371));
  NAND2_X1  g0171(.A1(G33), .A2(G97), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n325), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n371), .B(new_n372), .C1(new_n373), .C2(new_n324), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n331), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n336), .B1(new_n337), .B2(G238), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n369), .A3(new_n376), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT14), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n380), .A2(new_n381), .A3(G169), .ZN(new_n382));
  INV_X1    g0182(.A(new_n379), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n383), .A2(new_n377), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G179), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n382), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g0186(.A(new_n381), .B1(new_n380), .B2(G169), .ZN(new_n387));
  OAI21_X1  g0187(.A(new_n368), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n384), .A2(G190), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n380), .A2(G200), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n389), .A2(new_n390), .A3(new_n367), .ZN(new_n391));
  AOI21_X1  g0191(.A(KEYINPUT72), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n322), .A2(G222), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT68), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n393), .B(new_n394), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n326), .A2(G223), .B1(G77), .B2(new_n265), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n330), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n337), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n335), .B1(new_n398), .B2(new_n324), .ZN(new_n399));
  OR2_X1    g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n309), .A2(new_n359), .ZN(new_n401));
  INV_X1    g0201(.A(G150), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n401), .B1(new_n402), .B2(new_n257), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n220), .B1(new_n216), .B2(new_n217), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n273), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NOR2_X1   g0205(.A1(new_n311), .A2(G50), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n406), .B1(G50), .B2(new_n305), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n408), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n400), .A2(G200), .B1(KEYINPUT9), .B2(new_n409), .ZN(new_n410));
  NOR2_X1   g0210(.A1(new_n397), .A2(new_n399), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT9), .ZN(new_n412));
  AOI22_X1  g0212(.A1(new_n411), .A2(G190), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  XNOR2_X1  g0214(.A(new_n414), .B(KEYINPUT10), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n408), .B1(new_n411), .B2(G169), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n416), .A2(KEYINPUT70), .B1(new_n341), .B2(new_n411), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n417), .B1(KEYINPUT70), .B2(new_n416), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n415), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n388), .A2(new_n391), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT72), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n305), .A2(G77), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G77), .B2(new_n311), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT8), .B(G58), .ZN(new_n425));
  OAI22_X1  g0225(.A1(new_n425), .A2(new_n257), .B1(new_n220), .B2(new_n361), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  NOR2_X1   g0227(.A1(new_n427), .A2(new_n360), .ZN(new_n428));
  OAI21_X1  g0228(.A(new_n273), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  OR2_X1    g0230(.A1(new_n424), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n370), .A2(G232), .A3(new_n325), .ZN(new_n432));
  INV_X1    g0232(.A(G107), .ZN(new_n433));
  OAI221_X1 g0233(.A(new_n432), .B1(new_n433), .B2(new_n370), .C1(new_n327), .C2(new_n223), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n434), .A2(new_n331), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n336), .B1(new_n337), .B2(G244), .ZN(new_n436));
  NAND2_X1  g0236(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(G200), .ZN(new_n438));
  INV_X1    g0238(.A(G190), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n438), .B1(new_n439), .B2(new_n437), .ZN(new_n440));
  NOR2_X1   g0240(.A1(new_n424), .A2(new_n430), .ZN(new_n441));
  INV_X1    g0241(.A(G169), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n441), .B1(new_n437), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n435), .A2(new_n341), .A3(new_n436), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n440), .A2(new_n445), .ZN(new_n446));
  NOR4_X1   g0246(.A1(new_n392), .A2(new_n419), .A3(new_n422), .A4(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n356), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G33), .A2(G283), .ZN(new_n450));
  INV_X1    g0250(.A(G97), .ZN(new_n451));
  OAI211_X1 g0251(.A(new_n450), .B(new_n220), .C1(G33), .C2(new_n451), .ZN(new_n452));
  OAI211_X1 g0252(.A(new_n452), .B(new_n273), .C1(new_n220), .C2(G116), .ZN(new_n453));
  XOR2_X1   g0253(.A(new_n453), .B(KEYINPUT20), .Z(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n312), .A2(new_n455), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n304), .A2(G33), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n311), .A2(new_n316), .A3(new_n457), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n454), .B(new_n456), .C1(new_n455), .C2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT5), .ZN(new_n460));
  OAI211_X1 g0260(.A(new_n330), .B(G274), .C1(new_n460), .C2(G41), .ZN(new_n461));
  AND3_X1   g0261(.A1(new_n301), .A2(new_n303), .A3(G45), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(KEYINPUT5), .B2(new_n329), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n461), .B1(new_n463), .B2(KEYINPUT82), .ZN(new_n464));
  OAI21_X1  g0264(.A(new_n464), .B1(KEYINPUT82), .B2(new_n463), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n326), .A2(G264), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n370), .A2(G257), .A3(new_n325), .ZN(new_n467));
  INV_X1    g0267(.A(G303), .ZN(new_n468));
  OAI211_X1 g0268(.A(new_n466), .B(new_n467), .C1(new_n468), .C2(new_n370), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(new_n331), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n460), .A2(G41), .ZN(new_n471));
  OAI211_X1 g0271(.A(G270), .B(new_n330), .C1(new_n463), .C2(new_n471), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n465), .A2(new_n470), .A3(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n459), .A2(new_n473), .A3(G169), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT21), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(KEYINPUT83), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n474), .A2(new_n475), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT83), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n473), .A2(KEYINPUT21), .A3(G169), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n465), .A2(new_n470), .A3(G179), .A4(new_n472), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(new_n459), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n459), .B1(new_n473), .B2(G200), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n484), .B1(new_n439), .B2(new_n473), .ZN(new_n485));
  AND4_X1   g0285(.A1(new_n476), .A2(new_n479), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n433), .A2(KEYINPUT6), .A3(G97), .ZN(new_n487));
  NOR2_X1   g0287(.A1(new_n451), .A2(new_n433), .ZN(new_n488));
  NOR2_X1   g0288(.A1(new_n488), .A2(new_n208), .ZN(new_n489));
  OAI21_X1  g0289(.A(new_n487), .B1(new_n489), .B2(KEYINPUT6), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(G20), .B1(G77), .B2(new_n256), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n269), .B2(new_n433), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n492), .A2(new_n273), .B1(new_n451), .B2(new_n312), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n458), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g0295(.A1(new_n311), .A2(new_n457), .A3(KEYINPUT79), .A4(new_n316), .ZN(new_n496));
  AND2_X1   g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(G97), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n500));
  INV_X1    g0300(.A(G244), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n500), .B1(new_n373), .B2(new_n501), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n322), .B(G244), .C1(KEYINPUT80), .C2(KEYINPUT4), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n326), .A2(G250), .ZN(new_n504));
  NAND4_X1  g0304(.A1(new_n502), .A2(new_n503), .A3(new_n450), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n331), .ZN(new_n506));
  OAI211_X1 g0306(.A(G257), .B(new_n330), .C1(new_n463), .C2(new_n471), .ZN(new_n507));
  AND3_X1   g0307(.A1(new_n506), .A2(new_n465), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n499), .B1(new_n508), .B2(G190), .ZN(new_n509));
  AND2_X1   g0309(.A1(new_n465), .A2(new_n507), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n506), .A2(KEYINPUT81), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n512), .B1(new_n505), .B2(new_n331), .ZN(new_n513));
  OAI21_X1  g0313(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n514), .A2(G200), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n509), .A2(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n510), .A2(new_n506), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n517), .A2(new_n442), .B1(new_n498), .B2(new_n493), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n341), .B(new_n510), .C1(new_n511), .C2(new_n513), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AND2_X1   g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n322), .A2(G238), .B1(G33), .B2(G116), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n522), .B1(new_n501), .B2(new_n327), .ZN(new_n523));
  INV_X1    g0323(.A(G274), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n462), .A2(new_n524), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n462), .A2(G250), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(new_n331), .ZN(new_n527));
  AOI22_X1  g0327(.A1(new_n523), .A2(new_n331), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(new_n427), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n495), .A2(new_n529), .A3(new_n496), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n370), .A2(new_n220), .A3(G68), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT19), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n220), .B1(new_n372), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(G87), .B2(new_n209), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n532), .B1(new_n360), .B2(new_n451), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(new_n534), .A3(new_n535), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n536), .A2(new_n273), .B1(new_n312), .B2(new_n427), .ZN(new_n537));
  AOI22_X1  g0337(.A1(new_n528), .A2(new_n341), .B1(new_n530), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n523), .A2(new_n331), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n525), .B(new_n330), .C1(G250), .C2(new_n462), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n442), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n541), .A2(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n528), .A2(G190), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n495), .A2(G87), .A3(new_n496), .ZN(new_n546));
  AND2_X1   g0346(.A1(new_n546), .A2(new_n537), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n544), .A2(new_n545), .A3(new_n547), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n370), .A2(new_n220), .A3(G87), .ZN(new_n550));
  XNOR2_X1  g0350(.A(new_n550), .B(KEYINPUT22), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT23), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n220), .B2(G107), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n433), .A2(KEYINPUT23), .A3(G20), .ZN(new_n554));
  AOI22_X1  g0354(.A1(new_n553), .A2(new_n554), .B1(new_n359), .B2(G116), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n551), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(KEYINPUT24), .ZN(new_n557));
  INV_X1    g0357(.A(KEYINPUT24), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n551), .A2(new_n558), .A3(new_n555), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n557), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n273), .ZN(new_n561));
  AOI22_X1  g0361(.A1(new_n322), .A2(G250), .B1(G33), .B2(G294), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n370), .A2(G257), .A3(G1698), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n330), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n463), .A2(new_n471), .ZN(new_n565));
  NOR2_X1   g0365(.A1(new_n565), .A2(new_n331), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n564), .B1(new_n566), .B2(G264), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n567), .A2(new_n465), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n568), .A2(G200), .ZN(new_n569));
  NOR2_X1   g0369(.A1(new_n311), .A2(G107), .ZN(new_n570));
  OR2_X1    g0370(.A1(new_n570), .A2(KEYINPUT25), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n570), .A2(KEYINPUT25), .ZN(new_n572));
  AOI22_X1  g0372(.A1(new_n497), .A2(G107), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n567), .A2(G190), .A3(new_n465), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n561), .A2(new_n569), .A3(new_n573), .A4(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n568), .A2(new_n442), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n567), .A2(new_n341), .A3(new_n465), .ZN(new_n577));
  INV_X1    g0377(.A(new_n573), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n316), .B1(new_n557), .B2(new_n559), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n576), .B(new_n577), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  AND3_X1   g0380(.A1(new_n549), .A2(new_n575), .A3(new_n580), .ZN(new_n581));
  AND4_X1   g0381(.A1(new_n449), .A2(new_n486), .A3(new_n521), .A4(new_n581), .ZN(G372));
  NAND2_X1  g0382(.A1(new_n543), .A2(new_n548), .ZN(new_n583));
  OAI21_X1  g0383(.A(KEYINPUT26), .B1(new_n520), .B2(new_n583), .ZN(new_n584));
  AND2_X1   g0384(.A1(new_n547), .A2(new_n545), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n540), .A2(KEYINPUT84), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n539), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n588), .A2(G200), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n588), .A2(new_n442), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n585), .A2(new_n589), .B1(new_n590), .B2(new_n538), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT26), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n591), .A2(new_n592), .A3(new_n519), .A4(new_n518), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n590), .A2(new_n538), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n584), .A2(new_n593), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(KEYINPUT85), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT85), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n584), .A2(new_n593), .A3(new_n597), .A4(new_n594), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n516), .A2(new_n520), .A3(new_n575), .A4(new_n591), .ZN(new_n599));
  INV_X1    g0399(.A(new_n599), .ZN(new_n600));
  AOI22_X1  g0400(.A1(new_n478), .A2(new_n477), .B1(new_n482), .B2(new_n459), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(new_n476), .A3(new_n580), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n596), .A2(new_n598), .A3(new_n603), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n449), .A2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n445), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n391), .A2(new_n606), .ZN(new_n607));
  AOI21_X1  g0407(.A(new_n352), .B1(new_n388), .B2(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n342), .B1(new_n299), .B2(new_n314), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(KEYINPUT18), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n415), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n611), .A2(new_n418), .ZN(new_n612));
  XNOR2_X1  g0412(.A(new_n612), .B(KEYINPUT86), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n605), .A2(new_n613), .ZN(G369));
  AND2_X1   g0414(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n486), .A2(KEYINPUT87), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n220), .A2(G13), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n304), .A2(new_n617), .ZN(new_n618));
  OR2_X1    g0418(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n618), .A2(KEYINPUT27), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n619), .A2(G213), .A3(new_n620), .ZN(new_n621));
  INV_X1    g0421(.A(G343), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n459), .A2(new_n623), .ZN(new_n624));
  OR3_X1    g0424(.A1(new_n615), .A2(new_n616), .A3(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n601), .A2(new_n476), .A3(new_n624), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n580), .A2(new_n623), .ZN(new_n627));
  INV_X1    g0427(.A(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n623), .B1(new_n579), .B2(new_n578), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n575), .A2(new_n629), .ZN(new_n630));
  INV_X1    g0430(.A(new_n580), .ZN(new_n631));
  OAI21_X1  g0431(.A(new_n628), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n632), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n625), .A2(G330), .A3(new_n626), .A4(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n601), .A2(new_n476), .ZN(new_n635));
  INV_X1    g0435(.A(new_n623), .ZN(new_n636));
  NAND4_X1  g0436(.A1(new_n635), .A2(new_n630), .A3(new_n580), .A4(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n637), .A2(new_n628), .ZN(new_n638));
  INV_X1    g0438(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n634), .A2(new_n639), .ZN(G399));
  INV_X1    g0440(.A(new_n213), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(G41), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR3_X1   g0443(.A1(new_n209), .A2(G87), .A3(G116), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n643), .A2(G1), .A3(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n218), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n645), .B1(new_n646), .B2(new_n643), .ZN(new_n647));
  XNOR2_X1  g0447(.A(new_n647), .B(KEYINPUT28), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT88), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n602), .A2(new_n649), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n601), .A2(KEYINPUT88), .A3(new_n476), .A4(new_n580), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n599), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(new_n591), .ZN(new_n653));
  OAI21_X1  g0453(.A(KEYINPUT26), .B1(new_n653), .B2(new_n520), .ZN(new_n654));
  NAND4_X1  g0454(.A1(new_n549), .A2(new_n592), .A3(new_n519), .A4(new_n518), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(new_n594), .A3(new_n655), .ZN(new_n656));
  OAI211_X1 g0456(.A(KEYINPUT29), .B(new_n636), .C1(new_n652), .C2(new_n656), .ZN(new_n657));
  AOI22_X1  g0457(.A1(new_n595), .A2(KEYINPUT85), .B1(new_n600), .B2(new_n602), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n623), .B1(new_n658), .B2(new_n598), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n657), .B1(new_n659), .B2(KEYINPUT29), .ZN(new_n660));
  INV_X1    g0460(.A(G330), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n567), .A2(new_n528), .ZN(new_n662));
  INV_X1    g0462(.A(new_n481), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n508), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT30), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  AOI21_X1  g0466(.A(G179), .B1(new_n567), .B2(new_n465), .ZN(new_n667));
  NAND4_X1  g0467(.A1(new_n514), .A2(new_n473), .A3(new_n588), .A4(new_n667), .ZN(new_n668));
  NAND4_X1  g0468(.A1(new_n662), .A2(new_n663), .A3(new_n508), .A4(KEYINPUT30), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n666), .A2(new_n668), .A3(new_n669), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n671));
  AOI21_X1  g0471(.A(KEYINPUT31), .B1(new_n670), .B2(new_n623), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n521), .A2(new_n486), .A3(new_n581), .A4(new_n636), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n661), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n660), .A2(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(KEYINPUT89), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n660), .A2(KEYINPUT89), .A3(new_n676), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n648), .B1(new_n681), .B2(G1), .ZN(G364));
  AND2_X1   g0482(.A1(new_n625), .A2(new_n626), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(G330), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n625), .A2(G330), .A3(new_n626), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n300), .B1(new_n617), .B2(G45), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n643), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n684), .A2(new_n688), .ZN(new_n689));
  NOR2_X1   g0489(.A1(G13), .A2(G33), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G20), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  OR2_X1    g0493(.A1(new_n683), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n219), .B1(G20), .B2(new_n442), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n220), .A2(G179), .ZN(new_n697));
  NOR2_X1   g0497(.A1(G190), .A2(G200), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g0499(.A1(new_n699), .A2(KEYINPUT92), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(KEYINPUT92), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  INV_X1    g0502(.A(new_n702), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G159), .ZN(new_n704));
  XNOR2_X1  g0504(.A(new_n704), .B(KEYINPUT32), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n220), .A2(new_n341), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n706), .A2(G200), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n707), .A2(G190), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n439), .A2(G200), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n709), .A2(new_n341), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(G20), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n708), .A2(G68), .B1(new_n711), .B2(G97), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n697), .A2(new_n439), .A3(G200), .ZN(new_n713));
  INV_X1    g0513(.A(new_n713), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n714), .A2(G107), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n697), .A2(G190), .A3(G200), .ZN(new_n716));
  INV_X1    g0516(.A(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n717), .A2(G87), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n712), .A2(new_n715), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n707), .A2(new_n439), .ZN(new_n720));
  AOI21_X1  g0520(.A(new_n265), .B1(new_n720), .B2(G50), .ZN(new_n721));
  XNOR2_X1  g0521(.A(new_n706), .B(KEYINPUT91), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(new_n698), .ZN(new_n723));
  INV_X1    g0523(.A(new_n308), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n722), .A2(new_n709), .ZN(new_n725));
  OAI221_X1 g0525(.A(new_n721), .B1(new_n723), .B2(new_n361), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  OR3_X1    g0526(.A1(new_n705), .A2(new_n719), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G283), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n265), .B1(new_n713), .B2(new_n728), .ZN(new_n729));
  AOI22_X1  g0529(.A1(new_n720), .A2(G326), .B1(new_n711), .B2(G294), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n468), .B2(new_n716), .ZN(new_n731));
  INV_X1    g0531(.A(new_n725), .ZN(new_n732));
  AOI211_X1 g0532(.A(new_n729), .B(new_n731), .C1(G322), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(new_n723), .ZN(new_n734));
  AOI22_X1  g0534(.A1(G311), .A2(new_n734), .B1(new_n703), .B2(G329), .ZN(new_n735));
  XNOR2_X1  g0535(.A(KEYINPUT33), .B(G317), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(KEYINPUT93), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n708), .B1(new_n736), .B2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n733), .B(new_n735), .C1(new_n738), .C2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n696), .B1(new_n727), .B2(new_n741), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n692), .A2(new_n695), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n248), .A2(new_n333), .ZN(new_n744));
  INV_X1    g0544(.A(new_n277), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n641), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n747), .B1(new_n333), .B2(new_n218), .ZN(new_n748));
  INV_X1    g0548(.A(KEYINPUT90), .ZN(new_n749));
  AOI21_X1  g0549(.A(new_n744), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n750), .B1(new_n749), .B2(new_n748), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n641), .A2(new_n265), .ZN(new_n752));
  AOI22_X1  g0552(.A1(G355), .A2(new_n752), .B1(new_n455), .B2(new_n641), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  AOI211_X1 g0554(.A(new_n687), .B(new_n742), .C1(new_n743), .C2(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n689), .B1(new_n694), .B2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(G396));
  INV_X1    g0557(.A(new_n687), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n431), .A2(new_n623), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT95), .ZN(new_n760));
  OAI21_X1  g0560(.A(KEYINPUT96), .B1(new_n446), .B2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(KEYINPUT95), .ZN(new_n762));
  XNOR2_X1  g0562(.A(new_n759), .B(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(KEYINPUT96), .ZN(new_n764));
  NAND4_X1  g0564(.A1(new_n763), .A2(new_n764), .A3(new_n445), .A4(new_n440), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n604), .A2(new_n636), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n606), .A2(new_n623), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n761), .A2(new_n768), .A3(new_n765), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n767), .B1(new_n659), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n758), .B1(new_n771), .B2(new_n676), .ZN(new_n772));
  OAI21_X1  g0572(.A(new_n772), .B1(new_n676), .B2(new_n771), .ZN(new_n773));
  AOI22_X1  g0573(.A1(new_n708), .A2(G150), .B1(new_n720), .B2(G137), .ZN(new_n774));
  INV_X1    g0574(.A(G143), .ZN(new_n775));
  OAI221_X1 g0575(.A(new_n774), .B1(new_n723), .B2(new_n258), .C1(new_n775), .C2(new_n725), .ZN(new_n776));
  INV_X1    g0576(.A(KEYINPUT34), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n776), .A2(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n776), .A2(new_n777), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n703), .A2(G132), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n714), .A2(G68), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n781), .B1(new_n217), .B2(new_n716), .ZN(new_n782));
  AOI211_X1 g0582(.A(new_n277), .B(new_n782), .C1(new_n308), .C2(new_n711), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n778), .A2(new_n779), .A3(new_n780), .A4(new_n783), .ZN(new_n784));
  AOI22_X1  g0584(.A1(new_n708), .A2(G283), .B1(new_n720), .B2(G303), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n785), .B1(new_n455), .B2(new_n723), .ZN(new_n786));
  XNOR2_X1  g0586(.A(new_n786), .B(KEYINPUT94), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n370), .B1(new_n711), .B2(G97), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n717), .A2(G107), .B1(new_n714), .B2(G87), .ZN(new_n789));
  AOI22_X1  g0589(.A1(G294), .A2(new_n732), .B1(new_n703), .B2(G311), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n787), .A2(new_n788), .A3(new_n789), .A4(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n696), .B1(new_n784), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n695), .A2(new_n690), .ZN(new_n793));
  AOI211_X1 g0593(.A(new_n687), .B(new_n792), .C1(new_n361), .C2(new_n793), .ZN(new_n794));
  OAI21_X1  g0594(.A(new_n794), .B1(new_n770), .B2(new_n691), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n773), .A2(new_n795), .ZN(G384));
  OR2_X1    g0596(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n490), .A2(KEYINPUT35), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n797), .A2(G116), .A3(new_n221), .A4(new_n798), .ZN(new_n799));
  XOR2_X1   g0599(.A(new_n799), .B(KEYINPUT36), .Z(new_n800));
  NAND3_X1  g0600(.A1(new_n218), .A2(G77), .A3(new_n254), .ZN(new_n801));
  AOI211_X1 g0601(.A(G13), .B(new_n304), .C1(new_n801), .C2(new_n244), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT39), .ZN(new_n804));
  XOR2_X1   g0604(.A(new_n621), .B(KEYINPUT98), .Z(new_n805));
  NAND3_X1  g0605(.A1(new_n315), .A2(new_n321), .A3(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n299), .A2(new_n314), .ZN(new_n807));
  AOI21_X1  g0607(.A(KEYINPUT37), .B1(new_n807), .B2(new_n347), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n343), .A2(new_n806), .A3(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(KEYINPUT99), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g0611(.A1(new_n343), .A2(new_n806), .A3(new_n808), .A4(KEYINPUT99), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n806), .A2(new_n348), .A3(new_n609), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n814), .A2(KEYINPUT37), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n610), .A2(new_n352), .ZN(new_n817));
  OR2_X1    g0617(.A1(new_n817), .A2(new_n806), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT38), .B1(new_n816), .B2(new_n818), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n297), .A2(KEYINPUT16), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n820), .A2(new_n316), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n294), .A2(new_n298), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n314), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(KEYINPUT97), .ZN(new_n825));
  INV_X1    g0625(.A(new_n621), .ZN(new_n826));
  NAND3_X1  g0626(.A1(new_n824), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n824), .A2(new_n342), .ZN(new_n828));
  OAI21_X1  g0628(.A(KEYINPUT97), .B1(new_n823), .B2(new_n621), .ZN(new_n829));
  NAND4_X1  g0629(.A1(new_n827), .A2(new_n828), .A3(new_n348), .A4(new_n829), .ZN(new_n830));
  AOI22_X1  g0630(.A1(new_n811), .A2(new_n812), .B1(new_n830), .B2(KEYINPUT37), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n827), .A2(new_n829), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n352), .B1(KEYINPUT18), .B2(new_n343), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n832), .B1(new_n833), .B2(new_n344), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT38), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n831), .A2(new_n834), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n804), .B1(new_n819), .B2(new_n836), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n386), .A2(new_n387), .ZN(new_n838));
  NAND3_X1  g0638(.A1(new_n838), .A2(new_n368), .A3(new_n636), .ZN(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n830), .A2(KEYINPUT37), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n813), .A2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(new_n832), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n355), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n842), .A2(KEYINPUT38), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n835), .B1(new_n831), .B2(new_n834), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT39), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n837), .A2(new_n840), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  INV_X1    g0649(.A(new_n391), .ZN(new_n850));
  OAI211_X1 g0650(.A(new_n368), .B(new_n623), .C1(new_n838), .C2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n368), .A2(new_n623), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n388), .A2(new_n391), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n606), .A2(new_n636), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n855), .B1(new_n767), .B2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n805), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n849), .A2(new_n857), .B1(new_n610), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n848), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n604), .A2(new_n636), .ZN(new_n861));
  INV_X1    g0661(.A(KEYINPUT29), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g0663(.A1(new_n356), .A2(new_n447), .A3(new_n863), .A4(new_n657), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n613), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n860), .B(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n849), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n769), .B1(new_n853), .B2(new_n851), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  INV_X1    g0669(.A(new_n672), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n670), .A2(KEYINPUT31), .A3(new_n623), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n674), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n868), .A2(new_n869), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n868), .A2(new_n872), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n811), .A2(new_n812), .B1(KEYINPUT37), .B2(new_n814), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n817), .A2(new_n806), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n835), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n874), .B1(new_n845), .B2(new_n877), .ZN(new_n878));
  OAI22_X1  g0678(.A1(new_n867), .A2(new_n873), .B1(new_n878), .B2(new_n869), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n879), .A2(new_n449), .A3(new_n872), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n873), .B1(new_n845), .B2(new_n846), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n845), .A2(new_n877), .ZN(new_n882));
  INV_X1    g0682(.A(new_n874), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n881), .B1(new_n884), .B2(KEYINPUT40), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n449), .A2(new_n872), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n880), .A2(G330), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n866), .A2(new_n888), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n304), .B2(new_n617), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n866), .A2(new_n888), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n803), .B1(new_n890), .B2(new_n891), .ZN(G367));
  OAI221_X1 g0692(.A(new_n743), .B1(new_n213), .B2(new_n427), .C1(new_n747), .C2(new_n239), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n758), .ZN(new_n894));
  INV_X1    g0694(.A(new_n708), .ZN(new_n895));
  INV_X1    g0695(.A(new_n720), .ZN(new_n896));
  OAI22_X1  g0696(.A1(new_n895), .A2(new_n258), .B1(new_n896), .B2(new_n775), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n732), .A2(G150), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n703), .A2(G137), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n711), .ZN(new_n901));
  OAI22_X1  g0701(.A1(new_n901), .A2(new_n202), .B1(new_n713), .B2(new_n361), .ZN(new_n902));
  OAI221_X1 g0702(.A(new_n370), .B1(new_n724), .B2(new_n716), .C1(new_n723), .C2(new_n217), .ZN(new_n903));
  OR4_X1    g0703(.A1(new_n897), .A2(new_n900), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n713), .A2(new_n451), .ZN(new_n905));
  INV_X1    g0705(.A(G294), .ZN(new_n906));
  OAI21_X1  g0706(.A(new_n277), .B1(new_n895), .B2(new_n906), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n905), .B(new_n907), .C1(G107), .C2(new_n711), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT46), .ZN(new_n909));
  NOR3_X1   g0709(.A1(new_n716), .A2(new_n909), .A3(new_n455), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n910), .B1(new_n734), .B2(G283), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n909), .B1(new_n716), .B2(new_n455), .ZN(new_n912));
  XOR2_X1   g0712(.A(KEYINPUT105), .B(G317), .Z(new_n913));
  OR2_X1    g0713(.A1(new_n702), .A2(new_n913), .ZN(new_n914));
  NAND4_X1  g0714(.A1(new_n908), .A2(new_n911), .A3(new_n912), .A4(new_n914), .ZN(new_n915));
  AOI22_X1  g0715(.A1(new_n732), .A2(G303), .B1(G311), .B2(new_n720), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n916), .B(KEYINPUT104), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n904), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT47), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n894), .B1(new_n919), .B2(new_n695), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n591), .B1(new_n547), .B2(new_n636), .ZN(new_n921));
  OR3_X1    g0721(.A1(new_n594), .A2(new_n547), .A3(new_n636), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n921), .A2(new_n692), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  XNOR2_X1  g0724(.A(new_n686), .B(KEYINPUT103), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT44), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n518), .A2(new_n519), .A3(new_n623), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n516), .A2(new_n520), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n499), .A2(new_n623), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n928), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n927), .B1(new_n639), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n521), .A2(new_n930), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n638), .A2(KEYINPUT44), .A3(new_n934), .A4(new_n928), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n637), .A2(new_n932), .A3(new_n628), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT45), .Z(new_n938));
  AOI211_X1 g0738(.A(KEYINPUT101), .B(new_n634), .C1(new_n936), .C2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n634), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n936), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT101), .ZN(new_n942));
  AOI21_X1  g0742(.A(new_n940), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n635), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n632), .B1(new_n945), .B2(new_n623), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n946), .A2(new_n637), .ZN(new_n947));
  XNOR2_X1  g0747(.A(new_n685), .B(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n679), .B2(new_n680), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT102), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n944), .A2(new_n949), .A3(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n950), .B1(new_n944), .B2(new_n949), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n681), .B1(new_n952), .B2(new_n953), .ZN(new_n954));
  XOR2_X1   g0754(.A(new_n642), .B(KEYINPUT41), .Z(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n926), .B1(new_n954), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n940), .A2(new_n932), .ZN(new_n958));
  XNOR2_X1  g0758(.A(new_n958), .B(KEYINPUT100), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n921), .A2(new_n922), .ZN(new_n960));
  NOR2_X1   g0760(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n961));
  NOR2_X1   g0761(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g0762(.A(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n959), .A2(new_n961), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n631), .A2(new_n516), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n623), .B1(new_n965), .B2(new_n520), .ZN(new_n966));
  INV_X1    g0766(.A(new_n637), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n967), .A2(new_n932), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n966), .B1(new_n968), .B2(KEYINPUT42), .ZN(new_n969));
  OAI21_X1  g0769(.A(new_n969), .B1(KEYINPUT42), .B2(new_n968), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n960), .A2(KEYINPUT43), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g0772(.A1(new_n963), .A2(new_n964), .A3(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(new_n972), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n959), .A2(new_n961), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n974), .B1(new_n975), .B2(new_n962), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n973), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n924), .B1(new_n957), .B2(new_n977), .ZN(G387));
  AND2_X1   g0778(.A1(new_n679), .A2(new_n680), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n948), .ZN(new_n980));
  INV_X1    g0780(.A(new_n949), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n642), .A3(new_n981), .ZN(new_n982));
  OAI22_X1  g0782(.A1(new_n217), .A2(new_n725), .B1(new_n702), .B2(new_n402), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n983), .B1(G68), .B2(new_n734), .ZN(new_n984));
  NOR2_X1   g0784(.A1(new_n716), .A2(new_n361), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n901), .A2(new_n427), .ZN(new_n986));
  AOI211_X1 g0786(.A(new_n985), .B(new_n986), .C1(G159), .C2(new_n720), .ZN(new_n987));
  AOI211_X1 g0787(.A(new_n905), .B(new_n277), .C1(new_n309), .C2(new_n708), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n984), .A2(new_n987), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n703), .A2(G326), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n745), .B1(G116), .B2(new_n714), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n901), .A2(new_n728), .B1(new_n716), .B2(new_n906), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n708), .A2(G311), .B1(new_n720), .B2(G322), .ZN(new_n993));
  OAI221_X1 g0793(.A(new_n993), .B1(new_n723), .B2(new_n468), .C1(new_n725), .C2(new_n913), .ZN(new_n994));
  INV_X1    g0794(.A(KEYINPUT48), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n995), .B2(new_n994), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT49), .ZN(new_n998));
  OAI211_X1 g0798(.A(new_n990), .B(new_n991), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n997), .A2(new_n998), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n989), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1001), .A2(new_n695), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n236), .A2(G45), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT106), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n644), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1005), .A2(KEYINPUT107), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1005), .A2(KEYINPUT107), .ZN(new_n1007));
  AOI21_X1  g0807(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1009), .A2(KEYINPUT108), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n425), .A2(G50), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT50), .ZN(new_n1013));
  NAND3_X1  g0813(.A1(new_n1010), .A2(new_n1011), .A3(new_n1013), .ZN(new_n1014));
  NAND3_X1  g0814(.A1(new_n1004), .A2(new_n746), .A3(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(new_n1005), .A2(new_n752), .B1(new_n433), .B2(new_n641), .ZN(new_n1016));
  NAND2_X1  g0816(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n687), .B1(new_n1017), .B2(new_n743), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1002), .A2(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1019), .B1(new_n632), .B2(new_n692), .ZN(new_n1020));
  INV_X1    g0820(.A(new_n948), .ZN(new_n1021));
  AOI21_X1  g0821(.A(new_n1020), .B1(new_n1021), .B2(new_n926), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n982), .A2(new_n1022), .ZN(G393));
  XNOR2_X1  g0823(.A(new_n941), .B(new_n634), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n1024), .A2(new_n926), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n743), .B1(new_n451), .B2(new_n213), .C1(new_n747), .C2(new_n243), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(new_n758), .ZN(new_n1027));
  XOR2_X1   g0827(.A(new_n1027), .B(KEYINPUT109), .Z(new_n1028));
  INV_X1    g0828(.A(G87), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n745), .B1(new_n1029), .B2(new_n713), .ZN(new_n1030));
  NOR2_X1   g0830(.A1(new_n723), .A2(new_n425), .ZN(new_n1031));
  AOI211_X1 g0831(.A(new_n1030), .B(new_n1031), .C1(G143), .C2(new_n703), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n711), .A2(G77), .ZN(new_n1033));
  AOI22_X1  g0833(.A1(new_n708), .A2(G50), .B1(new_n717), .B2(G68), .ZN(new_n1034));
  NAND3_X1  g0834(.A1(new_n1032), .A2(new_n1033), .A3(new_n1034), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n725), .A2(new_n258), .B1(new_n402), .B2(new_n896), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT51), .Z(new_n1037));
  NOR2_X1   g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  AND2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT110), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(KEYINPUT110), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n732), .A2(G311), .B1(G317), .B2(new_n720), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT52), .Z(new_n1043));
  OAI211_X1 g0843(.A(new_n265), .B(new_n715), .C1(new_n723), .C2(new_n906), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(G322), .B2(new_n703), .ZN(new_n1045));
  OAI22_X1  g0845(.A1(new_n895), .A2(new_n468), .B1(new_n716), .B2(new_n728), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1046), .B1(G116), .B2(new_n711), .ZN(new_n1047));
  AND3_X1   g0847(.A1(new_n1043), .A2(new_n1045), .A3(new_n1047), .ZN(new_n1048));
  NOR3_X1   g0848(.A1(new_n1040), .A2(new_n1041), .A3(new_n1048), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n1028), .B1(new_n932), .B2(new_n693), .C1(new_n1049), .C2(new_n696), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1025), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n944), .A2(new_n949), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT102), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1053), .A2(new_n951), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n1024), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n643), .B1(new_n981), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1051), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n1057), .ZN(G390));
  AND3_X1   g0858(.A1(new_n868), .A2(G330), .A3(new_n872), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n767), .A2(new_n856), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n840), .B1(new_n1060), .B2(new_n854), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n1061), .B1(new_n837), .B2(new_n847), .ZN(new_n1062));
  OAI211_X1 g0862(.A(new_n636), .B(new_n766), .C1(new_n652), .C2(new_n656), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1063), .A2(new_n856), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n840), .B1(new_n1064), .B2(new_n854), .ZN(new_n1065));
  NAND2_X1  g0865(.A1(new_n1065), .A2(new_n882), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1059), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n845), .A2(new_n846), .A3(KEYINPUT39), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n845), .B2(new_n877), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1069), .A2(new_n1070), .B1(new_n840), .B2(new_n857), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n675), .A2(new_n868), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1072), .A3(new_n1066), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n356), .A2(new_n447), .A3(new_n675), .ZN(new_n1074));
  NAND3_X1  g0874(.A1(new_n864), .A2(new_n613), .A3(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n854), .B1(new_n675), .B2(new_n770), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1060), .B1(new_n1076), .B2(new_n1059), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n872), .A2(G330), .A3(new_n770), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1078), .A2(new_n855), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n1079), .A2(new_n856), .A3(new_n1072), .A4(new_n1063), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1077), .A2(new_n1080), .ZN(new_n1081));
  INV_X1    g0881(.A(new_n1081), .ZN(new_n1082));
  NOR2_X1   g0882(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1068), .A2(new_n1073), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1084), .A2(KEYINPUT111), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT111), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1068), .A2(new_n1073), .A3(new_n1083), .A4(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1085), .A2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1083), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n643), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1088), .A2(new_n1091), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n1089), .A2(new_n925), .ZN(new_n1093));
  INV_X1    g0893(.A(new_n793), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n723), .A2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n717), .A2(G150), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1096), .B(new_n1098), .C1(G125), .C2(new_n703), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n901), .A2(new_n258), .B1(new_n713), .B2(new_n217), .ZN(new_n1100));
  INV_X1    g0900(.A(G128), .ZN(new_n1101));
  INV_X1    g0901(.A(G132), .ZN(new_n1102));
  OAI221_X1 g0902(.A(new_n370), .B1(new_n896), .B2(new_n1101), .C1(new_n725), .C2(new_n1102), .ZN(new_n1103));
  AOI211_X1 g0903(.A(new_n1100), .B(new_n1103), .C1(G137), .C2(new_n708), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n708), .A2(G107), .B1(new_n720), .B2(G283), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n451), .B2(new_n723), .ZN(new_n1106));
  XOR2_X1   g0906(.A(new_n1106), .B(KEYINPUT112), .Z(new_n1107));
  OAI22_X1  g0907(.A1(new_n455), .A2(new_n725), .B1(new_n702), .B2(new_n906), .ZN(new_n1108));
  NAND4_X1  g0908(.A1(new_n718), .A2(new_n781), .A3(new_n1033), .A4(new_n265), .ZN(new_n1109));
  NOR2_X1   g0909(.A1(new_n1108), .A2(new_n1109), .ZN(new_n1110));
  AOI22_X1  g0910(.A1(new_n1099), .A2(new_n1104), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  OAI221_X1 g0911(.A(new_n758), .B1(new_n309), .B2(new_n1094), .C1(new_n1111), .C2(new_n696), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n837), .A2(new_n847), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1112), .B1(new_n1113), .B2(new_n690), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n1114), .B(KEYINPUT113), .ZN(new_n1115));
  NOR2_X1   g0915(.A1(new_n1093), .A2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1092), .A2(new_n1116), .ZN(G378));
  INV_X1    g0917(.A(KEYINPUT57), .ZN(new_n1118));
  XNOR2_X1  g0918(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1119), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n409), .A2(new_n621), .ZN(new_n1121));
  INV_X1    g0921(.A(new_n1121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n415), .A2(new_n418), .A3(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1122), .B1(new_n415), .B2(new_n418), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1120), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n1125), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1127), .A2(new_n1123), .A3(new_n1119), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1126), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1130), .B1(new_n885), .B2(new_n661), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT116), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1129), .A2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1126), .A2(new_n1128), .A3(KEYINPUT116), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n869), .B1(new_n882), .B2(new_n883), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1135), .B(G330), .C1(new_n1136), .C2(new_n881), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1131), .A2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n860), .A2(KEYINPUT117), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT117), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n848), .A2(new_n1140), .A3(new_n859), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1138), .A2(KEYINPUT118), .A3(new_n1139), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g0942(.A(new_n1137), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n1129), .B1(new_n879), .B2(G330), .ZN(new_n1144));
  NOR2_X1   g0944(.A1(new_n1143), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1146));
  NOR2_X1   g0946(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n860), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1131), .A2(new_n1148), .A3(new_n1137), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT118), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1142), .B1(new_n1147), .B2(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1075), .B1(new_n1085), .B2(new_n1087), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1118), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n1075), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1088), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT119), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1148), .B1(new_n1131), .B2(new_n1137), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n1118), .B1(new_n1159), .B2(new_n1149), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1156), .A2(new_n1157), .A3(new_n1160), .ZN(new_n1161));
  NOR3_X1   g0961(.A1(new_n1143), .A2(new_n1144), .A3(new_n860), .ZN(new_n1162));
  OAI21_X1  g0962(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1158), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT119), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1154), .A2(new_n1161), .A3(new_n642), .A4(new_n1164), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n926), .B(new_n1142), .C1(new_n1147), .C2(new_n1151), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n687), .B1(new_n217), .B2(new_n793), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(G128), .A2(new_n732), .B1(new_n734), .B2(G137), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n720), .A2(G125), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n708), .A2(G132), .B1(new_n711), .B2(G150), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  NOR2_X1   g0971(.A1(new_n716), .A2(new_n1095), .ZN(new_n1172));
  XOR2_X1   g0972(.A(new_n1172), .B(KEYINPUT115), .Z(new_n1173));
  NOR2_X1   g0973(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1175), .A2(KEYINPUT59), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n703), .A2(G124), .ZN(new_n1178));
  AOI211_X1 g0978(.A(G33), .B(G41), .C1(new_n714), .C2(G159), .ZN(new_n1179));
  NAND4_X1  g0979(.A1(new_n1176), .A2(new_n1177), .A3(new_n1178), .A4(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n277), .A2(new_n329), .ZN(new_n1181));
  NOR2_X1   g0981(.A1(new_n702), .A2(new_n728), .ZN(new_n1182));
  AOI211_X1 g0982(.A(new_n1181), .B(new_n1182), .C1(G107), .C2(new_n732), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n985), .B1(G68), .B2(new_n711), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(new_n720), .A2(G116), .B1(new_n714), .B2(new_n308), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1183), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n723), .A2(new_n427), .B1(new_n451), .B2(new_n895), .ZN(new_n1187));
  XOR2_X1   g0987(.A(new_n1187), .B(KEYINPUT114), .Z(new_n1188));
  NOR2_X1   g0988(.A1(new_n1186), .A2(new_n1188), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1189), .A2(KEYINPUT58), .ZN(new_n1191));
  OAI211_X1 g0991(.A(new_n1181), .B(new_n217), .C1(G33), .C2(G41), .ZN(new_n1192));
  AND4_X1   g0992(.A1(new_n1180), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1167), .B1(new_n696), .B2(new_n1193), .C1(new_n1135), .C2(new_n691), .ZN(new_n1194));
  AND2_X1   g0994(.A1(new_n1166), .A2(new_n1194), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1165), .A2(new_n1195), .ZN(G375));
  NAND2_X1  g0996(.A1(new_n1075), .A2(new_n1082), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1197), .ZN(new_n1198));
  XOR2_X1   g0998(.A(new_n955), .B(KEYINPUT120), .Z(new_n1199));
  NOR3_X1   g0999(.A1(new_n1198), .A2(new_n1083), .A3(new_n1199), .ZN(new_n1200));
  XNOR2_X1  g1000(.A(new_n1200), .B(KEYINPUT121), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1081), .A2(new_n926), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n855), .A2(new_n690), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1203), .B(KEYINPUT122), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n687), .B1(new_n202), .B2(new_n793), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(G107), .A2(new_n734), .B1(new_n732), .B2(G283), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n370), .B1(new_n714), .B2(G77), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1206), .B(new_n1207), .C1(new_n468), .C2(new_n702), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n896), .A2(new_n906), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n895), .A2(new_n455), .B1(new_n716), .B2(new_n451), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(new_n986), .A3(new_n1209), .A4(new_n1210), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n901), .A2(new_n217), .B1(new_n716), .B2(new_n258), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n277), .B(new_n1212), .C1(new_n308), .C2(new_n714), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n1101), .B2(new_n702), .C1(new_n402), .C2(new_n723), .ZN(new_n1214));
  XOR2_X1   g1014(.A(new_n1214), .B(KEYINPUT123), .Z(new_n1215));
  OAI22_X1  g1015(.A1(new_n1102), .A2(new_n896), .B1(new_n895), .B2(new_n1095), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1216), .B1(new_n732), .B2(G137), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1211), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1218));
  OAI211_X1 g1018(.A(new_n1204), .B(new_n1205), .C1(new_n696), .C2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1202), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1201), .A2(new_n1221), .ZN(G381));
  NAND3_X1  g1022(.A1(new_n982), .A2(new_n756), .A3(new_n1022), .ZN(new_n1223));
  OR4_X1    g1023(.A1(G384), .A2(G381), .A3(G390), .A4(new_n1223), .ZN(new_n1224));
  OR4_X1    g1024(.A1(G387), .A2(new_n1224), .A3(G375), .A4(G378), .ZN(G407));
  INV_X1    g1025(.A(G378), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n622), .A2(G213), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  OAI211_X1 g1029(.A(G407), .B(G213), .C1(G375), .C2(new_n1229), .ZN(G409));
  NAND2_X1  g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1231), .A2(new_n1223), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(KEYINPUT126), .ZN(new_n1233));
  INV_X1    g1033(.A(KEYINPUT126), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1231), .A2(new_n1234), .A3(new_n1223), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1233), .A2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n979), .B1(new_n1053), .B2(new_n951), .ZN(new_n1237));
  OAI21_X1  g1037(.A(new_n925), .B1(new_n1237), .B2(new_n955), .ZN(new_n1238));
  AND2_X1   g1038(.A1(new_n973), .A2(new_n976), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI21_X1  g1040(.A(G390), .B1(new_n1240), .B2(new_n924), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n924), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n1242), .B(new_n1057), .C1(new_n1238), .C2(new_n1239), .ZN(new_n1243));
  OAI21_X1  g1043(.A(new_n1236), .B1(new_n1241), .B2(new_n1243), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(G387), .A2(new_n1057), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n924), .A3(G390), .ZN(new_n1246));
  NAND4_X1  g1046(.A1(new_n1245), .A2(new_n1246), .A3(new_n1235), .A4(new_n1233), .ZN(new_n1247));
  INV_X1    g1047(.A(KEYINPUT61), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1244), .A2(new_n1247), .A3(new_n1248), .ZN(new_n1249));
  INV_X1    g1049(.A(KEYINPUT127), .ZN(new_n1250));
  XNOR2_X1  g1050(.A(new_n1249), .B(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT63), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1165), .A2(G378), .A3(new_n1195), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1152), .A2(new_n1153), .A3(new_n1199), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n926), .B1(new_n1162), .B2(new_n1158), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1194), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1226), .B1(new_n1254), .B2(new_n1256), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1258), .A2(new_n1227), .ZN(new_n1259));
  NOR2_X1   g1059(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1260));
  AND2_X1   g1060(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT60), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n1262), .B1(new_n1090), .B2(new_n1197), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n643), .B1(new_n1197), .B2(new_n1262), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1221), .B1(new_n1260), .B2(new_n1261), .C1(new_n1263), .C2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1267), .A2(new_n1220), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1268), .B2(new_n1261), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n1252), .B1(new_n1259), .B2(new_n1269), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1269), .A2(G2897), .A3(new_n1228), .ZN(new_n1271));
  INV_X1    g1071(.A(G2897), .ZN(new_n1272));
  OAI221_X1 g1072(.A(new_n1266), .B1(new_n1272), .B2(new_n1227), .C1(new_n1268), .C2(new_n1261), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n1271), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT125), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1274), .B(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1276), .A2(new_n1259), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1228), .B1(new_n1253), .B2(new_n1257), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1269), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1251), .A2(new_n1270), .A3(new_n1277), .A4(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  AND3_X1   g1082(.A1(new_n1278), .A2(new_n1282), .A3(new_n1279), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1248), .B1(new_n1278), .B2(new_n1274), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1282), .B1(new_n1278), .B2(new_n1279), .ZN(new_n1285));
  NOR3_X1   g1085(.A1(new_n1283), .A2(new_n1284), .A3(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1244), .A2(new_n1247), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1287), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1281), .B1(new_n1286), .B2(new_n1288), .ZN(G405));
  INV_X1    g1089(.A(new_n1253), .ZN(new_n1290));
  AOI21_X1  g1090(.A(G378), .B1(new_n1165), .B2(new_n1195), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1279), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1291), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1293), .A2(new_n1253), .A3(new_n1269), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1292), .A2(new_n1294), .ZN(new_n1295));
  XNOR2_X1  g1095(.A(new_n1295), .B(new_n1287), .ZN(G402));
endmodule


