//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 1 1 0 0 1 0 0 0 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1 1 0 1 1 0 0 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:15 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n710, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n750, new_n751, new_n752,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n762,
    new_n763, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n784, new_n785,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n798, new_n799, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n994, new_n995, new_n996,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1023,
    new_n1024, new_n1025, new_n1026, new_n1027, new_n1028, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1054,
    new_n1055, new_n1056, new_n1057, new_n1058, new_n1059, new_n1060,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069, new_n1070, new_n1071, new_n1072;
  INV_X1    g000(.A(G221), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT9), .B(G234), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G902), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(G469), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT83), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  OAI21_X1  g009(.A(KEYINPUT67), .B1(new_n195), .B2(G143), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT67), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n197), .A2(new_n198), .A3(G146), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(KEYINPUT66), .A3(G143), .ZN(new_n200));
  AOI21_X1  g014(.A(KEYINPUT66), .B1(new_n195), .B2(G143), .ZN(new_n201));
  OAI211_X1 g015(.A(new_n196), .B(new_n199), .C1(new_n200), .C2(new_n201), .ZN(new_n202));
  INV_X1    g016(.A(G128), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n195), .A2(G143), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n203), .B1(new_n204), .B2(KEYINPUT1), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n202), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(KEYINPUT1), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n198), .A2(G146), .ZN(new_n209));
  AND4_X1   g023(.A1(new_n208), .A2(new_n204), .A3(new_n209), .A4(G128), .ZN(new_n210));
  INV_X1    g024(.A(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G104), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT3), .B1(new_n212), .B2(G107), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT3), .ZN(new_n214));
  INV_X1    g028(.A(G107), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G104), .ZN(new_n216));
  INV_X1    g030(.A(G101), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n212), .A2(G107), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n213), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NOR2_X1   g033(.A1(new_n212), .A2(G107), .ZN(new_n220));
  NOR2_X1   g034(.A1(new_n215), .A2(G104), .ZN(new_n221));
  OAI21_X1  g035(.A(G101), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n219), .A2(new_n222), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n207), .A2(new_n211), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g038(.A(KEYINPUT1), .B1(new_n198), .B2(G146), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT84), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT84), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n204), .A2(new_n227), .A3(KEYINPUT1), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n226), .A2(G128), .A3(new_n228), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n204), .A2(new_n209), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n210), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n224), .B1(new_n223), .B2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT11), .ZN(new_n233));
  INV_X1    g047(.A(G134), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n233), .B1(new_n234), .B2(G137), .ZN(new_n235));
  INV_X1    g049(.A(G137), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT11), .A3(G134), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(G137), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT68), .B(G131), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n235), .A2(new_n237), .A3(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT69), .ZN(new_n244));
  AND2_X1   g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND4_X1  g059(.A1(new_n235), .A2(new_n237), .A3(KEYINPUT69), .A4(new_n238), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G131), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n242), .B1(new_n245), .B2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n232), .A2(KEYINPUT12), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(KEYINPUT73), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT73), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n251), .B(new_n242), .C1(new_n245), .C2(new_n247), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n232), .A2(new_n250), .A3(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT12), .ZN(new_n254));
  AND3_X1   g068(.A1(new_n253), .A2(KEYINPUT86), .A3(new_n254), .ZN(new_n255));
  AOI21_X1  g069(.A(KEYINPUT86), .B1(new_n253), .B2(new_n254), .ZN(new_n256));
  OAI21_X1  g070(.A(new_n249), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT10), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n258), .B1(new_n231), .B2(new_n223), .ZN(new_n259));
  INV_X1    g073(.A(new_n223), .ZN(new_n260));
  AND2_X1   g074(.A1(new_n196), .A2(new_n199), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT66), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n204), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n195), .A2(KEYINPUT66), .A3(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n205), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n260), .B(KEYINPUT10), .C1(new_n266), .C2(new_n210), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT0), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n268), .A2(new_n203), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(KEYINPUT0), .B2(G128), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT65), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n271), .A2(new_n268), .A3(new_n203), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n230), .ZN(new_n274));
  AOI22_X1  g088(.A1(new_n202), .A2(new_n273), .B1(new_n269), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n213), .A2(new_n216), .A3(new_n218), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G101), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n277), .A2(KEYINPUT4), .A3(new_n219), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT4), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n276), .A2(new_n279), .A3(G101), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n275), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n259), .A2(new_n267), .A3(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n252), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n243), .A2(new_n244), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(G131), .A3(new_n246), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n251), .B1(new_n285), .B2(new_n242), .ZN(new_n286));
  OAI21_X1  g100(.A(KEYINPUT85), .B1(new_n283), .B2(new_n286), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT85), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n250), .A2(new_n288), .A3(new_n252), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n282), .B1(new_n287), .B2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n194), .B1(new_n257), .B2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  XNOR2_X1  g107(.A(G110), .B(G140), .ZN(new_n294));
  INV_X1    g108(.A(G953), .ZN(new_n295));
  AND2_X1   g109(.A1(new_n295), .A2(G227), .ZN(new_n296));
  XNOR2_X1  g110(.A(new_n294), .B(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(new_n249), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n253), .A2(new_n254), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT86), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n253), .A2(KEYINPUT86), .A3(new_n254), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n298), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n194), .B1(new_n303), .B2(new_n290), .ZN(new_n304));
  INV_X1    g118(.A(new_n297), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n283), .A2(new_n286), .ZN(new_n306));
  AND2_X1   g120(.A1(new_n306), .A2(new_n282), .ZN(new_n307));
  OAI21_X1  g121(.A(new_n305), .B1(new_n290), .B2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  AOI22_X1  g123(.A1(new_n293), .A2(new_n297), .B1(new_n304), .B2(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n193), .B1(new_n310), .B2(new_n190), .ZN(new_n311));
  OAI21_X1  g125(.A(new_n297), .B1(new_n290), .B2(new_n307), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT88), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  OAI211_X1 g128(.A(KEYINPUT88), .B(new_n297), .C1(new_n290), .C2(new_n307), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n290), .A2(new_n297), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  AOI21_X1  g132(.A(new_n318), .B1(new_n257), .B2(KEYINPUT87), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT87), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n249), .C1(new_n255), .C2(new_n256), .ZN(new_n321));
  AOI21_X1  g135(.A(new_n316), .B1(new_n319), .B2(new_n321), .ZN(new_n322));
  NOR3_X1   g136(.A1(new_n322), .A2(G469), .A3(G902), .ZN(new_n323));
  OAI21_X1  g137(.A(new_n192), .B1(new_n311), .B2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(G214), .B1(G237), .B2(G902), .ZN(new_n325));
  INV_X1    g139(.A(G113), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(KEYINPUT2), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT2), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G113), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n331));
  INV_X1    g145(.A(G116), .ZN(new_n332));
  OAI21_X1  g146(.A(new_n331), .B1(new_n332), .B2(G119), .ZN(new_n333));
  INV_X1    g147(.A(G119), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n334), .A2(KEYINPUT72), .A3(G116), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(G119), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n330), .A2(new_n333), .A3(new_n335), .A4(new_n336), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n337), .A2(new_n219), .A3(new_n222), .ZN(new_n338));
  XOR2_X1   g152(.A(KEYINPUT90), .B(KEYINPUT5), .Z(new_n339));
  NOR2_X1   g153(.A1(new_n332), .A2(G119), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n326), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n333), .A2(new_n335), .A3(new_n336), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(new_n339), .ZN(new_n343));
  AND2_X1   g157(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n342), .A2(new_n327), .A3(new_n329), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(new_n337), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n278), .A2(new_n346), .A3(new_n280), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n347), .A2(KEYINPUT89), .ZN(new_n348));
  INV_X1    g162(.A(KEYINPUT89), .ZN(new_n349));
  NAND4_X1  g163(.A1(new_n278), .A2(new_n346), .A3(new_n349), .A4(new_n280), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n344), .B1(new_n348), .B2(new_n350), .ZN(new_n351));
  XNOR2_X1  g165(.A(G110), .B(G122), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n210), .B1(new_n202), .B2(new_n206), .ZN(new_n354));
  INV_X1    g168(.A(G125), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  OAI21_X1  g170(.A(new_n356), .B1(new_n355), .B2(new_n275), .ZN(new_n357));
  INV_X1    g171(.A(G224), .ZN(new_n358));
  NOR2_X1   g172(.A1(new_n358), .A2(G953), .ZN(new_n359));
  XOR2_X1   g173(.A(new_n357), .B(new_n359), .Z(new_n360));
  INV_X1    g174(.A(KEYINPUT91), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n351), .B2(new_n352), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT6), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n363), .B1(new_n351), .B2(new_n352), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n338), .A2(new_n343), .ZN(new_n365));
  AND2_X1   g179(.A1(new_n276), .A2(G101), .ZN(new_n366));
  AOI22_X1  g180(.A1(new_n366), .A2(new_n279), .B1(new_n345), .B2(new_n337), .ZN(new_n367));
  AOI21_X1  g181(.A(new_n349), .B1(new_n367), .B2(new_n278), .ZN(new_n368));
  AND4_X1   g182(.A1(new_n349), .A2(new_n278), .A3(new_n346), .A4(new_n280), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n365), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(new_n352), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(KEYINPUT91), .A3(new_n371), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n362), .A2(new_n364), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(KEYINPUT92), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g189(.A1(new_n362), .A2(new_n364), .A3(new_n372), .A4(KEYINPUT92), .ZN(new_n376));
  AOI211_X1 g190(.A(new_n353), .B(new_n360), .C1(new_n375), .C2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(KEYINPUT7), .ZN(new_n378));
  OR3_X1    g192(.A1(new_n357), .A2(new_n378), .A3(new_n359), .ZN(new_n379));
  XNOR2_X1  g193(.A(new_n352), .B(KEYINPUT8), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT5), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n341), .B1(new_n381), .B2(new_n342), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n338), .A2(new_n382), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n260), .B1(new_n343), .B2(new_n337), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n380), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n357), .B1(new_n378), .B2(new_n359), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n379), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n370), .A2(new_n371), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(G902), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  OAI21_X1  g205(.A(G210), .B1(G237), .B2(G902), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n377), .A2(new_n391), .A3(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n375), .A2(new_n376), .ZN(new_n395));
  INV_X1    g209(.A(new_n353), .ZN(new_n396));
  INV_X1    g210(.A(new_n360), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(new_n392), .B1(new_n398), .B2(new_n390), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n325), .B1(new_n394), .B2(new_n399), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n324), .A2(new_n400), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n207), .A2(new_n211), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT74), .ZN(new_n403));
  INV_X1    g217(.A(G131), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n236), .A2(G134), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(new_n238), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n406), .B1(new_n239), .B2(new_n241), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n402), .A2(new_n403), .A3(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(new_n406), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n243), .B2(new_n240), .ZN(new_n410));
  OAI21_X1  g224(.A(KEYINPUT74), .B1(new_n354), .B2(new_n410), .ZN(new_n411));
  AND2_X1   g225(.A1(new_n408), .A2(new_n411), .ZN(new_n412));
  INV_X1    g226(.A(new_n346), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n250), .A2(new_n275), .A3(new_n252), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT70), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n417), .B1(new_n354), .B2(new_n410), .ZN(new_n418));
  OAI211_X1 g232(.A(new_n407), .B(KEYINPUT70), .C1(new_n266), .C2(new_n210), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n418), .A2(new_n419), .B1(new_n275), .B2(new_n248), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n420), .A2(new_n413), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT28), .B1(new_n416), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n346), .B1(new_n402), .B2(new_n407), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n414), .A2(new_n423), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT28), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  NOR2_X1   g241(.A1(G237), .A2(G953), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n428), .A2(G210), .ZN(new_n429));
  XOR2_X1   g243(.A(new_n429), .B(KEYINPUT27), .Z(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT26), .B(G101), .ZN(new_n431));
  XNOR2_X1  g245(.A(new_n430), .B(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n427), .A2(new_n432), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n412), .A2(KEYINPUT30), .A3(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n418), .A2(new_n419), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n248), .A2(new_n275), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  XNOR2_X1  g251(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(KEYINPUT71), .B1(new_n437), .B2(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT71), .ZN(new_n441));
  NOR3_X1   g255(.A1(new_n420), .A2(new_n441), .A3(new_n438), .ZN(new_n442));
  OAI211_X1 g256(.A(new_n346), .B(new_n434), .C1(new_n440), .C2(new_n442), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n416), .A2(new_n432), .ZN(new_n444));
  AND3_X1   g258(.A1(new_n443), .A2(KEYINPUT31), .A3(new_n444), .ZN(new_n445));
  AOI21_X1  g259(.A(KEYINPUT31), .B1(new_n443), .B2(new_n444), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n433), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(G472), .A2(G902), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n448), .B(KEYINPUT75), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(KEYINPUT32), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(KEYINPUT32), .ZN(new_n454));
  INV_X1    g268(.A(new_n432), .ZN(new_n455));
  AOI21_X1  g269(.A(new_n455), .B1(new_n422), .B2(new_n426), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n443), .A2(new_n444), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT31), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n443), .A2(KEYINPUT31), .A3(new_n444), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n456), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n454), .B1(new_n461), .B2(new_n449), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n422), .A2(new_n426), .A3(new_n455), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT29), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n437), .A2(KEYINPUT71), .A3(new_n439), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n441), .B1(new_n420), .B2(new_n438), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n408), .A2(new_n411), .ZN(new_n467));
  AOI21_X1  g281(.A(new_n467), .B1(new_n306), .B2(new_n275), .ZN(new_n468));
  AOI22_X1  g282(.A1(new_n465), .A2(new_n466), .B1(new_n468), .B2(KEYINPUT30), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n416), .B1(new_n469), .B2(new_n346), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n463), .B(new_n464), .C1(new_n470), .C2(new_n455), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n412), .A2(new_n414), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n346), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n425), .B1(new_n473), .B2(new_n415), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT77), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n424), .A2(new_n475), .A3(new_n425), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n426), .A2(KEYINPUT77), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n474), .A2(KEYINPUT76), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n413), .B1(new_n412), .B2(new_n414), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n416), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT76), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n432), .A2(new_n464), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n478), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n471), .A2(new_n484), .A3(new_n190), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G472), .ZN(new_n486));
  NAND4_X1  g300(.A1(new_n447), .A2(KEYINPUT78), .A3(KEYINPUT32), .A4(new_n450), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n453), .A2(new_n462), .A3(new_n486), .A4(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(G234), .ZN(new_n489));
  OAI21_X1  g303(.A(G217), .B1(new_n489), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT23), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n491), .B1(new_n334), .B2(G128), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n334), .A2(G128), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n203), .A2(KEYINPUT23), .A3(G119), .ZN(new_n494));
  AND3_X1   g308(.A1(new_n492), .A2(new_n493), .A3(new_n494), .ZN(new_n495));
  XNOR2_X1  g309(.A(KEYINPUT80), .B(G110), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT79), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n498), .B1(new_n334), .B2(G128), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n203), .A2(KEYINPUT79), .A3(G119), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n499), .A2(new_n500), .A3(new_n493), .ZN(new_n501));
  XNOR2_X1  g315(.A(KEYINPUT24), .B(G110), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n497), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT81), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  NOR3_X1   g320(.A1(new_n355), .A2(KEYINPUT16), .A3(G140), .ZN(new_n507));
  XNOR2_X1  g321(.A(G125), .B(G140), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n507), .B1(KEYINPUT16), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(G146), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n195), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n506), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n509), .A2(G146), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n513), .A2(new_n510), .ZN(new_n514));
  INV_X1    g328(.A(G110), .ZN(new_n515));
  OAI221_X1 g329(.A(new_n514), .B1(new_n515), .B2(new_n495), .C1(new_n502), .C2(new_n501), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g331(.A(KEYINPUT22), .B(G137), .ZN(new_n518));
  NOR3_X1   g332(.A1(new_n187), .A2(new_n489), .A3(G953), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n518), .B(new_n519), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n512), .A2(new_n516), .A3(new_n520), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n190), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n490), .B1(new_n524), .B2(KEYINPUT25), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(KEYINPUT25), .B2(new_n524), .ZN(new_n526));
  AOI21_X1  g340(.A(G902), .B1(new_n489), .B2(G217), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n522), .A2(new_n523), .A3(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT82), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  OR2_X1    g344(.A1(new_n528), .A2(new_n529), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n526), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT102), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT101), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT99), .ZN(new_n536));
  OAI21_X1  g350(.A(new_n536), .B1(new_n198), .B2(G128), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n203), .A2(KEYINPUT99), .A3(G143), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n198), .A2(G128), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT13), .ZN(new_n540));
  AOI22_X1  g354(.A1(new_n537), .A2(new_n538), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OR2_X1    g355(.A1(new_n541), .A2(KEYINPUT100), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n539), .A2(new_n540), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n543), .B1(new_n541), .B2(KEYINPUT100), .ZN(new_n544));
  AOI21_X1  g358(.A(new_n234), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n537), .A2(new_n538), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n546), .A2(new_n234), .A3(new_n539), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT98), .ZN(new_n548));
  INV_X1    g362(.A(G122), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(new_n549), .B2(G116), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n332), .A2(KEYINPUT98), .A3(G122), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AND2_X1   g366(.A1(KEYINPUT97), .A2(G122), .ZN(new_n553));
  NOR2_X1   g367(.A1(KEYINPUT97), .A2(G122), .ZN(new_n554));
  OAI21_X1  g368(.A(G116), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n555), .A3(new_n215), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n215), .B1(new_n552), .B2(new_n555), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n547), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n547), .ZN(new_n560));
  AOI21_X1  g374(.A(new_n234), .B1(new_n546), .B2(new_n539), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n556), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OR2_X1    g376(.A1(KEYINPUT97), .A2(G122), .ZN(new_n563));
  NAND2_X1  g377(.A1(KEYINPUT97), .A2(G122), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n332), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(KEYINPUT14), .B2(new_n552), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT14), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n550), .A2(new_n567), .A3(new_n551), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n215), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  OAI22_X1  g383(.A1(new_n545), .A2(new_n559), .B1(new_n562), .B2(new_n569), .ZN(new_n570));
  INV_X1    g384(.A(G217), .ZN(new_n571));
  NOR3_X1   g385(.A1(new_n188), .A2(new_n571), .A3(G953), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n535), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n542), .A2(new_n544), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(G134), .ZN(new_n576));
  INV_X1    g390(.A(new_n559), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n552), .A2(KEYINPUT14), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n579), .A2(new_n555), .A3(new_n568), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(G107), .ZN(new_n581));
  OAI211_X1 g395(.A(new_n581), .B(new_n556), .C1(new_n560), .C2(new_n561), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n578), .A2(KEYINPUT101), .A3(new_n582), .A4(new_n572), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n570), .A2(new_n573), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n574), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n534), .B1(new_n585), .B2(new_n190), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(G478), .ZN(new_n588));
  NOR2_X1   g402(.A1(new_n588), .A2(KEYINPUT15), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n534), .A3(new_n190), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n587), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n585), .A2(new_n190), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n591), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(G475), .ZN(new_n597));
  INV_X1    g411(.A(G237), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n295), .A3(G214), .ZN(new_n599));
  NOR2_X1   g413(.A1(new_n599), .A2(new_n198), .ZN(new_n600));
  AOI21_X1  g414(.A(G143), .B1(new_n428), .B2(G214), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT18), .ZN(new_n603));
  OAI21_X1  g417(.A(new_n602), .B1(new_n603), .B2(new_n404), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n599), .A2(new_n198), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n428), .A2(G143), .A3(G214), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(KEYINPUT18), .A3(G131), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n508), .B(new_n195), .ZN(new_n609));
  NAND3_X1  g423(.A1(new_n604), .A2(new_n608), .A3(new_n609), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n241), .B1(new_n605), .B2(new_n606), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n611), .A2(KEYINPUT17), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(new_n513), .A3(new_n510), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n607), .A2(new_n240), .ZN(new_n614));
  NOR3_X1   g428(.A1(new_n614), .A2(new_n611), .A3(KEYINPUT17), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n610), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(G113), .B(G122), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n617), .B(new_n212), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n616), .B(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n597), .B1(new_n620), .B2(new_n190), .ZN(new_n621));
  OR2_X1    g435(.A1(new_n616), .A2(new_n619), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT93), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n623), .B1(new_n614), .B2(new_n611), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n602), .A2(new_n241), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n607), .A2(new_n240), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(KEYINPUT93), .A3(new_n626), .ZN(new_n627));
  XNOR2_X1  g441(.A(new_n508), .B(KEYINPUT19), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n628), .A2(new_n195), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n624), .A2(new_n627), .A3(new_n510), .A4(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n630), .A2(KEYINPUT94), .A3(new_n610), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(new_n619), .ZN(new_n632));
  AOI21_X1  g446(.A(KEYINPUT94), .B1(new_n630), .B2(new_n610), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n622), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(KEYINPUT20), .ZN(new_n635));
  NOR2_X1   g449(.A1(G475), .A2(G902), .ZN(new_n636));
  XOR2_X1   g450(.A(new_n636), .B(KEYINPUT95), .Z(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g453(.A(new_n635), .B1(new_n634), .B2(new_n638), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT96), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND4_X1  g456(.A1(new_n634), .A2(KEYINPUT96), .A3(new_n635), .A4(new_n638), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n621), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(G952), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n645), .A2(G953), .ZN(new_n646));
  OAI21_X1  g460(.A(new_n646), .B1(new_n489), .B2(new_n598), .ZN(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT21), .B(G898), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT103), .ZN(new_n649));
  AOI211_X1 g463(.A(new_n190), .B(new_n295), .C1(G234), .C2(G237), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND3_X1  g466(.A1(new_n596), .A2(new_n644), .A3(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n653), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n401), .A2(new_n488), .A3(new_n533), .A4(new_n654), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n655), .B(G101), .ZN(G3));
  NOR2_X1   g470(.A1(new_n324), .A2(new_n532), .ZN(new_n657));
  OAI211_X1 g471(.A(new_n325), .B(new_n652), .C1(new_n394), .C2(new_n399), .ZN(new_n658));
  INV_X1    g472(.A(new_n644), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n587), .A2(new_n588), .A3(new_n590), .ZN(new_n660));
  INV_X1    g474(.A(KEYINPUT105), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT33), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n585), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n578), .A2(new_n582), .A3(new_n572), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n584), .A3(KEYINPUT33), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n588), .A2(G902), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  OAI21_X1  g482(.A(new_n661), .B1(new_n666), .B2(new_n668), .ZN(new_n669));
  NAND4_X1  g483(.A1(new_n663), .A2(KEYINPUT105), .A3(new_n665), .A4(new_n667), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n660), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n659), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n658), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(G472), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n447), .B2(new_n190), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT104), .ZN(new_n676));
  OAI22_X1  g490(.A1(new_n675), .A2(new_n676), .B1(new_n449), .B2(new_n461), .ZN(new_n677));
  OAI21_X1  g491(.A(G472), .B1(new_n461), .B2(G902), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n678), .A2(KEYINPUT104), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n677), .A2(new_n679), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n657), .A2(new_n673), .A3(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(KEYINPUT34), .B(G104), .Z(new_n682));
  XNOR2_X1  g496(.A(new_n681), .B(new_n682), .ZN(G6));
  NOR2_X1   g497(.A1(new_n461), .A2(new_n449), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n678), .B2(KEYINPUT104), .ZN(new_n685));
  NOR2_X1   g499(.A1(new_n193), .A2(new_n190), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT83), .B1(new_n257), .B2(new_n291), .ZN(new_n687));
  OAI22_X1  g501(.A1(new_n305), .A2(new_n292), .B1(new_n687), .B2(new_n308), .ZN(new_n688));
  AOI21_X1  g502(.A(new_n686), .B1(new_n688), .B2(G469), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n257), .A2(KEYINPUT87), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n690), .A2(new_n321), .A3(new_n317), .ZN(new_n691));
  AND2_X1   g505(.A1(new_n314), .A2(new_n315), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n693), .A2(new_n193), .A3(new_n190), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n191), .B1(new_n689), .B2(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n675), .A2(new_n676), .ZN(new_n696));
  NAND4_X1  g510(.A1(new_n685), .A2(new_n533), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n621), .ZN(new_n699));
  INV_X1    g513(.A(new_n640), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT106), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n639), .ZN(new_n702));
  INV_X1    g516(.A(new_n634), .ZN(new_n703));
  OAI211_X1 g517(.A(KEYINPUT106), .B(KEYINPUT20), .C1(new_n703), .C2(new_n637), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n595), .A2(new_n699), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  NOR2_X1   g519(.A1(new_n658), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n698), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT35), .B(G107), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n707), .B(new_n708), .ZN(G9));
  NOR2_X1   g523(.A1(new_n521), .A2(KEYINPUT36), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n517), .B(new_n710), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n711), .A2(new_n527), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n526), .A2(new_n712), .ZN(new_n713));
  NAND3_X1  g527(.A1(new_n685), .A2(new_n696), .A3(new_n713), .ZN(new_n714));
  INV_X1    g528(.A(new_n325), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n393), .B1(new_n377), .B2(new_n391), .ZN(new_n716));
  NAND3_X1  g530(.A1(new_n398), .A2(new_n390), .A3(new_n392), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n715), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n654), .A2(new_n718), .A3(new_n695), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT37), .B(G110), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n720), .B(new_n721), .ZN(G12));
  NAND4_X1  g536(.A1(new_n488), .A2(new_n718), .A3(new_n695), .A4(new_n713), .ZN(new_n723));
  INV_X1    g537(.A(new_n647), .ZN(new_n724));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n724), .B1(new_n650), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n702), .A2(new_n699), .A3(new_n704), .A4(new_n727), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n728), .A2(new_n596), .ZN(new_n729));
  INV_X1    g543(.A(new_n729), .ZN(new_n730));
  NOR2_X1   g544(.A1(new_n723), .A2(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n203), .ZN(G30));
  XOR2_X1   g546(.A(new_n726), .B(KEYINPUT39), .Z(new_n733));
  NAND2_X1  g547(.A1(new_n695), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g548(.A(new_n734), .B(KEYINPUT40), .Z(new_n735));
  INV_X1    g549(.A(new_n713), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n416), .A2(new_n479), .ZN(new_n737));
  INV_X1    g551(.A(new_n737), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n738), .A2(new_n432), .B1(new_n443), .B2(new_n444), .ZN(new_n739));
  OAI21_X1  g553(.A(G472), .B1(new_n739), .B2(G902), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n453), .A2(new_n462), .A3(new_n487), .A4(new_n740), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n716), .A2(new_n717), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT38), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n596), .A2(new_n644), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n744), .A2(new_n715), .A3(new_n746), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n735), .A2(new_n736), .A3(new_n741), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G143), .ZN(G45));
  INV_X1    g563(.A(new_n671), .ZN(new_n750));
  NOR3_X1   g564(.A1(new_n750), .A2(new_n644), .A3(new_n726), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n401), .A2(new_n488), .A3(new_n713), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G146), .ZN(G48));
  OAI21_X1  g567(.A(G469), .B1(new_n322), .B2(G902), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n754), .A2(new_n192), .A3(new_n694), .ZN(new_n755));
  INV_X1    g569(.A(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n673), .A2(new_n488), .A3(new_n533), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(KEYINPUT41), .B(G113), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n757), .B(new_n758), .ZN(G15));
  NAND4_X1  g573(.A1(new_n706), .A2(new_n488), .A3(new_n533), .A4(new_n756), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G116), .ZN(G18));
  NOR2_X1   g575(.A1(new_n400), .A2(new_n755), .ZN(new_n762));
  NAND4_X1  g576(.A1(new_n762), .A2(new_n488), .A3(new_n654), .A4(new_n713), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(G119), .ZN(G21));
  NAND4_X1  g578(.A1(new_n754), .A2(new_n192), .A3(new_n694), .A4(new_n652), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n459), .A2(new_n460), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n477), .A2(new_n476), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n480), .B2(new_n481), .ZN(new_n769));
  NOR2_X1   g583(.A1(new_n474), .A2(KEYINPUT76), .ZN(new_n770));
  OAI21_X1  g584(.A(new_n432), .B1(new_n769), .B2(new_n770), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n449), .B1(new_n767), .B2(new_n771), .ZN(new_n772));
  NOR3_X1   g586(.A1(new_n675), .A2(new_n772), .A3(new_n532), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n766), .A2(new_n773), .A3(new_n718), .A4(new_n745), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT107), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n767), .A2(new_n771), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(new_n450), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n533), .A2(new_n778), .A3(new_n678), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n779), .A2(new_n765), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n780), .A2(KEYINPUT107), .A3(new_n718), .A4(new_n745), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n776), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g596(.A(new_n782), .B(G122), .ZN(G24));
  NOR3_X1   g597(.A1(new_n736), .A2(new_n675), .A3(new_n772), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n762), .A2(new_n751), .A3(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G125), .ZN(G27));
  NOR3_X1   g600(.A1(new_n394), .A2(new_n399), .A3(new_n715), .ZN(new_n787));
  NAND3_X1  g601(.A1(new_n787), .A2(new_n695), .A3(new_n751), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n486), .A2(new_n462), .A3(new_n451), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n533), .ZN(new_n790));
  OAI21_X1  g604(.A(KEYINPUT42), .B1(new_n788), .B2(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n716), .A2(new_n325), .A3(new_n717), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n324), .A2(new_n792), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n672), .A2(KEYINPUT42), .A3(new_n726), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n793), .A2(new_n488), .A3(new_n533), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n791), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(new_n404), .ZN(G33));
  AND4_X1   g611(.A1(new_n488), .A2(new_n533), .A3(new_n695), .A4(new_n787), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(new_n729), .ZN(new_n799));
  XNOR2_X1  g613(.A(new_n799), .B(G134), .ZN(G36));
  NAND2_X1  g614(.A1(new_n644), .A2(new_n671), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n801), .A2(KEYINPUT43), .ZN(new_n803));
  OR4_X1    g617(.A1(new_n680), .A2(new_n736), .A3(new_n802), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT44), .ZN(new_n805));
  OR2_X1    g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n792), .B1(new_n804), .B2(new_n805), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n193), .B1(new_n688), .B2(KEYINPUT45), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n808), .B1(KEYINPUT45), .B2(new_n688), .ZN(new_n809));
  INV_X1    g623(.A(new_n686), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT46), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n694), .ZN(new_n814));
  NOR2_X1   g628(.A1(new_n811), .A2(new_n812), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n192), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n806), .A2(new_n807), .A3(new_n733), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g632(.A(new_n818), .B(G137), .ZN(G39));
  INV_X1    g633(.A(KEYINPUT47), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  OAI211_X1 g635(.A(KEYINPUT47), .B(new_n192), .C1(new_n814), .C2(new_n815), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n751), .A2(new_n532), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n825), .A2(new_n488), .A3(new_n792), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(KEYINPUT108), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n824), .A2(new_n827), .ZN(new_n828));
  XOR2_X1   g642(.A(new_n828), .B(G140), .Z(G42));
  NAND2_X1  g643(.A1(new_n645), .A2(new_n295), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT121), .ZN(new_n831));
  NOR3_X1   g645(.A1(new_n802), .A2(new_n803), .A3(new_n647), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n762), .A3(new_n773), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n646), .ZN(new_n834));
  NOR2_X1   g648(.A1(new_n792), .A2(new_n755), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n790), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g652(.A(KEYINPUT120), .B(KEYINPUT48), .ZN(new_n839));
  XNOR2_X1  g653(.A(new_n838), .B(new_n839), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n750), .A2(new_n644), .ZN(new_n841));
  INV_X1    g655(.A(new_n741), .ZN(new_n842));
  AND4_X1   g656(.A1(new_n533), .A2(new_n842), .A3(new_n724), .A4(new_n835), .ZN(new_n843));
  AOI211_X1 g657(.A(new_n834), .B(new_n840), .C1(new_n841), .C2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n744), .A2(new_n715), .A3(new_n756), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n832), .A2(new_n773), .ZN(new_n846));
  OAI21_X1  g660(.A(KEYINPUT118), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n659), .A2(new_n671), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n843), .A2(new_n850), .B1(new_n836), .B2(new_n784), .ZN(new_n851));
  OAI211_X1 g665(.A(KEYINPUT118), .B(KEYINPUT50), .C1(new_n845), .C2(new_n846), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n849), .A2(new_n851), .A3(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT51), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT119), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n832), .A2(new_n773), .A3(new_n787), .ZN(new_n857));
  XOR2_X1   g671(.A(new_n857), .B(KEYINPUT116), .Z(new_n858));
  AND2_X1   g672(.A1(new_n754), .A2(new_n694), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n859), .A2(new_n191), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(new_n858), .B1(new_n823), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n855), .A2(new_n856), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n856), .B1(new_n855), .B2(new_n862), .ZN(new_n865));
  OAI21_X1  g679(.A(new_n844), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n858), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n824), .A2(KEYINPUT117), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT117), .ZN(new_n869));
  AOI21_X1  g683(.A(new_n861), .B1(new_n823), .B2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(new_n867), .B1(new_n868), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n854), .B1(new_n871), .B2(new_n853), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n831), .B1(new_n866), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(new_n865), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n863), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n876), .A2(new_n872), .A3(KEYINPUT121), .A4(new_n844), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  AND3_X1   g692(.A1(new_n757), .A2(new_n760), .A3(new_n763), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT111), .ZN(new_n880));
  AND3_X1   g694(.A1(new_n585), .A2(new_n534), .A3(new_n190), .ZN(new_n881));
  INV_X1    g695(.A(new_n589), .ZN(new_n882));
  NOR3_X1   g696(.A1(new_n881), .A2(new_n586), .A3(new_n882), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n880), .B1(new_n883), .B2(new_n593), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n591), .A2(KEYINPUT111), .A3(new_n594), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n728), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n488), .A2(new_n713), .A3(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n784), .A2(new_n751), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n793), .A2(new_n890), .B1(new_n798), .B2(new_n729), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n791), .A2(new_n795), .ZN(new_n892));
  NAND4_X1  g706(.A1(new_n879), .A2(new_n891), .A3(new_n892), .A4(new_n782), .ZN(new_n893));
  INV_X1    g707(.A(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n785), .B1(new_n723), .B2(new_n730), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n746), .A2(new_n726), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n401), .A2(new_n736), .A3(new_n741), .A4(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(KEYINPUT52), .A3(new_n752), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n752), .A2(new_n898), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n900), .B1(new_n901), .B2(new_n895), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n902), .ZN(new_n903));
  INV_X1    g717(.A(KEYINPUT112), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n883), .A2(new_n880), .A3(new_n593), .ZN(new_n905));
  AOI21_X1  g719(.A(KEYINPUT111), .B1(new_n591), .B2(new_n594), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n904), .B(new_n644), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n886), .B2(new_n644), .ZN(new_n909));
  OAI211_X1 g723(.A(new_n718), .B(new_n652), .C1(new_n908), .C2(new_n909), .ZN(new_n910));
  OAI22_X1  g724(.A1(new_n910), .A2(new_n697), .B1(new_n719), .B2(new_n714), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n488), .A2(new_n533), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n718), .A2(new_n652), .A3(new_n841), .ZN(new_n913));
  OAI22_X1  g727(.A1(new_n912), .A2(new_n719), .B1(new_n697), .B2(new_n913), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n911), .B1(KEYINPUT110), .B2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT110), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n655), .A2(new_n681), .A3(new_n916), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT113), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n914), .A2(KEYINPUT110), .ZN(new_n919));
  INV_X1    g733(.A(new_n909), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n658), .B1(new_n920), .B2(new_n907), .ZN(new_n921));
  INV_X1    g735(.A(new_n719), .ZN(new_n922));
  NOR3_X1   g736(.A1(new_n677), .A2(new_n679), .A3(new_n736), .ZN(new_n923));
  AOI22_X1  g737(.A1(new_n698), .A2(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n919), .A2(new_n917), .A3(new_n924), .A4(KEYINPUT113), .ZN(new_n925));
  INV_X1    g739(.A(new_n925), .ZN(new_n926));
  OAI211_X1 g740(.A(new_n894), .B(new_n903), .C1(new_n918), .C2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n919), .A2(new_n917), .A3(new_n924), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT113), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g744(.A(new_n893), .B1(new_n930), .B2(new_n925), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n752), .A2(new_n898), .A3(KEYINPUT52), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n895), .A2(KEYINPUT114), .ZN(new_n933));
  INV_X1    g747(.A(KEYINPUT114), .ZN(new_n934));
  OAI211_X1 g748(.A(new_n785), .B(new_n934), .C1(new_n723), .C2(new_n730), .ZN(new_n935));
  NAND3_X1  g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n936), .B2(new_n902), .ZN(new_n937));
  AOI22_X1  g751(.A1(new_n927), .A2(KEYINPUT53), .B1(new_n931), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n938), .A2(KEYINPUT54), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT53), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n927), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n879), .A2(new_n782), .A3(new_n892), .ZN(new_n942));
  AOI22_X1  g756(.A1(new_n902), .A2(new_n936), .B1(new_n942), .B2(KEYINPUT115), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n930), .A2(new_n925), .ZN(new_n944));
  AND2_X1   g758(.A1(new_n891), .A2(KEYINPUT53), .ZN(new_n945));
  INV_X1    g759(.A(KEYINPUT115), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n879), .A2(new_n892), .A3(new_n946), .A4(new_n782), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n943), .A2(new_n944), .A3(new_n945), .A4(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(KEYINPUT54), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n941), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n830), .B1(new_n878), .B2(new_n951), .ZN(new_n952));
  INV_X1    g766(.A(KEYINPUT49), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n859), .A2(new_n953), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n859), .A2(new_n953), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n533), .A2(new_n325), .A3(new_n192), .ZN(new_n956));
  NOR4_X1   g770(.A1(new_n954), .A2(new_n955), .A3(new_n801), .A4(new_n956), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n957), .A2(new_n842), .A3(new_n744), .ZN(new_n958));
  XNOR2_X1  g772(.A(new_n958), .B(KEYINPUT109), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n952), .A2(new_n959), .ZN(G75));
  NAND2_X1  g774(.A1(new_n936), .A2(new_n902), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n782), .A2(new_n757), .A3(new_n760), .A4(new_n763), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT115), .B1(new_n962), .B2(new_n796), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n961), .A2(new_n963), .A3(new_n947), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n945), .B1(new_n918), .B2(new_n926), .ZN(new_n966));
  INV_X1    g780(.A(new_n966), .ZN(new_n967));
  AOI22_X1  g781(.A1(new_n965), .A2(new_n967), .B1(new_n927), .B2(new_n940), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n968), .A2(new_n190), .ZN(new_n969));
  AOI21_X1  g783(.A(KEYINPUT56), .B1(new_n969), .B2(G210), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n353), .B1(new_n375), .B2(new_n376), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n971), .A2(new_n397), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n972), .A2(new_n377), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n973), .B(KEYINPUT55), .Z(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n970), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n295), .A2(G952), .ZN(new_n977));
  INV_X1    g791(.A(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n978), .B1(new_n970), .B2(new_n975), .ZN(new_n979));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n979), .ZN(G51));
  NOR3_X1   g794(.A1(new_n968), .A2(new_n190), .A3(new_n809), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n964), .A2(new_n966), .ZN(new_n982));
  AOI21_X1  g796(.A(KEYINPUT53), .B1(new_n931), .B2(new_n903), .ZN(new_n983));
  OAI21_X1  g797(.A(KEYINPUT54), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(new_n950), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n686), .B(KEYINPUT57), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n322), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n981), .B1(new_n987), .B2(KEYINPUT122), .ZN(new_n988));
  INV_X1    g802(.A(KEYINPUT122), .ZN(new_n989));
  INV_X1    g803(.A(new_n986), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n990), .B1(new_n984), .B2(new_n950), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n989), .B1(new_n991), .B2(new_n322), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n977), .B1(new_n988), .B2(new_n992), .ZN(G54));
  NAND3_X1  g807(.A1(new_n969), .A2(KEYINPUT58), .A3(G475), .ZN(new_n994));
  AND2_X1   g808(.A1(new_n994), .A2(new_n703), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n703), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n977), .ZN(G60));
  INV_X1    g811(.A(new_n666), .ZN(new_n998));
  NAND2_X1  g812(.A1(G478), .A2(G902), .ZN(new_n999));
  XNOR2_X1  g813(.A(new_n999), .B(KEYINPUT59), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n985), .A2(new_n998), .A3(new_n1000), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n998), .B1(new_n951), .B2(new_n1000), .ZN(new_n1002));
  NOR3_X1   g816(.A1(new_n1001), .A2(new_n1002), .A3(new_n977), .ZN(G63));
  XNOR2_X1  g817(.A(KEYINPUT125), .B(KEYINPUT61), .ZN(new_n1004));
  INV_X1    g818(.A(new_n1004), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n522), .A2(new_n523), .ZN(new_n1006));
  XNOR2_X1  g820(.A(KEYINPUT123), .B(KEYINPUT60), .ZN(new_n1007));
  NOR2_X1   g821(.A1(new_n571), .A2(new_n190), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1009), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1006), .B1(new_n968), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n941), .A2(new_n948), .ZN(new_n1012));
  NAND4_X1  g826(.A1(new_n1012), .A2(KEYINPUT124), .A3(new_n711), .A4(new_n1009), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1011), .A2(new_n1013), .A3(new_n978), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n1010), .B1(new_n941), .B2(new_n948), .ZN(new_n1015));
  AOI21_X1  g829(.A(KEYINPUT124), .B1(new_n1015), .B2(new_n711), .ZN(new_n1016));
  OAI21_X1  g830(.A(new_n1005), .B1(new_n1014), .B2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1015), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n977), .B1(new_n1018), .B2(new_n1006), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1016), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1019), .A2(new_n1020), .A3(new_n1013), .A4(new_n1004), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n1017), .A2(new_n1021), .ZN(G66));
  INV_X1    g836(.A(new_n649), .ZN(new_n1023));
  OAI21_X1  g837(.A(G953), .B1(new_n1023), .B2(new_n358), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n962), .B1(new_n930), .B2(new_n925), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(G953), .ZN(new_n1026));
  INV_X1    g840(.A(new_n971), .ZN(new_n1027));
  OAI21_X1  g841(.A(new_n1027), .B1(G898), .B2(new_n295), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n1026), .B(new_n1028), .ZN(G69));
  AOI21_X1  g843(.A(new_n295), .B1(G227), .B2(G900), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1030), .A2(KEYINPUT127), .ZN(new_n1031));
  OR2_X1    g845(.A1(new_n1030), .A2(KEYINPUT127), .ZN(new_n1032));
  AND3_X1   g846(.A1(new_n933), .A2(new_n752), .A3(new_n935), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n818), .A2(new_n1033), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT126), .ZN(new_n1035));
  NAND2_X1  g849(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n818), .A2(KEYINPUT126), .A3(new_n1033), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n817), .A2(new_n733), .ZN(new_n1039));
  NAND3_X1  g853(.A1(new_n837), .A2(new_n718), .A3(new_n745), .ZN(new_n1040));
  OAI211_X1 g854(.A(new_n892), .B(new_n799), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NOR2_X1   g855(.A1(new_n828), .A2(new_n1041), .ZN(new_n1042));
  NAND2_X1  g856(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n469), .B(new_n628), .ZN(new_n1044));
  INV_X1    g858(.A(new_n1044), .ZN(new_n1045));
  NOR2_X1   g859(.A1(new_n1045), .A2(G953), .ZN(new_n1046));
  AOI22_X1  g860(.A1(new_n1043), .A2(new_n1046), .B1(new_n725), .B2(G953), .ZN(new_n1047));
  INV_X1    g861(.A(new_n1047), .ZN(new_n1048));
  INV_X1    g862(.A(new_n818), .ZN(new_n1049));
  NAND3_X1  g863(.A1(new_n920), .A2(new_n672), .A3(new_n907), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n798), .A2(new_n733), .A3(new_n1050), .ZN(new_n1051));
  NOR3_X1   g865(.A1(new_n828), .A2(new_n1049), .A3(new_n1051), .ZN(new_n1052));
  NAND2_X1  g866(.A1(new_n1033), .A2(new_n748), .ZN(new_n1053));
  OR2_X1    g867(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1053), .A2(KEYINPUT62), .ZN(new_n1055));
  NAND3_X1  g869(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .ZN(new_n1056));
  AOI21_X1  g870(.A(new_n1044), .B1(new_n1056), .B2(new_n295), .ZN(new_n1057));
  OAI211_X1 g871(.A(new_n1031), .B(new_n1032), .C1(new_n1048), .C2(new_n1057), .ZN(new_n1058));
  INV_X1    g872(.A(new_n1057), .ZN(new_n1059));
  NAND4_X1  g873(.A1(new_n1059), .A2(new_n1047), .A3(KEYINPUT127), .A4(new_n1030), .ZN(new_n1060));
  AND2_X1   g874(.A1(new_n1058), .A2(new_n1060), .ZN(G72));
  NAND2_X1  g875(.A1(G472), .A2(G902), .ZN(new_n1062));
  XNOR2_X1  g876(.A(new_n1062), .B(KEYINPUT63), .ZN(new_n1063));
  OR2_X1    g877(.A1(new_n470), .A2(new_n455), .ZN(new_n1064));
  AOI21_X1  g878(.A(new_n1063), .B1(new_n1064), .B2(new_n457), .ZN(new_n1065));
  NAND2_X1  g879(.A1(new_n938), .A2(new_n1065), .ZN(new_n1066));
  NAND2_X1  g880(.A1(new_n1066), .A2(new_n978), .ZN(new_n1067));
  INV_X1    g881(.A(new_n1056), .ZN(new_n1068));
  AOI21_X1  g882(.A(new_n1063), .B1(new_n1068), .B2(new_n1025), .ZN(new_n1069));
  INV_X1    g883(.A(new_n1043), .ZN(new_n1070));
  AOI21_X1  g884(.A(new_n1063), .B1(new_n1070), .B2(new_n1025), .ZN(new_n1071));
  OAI22_X1  g885(.A1(new_n470), .A2(new_n1069), .B1(new_n1071), .B2(new_n455), .ZN(new_n1072));
  AOI21_X1  g886(.A(new_n1067), .B1(new_n1072), .B2(new_n1064), .ZN(G57));
endmodule


