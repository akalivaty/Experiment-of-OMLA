//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 0 1 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 1 1 0 1 0 1 0 0 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n693, new_n694,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n757, new_n758, new_n759, new_n761, new_n762, new_n763, new_n765,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n856, new_n857, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n921, new_n922, new_n923, new_n924, new_n925, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  XOR2_X1   g005(.A(G43gat), .B(G50gat), .Z(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  OR2_X1    g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G29gat), .A2(G36gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n207), .A2(new_n208), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  INV_X1    g012(.A(new_n213), .ZN(new_n214));
  NOR3_X1   g013(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n215));
  OR2_X1    g014(.A1(new_n215), .A2(KEYINPUT104), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT104), .ZN(new_n217));
  AOI21_X1  g016(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(new_n215), .ZN(new_n219));
  AOI22_X1  g018(.A1(new_n219), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n220));
  OAI22_X1  g019(.A1(new_n212), .A2(new_n218), .B1(new_n220), .B2(new_n209), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n206), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n222), .B(KEYINPUT106), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n223), .B1(new_n221), .B2(new_n206), .ZN(new_n224));
  NAND2_X1  g023(.A1(G229gat), .A2(G233gat), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n225), .B(KEYINPUT105), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(KEYINPUT13), .Z(new_n227));
  NAND2_X1  g026(.A1(new_n224), .A2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT107), .ZN(new_n229));
  XNOR2_X1  g028(.A(new_n228), .B(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT17), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n221), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n206), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n221), .A2(new_n231), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n232), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  AND2_X1   g034(.A1(new_n223), .A2(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n226), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT18), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n236), .A2(KEYINPUT18), .A3(new_n226), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n230), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XOR2_X1   g040(.A(KEYINPUT102), .B(KEYINPUT11), .Z(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT103), .ZN(new_n243));
  XOR2_X1   g042(.A(G113gat), .B(G141gat), .Z(new_n244));
  XNOR2_X1  g043(.A(new_n243), .B(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT12), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n241), .A2(new_n249), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n230), .A2(new_n248), .A3(new_n239), .A4(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  XOR2_X1   g052(.A(KEYINPUT65), .B(KEYINPUT25), .Z(new_n254));
  NAND2_X1  g053(.A1(G169gat), .A2(G176gat), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT23), .ZN(new_n257));
  NOR2_X1   g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(G169gat), .A2(G176gat), .ZN(new_n259));
  XNOR2_X1  g058(.A(KEYINPUT67), .B(G176gat), .ZN(new_n260));
  INV_X1    g059(.A(G169gat), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(KEYINPUT23), .ZN(new_n262));
  OAI22_X1  g061(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(G183gat), .A2(G190gat), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND4_X1  g065(.A1(KEYINPUT66), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AND3_X1   g069(.A1(new_n266), .A2(new_n267), .A3(new_n270), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n254), .B1(new_n263), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(KEYINPUT25), .B1(new_n262), .B2(G176gat), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n259), .B1(KEYINPUT23), .B2(new_n255), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n276));
  OR2_X1    g075(.A1(KEYINPUT69), .A2(KEYINPUT24), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT69), .A2(KEYINPUT24), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n265), .A2(KEYINPUT68), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT70), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(KEYINPUT70), .A2(G190gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  OAI21_X1  g085(.A(new_n268), .B1(new_n286), .B2(G183gat), .ZN(new_n287));
  OAI21_X1  g086(.A(new_n275), .B1(new_n281), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n272), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT72), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT71), .A2(G183gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n291), .A2(KEYINPUT27), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT27), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n293), .A2(KEYINPUT71), .A3(G183gat), .ZN(new_n294));
  NAND4_X1  g093(.A1(new_n292), .A2(new_n294), .A3(new_n284), .A4(new_n285), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT28), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(KEYINPUT70), .A2(G190gat), .ZN(new_n298));
  NOR2_X1   g097(.A1(KEYINPUT70), .A2(G190gat), .ZN(new_n299));
  NOR3_X1   g098(.A1(new_n298), .A2(new_n299), .A3(new_n296), .ZN(new_n300));
  XNOR2_X1  g099(.A(KEYINPUT27), .B(G183gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(G176gat), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n261), .A2(new_n304), .A3(KEYINPUT26), .ZN(new_n305));
  INV_X1    g104(.A(KEYINPUT26), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n306), .B1(G169gat), .B2(G176gat), .ZN(new_n307));
  OAI211_X1 g106(.A(new_n305), .B(new_n265), .C1(new_n307), .C2(new_n256), .ZN(new_n308));
  INV_X1    g107(.A(new_n308), .ZN(new_n309));
  AOI21_X1  g108(.A(new_n290), .B1(new_n303), .B2(new_n309), .ZN(new_n310));
  AOI211_X1 g109(.A(KEYINPUT72), .B(new_n308), .C1(new_n297), .C2(new_n302), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n289), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(G127gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G134gat), .ZN(new_n314));
  INV_X1    g113(.A(G134gat), .ZN(new_n315));
  NOR2_X1   g114(.A1(new_n315), .A2(G127gat), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT73), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n315), .A2(G127gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n313), .A2(G134gat), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(G113gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  AOI21_X1  g122(.A(KEYINPUT1), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(G113gat), .A2(G120gat), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n317), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n318), .A2(new_n319), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n328), .A2(KEYINPUT73), .A3(new_n325), .A4(new_n324), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n327), .A2(KEYINPUT74), .A3(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(KEYINPUT74), .B1(new_n327), .B2(new_n329), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT75), .ZN(new_n332));
  NOR3_X1   g131(.A1(new_n330), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n327), .A2(new_n329), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT74), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT74), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT75), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n312), .B1(new_n333), .B2(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n336), .A2(KEYINPUT75), .A3(new_n337), .ZN(new_n340));
  AOI22_X1  g139(.A1(new_n296), .A2(new_n295), .B1(new_n300), .B2(new_n301), .ZN(new_n341));
  OAI21_X1  g140(.A(KEYINPUT72), .B1(new_n341), .B2(new_n308), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n303), .A2(new_n290), .A3(new_n309), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n340), .A2(new_n344), .A3(new_n289), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(G227gat), .A2(G233gat), .ZN(new_n347));
  XOR2_X1   g146(.A(new_n347), .B(KEYINPUT64), .Z(new_n348));
  AOI21_X1  g147(.A(KEYINPUT76), .B1(new_n346), .B2(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT76), .ZN(new_n350));
  INV_X1    g149(.A(new_n348), .ZN(new_n351));
  AOI211_X1 g150(.A(new_n350), .B(new_n351), .C1(new_n339), .C2(new_n345), .ZN(new_n352));
  OAI21_X1  g151(.A(KEYINPUT32), .B1(new_n349), .B2(new_n352), .ZN(new_n353));
  XOR2_X1   g152(.A(G15gat), .B(G43gat), .Z(new_n354));
  XNOR2_X1  g153(.A(new_n354), .B(KEYINPUT78), .ZN(new_n355));
  XNOR2_X1  g154(.A(G71gat), .B(G99gat), .ZN(new_n356));
  XOR2_X1   g155(.A(new_n355), .B(new_n356), .Z(new_n357));
  AOI21_X1  g156(.A(new_n353), .B1(KEYINPUT33), .B2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(new_n358), .ZN(new_n359));
  OR3_X1    g158(.A1(new_n346), .A2(KEYINPUT34), .A3(new_n348), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT81), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  XOR2_X1   g161(.A(KEYINPUT80), .B(KEYINPUT34), .Z(new_n363));
  INV_X1    g162(.A(new_n347), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n363), .B1(new_n346), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n360), .A2(new_n361), .ZN(new_n366));
  AND3_X1   g165(.A1(new_n362), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT79), .ZN(new_n368));
  INV_X1    g167(.A(new_n357), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n332), .B1(new_n330), .B2(new_n331), .ZN(new_n370));
  AOI22_X1  g169(.A1(new_n370), .A2(new_n340), .B1(new_n344), .B2(new_n289), .ZN(new_n371));
  NOR2_X1   g170(.A1(new_n312), .A2(new_n333), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n348), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(new_n350), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n346), .A2(KEYINPUT76), .A3(new_n348), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT33), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n369), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n379), .B1(new_n376), .B2(KEYINPUT32), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT32), .ZN(new_n381));
  AOI211_X1 g180(.A(KEYINPUT77), .B(new_n381), .C1(new_n374), .C2(new_n375), .ZN(new_n382));
  OAI211_X1 g181(.A(new_n368), .B(new_n378), .C1(new_n380), .C2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n353), .A2(KEYINPUT77), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n379), .A3(KEYINPUT32), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n368), .B1(new_n387), .B2(new_n378), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n359), .B(new_n367), .C1(new_n384), .C2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n378), .B1(new_n380), .B2(new_n382), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n391), .A2(KEYINPUT79), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n358), .B1(new_n392), .B2(new_n383), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT83), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n393), .A2(new_n394), .A3(new_n367), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n390), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(G228gat), .A2(G233gat), .ZN(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT22), .ZN(new_n399));
  XNOR2_X1  g198(.A(KEYINPUT84), .B(G211gat), .ZN(new_n400));
  INV_X1    g199(.A(G218gat), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n399), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g201(.A(G197gat), .B(G204gat), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(G211gat), .B(G218gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n404), .A2(new_n405), .ZN(new_n408));
  OR2_X1    g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT3), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  XOR2_X1   g210(.A(G155gat), .B(G162gat), .Z(new_n412));
  INV_X1    g211(.A(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G155gat), .ZN(new_n414));
  INV_X1    g213(.A(G162gat), .ZN(new_n415));
  OAI21_X1  g214(.A(KEYINPUT2), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  XOR2_X1   g215(.A(G141gat), .B(G148gat), .Z(new_n417));
  AND3_X1   g216(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n416), .A2(KEYINPUT88), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT88), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n420), .B(KEYINPUT2), .C1(new_n414), .C2(new_n415), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n419), .A2(new_n417), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n412), .ZN(new_n423));
  OR2_X1    g222(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n423), .A2(KEYINPUT89), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n418), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  OAI21_X1  g225(.A(new_n398), .B1(new_n411), .B2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  XOR2_X1   g228(.A(KEYINPUT85), .B(KEYINPUT29), .Z(new_n430));
  NAND2_X1  g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n409), .B1(new_n431), .B2(KEYINPUT97), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT97), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n433), .A3(new_n430), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n427), .B1(new_n432), .B2(new_n434), .ZN(new_n435));
  XOR2_X1   g234(.A(new_n397), .B(KEYINPUT95), .Z(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n406), .A2(KEYINPUT96), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n438), .A2(new_n408), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n430), .B1(new_n406), .B2(KEYINPUT96), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n428), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n426), .A2(KEYINPUT92), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n426), .A2(KEYINPUT92), .ZN(new_n444));
  OAI21_X1  g243(.A(new_n441), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n409), .B1(new_n429), .B2(new_n430), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n437), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(G22gat), .B1(new_n435), .B2(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n424), .A2(new_n425), .ZN(new_n451));
  INV_X1    g250(.A(new_n418), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT92), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  OR2_X1    g254(.A1(new_n406), .A2(KEYINPUT96), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n456), .B(new_n430), .C1(new_n408), .C2(new_n438), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n455), .A2(new_n442), .B1(new_n457), .B2(new_n428), .ZN(new_n458));
  OAI21_X1  g257(.A(new_n436), .B1(new_n458), .B2(new_n446), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n431), .A2(KEYINPUT97), .ZN(new_n460));
  INV_X1    g259(.A(new_n409), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n460), .A2(new_n461), .A3(new_n434), .ZN(new_n462));
  OAI211_X1 g261(.A(new_n450), .B(new_n459), .C1(new_n462), .C2(new_n427), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n449), .A2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT98), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n462), .B2(new_n427), .ZN(new_n466));
  AOI21_X1  g265(.A(new_n465), .B1(new_n466), .B2(G22gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(G78gat), .B(G106gat), .ZN(new_n468));
  XNOR2_X1  g267(.A(KEYINPUT31), .B(G50gat), .ZN(new_n469));
  XNOR2_X1  g268(.A(new_n468), .B(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(new_n470), .ZN(new_n471));
  OAI21_X1  g270(.A(new_n464), .B1(new_n467), .B2(new_n471), .ZN(new_n472));
  NAND4_X1  g271(.A1(new_n449), .A2(new_n463), .A3(new_n465), .A4(new_n470), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n392), .A2(new_n383), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n367), .B1(new_n475), .B2(new_n359), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G8gat), .B(G36gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(KEYINPUT86), .ZN(new_n479));
  XOR2_X1   g278(.A(G64gat), .B(G92gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(G226gat), .A2(G233gat), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n312), .A2(new_n482), .ZN(new_n483));
  AOI22_X1  g282(.A1(new_n272), .A2(new_n288), .B1(new_n303), .B2(new_n309), .ZN(new_n484));
  INV_X1    g283(.A(new_n482), .ZN(new_n485));
  NOR3_X1   g284(.A1(new_n484), .A2(KEYINPUT29), .A3(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n409), .B1(new_n483), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n312), .A2(new_n482), .A3(new_n430), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n484), .A2(new_n485), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n461), .A2(new_n488), .A3(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n481), .B1(new_n487), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT30), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n487), .A2(new_n490), .A3(new_n481), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n487), .A2(new_n490), .A3(KEYINPUT30), .A4(new_n481), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT87), .ZN(new_n496));
  AND2_X1   g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g296(.A1(new_n495), .A2(new_n496), .ZN(new_n498));
  OAI21_X1  g297(.A(new_n494), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(new_n429), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n334), .B(KEYINPUT90), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n501), .B1(new_n426), .B2(new_n428), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n336), .A2(new_n337), .ZN(new_n504));
  NAND4_X1  g303(.A1(new_n455), .A2(KEYINPUT4), .A3(new_n442), .A4(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(G225gat), .A2(G233gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT91), .ZN(new_n507));
  INV_X1    g306(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n426), .A2(new_n334), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT4), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n503), .A2(new_n505), .A3(new_n508), .A4(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT5), .ZN(new_n513));
  INV_X1    g312(.A(new_n501), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n509), .B1(new_n426), .B2(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n513), .B1(new_n515), .B2(new_n507), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n500), .A2(new_n502), .ZN(new_n518));
  NOR3_X1   g317(.A1(new_n518), .A2(KEYINPUT5), .A3(new_n507), .ZN(new_n519));
  INV_X1    g318(.A(new_n509), .ZN(new_n520));
  OAI21_X1  g319(.A(KEYINPUT94), .B1(new_n520), .B2(new_n510), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n455), .A2(new_n510), .A3(new_n442), .A4(new_n504), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n509), .A2(new_n523), .A3(KEYINPUT4), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n521), .A2(new_n522), .A3(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n519), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n517), .A2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G1gat), .B(G29gat), .Z(new_n528));
  XNOR2_X1  g327(.A(G57gat), .B(G85gat), .ZN(new_n529));
  XNOR2_X1  g328(.A(new_n528), .B(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(KEYINPUT93), .B(KEYINPUT0), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n527), .A2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(KEYINPUT6), .ZN(new_n534));
  INV_X1    g333(.A(new_n532), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n517), .A2(new_n526), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n533), .A2(new_n534), .A3(new_n536), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n527), .A2(KEYINPUT6), .A3(new_n532), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n499), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT35), .ZN(new_n540));
  AND2_X1   g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND4_X1  g340(.A1(new_n396), .A2(new_n474), .A3(new_n477), .A4(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n449), .A2(KEYINPUT98), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n543), .A2(new_n470), .B1(new_n463), .B2(new_n449), .ZN(new_n544));
  INV_X1    g343(.A(new_n473), .ZN(new_n545));
  NOR2_X1   g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n359), .B1(new_n384), .B2(new_n388), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n367), .B(KEYINPUT82), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n546), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NOR2_X1   g348(.A1(new_n389), .A2(KEYINPUT83), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n394), .B1(new_n393), .B2(new_n367), .ZN(new_n551));
  OAI211_X1 g350(.A(new_n549), .B(new_n539), .C1(new_n550), .C2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n542), .B1(new_n553), .B2(new_n540), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT36), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n477), .C1(new_n550), .C2(new_n551), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n539), .A2(new_n474), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n537), .A2(new_n538), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT37), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n487), .A2(new_n490), .A3(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n461), .B1(new_n483), .B2(new_n486), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n488), .A2(new_n409), .A3(new_n489), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(new_n562), .A3(KEYINPUT37), .ZN(new_n563));
  XOR2_X1   g362(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n564));
  NOR2_X1   g363(.A1(new_n481), .A2(new_n564), .ZN(new_n565));
  NAND3_X1  g364(.A1(new_n560), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n566), .A2(new_n493), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n559), .B1(new_n487), .B2(new_n490), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT101), .ZN(new_n569));
  OR3_X1    g368(.A1(new_n568), .A2(new_n569), .A3(new_n481), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n569), .B1(new_n568), .B2(new_n481), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(new_n560), .A3(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n567), .B1(new_n572), .B2(new_n564), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n546), .B1(new_n558), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(KEYINPUT99), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n525), .A2(new_n503), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n507), .ZN(new_n577));
  OAI21_X1  g376(.A(new_n535), .B1(new_n577), .B2(KEYINPUT39), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT39), .B1(new_n515), .B2(new_n507), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n579), .B1(new_n576), .B2(new_n507), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n575), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n581), .A2(KEYINPUT40), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT40), .ZN(new_n583));
  OAI211_X1 g382(.A(new_n575), .B(new_n583), .C1(new_n578), .C2(new_n580), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n582), .A2(new_n533), .A3(new_n499), .A4(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n557), .B1(new_n574), .B2(new_n585), .ZN(new_n586));
  AOI22_X1  g385(.A1(new_n390), .A2(new_n395), .B1(new_n547), .B2(new_n548), .ZN(new_n587));
  OAI211_X1 g386(.A(new_n556), .B(new_n586), .C1(new_n555), .C2(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n253), .B1(new_n554), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT113), .ZN(new_n590));
  NAND2_X1  g389(.A1(G71gat), .A2(G78gat), .ZN(new_n591));
  OAI21_X1  g390(.A(KEYINPUT108), .B1(G71gat), .B2(G78gat), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NOR3_X1   g392(.A1(KEYINPUT108), .A2(G71gat), .A3(G78gat), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n591), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n595), .B(KEYINPUT109), .ZN(new_n596));
  XOR2_X1   g395(.A(G57gat), .B(G64gat), .Z(new_n597));
  INV_X1    g396(.A(new_n591), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(KEYINPUT9), .B2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  OR3_X1    g400(.A1(new_n599), .A2(new_n598), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(G85gat), .A2(G92gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n604), .B(KEYINPUT7), .ZN(new_n605));
  NAND2_X1  g404(.A1(G99gat), .A2(G106gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT8), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n605), .B(new_n607), .C1(G85gat), .C2(G92gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(G99gat), .B(G106gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n603), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT111), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n611), .A2(new_n612), .A3(KEYINPUT10), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n611), .B2(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n603), .A2(KEYINPUT10), .A3(new_n610), .ZN(new_n615));
  NAND3_X1  g414(.A1(new_n613), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(G230gat), .A2(G233gat), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n611), .A2(G230gat), .A3(G233gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(G120gat), .B(G148gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(G176gat), .B(G204gat), .ZN(new_n621));
  XOR2_X1   g420(.A(new_n620), .B(new_n621), .Z(new_n622));
  NAND3_X1  g421(.A1(new_n618), .A2(new_n619), .A3(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT112), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n616), .A2(new_n625), .A3(new_n617), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n625), .B1(new_n616), .B2(new_n617), .ZN(new_n628));
  OAI21_X1  g427(.A(new_n619), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n622), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n610), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n232), .A2(new_n234), .A3(new_n633), .ZN(new_n634));
  AND2_X1   g433(.A1(G232gat), .A2(G233gat), .ZN(new_n635));
  AOI22_X1  g434(.A1(new_n610), .A2(new_n221), .B1(KEYINPUT41), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT110), .ZN(new_n638));
  XNOR2_X1  g437(.A(G190gat), .B(G218gat), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n637), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G134gat), .B(G162gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n639), .A2(new_n638), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n635), .A2(KEYINPUT41), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n643), .B(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OR2_X1    g445(.A1(new_n642), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n642), .A2(new_n646), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n603), .A2(KEYINPUT21), .ZN(new_n650));
  NAND2_X1  g449(.A1(G231gat), .A2(G233gat), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n650), .B(new_n651), .Z(new_n652));
  XNOR2_X1  g451(.A(new_n652), .B(new_n313), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n206), .B1(new_n603), .B2(KEYINPUT21), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n652), .B(G127gat), .ZN(new_n656));
  INV_X1    g455(.A(new_n654), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(new_n414), .ZN(new_n660));
  XNOR2_X1  g459(.A(G183gat), .B(G211gat), .ZN(new_n661));
  XOR2_X1   g460(.A(new_n660), .B(new_n661), .Z(new_n662));
  NAND3_X1  g461(.A1(new_n655), .A2(new_n658), .A3(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  AOI21_X1  g463(.A(new_n662), .B1(new_n655), .B2(new_n658), .ZN(new_n665));
  OAI21_X1  g464(.A(new_n649), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n590), .B1(new_n632), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n665), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(new_n663), .ZN(new_n669));
  NAND4_X1  g468(.A1(new_n669), .A2(KEYINPUT113), .A3(new_n631), .A4(new_n649), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n589), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n558), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XOR2_X1   g473(.A(new_n674), .B(G1gat), .Z(G1324gat));
  INV_X1    g474(.A(new_n499), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT16), .B(G8gat), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(G8gat), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n679), .B1(new_n680), .B2(new_n677), .ZN(new_n681));
  MUX2_X1   g480(.A(new_n679), .B(new_n681), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g481(.A1(new_n548), .A2(new_n547), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n396), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n684), .A2(KEYINPUT36), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(new_n556), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(G15gat), .B1(new_n672), .B2(new_n687), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n396), .A2(new_n477), .ZN(new_n689));
  OR2_X1    g488(.A1(new_n689), .A2(G15gat), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n688), .B1(new_n672), .B2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(KEYINPUT114), .ZN(G1326gat));
  NOR2_X1   g491(.A1(new_n672), .A2(new_n474), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT43), .B(G22gat), .Z(new_n694));
  XNOR2_X1  g493(.A(new_n693), .B(new_n694), .ZN(G1327gat));
  INV_X1    g494(.A(new_n649), .ZN(new_n696));
  INV_X1    g495(.A(new_n588), .ZN(new_n697));
  AOI211_X1 g496(.A(new_n546), .B(new_n476), .C1(new_n390), .C2(new_n395), .ZN(new_n698));
  AOI22_X1  g497(.A1(new_n698), .A2(new_n541), .B1(new_n552), .B2(KEYINPUT35), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n696), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  INV_X1    g499(.A(new_n669), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n631), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n702), .A2(new_n253), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NOR4_X1   g503(.A1(new_n700), .A2(G29gat), .A3(new_n673), .A4(new_n704), .ZN(new_n705));
  XOR2_X1   g504(.A(new_n705), .B(KEYINPUT45), .Z(new_n706));
  AOI21_X1  g505(.A(new_n649), .B1(new_n554), .B2(new_n588), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n707), .A2(KEYINPUT44), .ZN(new_n708));
  OAI211_X1 g507(.A(KEYINPUT44), .B(new_n696), .C1(new_n697), .C2(new_n699), .ZN(new_n709));
  INV_X1    g508(.A(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n708), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n703), .ZN(new_n712));
  OAI21_X1  g511(.A(G29gat), .B1(new_n712), .B2(new_n673), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n706), .A2(new_n713), .ZN(G1328gat));
  NOR2_X1   g513(.A1(new_n700), .A2(new_n704), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n676), .A2(G36gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n715), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT115), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT46), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  OAI21_X1  g519(.A(G36gat), .B1(new_n712), .B2(new_n676), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n717), .A2(KEYINPUT115), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n717), .A2(KEYINPUT115), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(KEYINPUT46), .A3(new_n723), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n720), .A2(new_n721), .A3(new_n724), .ZN(G1329gat));
  INV_X1    g524(.A(KEYINPUT44), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n700), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n727), .A2(new_n686), .A3(new_n703), .A4(new_n709), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n728), .A2(G43gat), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT116), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT47), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(new_n689), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n702), .A2(G43gat), .A3(new_n649), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n589), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n729), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n731), .A2(new_n735), .ZN(new_n736));
  OAI211_X1 g535(.A(new_n729), .B(new_n734), .C1(new_n730), .C2(KEYINPUT47), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1330gat));
  NAND4_X1  g537(.A1(new_n727), .A2(new_n546), .A3(new_n703), .A4(new_n709), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n739), .A2(G50gat), .ZN(new_n740));
  NOR2_X1   g539(.A1(new_n474), .A2(G50gat), .ZN(new_n741));
  AND3_X1   g540(.A1(new_n707), .A2(new_n703), .A3(new_n741), .ZN(new_n742));
  INV_X1    g541(.A(new_n742), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT117), .ZN(new_n745));
  AOI21_X1  g544(.A(KEYINPUT48), .B1(new_n744), .B2(new_n745), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n742), .B1(new_n739), .B2(G50gat), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT48), .ZN(new_n748));
  NOR3_X1   g547(.A1(new_n747), .A2(KEYINPUT117), .A3(new_n748), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n746), .A2(new_n749), .ZN(G1331gat));
  NAND2_X1  g549(.A1(new_n554), .A2(new_n588), .ZN(new_n751));
  NOR3_X1   g550(.A1(new_n666), .A2(new_n252), .A3(new_n631), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(new_n558), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g555(.A(new_n676), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  XOR2_X1   g558(.A(new_n758), .B(new_n759), .Z(G1333gat));
  OR3_X1    g559(.A1(new_n753), .A2(G71gat), .A3(new_n689), .ZN(new_n761));
  OAI21_X1  g560(.A(G71gat), .B1(new_n753), .B2(new_n687), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  XOR2_X1   g562(.A(new_n763), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g563(.A1(new_n754), .A2(new_n546), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g565(.A1(new_n673), .A2(G85gat), .A3(new_n631), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n669), .A2(new_n252), .ZN(new_n768));
  AOI21_X1  g567(.A(KEYINPUT51), .B1(new_n707), .B2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT118), .ZN(new_n771));
  INV_X1    g570(.A(new_n768), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT51), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n707), .A2(new_n771), .A3(new_n774), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g575(.A(new_n771), .B1(new_n707), .B2(new_n774), .ZN(new_n777));
  OAI211_X1 g576(.A(new_n770), .B(KEYINPUT119), .C1(new_n776), .C2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n751), .A2(new_n696), .A3(new_n774), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n780), .A2(KEYINPUT118), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n769), .B1(new_n781), .B2(new_n775), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n782), .A2(KEYINPUT119), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n767), .B1(new_n779), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n772), .A2(new_n631), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n711), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(new_n558), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G85gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n784), .A2(new_n788), .ZN(G1336gat));
  OAI21_X1  g588(.A(new_n770), .B1(new_n776), .B2(new_n777), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n631), .A2(G92gat), .A3(new_n676), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n790), .A2(KEYINPUT121), .A3(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT121), .ZN(new_n793));
  INV_X1    g592(.A(new_n791), .ZN(new_n794));
  OAI21_X1  g593(.A(new_n793), .B1(new_n782), .B2(new_n794), .ZN(new_n795));
  NAND4_X1  g594(.A1(new_n727), .A2(new_n499), .A3(new_n709), .A4(new_n785), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT52), .B1(new_n796), .B2(G92gat), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n792), .A2(new_n795), .A3(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n796), .A2(G92gat), .ZN(new_n799));
  OAI211_X1 g598(.A(new_n696), .B(new_n768), .C1(new_n697), .C2(new_n699), .ZN(new_n800));
  AOI22_X1  g599(.A1(new_n800), .A2(new_n773), .B1(new_n707), .B2(new_n774), .ZN(new_n801));
  OAI21_X1  g600(.A(KEYINPUT120), .B1(new_n801), .B2(new_n794), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n799), .A2(new_n802), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n801), .A2(KEYINPUT120), .A3(new_n794), .ZN(new_n804));
  OAI21_X1  g603(.A(KEYINPUT52), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n798), .A2(new_n805), .ZN(G1337gat));
  NOR3_X1   g605(.A1(new_n689), .A2(G99gat), .A3(new_n631), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n807), .B1(new_n779), .B2(new_n783), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n786), .A2(new_n686), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G99gat), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(G1338gat));
  NAND4_X1  g610(.A1(new_n711), .A2(KEYINPUT122), .A3(new_n546), .A4(new_n785), .ZN(new_n812));
  NAND4_X1  g611(.A1(new_n727), .A2(new_n546), .A3(new_n709), .A4(new_n785), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n812), .A2(new_n815), .A3(G106gat), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n631), .A2(new_n474), .A3(G106gat), .ZN(new_n817));
  AOI21_X1  g616(.A(KEYINPUT53), .B1(new_n790), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n816), .A2(new_n818), .ZN(new_n819));
  NOR4_X1   g618(.A1(new_n801), .A2(G106gat), .A3(new_n474), .A4(new_n631), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n813), .A2(G106gat), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT53), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n819), .A2(new_n822), .ZN(G1339gat));
  NAND2_X1  g622(.A1(new_n618), .A2(KEYINPUT112), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(new_n825), .A3(new_n626), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n825), .B1(new_n616), .B2(new_n617), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(new_n617), .B2(new_n616), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n630), .A3(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND4_X1  g630(.A1(new_n826), .A2(KEYINPUT55), .A3(new_n630), .A4(new_n828), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n236), .A2(new_n226), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n224), .A2(new_n227), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n247), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n251), .A2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n831), .A2(new_n832), .A3(new_n623), .A4(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n669), .B1(new_n837), .B2(new_n696), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n696), .B1(new_n632), .B2(new_n836), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n831), .A2(new_n832), .A3(new_n252), .A4(new_n623), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n666), .A2(new_n252), .ZN(new_n842));
  AOI22_X1  g641(.A1(new_n838), .A2(new_n841), .B1(new_n631), .B2(new_n842), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n396), .A2(new_n549), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n673), .A2(new_n499), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(G113gat), .B1(new_n847), .B2(new_n252), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n838), .A2(new_n841), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n842), .A2(new_n631), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n851), .A2(new_n698), .A3(new_n845), .ZN(new_n852));
  INV_X1    g651(.A(new_n852), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n253), .A2(new_n322), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n848), .B1(new_n853), .B2(new_n854), .ZN(G1340gat));
  AOI21_X1  g654(.A(G120gat), .B1(new_n847), .B2(new_n632), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n631), .A2(new_n323), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n856), .B1(new_n853), .B2(new_n857), .ZN(G1341gat));
  NOR3_X1   g657(.A1(new_n852), .A2(new_n313), .A3(new_n701), .ZN(new_n859));
  INV_X1    g658(.A(new_n847), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n860), .A2(KEYINPUT123), .A3(new_n701), .ZN(new_n861));
  NOR2_X1   g660(.A1(new_n861), .A2(G127gat), .ZN(new_n862));
  OAI21_X1  g661(.A(KEYINPUT123), .B1(new_n860), .B2(new_n701), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n859), .B1(new_n862), .B2(new_n863), .ZN(G1342gat));
  NOR3_X1   g663(.A1(new_n860), .A2(G134gat), .A3(new_n649), .ZN(new_n865));
  INV_X1    g664(.A(new_n865), .ZN(new_n866));
  OR2_X1    g665(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n867));
  OAI21_X1  g666(.A(G134gat), .B1(new_n852), .B2(new_n649), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(KEYINPUT56), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(G1343gat));
  NAND2_X1  g669(.A1(new_n687), .A2(new_n845), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n851), .A2(new_n546), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(G141gat), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n873), .A2(new_n874), .A3(new_n252), .ZN(new_n875));
  AOI21_X1  g674(.A(KEYINPUT57), .B1(new_n851), .B2(new_n546), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT57), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n843), .A2(new_n877), .A3(new_n474), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NOR3_X1   g678(.A1(new_n879), .A2(new_n253), .A3(new_n871), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n875), .B1(new_n880), .B2(new_n874), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(KEYINPUT58), .ZN(G1344gat));
  INV_X1    g681(.A(KEYINPUT124), .ZN(new_n883));
  INV_X1    g682(.A(new_n871), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(new_n632), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n671), .A2(new_n253), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n849), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(KEYINPUT57), .B1(new_n887), .B2(new_n546), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(new_n878), .ZN(new_n889));
  OAI21_X1  g688(.A(G148gat), .B1(new_n885), .B2(new_n889), .ZN(new_n890));
  OAI211_X1 g689(.A(new_n884), .B(new_n632), .C1(new_n876), .C2(new_n878), .ZN(new_n891));
  INV_X1    g690(.A(G148gat), .ZN(new_n892));
  NOR2_X1   g691(.A1(new_n892), .A2(KEYINPUT59), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n890), .A2(KEYINPUT59), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n873), .A2(new_n892), .A3(new_n632), .ZN(new_n895));
  INV_X1    g694(.A(new_n895), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n883), .B1(new_n894), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT59), .ZN(new_n898));
  AOI22_X1  g697(.A1(new_n838), .A2(new_n841), .B1(new_n671), .B2(new_n253), .ZN(new_n899));
  OAI21_X1  g698(.A(new_n877), .B1(new_n899), .B2(new_n474), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n900), .B1(new_n872), .B2(new_n877), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n901), .A2(new_n632), .A3(new_n884), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n898), .B1(new_n902), .B2(G148gat), .ZN(new_n903));
  AND2_X1   g702(.A1(new_n891), .A2(new_n893), .ZN(new_n904));
  OAI211_X1 g703(.A(KEYINPUT124), .B(new_n895), .C1(new_n903), .C2(new_n904), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n897), .A2(new_n905), .ZN(G1345gat));
  NAND3_X1  g705(.A1(new_n873), .A2(new_n414), .A3(new_n669), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n879), .A2(new_n701), .A3(new_n871), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n907), .B1(new_n908), .B2(new_n414), .ZN(G1346gat));
  AOI21_X1  g708(.A(G162gat), .B1(new_n873), .B2(new_n696), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n879), .A2(new_n871), .ZN(new_n911));
  NOR2_X1   g710(.A1(new_n649), .A2(new_n415), .ZN(new_n912));
  AOI21_X1  g711(.A(new_n910), .B1(new_n911), .B2(new_n912), .ZN(G1347gat));
  NOR3_X1   g712(.A1(new_n843), .A2(new_n558), .A3(new_n676), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(new_n698), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n261), .A3(new_n253), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n844), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n252), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n261), .B2(new_n919), .ZN(G1348gat));
  AND4_X1   g719(.A1(new_n260), .A2(new_n914), .A3(new_n698), .A4(new_n632), .ZN(new_n921));
  OAI21_X1  g720(.A(new_n304), .B1(new_n917), .B2(new_n631), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT125), .ZN(new_n923));
  OR2_X1    g722(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n922), .A2(new_n923), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1349gat));
  OAI21_X1  g725(.A(G183gat), .B1(new_n915), .B2(new_n701), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n669), .A2(new_n301), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n927), .B1(new_n917), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g729(.A(G190gat), .B1(new_n915), .B2(new_n649), .ZN(new_n931));
  XNOR2_X1  g730(.A(new_n931), .B(KEYINPUT61), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n649), .A2(new_n286), .ZN(new_n933));
  OAI21_X1  g732(.A(new_n932), .B1(new_n917), .B2(new_n933), .ZN(G1351gat));
  INV_X1    g733(.A(KEYINPUT127), .ZN(new_n935));
  INV_X1    g734(.A(G197gat), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n901), .A2(KEYINPUT126), .ZN(new_n937));
  INV_X1    g736(.A(new_n878), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT126), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n938), .A2(new_n939), .A3(new_n900), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n558), .A2(new_n676), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n687), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(new_n253), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n936), .B1(new_n941), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n944), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n946), .A2(G197gat), .A3(new_n872), .ZN(new_n947));
  OAI21_X1  g746(.A(new_n935), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n939), .B1(new_n938), .B2(new_n900), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n888), .A2(new_n878), .A3(KEYINPUT126), .ZN(new_n950));
  NOR2_X1   g749(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g750(.A(G197gat), .B1(new_n951), .B2(new_n946), .ZN(new_n952));
  INV_X1    g751(.A(new_n947), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(KEYINPUT127), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n948), .A2(new_n954), .ZN(G1352gat));
  INV_X1    g754(.A(new_n943), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n632), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n957), .A2(G204gat), .A3(new_n872), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT62), .ZN(new_n959));
  OAI21_X1  g758(.A(G204gat), .B1(new_n951), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n959), .A2(new_n960), .ZN(G1353gat));
  OR2_X1    g760(.A1(new_n943), .A2(new_n872), .ZN(new_n962));
  INV_X1    g761(.A(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n400), .A3(new_n669), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n901), .A2(new_n669), .A3(new_n956), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g766(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n968));
  OAI21_X1  g767(.A(new_n964), .B1(new_n967), .B2(new_n968), .ZN(G1354gat));
  NAND2_X1  g768(.A1(new_n956), .A2(new_n696), .ZN(new_n970));
  OAI21_X1  g769(.A(G218gat), .B1(new_n951), .B2(new_n970), .ZN(new_n971));
  NAND3_X1  g770(.A1(new_n963), .A2(new_n401), .A3(new_n696), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(G1355gat));
endmodule


