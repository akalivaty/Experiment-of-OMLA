//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 0 1 1 1 1 0 1 0 1 0 0 0 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:08 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n717, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n764, new_n765, new_n766, new_n767, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n785, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n833, new_n834, new_n835, new_n836, new_n837, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n893, new_n894, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n987, new_n988, new_n989, new_n990, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1009, new_n1010;
  INV_X1    g000(.A(G22gat), .ZN(new_n202));
  NAND2_X1  g001(.A1(new_n202), .A2(G15gat), .ZN(new_n203));
  INV_X1    g002(.A(G15gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G1gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT16), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n203), .A2(new_n205), .A3(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(KEYINPUT89), .B(G8gat), .ZN(new_n209));
  XNOR2_X1  g008(.A(G15gat), .B(G22gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n208), .B(new_n209), .C1(G1gat), .C2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G8gat), .ZN(new_n212));
  AOI21_X1  g011(.A(G1gat), .B1(new_n203), .B2(new_n205), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT87), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI211_X1 g014(.A(new_n208), .B(KEYINPUT87), .C1(G1gat), .C2(new_n210), .ZN(new_n216));
  AND3_X1   g015(.A1(new_n215), .A2(new_n216), .A3(KEYINPUT88), .ZN(new_n217));
  AOI21_X1  g016(.A(KEYINPUT88), .B1(new_n215), .B2(new_n216), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n211), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT90), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT85), .ZN(new_n221));
  AND2_X1   g020(.A1(G43gat), .A2(G50gat), .ZN(new_n222));
  NOR2_X1   g021(.A1(G43gat), .A2(G50gat), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(G43gat), .ZN(new_n225));
  INV_X1    g024(.A(G50gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G43gat), .A2(G50gat), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(KEYINPUT85), .A3(new_n228), .ZN(new_n229));
  AND3_X1   g028(.A1(new_n224), .A2(new_n229), .A3(KEYINPUT15), .ZN(new_n230));
  OAI21_X1  g029(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n231), .A2(KEYINPUT86), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT86), .ZN(new_n233));
  OAI211_X1 g032(.A(new_n233), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n235));
  INV_X1    g034(.A(G29gat), .ZN(new_n236));
  INV_X1    g035(.A(G36gat), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n235), .A2(new_n236), .A3(new_n237), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n232), .A2(new_n234), .A3(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(G29gat), .A2(G36gat), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n230), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n229), .A3(KEYINPUT15), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n238), .A2(new_n231), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT15), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n227), .A2(new_n245), .A3(new_n228), .ZN(new_n246));
  NAND4_X1  g045(.A1(new_n243), .A2(new_n240), .A3(new_n244), .A4(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n242), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT17), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT17), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n242), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT90), .ZN(new_n253));
  OAI211_X1 g052(.A(new_n253), .B(new_n211), .C1(new_n217), .C2(new_n218), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n220), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(G229gat), .A2(G233gat), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n219), .A2(new_n248), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT18), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g059(.A1(new_n255), .A2(KEYINPUT18), .A3(new_n256), .A4(new_n257), .ZN(new_n261));
  XNOR2_X1  g060(.A(new_n219), .B(new_n248), .ZN(new_n262));
  XOR2_X1   g061(.A(new_n256), .B(KEYINPUT13), .Z(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n260), .A2(new_n261), .A3(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G113gat), .B(G141gat), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT83), .B(G197gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(new_n266), .B(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(KEYINPUT11), .B(G169gat), .ZN(new_n269));
  XNOR2_X1  g068(.A(new_n268), .B(new_n269), .ZN(new_n270));
  XOR2_X1   g069(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n271));
  XOR2_X1   g070(.A(new_n270), .B(new_n271), .Z(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND4_X1  g073(.A1(new_n260), .A2(new_n261), .A3(new_n264), .A4(new_n272), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT82), .ZN(new_n278));
  INV_X1    g077(.A(G134gat), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n279), .A2(G127gat), .ZN(new_n280));
  INV_X1    g079(.A(G127gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G134gat), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT1), .ZN(new_n283));
  AND3_X1   g082(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NOR2_X1   g083(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(KEYINPUT67), .A2(G120gat), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(KEYINPUT68), .A3(G113gat), .A4(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(new_n287), .ZN(new_n289));
  INV_X1    g088(.A(G113gat), .ZN(new_n290));
  NOR3_X1   g089(.A1(new_n289), .A2(new_n285), .A3(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT68), .ZN(new_n292));
  INV_X1    g091(.A(G120gat), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n292), .B1(new_n293), .B2(G113gat), .ZN(new_n294));
  OAI211_X1 g093(.A(new_n284), .B(new_n288), .C1(new_n291), .C2(new_n294), .ZN(new_n295));
  OR2_X1    g094(.A1(new_n280), .A2(KEYINPUT66), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n282), .A3(KEYINPUT66), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n297), .C1(KEYINPUT1), .C2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(G190gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n301), .A2(G183gat), .ZN(new_n302));
  INV_X1    g101(.A(G183gat), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(G190gat), .ZN(new_n304));
  OAI21_X1  g103(.A(KEYINPUT24), .B1(new_n302), .B2(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(G169gat), .A2(G176gat), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(G169gat), .A2(G176gat), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n308), .A2(KEYINPUT23), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n307), .A2(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT24), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(G183gat), .A3(G190gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT23), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(G176gat), .ZN(new_n314));
  INV_X1    g113(.A(G169gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n315), .A2(KEYINPUT65), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT65), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n317), .A2(G169gat), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n314), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n305), .A2(new_n310), .A3(new_n312), .A4(new_n319), .ZN(new_n320));
  XOR2_X1   g119(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n321));
  INV_X1    g120(.A(new_n312), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n303), .A2(G190gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n301), .A2(G183gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n322), .B1(new_n325), .B2(KEYINPUT24), .ZN(new_n326));
  INV_X1    g125(.A(G176gat), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n327), .A2(KEYINPUT23), .ZN(new_n328));
  OAI21_X1  g127(.A(KEYINPUT25), .B1(new_n328), .B2(G169gat), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n306), .B1(KEYINPUT23), .B2(new_n308), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI22_X1  g130(.A1(new_n320), .A2(new_n321), .B1(new_n326), .B2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT26), .ZN(new_n333));
  NAND3_X1  g132(.A1(new_n307), .A2(new_n333), .A3(new_n308), .ZN(new_n334));
  AOI22_X1  g133(.A1(new_n306), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  XNOR2_X1  g135(.A(KEYINPUT27), .B(G183gat), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT28), .B1(new_n337), .B2(new_n301), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n336), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI21_X1  g140(.A(new_n300), .B1(new_n332), .B2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G227gat), .ZN(new_n343));
  INV_X1    g142(.A(G233gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n295), .A2(new_n299), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n337), .A2(KEYINPUT28), .A3(new_n301), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n334), .B(new_n335), .C1(new_n347), .C2(new_n338), .ZN(new_n348));
  INV_X1    g147(.A(new_n321), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT65), .B(G169gat), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n350), .A2(new_n314), .B1(new_n309), .B2(new_n307), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n349), .B1(new_n326), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT25), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n353), .B1(new_n314), .B2(new_n315), .ZN(new_n354));
  AND4_X1   g153(.A1(new_n305), .A2(new_n354), .A3(new_n312), .A4(new_n310), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n346), .B(new_n348), .C1(new_n352), .C2(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n342), .A2(new_n345), .A3(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(KEYINPUT32), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT33), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n357), .A2(new_n359), .ZN(new_n360));
  XOR2_X1   g159(.A(G15gat), .B(G43gat), .Z(new_n361));
  XNOR2_X1  g160(.A(G71gat), .B(G99gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  NAND3_X1  g162(.A1(new_n358), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n363), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n357), .B(KEYINPUT32), .C1(new_n359), .C2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n364), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(KEYINPUT69), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT34), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n342), .A2(new_n356), .ZN(new_n370));
  INV_X1    g169(.A(new_n345), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g171(.A(KEYINPUT34), .B(new_n345), .C1(new_n342), .C2(new_n356), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  AND3_X1   g173(.A1(new_n374), .A2(new_n364), .A3(new_n366), .ZN(new_n375));
  INV_X1    g174(.A(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(new_n373), .ZN(new_n377));
  AOI22_X1  g176(.A1(new_n364), .A2(new_n366), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n368), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n367), .A2(KEYINPUT69), .A3(new_n374), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(G228gat), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n382), .A2(new_n344), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g183(.A1(G141gat), .A2(G148gat), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  NOR2_X1   g185(.A1(G141gat), .A2(G148gat), .ZN(new_n387));
  NOR3_X1   g186(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT2), .ZN(new_n388));
  XNOR2_X1  g187(.A(G155gat), .B(G162gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n384), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(G155gat), .B(G162gat), .Z(new_n391));
  INV_X1    g190(.A(G141gat), .ZN(new_n392));
  INV_X1    g191(.A(G148gat), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT2), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n394), .A2(new_n395), .A3(new_n385), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n391), .A2(new_n396), .A3(KEYINPUT73), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n394), .A2(new_n385), .ZN(new_n398));
  INV_X1    g197(.A(G155gat), .ZN(new_n399));
  INV_X1    g198(.A(G162gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n395), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G155gat), .A2(G162gat), .ZN(new_n402));
  AOI22_X1  g201(.A1(new_n398), .A2(KEYINPUT74), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  OR3_X1    g202(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT74), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n390), .A2(new_n397), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT3), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(G211gat), .A2(G218gat), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  AND2_X1   g210(.A1(G197gat), .A2(G204gat), .ZN(new_n412));
  NOR2_X1   g211(.A1(G197gat), .A2(G204gat), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT22), .ZN(new_n415));
  OAI211_X1 g214(.A(new_n408), .B(new_n411), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n411), .A2(new_n408), .ZN(new_n417));
  XNOR2_X1  g216(.A(G197gat), .B(G204gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n408), .A2(new_n415), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n417), .A2(new_n418), .A3(new_n419), .ZN(new_n420));
  AND3_X1   g219(.A1(new_n416), .A2(KEYINPUT70), .A3(new_n420), .ZN(new_n421));
  AOI21_X1  g220(.A(KEYINPUT70), .B1(new_n416), .B2(new_n420), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n383), .B1(new_n407), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT79), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT78), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n416), .A2(new_n420), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n427), .B1(new_n428), .B2(KEYINPUT29), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT29), .B1(new_n416), .B2(new_n420), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n430), .A2(KEYINPUT78), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n429), .A2(new_n406), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n398), .A2(KEYINPUT74), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n401), .A2(new_n402), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n404), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n388), .A2(new_n384), .A3(new_n389), .ZN(new_n436));
  AOI21_X1  g235(.A(KEYINPUT73), .B1(new_n391), .B2(new_n396), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  AOI21_X1  g237(.A(new_n426), .B1(new_n432), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n406), .B1(new_n430), .B2(KEYINPUT78), .ZN(new_n440));
  AOI211_X1 g239(.A(new_n427), .B(KEYINPUT29), .C1(new_n416), .C2(new_n420), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n426), .B(new_n438), .C1(new_n440), .C2(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n425), .B1(new_n439), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n405), .A2(new_n406), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT29), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n428), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n438), .B1(KEYINPUT3), .B2(new_n430), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  INV_X1    g249(.A(new_n383), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n444), .A2(new_n202), .A3(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n438), .B1(new_n440), .B2(new_n441), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT79), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n424), .B1(new_n455), .B2(new_n442), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n383), .B1(new_n448), .B2(new_n449), .ZN(new_n457));
  OAI21_X1  g256(.A(G22gat), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  XNOR2_X1  g257(.A(G78gat), .B(G106gat), .ZN(new_n459));
  XNOR2_X1  g258(.A(KEYINPUT31), .B(G50gat), .ZN(new_n460));
  XNOR2_X1  g259(.A(new_n459), .B(new_n460), .ZN(new_n461));
  AND3_X1   g260(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n461), .B1(new_n453), .B2(new_n458), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n278), .B1(new_n381), .B2(new_n464), .ZN(new_n465));
  NAND2_X1  g264(.A1(G225gat), .A2(G233gat), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  NOR2_X1   g266(.A1(new_n438), .A2(new_n346), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n390), .A2(new_n397), .ZN(new_n469));
  AOI22_X1  g268(.A1(new_n469), .A2(new_n435), .B1(new_n295), .B2(new_n299), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n468), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT75), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n471), .A2(new_n472), .A3(KEYINPUT5), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n438), .A2(new_n346), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n469), .A2(new_n295), .A3(new_n299), .A4(new_n435), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n466), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT75), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n438), .A2(KEYINPUT3), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n445), .A3(new_n346), .ZN(new_n480));
  INV_X1    g279(.A(KEYINPUT4), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n481), .B1(new_n438), .B2(new_n346), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n300), .A2(new_n405), .A3(KEYINPUT4), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n480), .A2(new_n466), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n473), .A2(new_n478), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g284(.A(new_n300), .B1(KEYINPUT3), .B2(new_n438), .ZN(new_n486));
  AOI21_X1  g285(.A(new_n467), .B1(new_n486), .B2(new_n445), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT76), .ZN(new_n488));
  AND3_X1   g287(.A1(new_n482), .A2(new_n483), .A3(new_n488), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n488), .B1(new_n482), .B2(new_n483), .ZN(new_n490));
  OAI211_X1 g289(.A(new_n487), .B(new_n477), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n485), .A2(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(G1gat), .B(G29gat), .ZN(new_n493));
  XNOR2_X1  g292(.A(new_n493), .B(KEYINPUT0), .ZN(new_n494));
  XNOR2_X1  g293(.A(G57gat), .B(G85gat), .ZN(new_n495));
  XOR2_X1   g294(.A(new_n494), .B(new_n495), .Z(new_n496));
  INV_X1    g295(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n492), .A2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT6), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n485), .A2(new_n491), .A3(new_n496), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n498), .A2(new_n499), .A3(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(KEYINPUT77), .A3(new_n499), .A4(new_n500), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n492), .A2(KEYINPUT6), .A3(new_n497), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n503), .A2(new_n504), .A3(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G8gat), .B(G36gat), .ZN(new_n507));
  XNOR2_X1  g306(.A(G64gat), .B(G92gat), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n507), .B(new_n508), .Z(new_n509));
  NAND2_X1  g308(.A1(G226gat), .A2(G233gat), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n510), .B(KEYINPUT71), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(KEYINPUT29), .ZN(new_n512));
  OAI21_X1  g311(.A(new_n512), .B1(new_n332), .B2(new_n341), .ZN(new_n513));
  OAI211_X1 g312(.A(new_n348), .B(new_n511), .C1(new_n352), .C2(new_n355), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(new_n423), .ZN(new_n516));
  NOR2_X1   g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n428), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n518), .B1(new_n513), .B2(new_n514), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n509), .B1(new_n517), .B2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT72), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT30), .ZN(new_n523));
  OAI211_X1 g322(.A(KEYINPUT72), .B(new_n509), .C1(new_n517), .C2(new_n519), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n522), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g324(.A(KEYINPUT30), .B(new_n509), .C1(new_n517), .C2(new_n519), .ZN(new_n526));
  INV_X1    g325(.A(new_n519), .ZN(new_n527));
  INV_X1    g326(.A(new_n509), .ZN(new_n528));
  OAI211_X1 g327(.A(new_n527), .B(new_n528), .C1(new_n515), .C2(new_n516), .ZN(new_n529));
  AND2_X1   g328(.A1(new_n526), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n525), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n461), .ZN(new_n533));
  AOI21_X1  g332(.A(new_n202), .B1(new_n444), .B2(new_n452), .ZN(new_n534));
  NOR3_X1   g333(.A1(new_n456), .A2(new_n457), .A3(G22gat), .ZN(new_n535));
  OAI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n453), .A2(new_n458), .A3(new_n461), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g337(.A1(new_n538), .A2(KEYINPUT82), .A3(new_n379), .A4(new_n380), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n465), .A2(new_n506), .A3(new_n532), .A4(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT35), .ZN(new_n541));
  INV_X1    g340(.A(new_n375), .ZN(new_n542));
  INV_X1    g341(.A(new_n378), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NOR3_X1   g343(.A1(new_n544), .A2(new_n531), .A3(KEYINPUT35), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n501), .A2(new_n505), .ZN(new_n546));
  AND3_X1   g345(.A1(new_n545), .A2(new_n546), .A3(new_n538), .ZN(new_n547));
  INV_X1    g346(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n541), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT37), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n550), .B1(new_n517), .B2(new_n519), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n515), .A2(new_n516), .ZN(new_n552));
  OAI211_X1 g351(.A(new_n552), .B(KEYINPUT37), .C1(new_n428), .C2(new_n515), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT38), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n551), .A2(new_n553), .A3(new_n554), .A4(new_n528), .ZN(new_n555));
  AND3_X1   g354(.A1(new_n555), .A2(new_n522), .A3(new_n524), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(new_n501), .A3(new_n505), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT81), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT81), .ZN(new_n559));
  NAND4_X1  g358(.A1(new_n556), .A2(new_n501), .A3(new_n559), .A4(new_n505), .ZN(new_n560));
  OAI211_X1 g359(.A(new_n527), .B(KEYINPUT37), .C1(new_n515), .C2(new_n516), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(new_n528), .A3(new_n551), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT38), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n558), .A2(new_n560), .A3(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n480), .B1(new_n489), .B2(new_n490), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT39), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n467), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n482), .A2(new_n483), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT76), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n482), .A2(new_n483), .A3(new_n488), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n466), .B1(new_n571), .B2(new_n480), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n474), .A2(new_n475), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT39), .B1(new_n573), .B2(new_n467), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(KEYINPUT80), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT80), .ZN(new_n576));
  OAI211_X1 g375(.A(new_n576), .B(KEYINPUT39), .C1(new_n573), .C2(new_n467), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n567), .B(new_n496), .C1(new_n572), .C2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT40), .ZN(new_n580));
  NAND2_X1  g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n467), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n582), .A2(new_n575), .A3(new_n577), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n583), .A2(KEYINPUT40), .A3(new_n496), .A4(new_n567), .ZN(new_n584));
  NAND4_X1  g383(.A1(new_n581), .A2(new_n584), .A3(new_n531), .A4(new_n498), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(new_n538), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n564), .A2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(new_n506), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n464), .B1(new_n589), .B2(new_n531), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n544), .A2(KEYINPUT36), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n591), .B1(new_n381), .B2(KEYINPUT36), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n588), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n277), .B1(new_n549), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g393(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n595), .B1(G57gat), .B2(G64gat), .ZN(new_n596));
  OR2_X1    g395(.A1(G71gat), .A2(G78gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(G71gat), .A2(G78gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  NOR2_X1   g398(.A1(new_n596), .A2(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(KEYINPUT91), .A2(G57gat), .ZN(new_n601));
  INV_X1    g400(.A(G64gat), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT9), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n606), .B1(new_n602), .B2(new_n601), .ZN(new_n607));
  OAI21_X1  g406(.A(KEYINPUT92), .B1(new_n604), .B2(new_n607), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n601), .A2(new_n602), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n605), .B2(new_n598), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT92), .ZN(new_n611));
  AOI22_X1  g410(.A1(new_n597), .A2(new_n598), .B1(new_n602), .B2(new_n601), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n610), .A2(new_n611), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n600), .B1(new_n608), .B2(new_n613), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n615));
  NAND2_X1  g414(.A1(G231gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n615), .B(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n281), .ZN(new_n618));
  AND2_X1   g417(.A1(new_n614), .A2(KEYINPUT21), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n619), .A2(new_n219), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n622));
  XNOR2_X1  g421(.A(new_n622), .B(new_n399), .ZN(new_n623));
  XOR2_X1   g422(.A(G183gat), .B(G211gat), .Z(new_n624));
  XNOR2_X1  g423(.A(new_n623), .B(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n621), .B(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G134gat), .B(G162gat), .Z(new_n627));
  AND2_X1   g426(.A1(G232gat), .A2(G233gat), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(KEYINPUT41), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n627), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(KEYINPUT97), .ZN(new_n631));
  NAND2_X1  g430(.A1(G99gat), .A2(G106gat), .ZN(new_n632));
  INV_X1    g431(.A(G85gat), .ZN(new_n633));
  INV_X1    g432(.A(G92gat), .ZN(new_n634));
  AOI22_X1  g433(.A1(KEYINPUT8), .A2(new_n632), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(G99gat), .B(G106gat), .ZN(new_n636));
  NAND4_X1  g435(.A1(KEYINPUT93), .A2(KEYINPUT7), .A3(G85gat), .A4(G92gat), .ZN(new_n637));
  NAND3_X1  g436(.A1(KEYINPUT93), .A2(G85gat), .A3(G92gat), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT7), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g439(.A1(new_n635), .A2(new_n636), .A3(new_n637), .A4(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT94), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n632), .A2(KEYINPUT8), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n633), .A2(new_n634), .ZN(new_n644));
  NAND4_X1  g443(.A1(new_n640), .A2(new_n637), .A3(new_n643), .A4(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n636), .ZN(new_n646));
  NAND2_X1  g445(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT95), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g448(.A1(new_n645), .A2(KEYINPUT95), .A3(new_n646), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT96), .B1(new_n642), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT94), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n641), .B(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT96), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n654), .A2(new_n655), .A3(new_n649), .A4(new_n650), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n657), .A2(new_n252), .B1(KEYINPUT41), .B2(new_n628), .ZN(new_n658));
  XOR2_X1   g457(.A(G190gat), .B(G218gat), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n652), .A2(new_n656), .A3(new_n248), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  AOI21_X1  g462(.A(new_n660), .B1(new_n658), .B2(new_n661), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n631), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n658), .A2(new_n661), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n666), .A2(new_n659), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n630), .B(KEYINPUT97), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n667), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n665), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g469(.A1(new_n626), .A2(new_n670), .ZN(new_n671));
  AOI21_X1  g470(.A(new_n611), .B1(new_n610), .B2(new_n612), .ZN(new_n672));
  NOR3_X1   g471(.A1(new_n604), .A2(new_n607), .A3(KEYINPUT92), .ZN(new_n673));
  OAI22_X1  g472(.A1(new_n672), .A2(new_n673), .B1(new_n599), .B2(new_n596), .ZN(new_n674));
  OAI21_X1  g473(.A(new_n674), .B1(new_n642), .B2(new_n651), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT10), .ZN(new_n676));
  AOI21_X1  g475(.A(new_n636), .B1(new_n645), .B2(KEYINPUT98), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(KEYINPUT98), .B2(new_n645), .ZN(new_n678));
  NAND3_X1  g477(.A1(new_n654), .A2(new_n614), .A3(new_n678), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n675), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  AOI211_X1 g479(.A(new_n676), .B(new_n600), .C1(new_n608), .C2(new_n613), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n652), .A2(new_n656), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT99), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n680), .A2(new_n682), .A3(KEYINPUT99), .ZN(new_n686));
  NAND2_X1  g485(.A1(G230gat), .A2(G233gat), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n685), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n687), .B1(new_n675), .B2(new_n679), .ZN(new_n689));
  XOR2_X1   g488(.A(G120gat), .B(G148gat), .Z(new_n690));
  XNOR2_X1  g489(.A(new_n690), .B(KEYINPUT100), .ZN(new_n691));
  XNOR2_X1  g490(.A(G176gat), .B(G204gat), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(new_n693));
  INV_X1    g492(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g493(.A1(new_n689), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n688), .A2(new_n695), .ZN(new_n696));
  XOR2_X1   g495(.A(new_n687), .B(KEYINPUT101), .Z(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n683), .A2(new_n698), .ZN(new_n699));
  INV_X1    g498(.A(new_n689), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n694), .ZN(new_n702));
  AOI21_X1  g501(.A(KEYINPUT102), .B1(new_n696), .B2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n695), .ZN(new_n704));
  INV_X1    g503(.A(new_n687), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n705), .B1(new_n683), .B2(new_n684), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n706), .B2(new_n686), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n693), .B1(new_n699), .B2(new_n700), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n707), .A2(new_n708), .A3(new_n709), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n703), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n671), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n594), .A2(new_n713), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n714), .A2(new_n506), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n206), .ZN(G1324gat));
  XOR2_X1   g515(.A(KEYINPUT16), .B(G8gat), .Z(new_n717));
  NAND4_X1  g516(.A1(new_n594), .A2(new_n531), .A3(new_n713), .A4(new_n717), .ZN(new_n718));
  OAI21_X1  g517(.A(G8gat), .B1(new_n714), .B2(new_n532), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(new_n718), .ZN(new_n720));
  MUX2_X1   g519(.A(new_n718), .B(new_n720), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g520(.A(G15gat), .B1(new_n714), .B2(new_n592), .ZN(new_n722));
  INV_X1    g521(.A(new_n544), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n723), .A2(new_n204), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n714), .B2(new_n724), .ZN(G1326gat));
  NAND2_X1  g524(.A1(new_n594), .A2(new_n464), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n726), .A2(new_n712), .ZN(new_n727));
  XOR2_X1   g526(.A(KEYINPUT43), .B(G22gat), .Z(new_n728));
  XNOR2_X1  g527(.A(new_n727), .B(new_n728), .ZN(G1327gat));
  INV_X1    g528(.A(new_n670), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n730), .B1(new_n549), .B2(new_n593), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n626), .A2(new_n711), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n277), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n731), .A2(new_n733), .ZN(new_n734));
  NOR3_X1   g533(.A1(new_n734), .A2(G29gat), .A3(new_n506), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT45), .Z(new_n736));
  NAND2_X1  g535(.A1(new_n549), .A2(new_n593), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n670), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT44), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n731), .A2(KEYINPUT44), .ZN(new_n741));
  AND2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n733), .B(KEYINPUT103), .Z(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744), .B2(new_n506), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n736), .A2(new_n745), .ZN(G1328gat));
  OAI21_X1  g545(.A(G36gat), .B1(new_n744), .B2(new_n532), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n734), .A2(G36gat), .A3(new_n532), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT46), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n747), .A2(new_n749), .ZN(G1329gat));
  NOR3_X1   g549(.A1(new_n734), .A2(G43gat), .A3(new_n544), .ZN(new_n751));
  INV_X1    g550(.A(new_n592), .ZN(new_n752));
  NAND4_X1  g551(.A1(new_n740), .A2(new_n752), .A3(new_n741), .A4(new_n743), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n751), .B1(new_n753), .B2(G43gat), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(KEYINPUT47), .ZN(G1330gat));
  OR4_X1    g554(.A1(G50gat), .A2(new_n726), .A3(new_n730), .A4(new_n732), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n740), .A2(new_n464), .A3(new_n741), .A4(new_n743), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G50gat), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT48), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n758), .A3(KEYINPUT48), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(G1331gat));
  INV_X1    g562(.A(new_n711), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n671), .A2(new_n277), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n765), .B1(new_n549), .B2(new_n593), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n589), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g567(.A(new_n531), .B(KEYINPUT104), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n771), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT49), .B(G64gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n772), .B1(new_n771), .B2(new_n773), .ZN(G1333gat));
  NAND3_X1  g573(.A1(new_n766), .A2(G71gat), .A3(new_n752), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT105), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n775), .A2(new_n776), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n766), .A2(new_n723), .ZN(new_n779));
  INV_X1    g578(.A(new_n779), .ZN(new_n780));
  OAI22_X1  g579(.A1(new_n777), .A2(new_n778), .B1(G71gat), .B2(new_n780), .ZN(new_n781));
  XNOR2_X1  g580(.A(KEYINPUT106), .B(KEYINPUT50), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n781), .B(new_n782), .Z(G1334gat));
  NAND2_X1  g582(.A1(new_n766), .A2(new_n464), .ZN(new_n784));
  XNOR2_X1  g583(.A(KEYINPUT107), .B(G78gat), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1335gat));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n787));
  INV_X1    g586(.A(new_n626), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n788), .A2(new_n276), .ZN(new_n789));
  INV_X1    g588(.A(new_n505), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n501), .B2(new_n502), .ZN(new_n791));
  AOI21_X1  g590(.A(new_n531), .B1(new_n791), .B2(new_n504), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n592), .B1(new_n792), .B2(new_n538), .ZN(new_n793));
  AOI22_X1  g592(.A1(new_n557), .A2(KEYINPUT81), .B1(KEYINPUT38), .B2(new_n562), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n586), .B1(new_n794), .B2(new_n560), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n547), .B1(new_n540), .B2(KEYINPUT35), .ZN(new_n797));
  OAI211_X1 g596(.A(new_n670), .B(new_n789), .C1(new_n796), .C2(new_n797), .ZN(new_n798));
  INV_X1    g597(.A(KEYINPUT51), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n787), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND4_X1  g599(.A1(new_n731), .A2(KEYINPUT108), .A3(KEYINPUT51), .A4(new_n789), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n798), .A2(new_n799), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT109), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g604(.A1(new_n800), .A2(new_n801), .A3(KEYINPUT109), .A4(new_n802), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NOR3_X1   g606(.A1(new_n506), .A2(new_n711), .A3(G85gat), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT110), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n788), .A2(new_n276), .A3(new_n711), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n740), .A2(new_n589), .A3(new_n741), .A4(new_n811), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n812), .A2(G85gat), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n809), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n808), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n815), .B1(new_n805), .B2(new_n806), .ZN(new_n816));
  INV_X1    g615(.A(new_n813), .ZN(new_n817));
  OAI21_X1  g616(.A(KEYINPUT110), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(G1336gat));
  NAND4_X1  g618(.A1(new_n740), .A2(new_n531), .A3(new_n741), .A4(new_n811), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n820), .A2(G92gat), .ZN(new_n821));
  XNOR2_X1  g620(.A(new_n798), .B(new_n799), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n769), .A2(G92gat), .A3(new_n711), .ZN(new_n823));
  AND2_X1   g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(KEYINPUT52), .B1(new_n821), .B2(new_n824), .ZN(new_n825));
  NAND4_X1  g624(.A1(new_n740), .A2(new_n741), .A3(new_n770), .A4(new_n811), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT52), .B1(new_n826), .B2(G92gat), .ZN(new_n827));
  INV_X1    g626(.A(KEYINPUT111), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n803), .A2(new_n823), .ZN(new_n829));
  AND3_X1   g628(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n828), .B1(new_n827), .B2(new_n829), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n825), .B1(new_n830), .B2(new_n831), .ZN(G1337gat));
  NOR3_X1   g631(.A1(new_n711), .A2(G99gat), .A3(new_n544), .ZN(new_n833));
  XNOR2_X1  g632(.A(new_n833), .B(KEYINPUT112), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n807), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n742), .A2(new_n752), .A3(new_n811), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G99gat), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n835), .A2(new_n837), .ZN(G1338gat));
  NAND3_X1  g637(.A1(new_n742), .A2(new_n464), .A3(new_n811), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(G106gat), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT53), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NOR3_X1   g641(.A1(new_n711), .A2(G106gat), .A3(new_n538), .ZN(new_n843));
  AND2_X1   g642(.A1(new_n803), .A2(new_n843), .ZN(new_n844));
  AOI22_X1  g643(.A1(new_n839), .A2(G106gat), .B1(new_n822), .B2(new_n843), .ZN(new_n845));
  OAI22_X1  g644(.A1(new_n842), .A2(new_n844), .B1(new_n845), .B2(new_n841), .ZN(G1339gat));
  NOR2_X1   g645(.A1(new_n262), .A2(new_n263), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n256), .B1(new_n255), .B2(new_n257), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n270), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AND2_X1   g648(.A1(new_n275), .A2(new_n849), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n850), .A2(new_n670), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n680), .A2(new_n682), .A3(new_n697), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(KEYINPUT54), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n853), .B1(new_n706), .B2(new_n686), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT54), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n683), .A2(new_n855), .A3(new_n698), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n694), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n707), .B1(new_n858), .B2(KEYINPUT55), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT55), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n854), .B2(new_n857), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n851), .A2(KEYINPUT113), .A3(new_n859), .A4(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n850), .A2(new_n670), .A3(new_n861), .ZN(new_n864));
  INV_X1    g663(.A(new_n853), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n688), .A2(new_n865), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n866), .A2(KEYINPUT55), .A3(new_n694), .A4(new_n856), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n696), .ZN(new_n868));
  OAI21_X1  g667(.A(new_n863), .B1(new_n864), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  NAND4_X1  g669(.A1(new_n276), .A2(new_n867), .A3(new_n696), .A4(new_n861), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n850), .B1(new_n703), .B2(new_n710), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n670), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n626), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n671), .A2(new_n277), .A3(new_n711), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n465), .A2(new_n539), .ZN(new_n877));
  AND2_X1   g676(.A1(new_n877), .A2(new_n589), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT115), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n876), .A2(KEYINPUT115), .A3(new_n878), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n770), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n290), .A3(new_n276), .ZN(new_n884));
  AOI211_X1 g683(.A(new_n464), .B(new_n544), .C1(new_n874), .C2(new_n875), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n770), .A2(new_n506), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(G113gat), .B1(new_n887), .B2(new_n277), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT114), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n888), .A2(new_n889), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n884), .B1(new_n890), .B2(new_n891), .ZN(G1340gat));
  NAND4_X1  g691(.A1(new_n883), .A2(new_n286), .A3(new_n287), .A4(new_n764), .ZN(new_n893));
  OAI21_X1  g692(.A(G120gat), .B1(new_n887), .B2(new_n711), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1341gat));
  NAND4_X1  g694(.A1(new_n885), .A2(G127gat), .A3(new_n788), .A4(new_n886), .ZN(new_n896));
  XNOR2_X1  g695(.A(new_n896), .B(KEYINPUT116), .ZN(new_n897));
  AOI21_X1  g696(.A(G127gat), .B1(new_n883), .B2(new_n788), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT117), .ZN(new_n899));
  OR3_X1    g698(.A1(new_n897), .A2(new_n898), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1342gat));
  NAND2_X1  g701(.A1(new_n881), .A2(new_n882), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n730), .A2(new_n531), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n903), .A2(new_n279), .A3(new_n904), .ZN(new_n905));
  OR2_X1    g704(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n906));
  OAI21_X1  g705(.A(G134gat), .B1(new_n887), .B2(new_n730), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(KEYINPUT56), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n906), .A2(new_n907), .A3(new_n908), .ZN(G1343gat));
  NAND2_X1  g708(.A1(new_n886), .A2(new_n592), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n871), .A2(new_n872), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n670), .B1(new_n911), .B2(KEYINPUT118), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT118), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n871), .A2(new_n872), .A3(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n870), .B1(new_n912), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT119), .B1(new_n915), .B2(new_n788), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT119), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n911), .A2(KEYINPUT118), .ZN(new_n918));
  AND3_X1   g717(.A1(new_n918), .A2(new_n730), .A3(new_n914), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n917), .B(new_n626), .C1(new_n919), .C2(new_n870), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n916), .A2(new_n920), .A3(new_n875), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT57), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n538), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n876), .A2(new_n464), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n922), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n910), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n392), .B1(new_n927), .B2(new_n276), .ZN(new_n928));
  NOR3_X1   g727(.A1(new_n925), .A2(new_n506), .A3(new_n752), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n769), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n276), .A2(new_n392), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(KEYINPUT58), .B1(new_n928), .B2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n932), .ZN(new_n934));
  INV_X1    g733(.A(KEYINPUT58), .ZN(new_n935));
  AOI211_X1 g734(.A(new_n277), .B(new_n910), .C1(new_n924), .C2(new_n926), .ZN(new_n936));
  OAI211_X1 g735(.A(new_n934), .B(new_n935), .C1(new_n936), .C2(new_n392), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n933), .A2(new_n937), .ZN(G1344gat));
  NAND4_X1  g737(.A1(new_n929), .A2(new_n393), .A3(new_n764), .A4(new_n769), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n864), .A2(new_n868), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n942), .B1(new_n912), .B2(new_n914), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n875), .B1(new_n943), .B2(new_n788), .ZN(new_n944));
  INV_X1    g743(.A(KEYINPUT122), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n538), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  OAI211_X1 g745(.A(new_n875), .B(KEYINPUT122), .C1(new_n943), .C2(new_n788), .ZN(new_n947));
  AOI21_X1  g746(.A(KEYINPUT57), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g747(.A1(new_n876), .A2(new_n923), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(new_n910), .ZN(new_n951));
  OR2_X1    g750(.A1(new_n951), .A2(KEYINPUT121), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n951), .A2(KEYINPUT121), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n952), .A2(new_n764), .A3(new_n953), .ZN(new_n954));
  OAI211_X1 g753(.A(KEYINPUT59), .B(G148gat), .C1(new_n950), .C2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n393), .B1(new_n927), .B2(new_n764), .ZN(new_n956));
  OAI211_X1 g755(.A(new_n941), .B(new_n955), .C1(KEYINPUT59), .C2(new_n956), .ZN(G1345gat));
  AND2_X1   g756(.A1(new_n927), .A2(new_n788), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n788), .A2(new_n399), .ZN(new_n959));
  OAI22_X1  g758(.A1(new_n958), .A2(new_n399), .B1(new_n930), .B2(new_n959), .ZN(G1346gat));
  NAND2_X1  g759(.A1(new_n924), .A2(new_n926), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(new_n670), .A3(new_n951), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT123), .ZN(new_n963));
  NAND2_X1  g762(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n927), .A2(KEYINPUT123), .A3(new_n670), .ZN(new_n965));
  NAND3_X1  g764(.A1(new_n964), .A2(G162gat), .A3(new_n965), .ZN(new_n966));
  NAND3_X1  g765(.A1(new_n929), .A2(new_n400), .A3(new_n904), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n966), .A2(new_n967), .ZN(G1347gat));
  NAND2_X1  g767(.A1(new_n506), .A2(new_n531), .ZN(new_n969));
  XOR2_X1   g768(.A(new_n969), .B(KEYINPUT125), .Z(new_n970));
  NAND2_X1  g769(.A1(new_n885), .A2(new_n970), .ZN(new_n971));
  OAI21_X1  g770(.A(G169gat), .B1(new_n971), .B2(new_n277), .ZN(new_n972));
  AOI21_X1  g771(.A(new_n589), .B1(new_n874), .B2(new_n875), .ZN(new_n973));
  AND2_X1   g772(.A1(new_n877), .A2(new_n770), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g774(.A(new_n975), .B(KEYINPUT124), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n276), .A2(new_n350), .ZN(new_n977));
  OAI21_X1  g776(.A(new_n972), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  XNOR2_X1  g777(.A(new_n978), .B(KEYINPUT126), .ZN(G1348gat));
  OAI21_X1  g778(.A(G176gat), .B1(new_n971), .B2(new_n711), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n764), .A2(new_n327), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n976), .B2(new_n981), .ZN(G1349gat));
  OAI21_X1  g781(.A(G183gat), .B1(new_n971), .B2(new_n626), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n788), .A2(new_n337), .ZN(new_n984));
  OAI21_X1  g783(.A(new_n983), .B1(new_n975), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g784(.A(new_n985), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g785(.A(G190gat), .B1(new_n971), .B2(new_n730), .ZN(new_n987));
  AND2_X1   g786(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n988));
  NOR2_X1   g787(.A1(new_n987), .A2(KEYINPUT61), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n670), .A2(new_n301), .ZN(new_n990));
  OAI22_X1  g789(.A1(new_n988), .A2(new_n989), .B1(new_n976), .B2(new_n990), .ZN(G1351gat));
  AND4_X1   g790(.A1(new_n464), .A2(new_n973), .A3(new_n592), .A4(new_n770), .ZN(new_n992));
  AOI21_X1  g791(.A(G197gat), .B1(new_n992), .B2(new_n276), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n970), .A2(new_n592), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n950), .A2(new_n995), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n276), .A2(G197gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n993), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  INV_X1    g797(.A(G204gat), .ZN(new_n999));
  NAND3_X1  g798(.A1(new_n992), .A2(new_n999), .A3(new_n764), .ZN(new_n1000));
  XOR2_X1   g799(.A(new_n1000), .B(KEYINPUT62), .Z(new_n1001));
  NOR3_X1   g800(.A1(new_n950), .A2(new_n711), .A3(new_n995), .ZN(new_n1002));
  OAI21_X1  g801(.A(new_n1001), .B1(new_n999), .B2(new_n1002), .ZN(G1353gat));
  NAND3_X1  g802(.A1(new_n992), .A2(new_n409), .A3(new_n788), .ZN(new_n1004));
  OAI211_X1 g803(.A(new_n788), .B(new_n994), .C1(new_n948), .C2(new_n949), .ZN(new_n1005));
  AND3_X1   g804(.A1(new_n1005), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1006));
  AOI21_X1  g805(.A(KEYINPUT63), .B1(new_n1005), .B2(G211gat), .ZN(new_n1007));
  OAI21_X1  g806(.A(new_n1004), .B1(new_n1006), .B2(new_n1007), .ZN(G1354gat));
  NAND3_X1  g807(.A1(new_n992), .A2(new_n410), .A3(new_n670), .ZN(new_n1009));
  NOR3_X1   g808(.A1(new_n950), .A2(new_n730), .A3(new_n995), .ZN(new_n1010));
  OAI21_X1  g809(.A(new_n1009), .B1(new_n1010), .B2(new_n410), .ZN(G1355gat));
endmodule


