//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 0 1 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:17 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n736, new_n737, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n763, new_n764, new_n765, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n775, new_n776, new_n777, new_n778,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n864, new_n865, new_n867, new_n868, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n876, new_n877, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n950, new_n951, new_n952, new_n954, new_n955,
    new_n956, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n986, new_n987, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT87), .ZN(new_n203));
  INV_X1    g002(.A(KEYINPUT16), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n203), .B1(new_n204), .B2(G1gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n202), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g005(.A1(new_n203), .A2(new_n204), .A3(G1gat), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n206), .A2(new_n207), .B1(G1gat), .B2(new_n202), .ZN(new_n208));
  OAI21_X1  g007(.A(KEYINPUT88), .B1(new_n202), .B2(G1gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(G8gat), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n208), .B(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n212));
  OR2_X1    g011(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n213));
  XOR2_X1   g012(.A(G57gat), .B(G64gat), .Z(new_n214));
  NAND2_X1  g013(.A1(new_n212), .A2(KEYINPUT92), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(G71gat), .B(G78gat), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(KEYINPUT93), .B1(new_n216), .B2(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n216), .A2(KEYINPUT93), .A3(new_n218), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  NAND4_X1  g021(.A1(new_n213), .A2(new_n214), .A3(new_n217), .A4(new_n215), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n223), .B(KEYINPUT94), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT21), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT95), .B(KEYINPUT19), .Z(new_n228));
  XNOR2_X1  g027(.A(new_n227), .B(new_n228), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G127gat), .B(G155gat), .ZN(new_n231));
  XOR2_X1   g030(.A(new_n231), .B(KEYINPUT20), .Z(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n225), .A2(new_n226), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(G231gat), .A3(G233gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(G231gat), .A2(G233gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n225), .A2(new_n226), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n233), .B1(new_n235), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n235), .A2(new_n233), .A3(new_n237), .ZN(new_n240));
  XOR2_X1   g039(.A(G183gat), .B(G211gat), .Z(new_n241));
  INV_X1    g040(.A(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n239), .A2(new_n240), .A3(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n242), .B1(new_n239), .B2(new_n240), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n230), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(new_n245), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n247), .A2(new_n229), .A3(new_n243), .ZN(new_n248));
  XOR2_X1   g047(.A(G190gat), .B(G218gat), .Z(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT14), .B(G29gat), .ZN(new_n251));
  INV_X1    g050(.A(G36gat), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(G29gat), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n254), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G50gat), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n258), .A2(G43gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT84), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n258), .A2(KEYINPUT84), .A3(G43gat), .ZN(new_n262));
  XNOR2_X1  g061(.A(KEYINPUT85), .B(G50gat), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n261), .B(new_n262), .C1(new_n263), .C2(G43gat), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT15), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT86), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OR2_X1    g067(.A1(new_n258), .A2(G43gat), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n269), .A2(new_n259), .A3(KEYINPUT15), .ZN(new_n270));
  AOI21_X1  g069(.A(new_n257), .B1(new_n268), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(new_n270), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n264), .A2(KEYINPUT86), .A3(new_n265), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n272), .B1(new_n273), .B2(new_n256), .ZN(new_n274));
  NOR2_X1   g073(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(G99gat), .A2(G106gat), .ZN(new_n276));
  INV_X1    g075(.A(G85gat), .ZN(new_n277));
  INV_X1    g076(.A(G92gat), .ZN(new_n278));
  AOI22_X1  g077(.A1(KEYINPUT8), .A2(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(KEYINPUT98), .A3(new_n281), .ZN(new_n282));
  AND2_X1   g081(.A1(new_n280), .A2(KEYINPUT98), .ZN(new_n283));
  OAI21_X1  g082(.A(KEYINPUT7), .B1(new_n280), .B2(KEYINPUT98), .ZN(new_n284));
  OAI211_X1 g083(.A(new_n279), .B(new_n282), .C1(new_n283), .C2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G99gat), .B(G106gat), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G232gat), .A2(G233gat), .ZN(new_n288));
  XOR2_X1   g087(.A(new_n288), .B(KEYINPUT96), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n275), .A2(new_n287), .B1(KEYINPUT41), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g090(.A(KEYINPUT17), .B1(new_n271), .B2(new_n274), .ZN(new_n292));
  INV_X1    g091(.A(new_n274), .ZN(new_n293));
  INV_X1    g092(.A(KEYINPUT17), .ZN(new_n294));
  AOI21_X1  g093(.A(KEYINPUT86), .B1(new_n264), .B2(new_n265), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n256), .B1(new_n295), .B2(new_n272), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n293), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n287), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n292), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n250), .B1(new_n291), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(new_n300), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n290), .A2(KEYINPUT41), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n302), .B(KEYINPUT97), .Z(new_n303));
  XOR2_X1   g102(.A(G134gat), .B(G162gat), .Z(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n291), .A2(new_n299), .A3(new_n250), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n301), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n305), .ZN(new_n308));
  INV_X1    g107(.A(new_n306), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n308), .B1(new_n309), .B2(new_n300), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n307), .A2(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(new_n311), .ZN(new_n312));
  AND3_X1   g111(.A1(new_n216), .A2(KEYINPUT93), .A3(new_n218), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n313), .A2(new_n219), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT94), .ZN(new_n315));
  XNOR2_X1  g114(.A(new_n223), .B(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n298), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n222), .A2(new_n224), .A3(new_n287), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT10), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n317), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND4_X1  g119(.A1(new_n222), .A2(new_n224), .A3(KEYINPUT10), .A4(new_n287), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G230gat), .A2(G233gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g123(.A(new_n323), .B1(new_n317), .B2(new_n318), .ZN(new_n325));
  OR2_X1    g124(.A1(new_n325), .A2(KEYINPUT99), .ZN(new_n326));
  XNOR2_X1  g125(.A(G120gat), .B(G148gat), .ZN(new_n327));
  XNOR2_X1  g126(.A(G176gat), .B(G204gat), .ZN(new_n328));
  XOR2_X1   g127(.A(new_n327), .B(new_n328), .Z(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  AOI21_X1  g129(.A(new_n330), .B1(new_n325), .B2(KEYINPUT99), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n324), .A2(new_n326), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(new_n323), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n333), .B1(new_n320), .B2(new_n321), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n330), .B1(new_n334), .B2(new_n325), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND4_X1  g136(.A1(new_n246), .A2(new_n248), .A3(new_n312), .A4(new_n337), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n292), .A2(new_n211), .A3(new_n297), .ZN(new_n339));
  NAND2_X1  g138(.A1(G229gat), .A2(G233gat), .ZN(new_n340));
  INV_X1    g139(.A(new_n211), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n275), .A2(new_n341), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n339), .A2(KEYINPUT18), .A3(new_n340), .A4(new_n342), .ZN(new_n343));
  XOR2_X1   g142(.A(new_n340), .B(KEYINPUT13), .Z(new_n344));
  NOR2_X1   g143(.A1(new_n275), .A2(new_n341), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n211), .A2(new_n271), .A3(new_n274), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n344), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G113gat), .B(G141gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(G197gat), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT11), .B(G169gat), .Z(new_n350));
  XNOR2_X1  g149(.A(new_n349), .B(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n351), .B(KEYINPUT12), .ZN(new_n352));
  AND3_X1   g151(.A1(new_n343), .A2(new_n347), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n339), .A2(new_n340), .A3(new_n342), .ZN(new_n354));
  XNOR2_X1  g153(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n355));
  AND3_X1   g154(.A1(new_n354), .A2(KEYINPUT90), .A3(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(KEYINPUT90), .B1(new_n354), .B2(new_n355), .ZN(new_n357));
  OAI21_X1  g156(.A(new_n353), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(new_n355), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n359), .A2(new_n347), .A3(new_n343), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n352), .B(KEYINPUT83), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n358), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G148gat), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(G155gat), .A2(G162gat), .ZN(new_n368));
  AOI22_X1  g167(.A1(new_n365), .A2(new_n367), .B1(KEYINPUT2), .B2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(new_n368), .ZN(new_n370));
  NOR2_X1   g169(.A1(G155gat), .A2(G162gat), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT73), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G155gat), .ZN(new_n373));
  INV_X1    g172(.A(G162gat), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT73), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n375), .A2(new_n376), .A3(new_n368), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n369), .A2(new_n372), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n375), .A2(new_n368), .ZN(new_n379));
  XNOR2_X1  g178(.A(G141gat), .B(G148gat), .ZN(new_n380));
  AND2_X1   g179(.A1(new_n368), .A2(KEYINPUT2), .ZN(new_n381));
  OAI211_X1 g180(.A(KEYINPUT73), .B(new_n379), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n378), .A2(new_n382), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT74), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n378), .A2(new_n382), .A3(KEYINPUT74), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n385), .A2(KEYINPUT3), .A3(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT65), .ZN(new_n388));
  INV_X1    g187(.A(G127gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n389), .A2(G134gat), .ZN(new_n390));
  INV_X1    g189(.A(G134gat), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n391), .A2(G127gat), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n388), .B1(new_n390), .B2(new_n392), .ZN(new_n393));
  INV_X1    g192(.A(G113gat), .ZN(new_n394));
  INV_X1    g193(.A(G120gat), .ZN(new_n395));
  NOR2_X1   g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT1), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(G113gat), .B2(G120gat), .ZN(new_n398));
  NOR2_X1   g197(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n391), .A2(G127gat), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n389), .A2(G134gat), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT65), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n393), .A2(new_n399), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G127gat), .B(G134gat), .ZN(new_n404));
  OAI211_X1 g203(.A(new_n404), .B(KEYINPUT65), .C1(new_n396), .C2(new_n398), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n403), .A2(new_n405), .ZN(new_n406));
  XOR2_X1   g205(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(new_n383), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n387), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g208(.A1(new_n406), .A2(new_n383), .A3(KEYINPUT4), .ZN(new_n410));
  AOI21_X1  g209(.A(KEYINPUT4), .B1(new_n406), .B2(new_n383), .ZN(new_n411));
  NOR2_X1   g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(G225gat), .A2(G233gat), .ZN(new_n413));
  NAND4_X1  g212(.A1(new_n409), .A2(new_n412), .A3(KEYINPUT5), .A4(new_n413), .ZN(new_n414));
  AND3_X1   g213(.A1(new_n409), .A2(new_n412), .A3(new_n413), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT5), .ZN(new_n416));
  AND2_X1   g215(.A1(new_n403), .A2(new_n405), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n385), .A2(new_n386), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n406), .A2(new_n383), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n413), .ZN(new_n421));
  AOI21_X1  g220(.A(new_n416), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n414), .B1(new_n415), .B2(new_n422), .ZN(new_n423));
  XOR2_X1   g222(.A(G1gat), .B(G29gat), .Z(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT76), .B(KEYINPUT0), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n424), .B(new_n425), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n423), .A2(new_n429), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT6), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n428), .B(new_n414), .C1(new_n415), .C2(new_n422), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  OR3_X1    g232(.A1(new_n423), .A2(new_n431), .A3(new_n429), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT22), .ZN(new_n436));
  INV_X1    g235(.A(G211gat), .ZN(new_n437));
  INV_X1    g236(.A(G218gat), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AND2_X1   g238(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n440));
  NOR2_X1   g239(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n441));
  INV_X1    g240(.A(G204gat), .ZN(new_n442));
  NOR3_X1   g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT67), .ZN(new_n444));
  INV_X1    g243(.A(G197gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(KEYINPUT67), .A2(G197gat), .ZN(new_n447));
  AOI21_X1  g246(.A(G204gat), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n439), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n437), .A2(new_n438), .ZN(new_n450));
  NOR2_X1   g249(.A1(G211gat), .A2(G218gat), .ZN(new_n451));
  OR2_X1    g250(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n442), .B1(new_n440), .B2(new_n441), .ZN(new_n455));
  NAND3_X1  g254(.A1(new_n446), .A2(G204gat), .A3(new_n447), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n452), .A3(new_n439), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(G226gat), .ZN(new_n460));
  INV_X1    g259(.A(G233gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT25), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT23), .ZN(new_n465));
  INV_X1    g264(.A(G169gat), .ZN(new_n466));
  INV_X1    g265(.A(G176gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G169gat), .A2(G176gat), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT64), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(KEYINPUT64), .A2(G169gat), .A3(G176gat), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g275(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT24), .ZN(new_n478));
  INV_X1    g277(.A(G183gat), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(G190gat), .ZN(new_n480));
  INV_X1    g279(.A(G190gat), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n481), .A2(G183gat), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n477), .B1(new_n480), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n464), .B1(new_n476), .B2(new_n483), .ZN(new_n484));
  AOI22_X1  g283(.A1(new_n469), .A2(new_n468), .B1(new_n473), .B2(new_n474), .ZN(new_n485));
  INV_X1    g284(.A(new_n477), .ZN(new_n486));
  OAI21_X1  g285(.A(KEYINPUT24), .B1(new_n481), .B2(G183gat), .ZN(new_n487));
  NOR2_X1   g286(.A1(new_n479), .A2(G190gat), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n485), .A2(KEYINPUT25), .A3(new_n489), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NOR3_X1   g291(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AOI22_X1  g293(.A1(new_n494), .A2(new_n475), .B1(G183gat), .B2(G190gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n479), .A2(KEYINPUT27), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT27), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(G183gat), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n496), .A2(new_n498), .A3(new_n481), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT28), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(KEYINPUT27), .B(G183gat), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n502), .A2(KEYINPUT28), .A3(new_n481), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n484), .A2(new_n490), .B1(new_n495), .B2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n463), .B1(new_n505), .B2(KEYINPUT29), .ZN(new_n506));
  INV_X1    g305(.A(new_n493), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n475), .A2(new_n507), .A3(new_n491), .ZN(new_n508));
  NAND2_X1  g307(.A1(G183gat), .A2(G190gat), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT28), .B1(new_n502), .B2(new_n481), .ZN(new_n510));
  AND4_X1   g309(.A1(KEYINPUT28), .A2(new_n496), .A3(new_n498), .A4(new_n481), .ZN(new_n511));
  OAI211_X1 g310(.A(new_n508), .B(new_n509), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n485), .A2(KEYINPUT25), .A3(new_n489), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT25), .B1(new_n485), .B2(new_n489), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n462), .ZN(new_n516));
  AOI211_X1 g315(.A(KEYINPUT68), .B(new_n459), .C1(new_n506), .C2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n506), .A2(new_n516), .ZN(new_n519));
  INV_X1    g318(.A(new_n459), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n518), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT69), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n522), .B1(new_n505), .B2(new_n463), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n515), .A2(KEYINPUT69), .A3(new_n462), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g324(.A1(new_n525), .A2(new_n459), .A3(new_n506), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n517), .B1(new_n521), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g326(.A(G8gat), .B(G36gat), .Z(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(KEYINPUT70), .ZN(new_n529));
  XNOR2_X1  g328(.A(G64gat), .B(G92gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(new_n531), .ZN(new_n532));
  OAI21_X1  g331(.A(KEYINPUT30), .B1(new_n527), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n519), .A2(new_n518), .A3(new_n520), .ZN(new_n534));
  AND3_X1   g333(.A1(new_n525), .A2(new_n459), .A3(new_n506), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT29), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n462), .B1(new_n515), .B2(new_n536), .ZN(new_n537));
  NOR2_X1   g336(.A1(new_n505), .A2(new_n463), .ZN(new_n538));
  OAI21_X1  g337(.A(new_n520), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(KEYINPUT68), .ZN(new_n540));
  OAI21_X1  g339(.A(new_n534), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT30), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n541), .A2(new_n542), .A3(new_n531), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n531), .B(KEYINPUT71), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n534), .B(new_n545), .C1(new_n535), .C2(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT72), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT72), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n527), .A2(new_n548), .A3(new_n545), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n435), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(G78gat), .B(G106gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(new_n552), .B(G22gat), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(KEYINPUT31), .B(G50gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n383), .A2(new_n407), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(new_n536), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n520), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(G228gat), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n560), .A2(new_n461), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(new_n563), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n454), .A2(KEYINPUT77), .A3(new_n458), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n452), .B1(new_n457), .B2(new_n439), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT77), .ZN(new_n567));
  AOI21_X1  g366(.A(KEYINPUT29), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n569));
  AND3_X1   g368(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n569), .B1(new_n565), .B2(new_n568), .ZN(new_n571));
  INV_X1    g370(.A(new_n407), .ZN(new_n572));
  NOR3_X1   g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OAI21_X1  g372(.A(new_n564), .B1(new_n573), .B2(new_n383), .ZN(new_n574));
  INV_X1    g373(.A(new_n559), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n385), .A2(new_n386), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n459), .A2(new_n536), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT3), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n576), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n561), .B1(new_n575), .B2(new_n579), .ZN(new_n580));
  AOI21_X1  g379(.A(new_n556), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n568), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT78), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n565), .A2(new_n568), .A3(new_n569), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n407), .A3(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n383), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n563), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n577), .A2(new_n578), .ZN(new_n588));
  INV_X1    g387(.A(new_n576), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n562), .B1(new_n590), .B2(new_n559), .ZN(new_n591));
  NOR3_X1   g390(.A1(new_n587), .A2(new_n591), .A3(new_n555), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n554), .B1(new_n581), .B2(new_n592), .ZN(new_n593));
  OAI21_X1  g392(.A(new_n555), .B1(new_n587), .B2(new_n591), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n571), .A2(new_n572), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n383), .B1(new_n595), .B2(new_n584), .ZN(new_n596));
  OAI211_X1 g395(.A(new_n580), .B(new_n556), .C1(new_n596), .C2(new_n563), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n594), .A2(new_n597), .A3(new_n553), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n593), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n551), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT66), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT36), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(KEYINPUT66), .A2(KEYINPUT36), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n515), .A2(new_n406), .ZN(new_n605));
  OAI211_X1 g404(.A(new_n417), .B(new_n512), .C1(new_n514), .C2(new_n513), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(G227gat), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n608), .A2(new_n461), .ZN(new_n609));
  INV_X1    g408(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT34), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT34), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n607), .A2(new_n613), .A3(new_n610), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n605), .A2(new_n609), .A3(new_n606), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT33), .ZN(new_n616));
  AND2_X1   g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XOR2_X1   g416(.A(G15gat), .B(G43gat), .Z(new_n618));
  XNOR2_X1  g417(.A(G71gat), .B(G99gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI211_X1 g420(.A(new_n612), .B(new_n614), .C1(new_n617), .C2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(KEYINPUT32), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n621), .B1(new_n615), .B2(new_n616), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n613), .B1(new_n607), .B2(new_n610), .ZN(new_n626));
  AOI211_X1 g425(.A(KEYINPUT34), .B(new_n609), .C1(new_n605), .C2(new_n606), .ZN(new_n627));
  OAI21_X1  g426(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n622), .A2(new_n624), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n624), .B1(new_n622), .B2(new_n628), .ZN(new_n630));
  OAI211_X1 g429(.A(new_n603), .B(new_n604), .C1(new_n629), .C2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n628), .ZN(new_n632));
  NOR3_X1   g431(.A1(new_n625), .A2(new_n626), .A3(new_n627), .ZN(new_n633));
  OAI21_X1  g432(.A(new_n623), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n622), .A2(new_n624), .A3(new_n628), .ZN(new_n635));
  NAND4_X1  g434(.A1(new_n634), .A2(new_n601), .A3(new_n602), .A4(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n631), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT38), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n638), .B(new_n545), .C1(new_n527), .C2(KEYINPUT37), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n459), .B1(new_n525), .B2(new_n506), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT80), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT37), .ZN(new_n643));
  OAI21_X1  g442(.A(KEYINPUT80), .B1(new_n519), .B2(new_n520), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n640), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT81), .B1(new_n643), .B2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT37), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n647), .B1(new_n640), .B2(new_n641), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT81), .ZN(new_n649));
  OAI211_X1 g448(.A(new_n648), .B(new_n649), .C1(new_n640), .C2(new_n644), .ZN(new_n650));
  AOI21_X1  g449(.A(new_n639), .B1(new_n646), .B2(new_n650), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n531), .B1(new_n541), .B2(new_n647), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n527), .A2(KEYINPUT37), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n638), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n541), .A2(new_n531), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n433), .A2(new_n434), .A3(new_n655), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n651), .A2(new_n654), .A3(new_n656), .ZN(new_n657));
  AND3_X1   g456(.A1(new_n594), .A2(new_n553), .A3(new_n597), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n553), .B1(new_n594), .B2(new_n597), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  AOI22_X1  g459(.A1(new_n533), .A2(new_n543), .B1(new_n547), .B2(new_n549), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n409), .A2(new_n412), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT79), .B(KEYINPUT39), .Z(new_n663));
  NAND3_X1  g462(.A1(new_n662), .A2(new_n421), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(new_n429), .ZN(new_n665));
  OAI21_X1  g464(.A(KEYINPUT39), .B1(new_n420), .B2(new_n421), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n666), .B1(new_n662), .B2(new_n421), .ZN(new_n667));
  INV_X1    g466(.A(KEYINPUT40), .ZN(new_n668));
  OR3_X1    g467(.A1(new_n665), .A2(new_n667), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g468(.A(new_n668), .B1(new_n665), .B2(new_n667), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n432), .A3(new_n670), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n660), .B1(new_n661), .B2(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n600), .B(new_n637), .C1(new_n657), .C2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n435), .A2(new_n544), .A3(new_n550), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n634), .A2(new_n635), .ZN(new_n675));
  NOR3_X1   g474(.A1(new_n675), .A2(new_n658), .A3(new_n659), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT35), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n593), .A2(new_n598), .A3(new_n635), .A4(new_n634), .ZN(new_n679));
  OAI21_X1  g478(.A(KEYINPUT35), .B1(new_n551), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT82), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n673), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n673), .B2(new_n681), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n363), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT91), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT91), .ZN(new_n687));
  OAI211_X1 g486(.A(new_n687), .B(new_n363), .C1(new_n683), .C2(new_n684), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n338), .B1(new_n686), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n435), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g491(.A1(new_n544), .A2(new_n550), .ZN(new_n693));
  XOR2_X1   g492(.A(KEYINPUT16), .B(G8gat), .Z(new_n694));
  AND3_X1   g493(.A1(new_n689), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(G8gat), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n689), .B2(new_n693), .ZN(new_n697));
  OAI21_X1  g496(.A(KEYINPUT42), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  INV_X1    g498(.A(G15gat), .ZN(new_n700));
  INV_X1    g499(.A(new_n675), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n689), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n637), .ZN(new_n703));
  AND2_X1   g502(.A1(new_n689), .A2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n704), .B2(new_n700), .ZN(G1326gat));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n599), .ZN(new_n706));
  XNOR2_X1  g505(.A(KEYINPUT43), .B(G22gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1327gat));
  NAND2_X1  g507(.A1(new_n686), .A2(new_n688), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n246), .A2(new_n248), .ZN(new_n710));
  INV_X1    g509(.A(new_n710), .ZN(new_n711));
  NOR2_X1   g510(.A1(new_n711), .A2(new_n336), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g512(.A1(new_n713), .A2(new_n312), .ZN(new_n714));
  AND2_X1   g513(.A1(new_n709), .A2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n435), .A2(G29gat), .ZN(new_n717));
  AND3_X1   g516(.A1(new_n715), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n716), .B1(new_n715), .B2(new_n717), .ZN(new_n719));
  OAI211_X1 g518(.A(KEYINPUT44), .B(new_n311), .C1(new_n683), .C2(new_n684), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n312), .B1(new_n673), .B2(new_n681), .ZN(new_n721));
  OR2_X1    g520(.A1(new_n721), .A2(KEYINPUT44), .ZN(new_n722));
  AND2_X1   g521(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g522(.A(KEYINPUT90), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n359), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n354), .A2(KEYINPUT90), .A3(new_n355), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AOI22_X1  g526(.A1(new_n727), .A2(new_n353), .B1(new_n360), .B2(new_n361), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n713), .A2(new_n728), .ZN(new_n729));
  AND2_X1   g528(.A1(new_n723), .A2(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n730), .A2(new_n690), .ZN(new_n731));
  OAI22_X1  g530(.A1(new_n718), .A2(new_n719), .B1(new_n731), .B2(new_n254), .ZN(G1328gat));
  NAND3_X1  g531(.A1(new_n715), .A2(new_n252), .A3(new_n693), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(KEYINPUT46), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT46), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n715), .A2(new_n735), .A3(new_n252), .A4(new_n693), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n730), .A2(new_n693), .ZN(new_n737));
  OAI211_X1 g536(.A(new_n734), .B(new_n736), .C1(new_n252), .C2(new_n737), .ZN(G1329gat));
  NOR2_X1   g537(.A1(new_n675), .A2(G43gat), .ZN(new_n739));
  NAND3_X1  g538(.A1(new_n709), .A2(new_n714), .A3(new_n739), .ZN(new_n740));
  NAND4_X1  g539(.A1(new_n720), .A2(new_n722), .A3(new_n703), .A4(new_n729), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(G43gat), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT47), .Z(G1330gat));
  NAND3_X1  g543(.A1(new_n723), .A2(new_n599), .A3(new_n729), .ZN(new_n745));
  INV_X1    g544(.A(new_n263), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n673), .A2(new_n681), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT82), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n673), .A2(new_n681), .A3(new_n682), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n687), .B1(new_n751), .B2(new_n363), .ZN(new_n752));
  INV_X1    g551(.A(new_n688), .ZN(new_n753));
  OAI211_X1 g552(.A(KEYINPUT100), .B(new_n714), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n660), .A2(new_n746), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(KEYINPUT100), .B1(new_n709), .B2(new_n714), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n747), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT48), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  OAI211_X1 g559(.A(new_n747), .B(KEYINPUT48), .C1(new_n756), .C2(new_n757), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(G1331gat));
  NAND4_X1  g561(.A1(new_n711), .A2(new_n728), .A3(new_n312), .A4(new_n336), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n673), .B2(new_n681), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n690), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(G57gat), .ZN(G1332gat));
  AND2_X1   g565(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n693), .A2(KEYINPUT101), .ZN(new_n768));
  OR2_X1    g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n764), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(KEYINPUT102), .ZN(new_n772));
  NOR2_X1   g571(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1333gat));
  INV_X1    g573(.A(G71gat), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n764), .A2(new_n775), .A3(new_n701), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n764), .A2(new_n703), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n776), .B1(new_n777), .B2(new_n775), .ZN(new_n778));
  XOR2_X1   g577(.A(new_n778), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g578(.A1(new_n764), .A2(new_n599), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g580(.A1(new_n711), .A2(new_n363), .ZN(new_n782));
  AND2_X1   g581(.A1(new_n721), .A2(new_n782), .ZN(new_n783));
  OR2_X1    g582(.A1(new_n783), .A2(KEYINPUT51), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n721), .A2(KEYINPUT51), .A3(new_n782), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT103), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n783), .A2(KEYINPUT103), .A3(KEYINPUT51), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n784), .A2(new_n787), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n789), .A2(new_n277), .A3(new_n690), .A4(new_n336), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n711), .A2(new_n363), .A3(new_n337), .ZN(new_n791));
  AND3_X1   g590(.A1(new_n723), .A2(new_n690), .A3(new_n791), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n277), .B2(new_n792), .ZN(G1336gat));
  NAND3_X1  g592(.A1(new_n769), .A2(new_n278), .A3(new_n336), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT104), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n789), .A2(new_n795), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT105), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n720), .A2(new_n722), .A3(new_n769), .A4(new_n791), .ZN(new_n798));
  AOI21_X1  g597(.A(KEYINPUT52), .B1(new_n798), .B2(G92gat), .ZN(new_n799));
  AND3_X1   g598(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n797), .B1(new_n796), .B2(new_n799), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT52), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n723), .A2(new_n693), .A3(new_n791), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n784), .A2(new_n785), .ZN(new_n804));
  AOI22_X1  g603(.A1(new_n803), .A2(G92gat), .B1(new_n804), .B2(new_n795), .ZN(new_n805));
  OAI22_X1  g604(.A1(new_n800), .A2(new_n801), .B1(new_n802), .B2(new_n805), .ZN(G1337gat));
  NAND3_X1  g605(.A1(new_n723), .A2(new_n703), .A3(new_n791), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(G99gat), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n675), .A2(G99gat), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n789), .A2(new_n336), .A3(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT106), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT106), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n808), .A2(new_n810), .A3(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n812), .A2(new_n814), .ZN(G1338gat));
  NAND3_X1  g614(.A1(new_n723), .A2(new_n599), .A3(new_n791), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G106gat), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT53), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR3_X1   g618(.A1(new_n660), .A2(G106gat), .A3(new_n337), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT107), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n789), .A2(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n816), .A2(G106gat), .B1(new_n804), .B2(new_n821), .ZN(new_n823));
  OAI22_X1  g622(.A1(new_n819), .A2(new_n822), .B1(new_n823), .B2(new_n818), .ZN(G1339gat));
  NOR2_X1   g623(.A1(new_n338), .A2(new_n363), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n340), .B1(new_n339), .B2(new_n342), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n345), .A2(new_n346), .A3(new_n344), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n351), .B1(new_n826), .B2(new_n827), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n358), .A2(new_n828), .A3(new_n336), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AND3_X1   g629(.A1(new_n320), .A2(new_n333), .A3(new_n321), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT54), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n831), .A2(new_n334), .A3(new_n832), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n322), .A2(new_n832), .A3(new_n323), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n330), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n830), .B1(new_n833), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n320), .A2(new_n333), .A3(new_n321), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n324), .A2(KEYINPUT54), .A3(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n329), .B1(new_n334), .B2(new_n832), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n838), .A2(KEYINPUT55), .A3(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n836), .A2(new_n332), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n829), .B1(new_n841), .B2(new_n728), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n312), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n311), .A2(new_n358), .A3(new_n828), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n843), .A2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n825), .B1(new_n847), .B2(new_n710), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n848), .A2(new_n599), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n675), .A2(new_n435), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT108), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND3_X1  g652(.A1(new_n849), .A2(KEYINPUT108), .A3(new_n850), .ZN(new_n854));
  AOI21_X1  g653(.A(new_n769), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  NOR2_X1   g654(.A1(new_n855), .A2(KEYINPUT109), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT109), .ZN(new_n857));
  AOI211_X1 g656(.A(new_n857), .B(new_n769), .C1(new_n853), .C2(new_n854), .ZN(new_n858));
  OAI211_X1 g657(.A(new_n394), .B(new_n363), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n769), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n849), .A2(new_n860), .A3(new_n850), .ZN(new_n861));
  OAI21_X1  g660(.A(G113gat), .B1(new_n861), .B2(new_n728), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n859), .A2(new_n862), .ZN(G1340gat));
  OAI211_X1 g662(.A(new_n395), .B(new_n336), .C1(new_n856), .C2(new_n858), .ZN(new_n864));
  OAI21_X1  g663(.A(G120gat), .B1(new_n861), .B2(new_n337), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n864), .A2(new_n865), .ZN(G1341gat));
  NAND3_X1  g665(.A1(new_n855), .A2(new_n389), .A3(new_n711), .ZN(new_n867));
  OAI21_X1  g666(.A(G127gat), .B1(new_n861), .B2(new_n710), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1342gat));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n661), .A2(new_n311), .ZN(new_n871));
  XNOR2_X1  g670(.A(new_n871), .B(KEYINPUT110), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n872), .A2(G134gat), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n870), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g673(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n875));
  OAI21_X1  g674(.A(G134gat), .B1(new_n861), .B2(new_n312), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n874), .A2(KEYINPUT56), .ZN(new_n877));
  NAND3_X1  g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1343gat));
  NAND4_X1  g677(.A1(new_n363), .A2(new_n332), .A3(new_n840), .A4(new_n836), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n311), .B1(new_n879), .B2(new_n829), .ZN(new_n880));
  OAI21_X1  g679(.A(new_n710), .B1(new_n880), .B2(new_n845), .ZN(new_n881));
  INV_X1    g680(.A(new_n825), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n660), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  XNOR2_X1  g682(.A(KEYINPUT111), .B(KEYINPUT57), .ZN(new_n884));
  INV_X1    g683(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(KEYINPUT112), .B1(new_n883), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT112), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n887), .B(new_n884), .C1(new_n848), .C2(new_n660), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n829), .A2(KEYINPUT113), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT113), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n358), .A2(new_n828), .A3(new_n890), .A4(new_n336), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n879), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n845), .B1(new_n892), .B2(new_n312), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n882), .B1(new_n893), .B2(new_n711), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n894), .A2(KEYINPUT57), .A3(new_n599), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n886), .A2(new_n888), .A3(new_n895), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n637), .A2(new_n690), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n769), .A2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n896), .A2(new_n363), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n899), .A2(G141gat), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT114), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n883), .A2(new_n898), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n902), .A2(new_n364), .A3(new_n363), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n900), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n901), .A2(new_n904), .A3(KEYINPUT58), .ZN(new_n905));
  INV_X1    g704(.A(KEYINPUT58), .ZN(new_n906));
  OAI211_X1 g705(.A(new_n900), .B(new_n903), .C1(KEYINPUT114), .C2(new_n906), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n905), .A2(new_n907), .ZN(G1344gat));
  INV_X1    g707(.A(KEYINPUT115), .ZN(new_n909));
  NOR3_X1   g708(.A1(new_n769), .A2(new_n337), .A3(new_n897), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n883), .A2(new_n366), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n896), .A2(new_n336), .A3(new_n898), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n366), .A2(KEYINPUT59), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g713(.A(KEYINPUT57), .B1(new_n894), .B2(new_n599), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n660), .B(new_n884), .C1(new_n881), .C2(new_n882), .ZN(new_n916));
  OAI21_X1  g715(.A(new_n910), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n917), .A2(G148gat), .ZN(new_n918));
  AND2_X1   g717(.A1(new_n918), .A2(KEYINPUT59), .ZN(new_n919));
  OAI211_X1 g718(.A(new_n909), .B(new_n911), .C1(new_n914), .C2(new_n919), .ZN(new_n920));
  AOI22_X1  g719(.A1(new_n912), .A2(new_n913), .B1(new_n918), .B2(KEYINPUT59), .ZN(new_n921));
  INV_X1    g720(.A(new_n911), .ZN(new_n922));
  OAI21_X1  g721(.A(KEYINPUT115), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n920), .A2(new_n923), .ZN(G1345gat));
  AOI21_X1  g723(.A(G155gat), .B1(new_n902), .B2(new_n711), .ZN(new_n925));
  AND2_X1   g724(.A1(new_n896), .A2(new_n898), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n710), .A2(new_n373), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n925), .B1(new_n926), .B2(new_n927), .ZN(G1346gat));
  NAND3_X1  g727(.A1(new_n896), .A2(new_n311), .A3(new_n898), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G162gat), .ZN(new_n930));
  NOR4_X1   g729(.A1(new_n872), .A2(G162gat), .A3(new_n435), .A4(new_n703), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n883), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT116), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n930), .A2(KEYINPUT116), .A3(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1347gat));
  NAND2_X1  g736(.A1(new_n693), .A2(new_n435), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT117), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n938), .B(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n940), .A2(new_n701), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n849), .A2(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n942), .A2(new_n466), .A3(new_n728), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n848), .A2(new_n690), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n860), .A2(new_n679), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  INV_X1    g745(.A(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(new_n363), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n943), .B1(new_n466), .B2(new_n948), .ZN(G1348gat));
  OAI21_X1  g748(.A(new_n467), .B1(new_n946), .B2(new_n337), .ZN(new_n950));
  XNOR2_X1  g749(.A(new_n950), .B(KEYINPUT118), .ZN(new_n951));
  NOR3_X1   g750(.A1(new_n942), .A2(new_n467), .A3(new_n337), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(G1349gat));
  NAND3_X1  g752(.A1(new_n947), .A2(new_n502), .A3(new_n711), .ZN(new_n954));
  OAI21_X1  g753(.A(G183gat), .B1(new_n942), .B2(new_n710), .ZN(new_n955));
  NAND3_X1  g754(.A1(new_n954), .A2(KEYINPUT119), .A3(new_n955), .ZN(new_n956));
  XNOR2_X1  g755(.A(new_n956), .B(KEYINPUT60), .ZN(G1350gat));
  NOR3_X1   g756(.A1(new_n946), .A2(G190gat), .A3(new_n312), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n849), .A2(new_n311), .A3(new_n941), .ZN(new_n959));
  AND2_X1   g758(.A1(new_n959), .A2(G190gat), .ZN(new_n960));
  NOR2_X1   g759(.A1(new_n960), .A2(KEYINPUT120), .ZN(new_n961));
  INV_X1    g760(.A(KEYINPUT61), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n958), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g762(.A1(new_n960), .A2(KEYINPUT120), .ZN(new_n964));
  OAI21_X1  g763(.A(KEYINPUT61), .B1(new_n960), .B2(KEYINPUT120), .ZN(new_n965));
  OAI21_X1  g764(.A(new_n963), .B1(new_n964), .B2(new_n965), .ZN(G1351gat));
  NAND2_X1  g765(.A1(new_n940), .A2(new_n637), .ZN(new_n967));
  INV_X1    g766(.A(KEYINPUT122), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n967), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n940), .A2(KEYINPUT122), .A3(new_n637), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n969), .A2(KEYINPUT123), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT123), .B1(new_n969), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n894), .A2(new_n599), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT57), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(new_n916), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n973), .A2(new_n978), .ZN(new_n979));
  OAI21_X1  g778(.A(G197gat), .B1(new_n979), .B2(new_n728), .ZN(new_n980));
  NOR3_X1   g779(.A1(new_n860), .A2(new_n660), .A3(new_n703), .ZN(new_n981));
  NAND4_X1  g780(.A1(new_n944), .A2(new_n445), .A3(new_n363), .A4(new_n981), .ZN(new_n982));
  XNOR2_X1  g781(.A(new_n982), .B(KEYINPUT121), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT124), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g785(.A1(new_n980), .A2(KEYINPUT124), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1352gat));
  NAND2_X1  g787(.A1(new_n944), .A2(new_n981), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n989), .A2(G204gat), .A3(new_n337), .ZN(new_n990));
  XNOR2_X1  g789(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  OAI21_X1  g791(.A(G204gat), .B1(new_n979), .B2(new_n337), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(G1353gat));
  NAND4_X1  g793(.A1(new_n944), .A2(new_n437), .A3(new_n711), .A4(new_n981), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n710), .B1(new_n969), .B2(new_n970), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n996), .B1(new_n915), .B2(new_n916), .ZN(new_n997));
  AND3_X1   g796(.A1(new_n997), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n998));
  AOI21_X1  g797(.A(KEYINPUT63), .B1(new_n997), .B2(G211gat), .ZN(new_n999));
  OAI21_X1  g798(.A(new_n995), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g799(.A(KEYINPUT126), .ZN(new_n1001));
  NAND2_X1  g800(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  OAI211_X1 g801(.A(KEYINPUT126), .B(new_n995), .C1(new_n998), .C2(new_n999), .ZN(new_n1003));
  NAND2_X1  g802(.A1(new_n1002), .A2(new_n1003), .ZN(G1354gat));
  NOR3_X1   g803(.A1(new_n989), .A2(G218gat), .A3(new_n312), .ZN(new_n1005));
  NAND3_X1  g804(.A1(new_n973), .A2(new_n978), .A3(new_n311), .ZN(new_n1006));
  AOI21_X1  g805(.A(new_n1005), .B1(new_n1006), .B2(G218gat), .ZN(new_n1007));
  XNOR2_X1  g806(.A(new_n1007), .B(KEYINPUT127), .ZN(G1355gat));
endmodule


