//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 1 1 1 0 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n724, new_n725, new_n726, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037;
  INV_X1    g000(.A(G217), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AOI21_X1  g002(.A(new_n187), .B1(G234), .B2(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G119), .ZN(new_n191));
  INV_X1    g005(.A(G119), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n191), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  XNOR2_X1  g009(.A(KEYINPUT24), .B(G110), .ZN(new_n196));
  INV_X1    g010(.A(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT70), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT23), .ZN(new_n200));
  OAI21_X1  g014(.A(new_n200), .B1(new_n192), .B2(G128), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n201), .A2(new_n193), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT69), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT69), .A4(new_n193), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  AOI21_X1  g021(.A(new_n199), .B1(new_n207), .B2(G110), .ZN(new_n208));
  INV_X1    g022(.A(G110), .ZN(new_n209));
  AOI211_X1 g023(.A(KEYINPUT70), .B(new_n209), .C1(new_n205), .C2(new_n206), .ZN(new_n210));
  OAI21_X1  g024(.A(new_n198), .B1(new_n208), .B2(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(G140), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G125), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n213), .A2(KEYINPUT16), .ZN(new_n214));
  INV_X1    g028(.A(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G125), .ZN(new_n216));
  NOR3_X1   g030(.A1(new_n216), .A2(KEYINPUT71), .A3(G140), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n216), .A2(G140), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n213), .A2(new_n219), .A3(KEYINPUT71), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  AOI21_X1  g035(.A(KEYINPUT72), .B1(new_n221), .B2(KEYINPUT16), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT72), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT16), .ZN(new_n224));
  AOI211_X1 g038(.A(new_n223), .B(new_n224), .C1(new_n218), .C2(new_n220), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n215), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(G146), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  XNOR2_X1  g042(.A(G125), .B(G140), .ZN(new_n229));
  AOI21_X1  g043(.A(new_n217), .B1(new_n229), .B2(KEYINPUT71), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n223), .B1(new_n230), .B2(new_n224), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n221), .A2(KEYINPUT72), .A3(KEYINPUT16), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n214), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(G146), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n211), .B1(new_n228), .B2(new_n234), .ZN(new_n235));
  AOI211_X1 g049(.A(new_n227), .B(new_n214), .C1(new_n231), .C2(new_n232), .ZN(new_n236));
  OAI22_X1  g050(.A1(new_n195), .A2(new_n197), .B1(new_n203), .B2(G110), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n229), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n236), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g054(.A(KEYINPUT22), .B(G137), .ZN(new_n241));
  INV_X1    g055(.A(G953), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(G221), .A3(G234), .ZN(new_n243));
  XNOR2_X1  g057(.A(new_n241), .B(new_n243), .ZN(new_n244));
  NOR3_X1   g058(.A1(new_n235), .A2(new_n240), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(new_n244), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n209), .B1(new_n205), .B2(new_n206), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n247), .B(new_n199), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n233), .A2(G146), .ZN(new_n249));
  OAI211_X1 g063(.A(new_n248), .B(new_n198), .C1(new_n249), .C2(new_n236), .ZN(new_n250));
  INV_X1    g064(.A(new_n240), .ZN(new_n251));
  AOI21_X1  g065(.A(new_n246), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n188), .B1(new_n245), .B2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(KEYINPUT73), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT25), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  OAI211_X1 g070(.A(KEYINPUT25), .B(new_n188), .C1(new_n245), .C2(new_n252), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n257), .A2(KEYINPUT73), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n244), .B1(new_n235), .B2(new_n240), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n250), .A2(new_n251), .A3(new_n246), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(KEYINPUT25), .B1(new_n261), .B2(new_n188), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n189), .B(new_n256), .C1(new_n258), .C2(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n189), .A2(G902), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(G472), .A2(G902), .ZN(new_n267));
  XOR2_X1   g081(.A(G116), .B(G119), .Z(new_n268));
  XNOR2_X1  g082(.A(KEYINPUT2), .B(G113), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT65), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  XOR2_X1   g084(.A(KEYINPUT2), .B(G113), .Z(new_n271));
  INV_X1    g085(.A(KEYINPUT65), .ZN(new_n272));
  XNOR2_X1  g086(.A(G116), .B(G119), .ZN(new_n273));
  NAND3_X1  g087(.A1(new_n271), .A2(new_n272), .A3(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n270), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n268), .A2(new_n269), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT11), .ZN(new_n278));
  INV_X1    g092(.A(G134), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n278), .B1(new_n279), .B2(G137), .ZN(new_n280));
  INV_X1    g094(.A(G137), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT11), .A3(G134), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(G137), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(G131), .ZN(new_n285));
  INV_X1    g099(.A(G131), .ZN(new_n286));
  NAND4_X1  g100(.A1(new_n280), .A2(new_n282), .A3(new_n286), .A4(new_n283), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n285), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n227), .A2(G143), .ZN(new_n289));
  INV_X1    g103(.A(G143), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G146), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  NOR2_X1   g106(.A1(KEYINPUT0), .A2(G128), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT0), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n294), .A2(new_n190), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n292), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  XNOR2_X1  g110(.A(G143), .B(G146), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n297), .B1(new_n294), .B2(new_n190), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(G128), .B1(new_n289), .B2(new_n291), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n290), .A2(KEYINPUT1), .A3(G146), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  OAI21_X1  g116(.A(KEYINPUT64), .B1(new_n300), .B2(new_n302), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT64), .ZN(new_n304));
  OAI211_X1 g118(.A(new_n304), .B(new_n301), .C1(new_n297), .C2(G128), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT1), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n297), .A2(new_n306), .A3(G128), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n283), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n279), .A2(G137), .ZN(new_n310));
  OAI21_X1  g124(.A(G131), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(new_n287), .ZN(new_n312));
  INV_X1    g126(.A(new_n312), .ZN(new_n313));
  AOI221_X4 g127(.A(KEYINPUT30), .B1(new_n288), .B2(new_n299), .C1(new_n308), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n308), .A2(new_n313), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n288), .A2(new_n299), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n315), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  OAI21_X1  g132(.A(new_n277), .B1(new_n314), .B2(new_n318), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT31), .ZN(new_n320));
  XNOR2_X1  g134(.A(KEYINPUT26), .B(G101), .ZN(new_n321));
  NOR2_X1   g135(.A1(G237), .A2(G953), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n322), .A2(G210), .ZN(new_n323));
  XNOR2_X1  g137(.A(new_n321), .B(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(KEYINPUT66), .B(KEYINPUT27), .ZN(new_n325));
  XOR2_X1   g139(.A(new_n324), .B(new_n325), .Z(new_n326));
  AOI22_X1  g140(.A1(new_n270), .A2(new_n274), .B1(new_n268), .B2(new_n269), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n316), .A2(new_n327), .A3(new_n317), .ZN(new_n328));
  NAND4_X1  g142(.A1(new_n319), .A2(new_n320), .A3(new_n326), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT67), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n319), .A2(new_n326), .A3(new_n328), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(KEYINPUT31), .ZN(new_n332));
  AND2_X1   g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n326), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT28), .ZN(new_n335));
  AND4_X1   g149(.A1(new_n306), .A2(new_n289), .A3(new_n291), .A4(G128), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n301), .B1(new_n297), .B2(G128), .ZN(new_n337));
  AOI21_X1  g151(.A(new_n336), .B1(new_n337), .B2(KEYINPUT64), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n312), .B1(new_n338), .B2(new_n305), .ZN(new_n339));
  AND2_X1   g153(.A1(new_n288), .A2(new_n299), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n277), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n335), .B1(new_n341), .B2(new_n328), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n328), .A2(new_n335), .ZN(new_n343));
  INV_X1    g157(.A(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n334), .B1(new_n342), .B2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT67), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n345), .B1(new_n332), .B2(new_n346), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n267), .B1(new_n333), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n348), .A2(KEYINPUT32), .ZN(new_n349));
  INV_X1    g163(.A(new_n328), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n327), .B1(new_n316), .B2(new_n317), .ZN(new_n351));
  OAI21_X1  g165(.A(KEYINPUT28), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n326), .B1(new_n352), .B2(new_n343), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT30), .B1(new_n339), .B2(new_n340), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n316), .A2(new_n315), .A3(new_n317), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n350), .B1(new_n356), .B2(new_n277), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n320), .B1(new_n357), .B2(new_n326), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n353), .B1(new_n358), .B2(KEYINPUT67), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n330), .A2(new_n332), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT32), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n361), .A2(new_n362), .A3(new_n267), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n349), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G472), .ZN(new_n365));
  NOR3_X1   g179(.A1(new_n342), .A2(new_n344), .A3(new_n334), .ZN(new_n366));
  AOI21_X1  g180(.A(G902), .B1(new_n366), .B2(KEYINPUT29), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n352), .A2(new_n326), .A3(new_n343), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n327), .B1(new_n354), .B2(new_n355), .ZN(new_n369));
  OAI21_X1  g183(.A(new_n334), .B1(new_n369), .B2(new_n350), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT29), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n368), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n365), .B1(new_n367), .B2(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(KEYINPUT68), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n266), .B1(new_n364), .B2(new_n374), .ZN(new_n375));
  XNOR2_X1  g189(.A(KEYINPUT9), .B(G234), .ZN(new_n376));
  OAI21_X1  g190(.A(G221), .B1(new_n376), .B2(G902), .ZN(new_n377));
  XOR2_X1   g191(.A(new_n377), .B(KEYINPUT74), .Z(new_n378));
  XNOR2_X1  g192(.A(G110), .B(G140), .ZN(new_n379));
  AND2_X1   g193(.A1(new_n242), .A2(G227), .ZN(new_n380));
  XNOR2_X1  g194(.A(new_n379), .B(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G104), .ZN(new_n383));
  OAI21_X1  g197(.A(KEYINPUT3), .B1(new_n383), .B2(G107), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT3), .ZN(new_n385));
  INV_X1    g199(.A(G107), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n385), .A2(new_n386), .A3(G104), .ZN(new_n387));
  INV_X1    g201(.A(G101), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(G107), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n384), .A2(new_n387), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n383), .A2(G107), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n386), .A2(G104), .ZN(new_n392));
  OAI21_X1  g206(.A(G101), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT10), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n308), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n384), .A2(new_n387), .A3(new_n389), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(G101), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n399), .A2(KEYINPUT4), .A3(new_n390), .ZN(new_n400));
  XOR2_X1   g214(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n401));
  NAND3_X1  g215(.A1(new_n398), .A2(G101), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n299), .A3(new_n402), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n390), .B(new_n393), .C1(new_n337), .C2(new_n336), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(new_n395), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n397), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n288), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT78), .ZN(new_n408));
  INV_X1    g222(.A(new_n288), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n397), .A2(new_n403), .A3(new_n405), .A4(new_n409), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(KEYINPUT78), .A3(new_n288), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n382), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND4_X1  g227(.A1(new_n303), .A2(new_n394), .A3(new_n305), .A4(new_n307), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(new_n404), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(new_n288), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT77), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT12), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n416), .A2(new_n417), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n409), .B1(new_n414), .B2(new_n404), .ZN(new_n420));
  OAI21_X1  g234(.A(KEYINPUT77), .B1(new_n420), .B2(KEYINPUT12), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(KEYINPUT12), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n423), .A2(new_n410), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n413), .B1(new_n424), .B2(new_n382), .ZN(new_n425));
  INV_X1    g239(.A(G469), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n425), .A2(KEYINPUT79), .A3(new_n426), .A4(new_n188), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n382), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n411), .A2(new_n412), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n381), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n428), .A2(new_n430), .A3(new_n426), .A4(new_n188), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT79), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n427), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n429), .A2(new_n382), .ZN(new_n435));
  INV_X1    g249(.A(new_n424), .ZN(new_n436));
  XOR2_X1   g250(.A(new_n381), .B(KEYINPUT75), .Z(new_n437));
  OAI21_X1  g251(.A(new_n435), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n188), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G469), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n378), .B1(new_n434), .B2(new_n440), .ZN(new_n441));
  AND3_X1   g255(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n442));
  AOI21_X1  g256(.A(G143), .B1(new_n322), .B2(G214), .ZN(new_n443));
  OAI21_X1  g257(.A(G131), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n322), .A2(G214), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(new_n290), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n322), .A2(G143), .A3(G214), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n446), .A2(new_n286), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n444), .A2(new_n448), .ZN(new_n449));
  MUX2_X1   g263(.A(new_n449), .B(new_n444), .S(KEYINPUT17), .Z(new_n450));
  NAND3_X1  g264(.A1(new_n228), .A2(new_n234), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G113), .B(G122), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n383), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n238), .B1(new_n221), .B2(new_n227), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT18), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n446), .B(new_n447), .C1(new_n455), .C2(new_n286), .ZN(new_n456));
  OAI211_X1 g270(.A(new_n454), .B(new_n456), .C1(new_n455), .C2(new_n444), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n451), .A2(new_n453), .A3(new_n457), .ZN(new_n458));
  MUX2_X1   g272(.A(new_n229), .B(new_n230), .S(KEYINPUT19), .Z(new_n459));
  OAI21_X1  g273(.A(new_n449), .B1(new_n459), .B2(G146), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n460), .B2(new_n236), .ZN(new_n461));
  INV_X1    g275(.A(new_n453), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n458), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g278(.A1(G475), .A2(G902), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT20), .ZN(new_n467));
  INV_X1    g281(.A(new_n465), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n468), .B1(new_n458), .B2(new_n463), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT20), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  INV_X1    g285(.A(new_n458), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n453), .B1(new_n451), .B2(new_n457), .ZN(new_n473));
  OAI21_X1  g287(.A(new_n188), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n467), .A2(new_n471), .B1(G475), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n290), .A2(KEYINPUT13), .A3(G128), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT13), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n477), .B1(new_n190), .B2(G143), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n190), .A2(G143), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n476), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(G134), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n290), .A2(G128), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n190), .A2(G143), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n279), .ZN(new_n484));
  INV_X1    g298(.A(G116), .ZN(new_n485));
  NOR2_X1   g299(.A1(new_n485), .A2(G122), .ZN(new_n486));
  INV_X1    g300(.A(G122), .ZN(new_n487));
  NOR2_X1   g301(.A1(new_n487), .A2(G116), .ZN(new_n488));
  OAI21_X1  g302(.A(G107), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n487), .A2(G116), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n485), .A2(G122), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n386), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  NAND3_X1  g307(.A1(new_n481), .A2(new_n484), .A3(new_n493), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT14), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n495), .A2(new_n485), .A3(G122), .ZN(new_n496));
  AOI21_X1  g310(.A(KEYINPUT14), .B1(new_n487), .B2(G116), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n488), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n498), .A2(G107), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n290), .A2(G128), .ZN(new_n500));
  OAI21_X1  g314(.A(G134), .B1(new_n479), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n484), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n502), .A3(new_n492), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n494), .A2(new_n503), .ZN(new_n504));
  NOR3_X1   g318(.A1(new_n376), .A2(new_n187), .A3(G953), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n505), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n494), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  AND2_X1   g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT15), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(G478), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n188), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n506), .A2(new_n188), .A3(new_n508), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n513), .A2(new_n510), .A3(G478), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(G234), .A2(G237), .ZN(new_n517));
  AND3_X1   g331(.A1(new_n517), .A2(G952), .A3(new_n242), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n517), .A2(G902), .A3(G953), .ZN(new_n519));
  XOR2_X1   g333(.A(new_n519), .B(KEYINPUT84), .Z(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(KEYINPUT21), .B(G898), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n518), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n475), .A2(new_n516), .A3(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n277), .A2(new_n400), .A3(new_n402), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n485), .A2(KEYINPUT5), .A3(G119), .ZN(new_n527));
  INV_X1    g341(.A(G113), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n273), .A2(KEYINPUT5), .ZN(new_n530));
  AOI22_X1  g344(.A1(new_n270), .A2(new_n274), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(new_n394), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n526), .A2(new_n533), .ZN(new_n534));
  XNOR2_X1  g348(.A(G110), .B(G122), .ZN(new_n535));
  INV_X1    g349(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n526), .A2(new_n533), .A3(new_n535), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n537), .A2(KEYINPUT6), .A3(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(new_n216), .B1(new_n296), .B2(new_n298), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n540), .B1(new_n308), .B2(new_n216), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n242), .A2(G224), .ZN(new_n542));
  XNOR2_X1  g356(.A(new_n542), .B(KEYINPUT81), .ZN(new_n543));
  XNOR2_X1  g357(.A(new_n541), .B(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT6), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n534), .A2(new_n545), .A3(new_n536), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n539), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT7), .ZN(new_n548));
  NOR2_X1   g362(.A1(new_n543), .A2(new_n548), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  OR2_X1    g364(.A1(new_n541), .A2(new_n550), .ZN(new_n551));
  AND2_X1   g365(.A1(new_n551), .A2(new_n538), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT83), .ZN(new_n553));
  OAI21_X1  g367(.A(new_n529), .B1(new_n530), .B2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n553), .B2(new_n530), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n275), .A2(new_n532), .ZN(new_n556));
  OAI22_X1  g370(.A1(new_n555), .A2(new_n556), .B1(new_n532), .B2(new_n531), .ZN(new_n557));
  XNOR2_X1  g371(.A(KEYINPUT82), .B(KEYINPUT8), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n535), .B(new_n558), .ZN(new_n559));
  AOI22_X1  g373(.A1(new_n557), .A2(new_n559), .B1(new_n541), .B2(new_n550), .ZN(new_n560));
  AOI21_X1  g374(.A(G902), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  OAI21_X1  g375(.A(G210), .B1(G237), .B2(G902), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n547), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(new_n562), .B1(new_n547), .B2(new_n561), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(G214), .B1(G237), .B2(G902), .ZN(new_n567));
  XNOR2_X1  g381(.A(new_n567), .B(KEYINPUT80), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n525), .A2(new_n566), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n375), .A2(new_n441), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g384(.A(new_n570), .B(G101), .ZN(G3));
  NAND2_X1  g385(.A1(new_n361), .A2(new_n188), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(KEYINPUT85), .A3(G472), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT85), .ZN(new_n574));
  AOI21_X1  g388(.A(G902), .B1(new_n359), .B2(new_n360), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n574), .B1(new_n575), .B2(new_n365), .ZN(new_n576));
  AOI22_X1  g390(.A1(new_n573), .A2(new_n576), .B1(new_n267), .B2(new_n361), .ZN(new_n577));
  INV_X1    g391(.A(new_n266), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n577), .A2(new_n578), .A3(new_n441), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT33), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT86), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n504), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n581), .B1(new_n583), .B2(new_n505), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT87), .ZN(new_n585));
  AOI211_X1 g399(.A(KEYINPUT86), .B(new_n505), .C1(new_n494), .C2(new_n503), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g402(.A(KEYINPUT86), .B1(new_n494), .B2(new_n503), .ZN(new_n589));
  OAI21_X1  g403(.A(KEYINPUT33), .B1(new_n589), .B2(new_n507), .ZN(new_n590));
  OAI21_X1  g404(.A(KEYINPUT87), .B1(new_n590), .B2(new_n586), .ZN(new_n591));
  AOI22_X1  g405(.A1(new_n588), .A2(new_n591), .B1(new_n581), .B2(new_n509), .ZN(new_n592));
  AOI21_X1  g406(.A(new_n580), .B1(new_n592), .B2(new_n188), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n513), .A2(G478), .ZN(new_n594));
  OAI21_X1  g408(.A(KEYINPUT88), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n509), .A2(new_n581), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n597));
  NOR3_X1   g411(.A1(new_n590), .A2(KEYINPUT87), .A3(new_n586), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n188), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G478), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT88), .ZN(new_n601));
  INV_X1    g415(.A(new_n594), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n474), .A2(G475), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n466), .A2(KEYINPUT20), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n469), .A2(new_n470), .ZN(new_n607));
  OAI21_X1  g421(.A(new_n605), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n567), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n547), .A2(new_n561), .ZN(new_n611));
  INV_X1    g425(.A(new_n562), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n610), .B1(new_n613), .B2(new_n563), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n524), .ZN(new_n615));
  NOR3_X1   g429(.A1(new_n579), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(KEYINPUT34), .B(G104), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n616), .B(new_n617), .ZN(G6));
  INV_X1    g432(.A(KEYINPUT89), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n467), .A2(new_n619), .A3(new_n471), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n469), .A2(KEYINPUT89), .A3(new_n470), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT90), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n451), .A2(new_n457), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n462), .ZN(new_n625));
  AOI21_X1  g439(.A(G902), .B1(new_n625), .B2(new_n458), .ZN(new_n626));
  INV_X1    g440(.A(G475), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n623), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n474), .A2(KEYINPUT90), .A3(G475), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n629), .A3(new_n515), .ZN(new_n630));
  NOR3_X1   g444(.A1(new_n615), .A2(new_n622), .A3(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n579), .A2(new_n632), .ZN(new_n633));
  XNOR2_X1  g447(.A(KEYINPUT35), .B(G107), .ZN(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G9));
  AND2_X1   g449(.A1(new_n569), .A2(new_n441), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n235), .A2(new_n240), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n246), .A2(KEYINPUT36), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n637), .B(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(new_n264), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n263), .A2(new_n642), .ZN(new_n643));
  AND3_X1   g457(.A1(new_n577), .A2(KEYINPUT91), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g458(.A(KEYINPUT91), .B1(new_n577), .B2(new_n643), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n636), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(KEYINPUT37), .B(G110), .Z(new_n647));
  XNOR2_X1  g461(.A(new_n646), .B(new_n647), .ZN(G12));
  AOI21_X1  g462(.A(new_n362), .B1(new_n361), .B2(new_n267), .ZN(new_n649));
  INV_X1    g463(.A(new_n267), .ZN(new_n650));
  AOI211_X1 g464(.A(KEYINPUT32), .B(new_n650), .C1(new_n359), .C2(new_n360), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n367), .A2(new_n372), .ZN(new_n652));
  AOI21_X1  g466(.A(KEYINPUT68), .B1(new_n652), .B2(G472), .ZN(new_n653));
  INV_X1    g467(.A(KEYINPUT68), .ZN(new_n654));
  AOI211_X1 g468(.A(new_n654), .B(new_n365), .C1(new_n367), .C2(new_n372), .ZN(new_n655));
  OAI22_X1  g469(.A1(new_n649), .A2(new_n651), .B1(new_n653), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n567), .B1(new_n564), .B2(new_n565), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n657), .B1(new_n263), .B2(new_n642), .ZN(new_n658));
  OR2_X1    g472(.A1(new_n520), .A2(G900), .ZN(new_n659));
  INV_X1    g473(.A(new_n518), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n661), .ZN(new_n662));
  NOR3_X1   g476(.A1(new_n622), .A2(new_n630), .A3(new_n662), .ZN(new_n663));
  NAND4_X1  g477(.A1(new_n656), .A2(new_n441), .A3(new_n658), .A4(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XNOR2_X1  g479(.A(new_n661), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n441), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g481(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n667), .A2(KEYINPUT40), .ZN(new_n669));
  OAI21_X1  g483(.A(new_n334), .B1(new_n350), .B2(new_n351), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n331), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n365), .B1(new_n671), .B2(new_n188), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n672), .B1(new_n349), .B2(new_n363), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  OAI21_X1  g488(.A(KEYINPUT38), .B1(new_n564), .B2(new_n565), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT38), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n613), .A2(new_n676), .A3(new_n563), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n675), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n608), .A2(new_n567), .A3(new_n515), .ZN(new_n680));
  NOR3_X1   g494(.A1(new_n679), .A2(new_n643), .A3(new_n680), .ZN(new_n681));
  NAND4_X1  g495(.A1(new_n668), .A2(new_n669), .A3(new_n674), .A4(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G143), .ZN(G45));
  AOI21_X1  g497(.A(new_n601), .B1(new_n600), .B2(new_n602), .ZN(new_n684));
  AOI211_X1 g498(.A(KEYINPUT88), .B(new_n594), .C1(new_n599), .C2(G478), .ZN(new_n685));
  OAI211_X1 g499(.A(new_n608), .B(new_n661), .C1(new_n684), .C2(new_n685), .ZN(new_n686));
  INV_X1    g500(.A(KEYINPUT92), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n604), .A2(KEYINPUT92), .A3(new_n608), .A4(new_n661), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n688), .A2(new_n658), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n656), .A2(new_n441), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(new_n227), .ZN(G48));
  NOR2_X1   g507(.A1(new_n609), .A2(new_n615), .ZN(new_n694));
  INV_X1    g508(.A(new_n378), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n425), .A2(new_n188), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n434), .A2(new_n695), .A3(new_n697), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n375), .A2(new_n694), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(KEYINPUT93), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT41), .B(G113), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G15));
  NAND3_X1  g516(.A1(new_n375), .A2(new_n631), .A3(new_n698), .ZN(new_n703));
  XNOR2_X1  g517(.A(new_n703), .B(G116), .ZN(G18));
  AND4_X1   g518(.A1(new_n695), .A2(new_n434), .A3(new_n614), .A4(new_n697), .ZN(new_n705));
  INV_X1    g519(.A(new_n189), .ZN(new_n706));
  AOI21_X1  g520(.A(new_n706), .B1(new_n262), .B2(new_n254), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n253), .A2(new_n255), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(KEYINPUT73), .A3(new_n257), .ZN(new_n709));
  AOI21_X1  g523(.A(new_n641), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  NOR2_X1   g524(.A1(new_n710), .A2(new_n525), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n705), .A2(new_n711), .A3(new_n656), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G119), .ZN(G21));
  NAND3_X1  g527(.A1(new_n332), .A2(new_n329), .A3(new_n345), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n267), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n715), .B1(new_n575), .B2(new_n365), .ZN(new_n716));
  NOR2_X1   g530(.A1(new_n266), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT94), .B1(new_n475), .B2(new_n516), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT94), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n608), .A2(new_n719), .A3(new_n515), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n657), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n717), .A2(new_n721), .A3(new_n698), .A4(new_n524), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G122), .ZN(G24));
  NOR2_X1   g537(.A1(new_n710), .A2(new_n716), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n705), .A2(new_n724), .A3(new_n688), .A4(new_n689), .ZN(new_n725));
  XNOR2_X1  g539(.A(KEYINPUT95), .B(G125), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n725), .B(new_n726), .ZN(G27));
  NAND4_X1  g541(.A1(new_n613), .A2(new_n695), .A3(new_n563), .A4(new_n567), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n426), .A2(new_n188), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT96), .B1(new_n429), .B2(new_n382), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT96), .ZN(new_n731));
  AOI211_X1 g545(.A(new_n731), .B(new_n381), .C1(new_n411), .C2(new_n412), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n437), .B1(new_n423), .B2(new_n410), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n730), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  AOI21_X1  g548(.A(new_n729), .B1(new_n734), .B2(G469), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n728), .B1(new_n735), .B2(new_n434), .ZN(new_n736));
  AND3_X1   g550(.A1(new_n656), .A2(new_n578), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g551(.A1(new_n688), .A2(new_n689), .ZN(new_n738));
  INV_X1    g552(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g553(.A(KEYINPUT42), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n653), .A2(new_n655), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT97), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n741), .B1(new_n364), .B2(new_n742), .ZN(new_n743));
  NAND3_X1  g557(.A1(new_n349), .A2(KEYINPUT97), .A3(new_n363), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n266), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n688), .A2(new_n736), .A3(KEYINPUT42), .A4(new_n689), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(KEYINPUT98), .A3(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT98), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n742), .B1(new_n649), .B2(new_n651), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n750), .A2(new_n744), .A3(new_n374), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n578), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n749), .B1(new_n752), .B2(new_n746), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n740), .B1(new_n748), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(new_n286), .ZN(G33));
  NAND4_X1  g569(.A1(new_n656), .A2(new_n736), .A3(new_n578), .A4(new_n663), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  INV_X1    g571(.A(KEYINPUT100), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n577), .A2(new_n758), .A3(new_n710), .ZN(new_n759));
  OAI21_X1  g573(.A(new_n758), .B1(new_n577), .B2(new_n710), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n604), .A2(new_n475), .ZN(new_n761));
  AOI21_X1  g575(.A(KEYINPUT43), .B1(new_n475), .B2(KEYINPUT99), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n604), .B(new_n475), .C1(KEYINPUT99), .C2(KEYINPUT43), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n759), .A2(new_n760), .A3(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT44), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND4_X1  g582(.A1(new_n759), .A2(KEYINPUT44), .A3(new_n760), .A4(new_n765), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n734), .A2(KEYINPUT45), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT45), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n426), .B1(new_n438), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n770), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n729), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(KEYINPUT46), .A3(new_n774), .ZN(new_n775));
  NAND2_X1  g589(.A1(new_n775), .A2(new_n434), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n729), .B1(new_n770), .B2(new_n772), .ZN(new_n777));
  NOR2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n695), .B1(new_n776), .B2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n666), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n613), .A2(new_n563), .A3(new_n567), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n768), .A2(new_n769), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  INV_X1    g598(.A(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n779), .A2(new_n785), .ZN(new_n786));
  OAI211_X1 g600(.A(KEYINPUT47), .B(new_n695), .C1(new_n776), .C2(new_n778), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n656), .A2(new_n578), .A3(new_n781), .ZN(new_n789));
  NAND3_X1  g603(.A1(new_n788), .A2(new_n739), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G140), .ZN(G42));
  INV_X1    g605(.A(KEYINPUT106), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n725), .B(new_n664), .C1(new_n691), .C2(new_n690), .ZN(new_n793));
  XOR2_X1   g607(.A(new_n661), .B(KEYINPUT105), .Z(new_n794));
  NOR3_X1   g608(.A1(new_n643), .A2(new_n378), .A3(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n735), .A2(new_n434), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n674), .A2(new_n795), .A3(new_n721), .A4(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n792), .B1(new_n793), .B2(new_n798), .ZN(new_n799));
  INV_X1    g613(.A(new_n691), .ZN(new_n800));
  OAI211_X1 g614(.A(new_n800), .B(new_n658), .C1(new_n739), .C2(new_n663), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n797), .A3(KEYINPUT106), .A4(new_n725), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n793), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(KEYINPUT52), .A3(new_n797), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n804), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n622), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n515), .A2(KEYINPUT103), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT103), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n512), .A2(new_n810), .A3(new_n514), .ZN(new_n811));
  AOI21_X1  g625(.A(new_n662), .B1(new_n809), .B2(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n628), .A2(new_n812), .A3(new_n629), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n813), .A2(new_n781), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n643), .A2(new_n808), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT104), .B1(new_n691), .B2(new_n815), .ZN(new_n816));
  AND3_X1   g630(.A1(new_n643), .A2(new_n808), .A3(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT104), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n818), .A3(new_n656), .A4(new_n441), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  AND2_X1   g634(.A1(new_n722), .A2(new_n712), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n724), .A2(new_n688), .A3(new_n689), .A4(new_n736), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n822), .A2(new_n756), .ZN(new_n823));
  OAI211_X1 g637(.A(new_n375), .B(new_n698), .C1(new_n631), .C2(new_n694), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n820), .A2(new_n821), .A3(new_n823), .A4(new_n824), .ZN(new_n825));
  INV_X1    g639(.A(new_n568), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(new_n524), .C1(new_n564), .C2(new_n565), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n475), .A2(new_n809), .A3(new_n811), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n827), .B1(new_n609), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n577), .A2(new_n829), .A3(new_n578), .A4(new_n441), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n830), .A2(new_n570), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n646), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n754), .A2(new_n825), .A3(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT53), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n807), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND4_X1   g649(.A1(new_n824), .A2(new_n820), .A3(new_n821), .A4(new_n823), .ZN(new_n836));
  INV_X1    g650(.A(new_n740), .ZN(new_n837));
  AOI21_X1  g651(.A(KEYINPUT98), .B1(new_n745), .B2(new_n747), .ZN(new_n838));
  NOR3_X1   g652(.A1(new_n752), .A2(new_n749), .A3(new_n746), .ZN(new_n839));
  OAI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n830), .A2(new_n570), .ZN(new_n841));
  INV_X1    g655(.A(new_n645), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n577), .A2(KEYINPUT91), .A3(new_n643), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g658(.A(new_n841), .B1(new_n844), .B2(new_n636), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n840), .A3(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n799), .A2(new_n802), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n847), .A2(KEYINPUT52), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n846), .B1(new_n804), .B2(new_n848), .ZN(new_n849));
  OAI211_X1 g663(.A(KEYINPUT54), .B(new_n835), .C1(new_n849), .C2(new_n834), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT54), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n807), .A2(new_n833), .A3(KEYINPUT53), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n851), .B(new_n852), .C1(new_n849), .C2(KEYINPUT53), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n266), .A2(new_n660), .ZN(new_n854));
  AND2_X1   g668(.A1(new_n854), .A2(new_n673), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n434), .A2(new_n697), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n856), .A2(new_n728), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n604), .A2(new_n608), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n855), .A2(KEYINPUT109), .A3(new_n857), .A4(new_n858), .ZN(new_n859));
  INV_X1    g673(.A(KEYINPUT109), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n857), .A2(new_n854), .A3(new_n673), .ZN(new_n861));
  INV_X1    g675(.A(new_n858), .ZN(new_n862));
  OAI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n765), .A2(new_n518), .A3(new_n857), .ZN(new_n864));
  AOI22_X1  g678(.A1(new_n859), .A2(new_n863), .B1(new_n864), .B2(new_n724), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n434), .A2(new_n695), .A3(new_n697), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n675), .A2(new_n610), .A3(new_n677), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n866), .A2(new_n867), .A3(KEYINPUT108), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT108), .B1(new_n866), .B2(new_n867), .ZN(new_n869));
  AND2_X1   g683(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT50), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n765), .A2(new_n518), .A3(new_n717), .ZN(new_n872));
  NOR3_X1   g686(.A1(new_n870), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n765), .A2(new_n518), .A3(new_n717), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n869), .ZN(new_n875));
  AOI21_X1  g689(.A(KEYINPUT50), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n865), .B1(new_n873), .B2(new_n876), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(KEYINPUT110), .ZN(new_n878));
  OAI21_X1  g692(.A(new_n871), .B1(new_n870), .B2(new_n872), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n874), .A2(KEYINPUT50), .A3(new_n875), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT110), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n881), .A2(new_n882), .A3(new_n865), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n872), .A2(new_n781), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT101), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n856), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n434), .A2(KEYINPUT101), .A3(new_n697), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT107), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n886), .A2(KEYINPUT107), .A3(new_n887), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n695), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n884), .B1(new_n788), .B2(new_n892), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n878), .A2(KEYINPUT51), .A3(new_n883), .A4(new_n893), .ZN(new_n894));
  OAI211_X1 g708(.A(G952), .B(new_n242), .C1(new_n861), .C2(new_n609), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n895), .B1(new_n705), .B2(new_n874), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n864), .A2(new_n745), .ZN(new_n897));
  AND2_X1   g711(.A1(new_n897), .A2(KEYINPUT48), .ZN(new_n898));
  NOR2_X1   g712(.A1(new_n897), .A2(KEYINPUT48), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n893), .A2(new_n881), .A3(new_n865), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT51), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g717(.A1(new_n894), .A2(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n850), .A2(new_n853), .A3(new_n904), .ZN(new_n905));
  NOR2_X1   g719(.A1(G952), .A2(G953), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT111), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n905), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n679), .A2(new_n695), .A3(new_n826), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n909), .A2(new_n266), .A3(new_n761), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n888), .A2(KEYINPUT49), .ZN(new_n912));
  OAI211_X1 g726(.A(new_n673), .B(new_n910), .C1(new_n911), .C2(new_n912), .ZN(new_n913));
  XOR2_X1   g727(.A(new_n913), .B(KEYINPUT102), .Z(new_n914));
  NAND2_X1  g728(.A1(new_n908), .A2(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT112), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n908), .A2(KEYINPUT112), .A3(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(G75));
  NAND2_X1  g733(.A1(new_n848), .A2(new_n804), .ZN(new_n920));
  AOI21_X1  g734(.A(KEYINPUT53), .B1(new_n920), .B2(new_n833), .ZN(new_n921));
  INV_X1    g735(.A(new_n852), .ZN(new_n922));
  OAI211_X1 g736(.A(G210), .B(G902), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT56), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n539), .A2(new_n546), .ZN(new_n925));
  XOR2_X1   g739(.A(new_n925), .B(new_n544), .Z(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(KEYINPUT55), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT114), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n923), .A2(new_n924), .A3(new_n928), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n242), .A2(G952), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(KEYINPUT115), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n929), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT113), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n923), .A2(new_n933), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n799), .A2(new_n802), .A3(new_n803), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n803), .B1(new_n799), .B2(new_n802), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n833), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n937), .A2(new_n834), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n188), .B1(new_n938), .B2(new_n852), .ZN(new_n939));
  AOI21_X1  g753(.A(KEYINPUT113), .B1(new_n939), .B2(G210), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n924), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n932), .B1(new_n941), .B2(new_n927), .ZN(G51));
  OAI21_X1  g756(.A(KEYINPUT54), .B1(new_n921), .B2(new_n922), .ZN(new_n943));
  AND2_X1   g757(.A1(new_n943), .A2(new_n853), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n729), .B(KEYINPUT57), .Z(new_n945));
  OAI21_X1  g759(.A(new_n425), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n939), .A2(new_n770), .A3(new_n772), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n930), .B1(new_n946), .B2(new_n947), .ZN(G54));
  INV_X1    g762(.A(KEYINPUT116), .ZN(new_n949));
  AND2_X1   g763(.A1(KEYINPUT58), .A2(G475), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n939), .A2(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(new_n464), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n949), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n930), .B1(new_n951), .B2(new_n952), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n939), .A2(KEYINPUT116), .A3(new_n464), .A4(new_n950), .ZN(new_n955));
  AND3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G60));
  INV_X1    g770(.A(new_n592), .ZN(new_n957));
  NAND2_X1  g771(.A1(G478), .A2(G902), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT59), .Z(new_n959));
  AOI211_X1 g773(.A(new_n957), .B(new_n959), .C1(new_n943), .C2(new_n853), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n850), .B2(new_n853), .ZN(new_n961));
  NOR2_X1   g775(.A1(new_n961), .A2(new_n592), .ZN(new_n962));
  INV_X1    g776(.A(new_n931), .ZN(new_n963));
  NOR3_X1   g777(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(G63));
  XOR2_X1   g778(.A(new_n261), .B(KEYINPUT118), .Z(new_n965));
  NOR2_X1   g779(.A1(new_n921), .A2(new_n922), .ZN(new_n966));
  NAND2_X1  g780(.A1(G217), .A2(G902), .ZN(new_n967));
  XNOR2_X1  g781(.A(new_n967), .B(KEYINPUT60), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n965), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n968), .B1(new_n938), .B2(new_n852), .ZN(new_n970));
  XNOR2_X1  g784(.A(new_n639), .B(KEYINPUT117), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n969), .A2(new_n931), .A3(new_n972), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND4_X1  g789(.A1(new_n969), .A2(new_n972), .A3(KEYINPUT61), .A4(new_n931), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(G66));
  AND3_X1   g791(.A1(new_n845), .A2(new_n824), .A3(new_n821), .ZN(new_n978));
  OR3_X1    g792(.A1(new_n978), .A2(KEYINPUT119), .A3(G953), .ZN(new_n979));
  OAI21_X1  g793(.A(KEYINPUT119), .B1(new_n978), .B2(G953), .ZN(new_n980));
  INV_X1    g794(.A(G224), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n522), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n979), .A2(new_n980), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n925), .B1(G898), .B2(new_n242), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  XNOR2_X1  g799(.A(new_n356), .B(new_n459), .ZN(new_n986));
  AOI21_X1  g800(.A(new_n986), .B1(G900), .B2(G953), .ZN(new_n987));
  INV_X1    g801(.A(new_n778), .ZN(new_n988));
  AOI22_X1  g802(.A1(new_n777), .A2(KEYINPUT46), .B1(new_n433), .B2(new_n427), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n378), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  NAND4_X1  g804(.A1(new_n990), .A2(new_n745), .A3(new_n666), .A4(new_n721), .ZN(new_n991));
  AND4_X1   g805(.A1(new_n840), .A2(new_n790), .A3(new_n991), .A4(new_n756), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT121), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n793), .B(new_n993), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n783), .A2(KEYINPUT123), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT123), .B1(new_n783), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n987), .B1(new_n997), .B2(G953), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n781), .B1(new_n609), .B2(new_n828), .ZN(new_n999));
  NAND4_X1  g813(.A1(new_n375), .A2(new_n441), .A3(new_n999), .A4(new_n666), .ZN(new_n1000));
  AND3_X1   g814(.A1(new_n783), .A2(new_n790), .A3(new_n1000), .ZN(new_n1001));
  AND3_X1   g815(.A1(new_n994), .A2(KEYINPUT62), .A3(new_n682), .ZN(new_n1002));
  AOI21_X1  g816(.A(KEYINPUT62), .B1(new_n994), .B2(new_n682), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  NAND2_X1  g818(.A1(new_n1004), .A2(KEYINPUT122), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT122), .ZN(new_n1006));
  OAI211_X1 g820(.A(new_n1001), .B(new_n1006), .C1(new_n1002), .C2(new_n1003), .ZN(new_n1007));
  AOI21_X1  g821(.A(G953), .B1(new_n1005), .B2(new_n1007), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n986), .B(KEYINPUT120), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n998), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1009), .A2(KEYINPUT124), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n242), .B1(G227), .B2(G900), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1014));
  OAI211_X1 g828(.A(new_n998), .B(new_n1014), .C1(new_n1008), .C2(new_n1009), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1013), .A2(new_n1015), .ZN(G72));
  NAND2_X1  g830(.A1(G472), .A2(G902), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT63), .Z(new_n1018));
  NAND3_X1  g832(.A1(new_n845), .A2(new_n824), .A3(new_n821), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1018), .B1(new_n997), .B2(new_n1019), .ZN(new_n1020));
  INV_X1    g834(.A(new_n357), .ZN(new_n1021));
  NOR2_X1   g835(.A1(new_n1021), .A2(new_n326), .ZN(new_n1022));
  AOI21_X1  g836(.A(new_n930), .B1(new_n1020), .B2(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1018), .ZN(new_n1024));
  XNOR2_X1  g838(.A(new_n370), .B(KEYINPUT126), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1024), .B1(new_n1025), .B2(new_n331), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n835), .B(new_n1026), .C1(new_n849), .C2(new_n834), .ZN(new_n1027));
  INV_X1    g841(.A(KEYINPUT127), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1023), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g845(.A1(new_n1021), .A2(new_n326), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1005), .A2(new_n978), .A3(new_n1007), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n1033), .A2(new_n1018), .ZN(new_n1034));
  INV_X1    g848(.A(KEYINPUT125), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1032), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  NAND3_X1  g850(.A1(new_n1033), .A2(KEYINPUT125), .A3(new_n1018), .ZN(new_n1037));
  AOI21_X1  g851(.A(new_n1031), .B1(new_n1036), .B2(new_n1037), .ZN(G57));
endmodule


