//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 0 1 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 0 1 0 1 1 1 0 0 0 0 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n772, new_n774, new_n775, new_n776,
    new_n777, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n801, new_n802, new_n803, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1014, new_n1015, new_n1016, new_n1017,
    new_n1018, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067,
    new_n1068, new_n1069;
  INV_X1    g000(.A(KEYINPUT99), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT95), .ZN(new_n189));
  INV_X1    g003(.A(G134), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT13), .B1(new_n191), .B2(G128), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n191), .A2(G128), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(new_n193), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n194), .A2(KEYINPUT93), .B1(KEYINPUT13), .B2(new_n195), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT93), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n192), .A2(new_n197), .A3(new_n193), .ZN(new_n198));
  AOI21_X1  g012(.A(new_n190), .B1(new_n196), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G128), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n193), .A2(new_n201), .A3(new_n190), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT94), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n193), .A2(new_n201), .A3(KEYINPUT94), .A4(new_n190), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G122), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G122), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n210), .A3(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n206), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n189), .B1(new_n199), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n194), .A2(KEYINPUT93), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n195), .A2(KEYINPUT13), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n198), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(G134), .ZN(new_n221));
  AOI22_X1  g035(.A1(new_n204), .A2(new_n205), .B1(new_n212), .B2(new_n214), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n221), .A2(KEYINPUT95), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n190), .B1(new_n193), .B2(new_n201), .ZN(new_n224));
  INV_X1    g038(.A(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n225), .A2(KEYINPUT96), .A3(new_n202), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT96), .ZN(new_n227));
  INV_X1    g041(.A(new_n202), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n228), .B2(new_n224), .ZN(new_n229));
  AND3_X1   g043(.A1(new_n226), .A2(new_n229), .A3(new_n214), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n209), .A2(KEYINPUT14), .A3(G122), .ZN(new_n231));
  AND2_X1   g045(.A1(new_n231), .A2(G107), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n232), .B1(KEYINPUT14), .B2(new_n211), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(KEYINPUT97), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n235));
  OAI211_X1 g049(.A(new_n232), .B(new_n235), .C1(KEYINPUT14), .C2(new_n211), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n234), .A2(new_n236), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n217), .A2(new_n223), .B1(new_n230), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT9), .B(G234), .ZN(new_n239));
  INV_X1    g053(.A(G217), .ZN(new_n240));
  NOR3_X1   g054(.A1(new_n239), .A2(new_n240), .A3(G953), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(KEYINPUT98), .A3(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n230), .A2(new_n237), .ZN(new_n243));
  NOR3_X1   g057(.A1(new_n199), .A2(new_n216), .A3(new_n189), .ZN(new_n244));
  AOI21_X1  g058(.A(KEYINPUT95), .B1(new_n221), .B2(new_n222), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  INV_X1    g060(.A(new_n241), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n242), .A2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(KEYINPUT98), .B1(new_n238), .B2(new_n241), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n188), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G478), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(KEYINPUT15), .ZN(new_n253));
  OR2_X1    g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n253), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(G221), .ZN(new_n258));
  INV_X1    g072(.A(new_n239), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n259), .B2(new_n188), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n261), .B1(new_n190), .B2(G137), .ZN(new_n262));
  INV_X1    g076(.A(G137), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT11), .A3(G134), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n190), .A2(G137), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(KEYINPUT67), .B1(new_n266), .B2(G131), .ZN(new_n267));
  INV_X1    g081(.A(new_n267), .ZN(new_n268));
  AND2_X1   g082(.A1(KEYINPUT66), .A2(G131), .ZN(new_n269));
  NOR2_X1   g083(.A1(KEYINPUT66), .A2(G131), .ZN(new_n270));
  NOR2_X1   g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n271), .A2(new_n262), .A3(new_n264), .A4(new_n265), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n264), .A2(new_n265), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT11), .B1(new_n263), .B2(G134), .ZN(new_n274));
  OAI211_X1 g088(.A(KEYINPUT67), .B(G131), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n268), .A2(new_n272), .A3(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n191), .A2(G146), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n278));
  OAI21_X1  g092(.A(G128), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G146), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(G143), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n191), .A2(G146), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  OAI21_X1  g098(.A(KEYINPUT65), .B1(new_n191), .B2(G146), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n286), .A2(new_n280), .A3(G143), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n200), .A2(KEYINPUT1), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n285), .A2(new_n287), .A3(new_n282), .A4(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n284), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G104), .ZN(new_n291));
  OAI21_X1  g105(.A(KEYINPUT3), .B1(new_n291), .B2(G107), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT3), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n293), .A2(new_n213), .A3(G104), .ZN(new_n294));
  INV_X1    g108(.A(G101), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(G107), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n292), .A2(new_n294), .A3(new_n295), .A4(new_n296), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n291), .A2(G107), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n213), .A2(G104), .ZN(new_n299));
  OAI21_X1  g113(.A(G101), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n297), .A2(new_n300), .ZN(new_n303));
  NAND3_X1  g117(.A1(new_n285), .A2(new_n287), .A3(new_n282), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(new_n279), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n303), .B1(new_n289), .B2(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n276), .B1(new_n302), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(KEYINPUT12), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n305), .A2(new_n289), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n301), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n292), .A2(new_n294), .A3(new_n296), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G101), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n314), .A2(KEYINPUT4), .A3(new_n297), .ZN(new_n315));
  AND3_X1   g129(.A1(new_n285), .A2(new_n287), .A3(new_n282), .ZN(new_n316));
  NAND2_X1  g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT64), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(KEYINPUT64), .A2(KEYINPUT0), .A3(G128), .ZN(new_n321));
  AND2_X1   g135(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT0), .ZN(new_n323));
  AOI22_X1  g137(.A1(new_n281), .A2(new_n282), .B1(new_n323), .B2(new_n200), .ZN(new_n324));
  AOI22_X1  g138(.A1(new_n316), .A2(new_n318), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g139(.A(KEYINPUT4), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n313), .A2(new_n326), .A3(G101), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n315), .A2(new_n325), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n275), .A2(new_n272), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(new_n267), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n311), .B1(new_n284), .B2(new_n289), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n301), .ZN(new_n332));
  NAND4_X1  g146(.A1(new_n312), .A2(new_n328), .A3(new_n330), .A4(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT12), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n276), .B(new_n334), .C1(new_n302), .C2(new_n306), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n308), .A2(new_n333), .A3(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(G110), .B(G140), .ZN(new_n337));
  INV_X1    g151(.A(G953), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G227), .ZN(new_n339));
  XNOR2_X1  g153(.A(new_n337), .B(new_n339), .ZN(new_n340));
  XNOR2_X1  g154(.A(KEYINPUT81), .B(KEYINPUT82), .ZN(new_n341));
  XNOR2_X1  g155(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n336), .A2(new_n343), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n332), .B1(new_n306), .B2(KEYINPUT10), .ZN(new_n345));
  INV_X1    g159(.A(new_n328), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n276), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(new_n342), .A3(new_n333), .ZN(new_n348));
  AND2_X1   g162(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g163(.A(G469), .B1(new_n349), .B2(G902), .ZN(new_n350));
  INV_X1    g164(.A(G469), .ZN(new_n351));
  INV_X1    g165(.A(new_n333), .ZN(new_n352));
  AOI22_X1  g166(.A1(new_n310), .A2(new_n311), .B1(new_n301), .B2(new_n331), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n330), .B1(new_n353), .B2(new_n328), .ZN(new_n354));
  OAI211_X1 g168(.A(KEYINPUT83), .B(new_n343), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n308), .A2(new_n333), .A3(new_n342), .A4(new_n335), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n347), .A2(new_n333), .ZN(new_n358));
  AOI21_X1  g172(.A(KEYINPUT83), .B1(new_n358), .B2(new_n343), .ZN(new_n359));
  OAI211_X1 g173(.A(new_n351), .B(new_n188), .C1(new_n357), .C2(new_n359), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n260), .B1(new_n350), .B2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(G475), .ZN(new_n362));
  INV_X1    g176(.A(G237), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n363), .A2(new_n338), .A3(G214), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n191), .ZN(new_n365));
  NOR2_X1   g179(.A1(G237), .A2(G953), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n366), .A2(G143), .A3(G214), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT90), .ZN(new_n369));
  AND3_X1   g183(.A1(new_n369), .A2(KEYINPUT18), .A3(G131), .ZN(new_n370));
  OR2_X1    g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n368), .A2(new_n370), .ZN(new_n372));
  INV_X1    g186(.A(G140), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G125), .ZN(new_n374));
  INV_X1    g188(.A(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G140), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G146), .ZN(new_n378));
  XNOR2_X1  g192(.A(G125), .B(G140), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n280), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n371), .A2(new_n372), .A3(new_n381), .ZN(new_n382));
  OR2_X1    g196(.A1(new_n269), .A2(new_n270), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n364), .A2(new_n191), .ZN(new_n384));
  AOI21_X1  g198(.A(G143), .B1(new_n366), .B2(G214), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n383), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g200(.A(KEYINPUT17), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n365), .A2(new_n271), .A3(new_n367), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n386), .A2(new_n387), .A3(new_n388), .ZN(new_n389));
  NAND3_X1  g203(.A1(new_n368), .A2(KEYINPUT17), .A3(new_n383), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT16), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n392), .A2(new_n373), .A3(G125), .ZN(new_n393));
  OAI211_X1 g207(.A(G146), .B(new_n393), .C1(new_n377), .C2(new_n392), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT77), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n393), .B1(new_n377), .B2(new_n392), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n280), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n379), .A2(KEYINPUT16), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT77), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G146), .A4(new_n393), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n395), .A2(new_n397), .A3(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n382), .B1(new_n391), .B2(new_n401), .ZN(new_n402));
  XNOR2_X1  g216(.A(G113), .B(G122), .ZN(new_n403));
  XNOR2_X1  g217(.A(new_n403), .B(new_n291), .ZN(new_n404));
  INV_X1    g218(.A(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n402), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g220(.A(new_n404), .B(new_n382), .C1(new_n391), .C2(new_n401), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(new_n188), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n362), .B1(new_n409), .B2(KEYINPUT92), .ZN(new_n410));
  INV_X1    g224(.A(KEYINPUT92), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n408), .A2(new_n411), .A3(new_n188), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n386), .A2(new_n388), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n414));
  XNOR2_X1  g228(.A(new_n379), .B(new_n414), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n413), .B(new_n394), .C1(G146), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n382), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n417), .A2(new_n405), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n418), .A2(new_n407), .ZN(new_n419));
  NOR2_X1   g233(.A1(G475), .A2(G902), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  AOI21_X1  g235(.A(KEYINPUT91), .B1(new_n418), .B2(new_n407), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(KEYINPUT20), .B2(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n419), .A2(KEYINPUT91), .A3(new_n424), .A4(new_n420), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n410), .A2(new_n412), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n338), .A2(G952), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n427), .B1(G234), .B2(G237), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n188), .B(new_n338), .C1(G234), .C2(G237), .ZN(new_n429));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(G898), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n428), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n257), .A2(new_n361), .A3(new_n426), .A4(new_n432), .ZN(new_n433));
  OAI21_X1  g247(.A(G210), .B1(G237), .B2(G902), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n323), .A2(new_n200), .ZN(new_n436));
  NAND4_X1  g250(.A1(new_n283), .A2(new_n436), .A3(new_n320), .A4(new_n321), .ZN(new_n437));
  NAND4_X1  g251(.A1(new_n285), .A2(new_n287), .A3(new_n318), .A4(new_n282), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(G125), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n284), .A2(new_n375), .A3(new_n289), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G224), .ZN(new_n443));
  NOR2_X1   g257(.A1(new_n443), .A2(G953), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n442), .B(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(KEYINPUT2), .B(G113), .Z(new_n446));
  XNOR2_X1  g260(.A(G116), .B(G119), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT69), .ZN(new_n448));
  XNOR2_X1  g262(.A(KEYINPUT2), .B(G113), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT69), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n209), .A2(G119), .ZN(new_n451));
  INV_X1    g265(.A(G119), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(G116), .ZN(new_n453));
  OAI211_X1 g267(.A(new_n449), .B(new_n450), .C1(new_n451), .C2(new_n453), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n448), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n315), .A2(new_n455), .A3(new_n327), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n447), .A2(KEYINPUT5), .ZN(new_n457));
  INV_X1    g271(.A(G113), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT5), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n458), .B1(new_n451), .B2(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n457), .A2(new_n460), .B1(new_n446), .B2(new_n447), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(new_n301), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n456), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT6), .ZN(new_n464));
  XNOR2_X1  g278(.A(G110), .B(G122), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n463), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g283(.A1(new_n463), .A2(KEYINPUT86), .A3(new_n464), .A4(new_n466), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n464), .B1(new_n463), .B2(new_n466), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n456), .A2(new_n462), .A3(new_n465), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n472), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n474));
  AOI21_X1  g288(.A(KEYINPUT85), .B1(new_n472), .B2(new_n473), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n445), .B(new_n471), .C1(new_n474), .C2(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT8), .ZN(new_n478));
  XNOR2_X1  g292(.A(new_n465), .B(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n461), .B2(new_n303), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT88), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n452), .A2(G116), .ZN(new_n482));
  OAI21_X1  g296(.A(G113), .B1(new_n482), .B2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT87), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  OAI211_X1 g299(.A(KEYINPUT87), .B(G113), .C1(new_n482), .C2(KEYINPUT5), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n457), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n446), .A2(new_n447), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n480), .B(new_n481), .C1(new_n489), .C2(new_n303), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n465), .B(KEYINPUT8), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n457), .A2(new_n460), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n492), .A2(new_n488), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n491), .B1(new_n493), .B2(new_n301), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n303), .B1(new_n487), .B2(new_n488), .ZN(new_n495));
  OAI21_X1  g309(.A(KEYINPUT88), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n490), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT89), .ZN(new_n498));
  OAI21_X1  g312(.A(KEYINPUT7), .B1(new_n443), .B2(G953), .ZN(new_n499));
  AND3_X1   g313(.A1(new_n284), .A2(new_n375), .A3(new_n289), .ZN(new_n500));
  AOI21_X1  g314(.A(new_n375), .B1(new_n437), .B2(new_n438), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g316(.A(new_n499), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n440), .A2(new_n441), .A3(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n497), .A2(new_n498), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(new_n473), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n505), .B1(new_n490), .B2(new_n496), .ZN(new_n509));
  NOR2_X1   g323(.A1(new_n509), .A2(new_n498), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n188), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n435), .B1(new_n477), .B2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n473), .ZN(new_n513));
  AOI21_X1  g327(.A(new_n513), .B1(new_n509), .B2(new_n498), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n497), .A2(new_n506), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(KEYINPUT89), .ZN(new_n516));
  AOI21_X1  g330(.A(G902), .B1(new_n514), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n517), .A2(new_n434), .A3(new_n476), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n512), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g333(.A(G214), .B1(G237), .B2(G902), .ZN(new_n520));
  XOR2_X1   g334(.A(new_n520), .B(KEYINPUT84), .Z(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n519), .A2(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n187), .B1(new_n433), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT73), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n200), .B2(G119), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n200), .A2(G119), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n452), .A2(KEYINPUT73), .A3(G128), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n527), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT74), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT74), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n526), .A2(new_n528), .A3(new_n531), .A4(new_n527), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n530), .A2(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(G110), .ZN(new_n534));
  AND2_X1   g348(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n535));
  NOR2_X1   g349(.A1(new_n534), .A2(KEYINPUT24), .ZN(new_n536));
  OAI21_X1  g350(.A(KEYINPUT75), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT24), .B(G110), .ZN(new_n538));
  INV_X1    g352(.A(KEYINPUT75), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AND2_X1   g354(.A1(new_n537), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT76), .B1(new_n452), .B2(G128), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT23), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT23), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n527), .A2(KEYINPUT76), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n452), .A2(G128), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n543), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI22_X1  g361(.A1(new_n533), .A2(new_n541), .B1(G110), .B2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n548), .A2(new_n401), .ZN(new_n549));
  AND2_X1   g363(.A1(new_n394), .A2(new_n380), .ZN(new_n550));
  AOI22_X1  g364(.A1(new_n530), .A2(new_n532), .B1(new_n540), .B2(new_n537), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n547), .A2(G110), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(KEYINPUT78), .ZN(new_n554));
  AND2_X1   g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI211_X1 g369(.A(new_n550), .B(KEYINPUT78), .C1(new_n551), .C2(new_n552), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  OAI21_X1  g371(.A(new_n549), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  INV_X1    g373(.A(G234), .ZN(new_n560));
  NOR3_X1   g374(.A1(new_n258), .A2(new_n560), .A3(G953), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n559), .B(new_n561), .Z(new_n562));
  INV_X1    g376(.A(new_n562), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n558), .A2(KEYINPUT79), .A3(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT79), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n553), .A2(new_n554), .ZN(new_n566));
  AOI22_X1  g380(.A1(new_n566), .A2(new_n556), .B1(new_n401), .B2(new_n548), .ZN(new_n567));
  OAI21_X1  g381(.A(new_n565), .B1(new_n567), .B2(new_n562), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  OAI211_X1 g383(.A(new_n549), .B(new_n562), .C1(new_n555), .C2(new_n557), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g385(.A(G217), .B1(new_n560), .B2(G902), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n188), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n571), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n188), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n576), .B1(new_n568), .B2(new_n564), .ZN(new_n577));
  OAI21_X1  g391(.A(KEYINPUT80), .B1(new_n577), .B2(KEYINPUT25), .ZN(new_n578));
  AOI21_X1  g392(.A(G902), .B1(new_n567), .B2(new_n562), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n569), .A2(KEYINPUT25), .A3(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  XOR2_X1   g396(.A(new_n572), .B(KEYINPUT72), .Z(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT79), .B1(new_n558), .B2(new_n563), .ZN(new_n585));
  NOR3_X1   g399(.A1(new_n567), .A2(new_n565), .A3(new_n562), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n579), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT25), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n584), .B1(new_n589), .B2(KEYINPUT80), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n575), .B1(new_n582), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n190), .A2(G137), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n263), .A2(G134), .ZN(new_n593));
  OAI21_X1  g407(.A(G131), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n594), .B1(new_n266), .B2(new_n383), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(KEYINPUT68), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT68), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n272), .A2(new_n597), .A3(new_n594), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n596), .A2(new_n290), .A3(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n325), .B1(new_n329), .B2(new_n267), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT30), .ZN(new_n601));
  NAND3_X1  g415(.A1(new_n599), .A2(new_n600), .A3(new_n601), .ZN(new_n602));
  INV_X1    g416(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n595), .A2(KEYINPUT70), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT70), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n272), .A2(new_n605), .A3(new_n594), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n290), .A3(new_n606), .ZN(new_n607));
  AOI21_X1  g421(.A(new_n601), .B1(new_n607), .B2(new_n600), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n455), .B1(new_n603), .B2(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n455), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n607), .A2(new_n600), .A3(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n366), .A2(G210), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n612), .B(KEYINPUT27), .ZN(new_n613));
  XNOR2_X1  g427(.A(KEYINPUT26), .B(G101), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n609), .A2(new_n611), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(KEYINPUT31), .ZN(new_n617));
  INV_X1    g431(.A(new_n611), .ZN(new_n618));
  AND2_X1   g432(.A1(new_n607), .A2(new_n600), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n602), .B1(new_n619), .B2(new_n601), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n618), .B1(new_n620), .B2(new_n455), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT31), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n621), .A2(new_n622), .A3(new_n615), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT71), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n611), .A2(KEYINPUT28), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT28), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n607), .A2(new_n600), .A3(new_n610), .A4(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n625), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(new_n610), .B1(new_n599), .B2(new_n600), .ZN(new_n629));
  INV_X1    g443(.A(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n615), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n624), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n629), .B1(new_n625), .B2(new_n627), .ZN(new_n634));
  NOR3_X1   g448(.A1(new_n634), .A2(KEYINPUT71), .A3(new_n615), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n617), .B(new_n623), .C1(new_n633), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(G472), .A2(G902), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT32), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT32), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n639), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT29), .ZN(new_n643));
  OAI21_X1  g457(.A(new_n643), .B1(new_n621), .B2(new_n615), .ZN(new_n644));
  AOI21_X1  g458(.A(new_n644), .B1(new_n615), .B2(new_n634), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n619), .A2(new_n610), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n625), .B2(new_n627), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT29), .A3(new_n615), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(new_n188), .ZN(new_n649));
  OAI21_X1  g463(.A(G472), .B1(new_n645), .B2(new_n649), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n591), .B1(new_n642), .B2(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(new_n523), .ZN(new_n652));
  INV_X1    g466(.A(new_n426), .ZN(new_n653));
  NOR3_X1   g467(.A1(new_n256), .A2(new_n653), .A3(new_n431), .ZN(new_n654));
  NAND4_X1  g468(.A1(new_n652), .A2(new_n654), .A3(KEYINPUT99), .A4(new_n361), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n524), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n656), .B(G101), .ZN(G3));
  NAND3_X1  g471(.A1(new_n589), .A2(KEYINPUT80), .A3(new_n580), .ZN(new_n658));
  AOI21_X1  g472(.A(KEYINPUT25), .B1(new_n569), .B2(new_n579), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT80), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n583), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI22_X1  g475(.A1(new_n658), .A2(new_n661), .B1(new_n574), .B2(new_n571), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n662), .A2(new_n361), .ZN(new_n663));
  AND3_X1   g477(.A1(new_n517), .A2(new_n434), .A3(new_n476), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n434), .B1(new_n517), .B2(new_n476), .ZN(new_n665));
  OAI211_X1 g479(.A(new_n520), .B(new_n432), .C1(new_n664), .C2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(KEYINPUT33), .B1(new_n238), .B2(new_n241), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n217), .A2(new_n223), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n668), .A2(new_n243), .A3(new_n241), .ZN(new_n669));
  OAI21_X1  g483(.A(KEYINPUT100), .B1(new_n667), .B2(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n238), .A2(new_n241), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT100), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n248), .A2(new_n671), .A3(new_n672), .A4(KEYINPUT33), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n670), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT33), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n675), .B1(new_n249), .B2(new_n250), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n252), .A2(G902), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n251), .A2(new_n252), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n680), .A2(new_n653), .ZN(new_n681));
  NOR2_X1   g495(.A1(new_n666), .A2(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n636), .A2(new_n188), .ZN(new_n683));
  AOI22_X1  g497(.A1(new_n683), .A2(G472), .B1(new_n637), .B2(new_n636), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n663), .A2(new_n682), .A3(new_n684), .ZN(new_n685));
  XOR2_X1   g499(.A(KEYINPUT34), .B(G104), .Z(new_n686));
  XNOR2_X1  g500(.A(new_n685), .B(new_n686), .ZN(G6));
  NAND2_X1  g501(.A1(new_n410), .A2(new_n412), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n421), .B(KEYINPUT20), .ZN(new_n689));
  AND2_X1   g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n256), .A2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n666), .A2(new_n691), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n663), .A2(new_n684), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(new_n213), .ZN(new_n694));
  XNOR2_X1  g508(.A(KEYINPUT101), .B(KEYINPUT35), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n694), .B(new_n695), .ZN(G9));
  NOR2_X1   g510(.A1(new_n563), .A2(KEYINPUT36), .ZN(new_n697));
  XNOR2_X1  g511(.A(new_n567), .B(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n698), .A2(new_n573), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n699), .B1(new_n658), .B2(new_n661), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT102), .ZN(new_n701));
  NOR2_X1   g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI211_X1 g516(.A(KEYINPUT102), .B(new_n699), .C1(new_n658), .C2(new_n661), .ZN(new_n703));
  NOR2_X1   g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n704), .A2(new_n684), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n524), .A2(new_n655), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  XOR2_X1   g521(.A(KEYINPUT37), .B(G110), .Z(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(KEYINPUT103), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n707), .B(new_n709), .ZN(G12));
  AND3_X1   g524(.A1(new_n636), .A2(new_n640), .A3(new_n637), .ZN(new_n711));
  AOI21_X1  g525(.A(new_n640), .B1(new_n636), .B2(new_n637), .ZN(new_n712));
  OAI21_X1  g526(.A(new_n650), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(new_n361), .ZN(new_n714));
  NOR3_X1   g528(.A1(new_n714), .A2(new_n702), .A3(new_n703), .ZN(new_n715));
  XOR2_X1   g529(.A(KEYINPUT104), .B(G900), .Z(new_n716));
  AOI21_X1  g530(.A(new_n428), .B1(new_n429), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n690), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n257), .A2(new_n719), .ZN(new_n720));
  INV_X1    g534(.A(new_n520), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n721), .B1(new_n512), .B2(new_n518), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n715), .A2(new_n724), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G128), .ZN(G30));
  AOI21_X1  g540(.A(new_n632), .B1(new_n609), .B2(new_n611), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n611), .A2(new_n632), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n188), .B1(new_n646), .B2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(G472), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  INV_X1    g544(.A(KEYINPUT105), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n730), .B(new_n731), .ZN(new_n732));
  AOI21_X1  g546(.A(new_n732), .B1(new_n639), .B2(new_n641), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(KEYINPUT106), .ZN(new_n734));
  INV_X1    g548(.A(new_n734), .ZN(new_n735));
  XOR2_X1   g549(.A(new_n519), .B(KEYINPUT38), .Z(new_n736));
  INV_X1    g550(.A(new_n699), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n582), .B2(new_n590), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n256), .A2(new_n653), .ZN(new_n739));
  NOR4_X1   g553(.A1(new_n736), .A2(new_n721), .A3(new_n738), .A4(new_n739), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n717), .B(KEYINPUT39), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n361), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(new_n742), .B(KEYINPUT107), .Z(new_n743));
  AND2_X1   g557(.A1(new_n743), .A2(KEYINPUT40), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n743), .A2(KEYINPUT40), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n735), .B(new_n740), .C1(new_n744), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G143), .ZN(G45));
  NAND2_X1  g561(.A1(new_n738), .A2(KEYINPUT102), .ZN(new_n748));
  OAI211_X1 g562(.A(new_n701), .B(new_n737), .C1(new_n582), .C2(new_n590), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n748), .A2(new_n361), .A3(new_n713), .A4(new_n749), .ZN(new_n750));
  NAND2_X1  g564(.A1(new_n423), .A2(new_n425), .ZN(new_n751));
  AOI221_X4 g565(.A(new_n717), .B1(new_n688), .B2(new_n751), .C1(new_n678), .C2(new_n679), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n752), .A2(KEYINPUT108), .A3(new_n722), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n680), .A2(new_n653), .A3(new_n718), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n520), .B1(new_n664), .B2(new_n665), .ZN(new_n756));
  OAI21_X1  g570(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n753), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n750), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(new_n280), .ZN(G48));
  OAI21_X1  g574(.A(new_n188), .B1(new_n357), .B2(new_n359), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(G469), .ZN(new_n762));
  INV_X1    g576(.A(new_n260), .ZN(new_n763));
  AND3_X1   g577(.A1(new_n762), .A2(new_n763), .A3(new_n360), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n651), .A2(KEYINPUT109), .A3(new_n682), .A4(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n682), .A2(new_n713), .A3(new_n662), .A4(new_n764), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT109), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n765), .A2(new_n768), .ZN(new_n769));
  XNOR2_X1  g583(.A(KEYINPUT41), .B(G113), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n769), .B(new_n770), .ZN(G15));
  NAND4_X1  g585(.A1(new_n692), .A2(new_n713), .A3(new_n662), .A4(new_n764), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(G116), .ZN(G18));
  AND2_X1   g587(.A1(new_n713), .A2(new_n654), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n762), .A2(new_n763), .A3(new_n360), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n756), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n704), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G119), .ZN(G21));
  OAI211_X1 g592(.A(new_n623), .B(new_n617), .C1(new_n615), .C2(new_n647), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n779), .A2(new_n637), .ZN(new_n780));
  AND2_X1   g594(.A1(new_n623), .A2(new_n617), .ZN(new_n781));
  INV_X1    g595(.A(new_n635), .ZN(new_n782));
  OAI21_X1  g596(.A(KEYINPUT71), .B1(new_n634), .B2(new_n615), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  AOI21_X1  g598(.A(G902), .B1(new_n781), .B2(new_n784), .ZN(new_n785));
  INV_X1    g599(.A(G472), .ZN(new_n786));
  OAI21_X1  g600(.A(new_n780), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n591), .A2(new_n787), .ZN(new_n788));
  INV_X1    g602(.A(KEYINPUT110), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n762), .A2(new_n763), .A3(new_n360), .A4(new_n432), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n739), .A2(new_n756), .A3(new_n790), .ZN(new_n791));
  NAND3_X1  g605(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AOI22_X1  g606(.A1(new_n683), .A2(G472), .B1(new_n637), .B2(new_n779), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n662), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n426), .B1(new_n254), .B2(new_n255), .ZN(new_n795));
  NAND4_X1  g609(.A1(new_n764), .A2(new_n722), .A3(new_n432), .A4(new_n795), .ZN(new_n796));
  OAI21_X1  g610(.A(KEYINPUT110), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n792), .A2(new_n797), .ZN(new_n798));
  XOR2_X1   g612(.A(KEYINPUT111), .B(G122), .Z(new_n799));
  XNOR2_X1  g613(.A(new_n798), .B(new_n799), .ZN(G24));
  NOR2_X1   g614(.A1(new_n787), .A2(new_n700), .ZN(new_n801));
  NOR3_X1   g615(.A1(new_n755), .A2(new_n756), .A3(new_n775), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  XNOR2_X1  g617(.A(new_n803), .B(G125), .ZN(G27));
  INV_X1    g618(.A(KEYINPUT42), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n713), .A2(new_n662), .ZN(new_n806));
  NAND2_X1  g620(.A1(G469), .A2(G902), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT112), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n344), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n336), .A2(KEYINPUT112), .A3(new_n343), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n809), .A2(G469), .A3(new_n348), .A4(new_n810), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n360), .A2(new_n807), .A3(new_n811), .ZN(new_n812));
  AND2_X1   g626(.A1(new_n812), .A2(new_n763), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n664), .A2(new_n665), .A3(new_n721), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n752), .A2(new_n813), .A3(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n805), .B1(new_n806), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n812), .A2(new_n763), .ZN(new_n817));
  NAND3_X1  g631(.A1(new_n512), .A2(new_n518), .A3(new_n520), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n755), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n819), .A2(KEYINPUT42), .A3(new_n662), .A4(new_n713), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n816), .A2(new_n820), .ZN(new_n821));
  XNOR2_X1  g635(.A(new_n821), .B(G131), .ZN(G33));
  NOR2_X1   g636(.A1(new_n817), .A2(new_n818), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n651), .A2(new_n720), .A3(new_n823), .ZN(new_n824));
  XNOR2_X1  g638(.A(new_n824), .B(G134), .ZN(G36));
  NAND4_X1  g639(.A1(new_n809), .A2(KEYINPUT45), .A3(new_n348), .A4(new_n810), .ZN(new_n826));
  OAI211_X1 g640(.A(new_n826), .B(G469), .C1(KEYINPUT45), .C2(new_n349), .ZN(new_n827));
  NAND2_X1  g641(.A1(new_n827), .A2(new_n807), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT46), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n360), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n828), .A2(new_n829), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND2_X1   g647(.A1(new_n814), .A2(new_n741), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n763), .A3(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n835), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n700), .A2(new_n684), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n680), .A2(new_n426), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT44), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  INV_X1    g657(.A(new_n841), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n844), .A2(KEYINPUT44), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n836), .A2(new_n843), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(G137), .ZN(G39));
  NAND3_X1  g661(.A1(new_n833), .A2(KEYINPUT47), .A3(new_n763), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n763), .B1(new_n831), .B2(new_n832), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT47), .ZN(new_n850));
  NAND2_X1  g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  NOR4_X1   g666(.A1(new_n713), .A2(new_n662), .A3(new_n755), .A4(new_n818), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  XNOR2_X1  g668(.A(new_n854), .B(G140), .ZN(G42));
  AND2_X1   g669(.A1(new_n762), .A2(new_n360), .ZN(new_n856));
  XOR2_X1   g670(.A(new_n856), .B(KEYINPUT113), .Z(new_n857));
  NOR2_X1   g671(.A1(new_n857), .A2(KEYINPUT49), .ZN(new_n858));
  XOR2_X1   g672(.A(new_n858), .B(KEYINPUT114), .Z(new_n859));
  NOR3_X1   g673(.A1(new_n838), .A2(new_n521), .A3(new_n260), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n736), .A2(new_n662), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n861), .B1(KEYINPUT49), .B2(new_n857), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n859), .A2(new_n734), .A3(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n818), .A2(new_n775), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n864), .A2(new_n662), .A3(new_n428), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n735), .A2(new_n681), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n840), .A2(new_n428), .A3(new_n839), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n794), .ZN(new_n868));
  AND2_X1   g682(.A1(new_n868), .A2(new_n776), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n866), .A2(new_n427), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT48), .ZN(new_n871));
  INV_X1    g685(.A(new_n867), .ZN(new_n872));
  INV_X1    g686(.A(KEYINPUT119), .ZN(new_n873));
  NAND3_X1  g687(.A1(new_n872), .A2(new_n873), .A3(new_n864), .ZN(new_n874));
  INV_X1    g688(.A(new_n864), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT119), .B1(new_n867), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n871), .B1(new_n877), .B2(new_n651), .ZN(new_n878));
  AOI211_X1 g692(.A(KEYINPUT48), .B(new_n806), .C1(new_n874), .C2(new_n876), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n870), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(KEYINPUT120), .ZN(new_n881));
  INV_X1    g695(.A(KEYINPUT120), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n870), .B(new_n882), .C1(new_n879), .C2(new_n878), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g698(.A1(new_n735), .A2(new_n865), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n680), .A2(new_n653), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n877), .A2(new_n801), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n764), .A2(KEYINPUT118), .A3(new_n721), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT118), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n890), .B1(new_n775), .B2(new_n520), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n736), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(KEYINPUT50), .B1(new_n893), .B2(new_n868), .ZN(new_n894));
  AND3_X1   g708(.A1(new_n893), .A2(KEYINPUT50), .A3(new_n868), .ZN(new_n895));
  OAI211_X1 g709(.A(new_n887), .B(new_n888), .C1(new_n894), .C2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n848), .B(new_n851), .C1(new_n763), .C2(new_n857), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT117), .ZN(new_n898));
  INV_X1    g712(.A(new_n868), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n898), .B1(new_n899), .B2(new_n818), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n868), .A2(KEYINPUT117), .A3(new_n814), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n897), .A2(new_n900), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(KEYINPUT51), .B1(new_n896), .B2(new_n903), .ZN(new_n904));
  AND2_X1   g718(.A1(new_n887), .A2(new_n888), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT51), .ZN(new_n906));
  OR2_X1    g720(.A1(new_n895), .A2(new_n894), .ZN(new_n907));
  NAND4_X1  g721(.A1(new_n905), .A2(new_n906), .A3(new_n902), .A4(new_n907), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n884), .A2(new_n909), .ZN(new_n910));
  AOI22_X1  g724(.A1(new_n715), .A2(new_n724), .B1(new_n801), .B2(new_n802), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n700), .A2(new_n718), .A3(new_n813), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n722), .A2(new_n795), .ZN(new_n913));
  NOR3_X1   g727(.A1(new_n912), .A2(new_n733), .A3(new_n913), .ZN(new_n914));
  INV_X1    g728(.A(new_n758), .ZN(new_n915));
  AOI21_X1  g729(.A(new_n914), .B1(new_n715), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n911), .A2(new_n916), .A3(KEYINPUT52), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT52), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n803), .B1(new_n750), .B2(new_n723), .ZN(new_n919));
  INV_X1    g733(.A(new_n732), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n642), .A2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n913), .ZN(new_n922));
  NOR2_X1   g736(.A1(new_n817), .A2(new_n717), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n921), .A2(new_n922), .A3(new_n700), .A4(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(new_n750), .B2(new_n758), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n918), .B1(new_n919), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n917), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n798), .A2(new_n777), .A3(new_n772), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n766), .B(KEYINPUT109), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT115), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n738), .A2(new_n793), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n931), .B1(new_n932), .B2(new_n815), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n801), .A2(new_n819), .A3(KEYINPUT115), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g749(.A(new_n714), .ZN(new_n936));
  NOR3_X1   g750(.A1(new_n719), .A2(new_n818), .A3(new_n256), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n704), .A2(new_n936), .A3(new_n937), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n821), .A2(new_n935), .A3(new_n938), .A4(new_n824), .ZN(new_n939));
  OAI21_X1  g753(.A(new_n681), .B1(new_n257), .B2(new_n653), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n523), .A2(new_n431), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n663), .A2(new_n684), .A3(new_n940), .A4(new_n941), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n656), .B(new_n942), .C1(new_n705), .C2(new_n706), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n939), .A2(new_n943), .ZN(new_n944));
  AND4_X1   g758(.A1(KEYINPUT53), .A2(new_n927), .A3(new_n930), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n748), .A2(new_n749), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n713), .A2(new_n776), .A3(new_n654), .ZN(new_n947));
  OAI21_X1  g761(.A(new_n772), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n769), .A3(new_n798), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n950), .A2(new_n939), .A3(new_n943), .ZN(new_n951));
  AOI21_X1  g765(.A(KEYINPUT53), .B1(new_n951), .B2(new_n927), .ZN(new_n952));
  OAI21_X1  g766(.A(KEYINPUT54), .B1(new_n945), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(KEYINPUT116), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT53), .ZN(new_n955));
  AND2_X1   g769(.A1(new_n917), .A2(new_n926), .ZN(new_n956));
  AND4_X1   g770(.A1(new_n821), .A2(new_n935), .A3(new_n824), .A4(new_n938), .ZN(new_n957));
  INV_X1    g771(.A(new_n943), .ZN(new_n958));
  NAND3_X1  g772(.A1(new_n930), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n956), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT54), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n951), .A2(KEYINPUT53), .A3(new_n927), .ZN(new_n962));
  NAND3_X1  g776(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n953), .A2(new_n954), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n961), .B1(new_n960), .B2(new_n962), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT116), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n910), .B1(new_n964), .B2(new_n966), .ZN(new_n967));
  NOR2_X1   g781(.A1(G952), .A2(G953), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n863), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n969), .A2(KEYINPUT121), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT121), .ZN(new_n971));
  OAI211_X1 g785(.A(new_n971), .B(new_n863), .C1(new_n967), .C2(new_n968), .ZN(new_n972));
  NAND2_X1  g786(.A1(new_n970), .A2(new_n972), .ZN(G75));
  NAND2_X1  g787(.A1(new_n960), .A2(new_n962), .ZN(new_n974));
  NAND3_X1  g788(.A1(new_n974), .A2(G210), .A3(G902), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT56), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n471), .B1(new_n474), .B2(new_n475), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n977), .B(new_n445), .ZN(new_n978));
  XNOR2_X1  g792(.A(new_n978), .B(KEYINPUT55), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n975), .A2(new_n976), .A3(new_n979), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n979), .B1(new_n975), .B2(new_n976), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n338), .A2(G952), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n980), .A2(new_n981), .A3(new_n982), .ZN(G51));
  XOR2_X1   g797(.A(new_n807), .B(KEYINPUT57), .Z(new_n984));
  INV_X1    g798(.A(new_n963), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n984), .B1(new_n985), .B2(new_n965), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n359), .B2(new_n357), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n974), .A2(G902), .ZN(new_n988));
  OR2_X1    g802(.A1(new_n988), .A2(new_n827), .ZN(new_n989));
  AOI21_X1  g803(.A(new_n982), .B1(new_n987), .B2(new_n989), .ZN(G54));
  INV_X1    g804(.A(new_n419), .ZN(new_n991));
  NAND2_X1  g805(.A1(KEYINPUT58), .A2(G475), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n991), .B1(new_n988), .B2(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n993), .B1(G952), .B2(new_n338), .ZN(new_n994));
  NOR3_X1   g808(.A1(new_n988), .A2(new_n991), .A3(new_n992), .ZN(new_n995));
  NOR2_X1   g809(.A1(new_n994), .A2(new_n995), .ZN(G60));
  AND2_X1   g810(.A1(new_n674), .A2(new_n676), .ZN(new_n997));
  NAND2_X1  g811(.A1(G478), .A2(G902), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n998), .B(KEYINPUT59), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  AOI21_X1  g814(.A(new_n1000), .B1(new_n953), .B2(new_n963), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n964), .A2(new_n966), .A3(new_n999), .ZN(new_n1002));
  INV_X1    g816(.A(new_n997), .ZN(new_n1003));
  AOI211_X1 g817(.A(new_n982), .B(new_n1001), .C1(new_n1002), .C2(new_n1003), .ZN(G63));
  NAND2_X1  g818(.A1(G217), .A2(G902), .ZN(new_n1005));
  XOR2_X1   g819(.A(new_n1005), .B(KEYINPUT60), .Z(new_n1006));
  OAI21_X1  g820(.A(new_n1006), .B1(new_n945), .B2(new_n952), .ZN(new_n1007));
  OR2_X1    g821(.A1(new_n1007), .A2(new_n698), .ZN(new_n1008));
  INV_X1    g822(.A(new_n571), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n982), .B1(new_n1007), .B2(new_n1009), .ZN(new_n1010));
  AOI22_X1  g824(.A1(new_n1008), .A2(new_n1010), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n1011));
  NOR2_X1   g825(.A1(KEYINPUT122), .A2(KEYINPUT61), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1011), .B(new_n1012), .ZN(G66));
  INV_X1    g827(.A(new_n430), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n338), .B1(new_n1014), .B2(G224), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n930), .A2(new_n958), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(new_n1016), .B2(new_n338), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n977), .B1(G898), .B2(new_n338), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1017), .B(new_n1018), .Z(G69));
  INV_X1    g833(.A(KEYINPUT123), .ZN(new_n1020));
  NOR2_X1   g834(.A1(new_n919), .A2(new_n759), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n746), .A2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g836(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1023));
  NAND4_X1  g837(.A1(new_n743), .A2(new_n651), .A3(new_n814), .A4(new_n940), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n846), .A2(new_n854), .A3(new_n1024), .ZN(new_n1025));
  NOR2_X1   g839(.A1(new_n1023), .A2(new_n1025), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1022), .A2(KEYINPUT62), .ZN(new_n1027));
  AOI21_X1  g841(.A(G953), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  XNOR2_X1  g842(.A(new_n620), .B(new_n415), .ZN(new_n1029));
  INV_X1    g843(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n1020), .B1(new_n1028), .B2(new_n1030), .ZN(new_n1031));
  AND2_X1   g845(.A1(new_n846), .A2(new_n854), .ZN(new_n1032));
  OAI211_X1 g846(.A(new_n1032), .B(new_n1024), .C1(KEYINPUT62), .C2(new_n1022), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1027), .ZN(new_n1034));
  OAI21_X1  g848(.A(new_n338), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NAND3_X1  g849(.A1(new_n1035), .A2(KEYINPUT123), .A3(new_n1029), .ZN(new_n1036));
  AOI21_X1  g850(.A(new_n338), .B1(G227), .B2(G900), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n720), .A2(new_n823), .ZN(new_n1038));
  NAND2_X1  g852(.A1(new_n922), .A2(new_n741), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1038), .B1(new_n849), .B2(new_n1039), .ZN(new_n1040));
  AOI22_X1  g854(.A1(new_n1040), .A2(new_n651), .B1(new_n816), .B2(new_n820), .ZN(new_n1041));
  NAND4_X1  g855(.A1(new_n1032), .A2(new_n338), .A3(new_n1021), .A4(new_n1041), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1029), .B1(G900), .B2(G953), .ZN(new_n1043));
  AOI21_X1  g857(.A(new_n1037), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g858(.A1(new_n1031), .A2(new_n1036), .A3(new_n1044), .ZN(new_n1045));
  AND3_X1   g859(.A1(new_n1042), .A2(KEYINPUT124), .A3(new_n1043), .ZN(new_n1046));
  AOI21_X1  g860(.A(KEYINPUT124), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1047));
  NOR2_X1   g861(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1031), .A2(new_n1048), .A3(new_n1036), .ZN(new_n1049));
  INV_X1    g863(.A(KEYINPUT125), .ZN(new_n1050));
  AND3_X1   g864(.A1(new_n1049), .A2(new_n1050), .A3(new_n1037), .ZN(new_n1051));
  AOI21_X1  g865(.A(new_n1050), .B1(new_n1049), .B2(new_n1037), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1045), .B1(new_n1051), .B2(new_n1052), .ZN(G72));
  NAND2_X1  g867(.A1(G472), .A2(G902), .ZN(new_n1054));
  XOR2_X1   g868(.A(new_n1054), .B(KEYINPUT63), .Z(new_n1055));
  NAND2_X1  g869(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1056));
  OAI21_X1  g870(.A(new_n1055), .B1(new_n1056), .B2(new_n1016), .ZN(new_n1057));
  NAND2_X1  g871(.A1(new_n1057), .A2(new_n727), .ZN(new_n1058));
  NAND3_X1  g872(.A1(new_n1032), .A2(new_n1021), .A3(new_n1041), .ZN(new_n1059));
  OAI21_X1  g873(.A(new_n1055), .B1(new_n1059), .B2(new_n1016), .ZN(new_n1060));
  AOI21_X1  g874(.A(new_n728), .B1(new_n620), .B2(new_n455), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n982), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1058), .A2(new_n1062), .ZN(new_n1063));
  INV_X1    g877(.A(new_n727), .ZN(new_n1064));
  INV_X1    g878(.A(new_n1061), .ZN(new_n1065));
  NAND4_X1  g879(.A1(new_n974), .A2(new_n1064), .A3(new_n1055), .A4(new_n1065), .ZN(new_n1066));
  INV_X1    g880(.A(KEYINPUT126), .ZN(new_n1067));
  OR2_X1    g881(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g882(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1069));
  AOI21_X1  g883(.A(new_n1063), .B1(new_n1068), .B2(new_n1069), .ZN(G57));
endmodule


