//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 1 0 0 1 1 1 1 0 0 0 1 1 0 0 0 1 0 1 0 1 0 0 0 0 1 0 1 0 1 0 1 0 0 1 0 0 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n710, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993;
  INV_X1    g000(.A(KEYINPUT15), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G478), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  INV_X1    g003(.A(G128), .ZN(new_n190));
  NOR2_X1   g004(.A1(new_n190), .A2(G143), .ZN(new_n191));
  INV_X1    g005(.A(KEYINPUT13), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n189), .B1(new_n191), .B2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT93), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G128), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(G143), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(KEYINPUT13), .ZN(new_n198));
  AND3_X1   g012(.A1(new_n193), .A2(new_n194), .A3(new_n198), .ZN(new_n199));
  AOI21_X1  g013(.A(new_n194), .B1(new_n193), .B2(new_n198), .ZN(new_n200));
  XNOR2_X1  g014(.A(G128), .B(G143), .ZN(new_n201));
  AND2_X1   g015(.A1(new_n201), .A2(new_n189), .ZN(new_n202));
  NOR3_X1   g016(.A1(new_n199), .A2(new_n200), .A3(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G116), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(KEYINPUT67), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT67), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G116), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n205), .A2(new_n207), .A3(G122), .ZN(new_n208));
  INV_X1    g022(.A(G122), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G116), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G107), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n208), .A2(new_n213), .A3(new_n210), .ZN(new_n214));
  AND3_X1   g028(.A1(new_n212), .A2(KEYINPUT92), .A3(new_n214), .ZN(new_n215));
  AOI21_X1  g029(.A(KEYINPUT92), .B1(new_n212), .B2(new_n214), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n203), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n201), .A2(new_n189), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n211), .A2(KEYINPUT14), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT14), .ZN(new_n220));
  OAI21_X1  g034(.A(G107), .B1(new_n208), .B2(new_n220), .ZN(new_n221));
  OAI221_X1 g035(.A(new_n214), .B1(new_n202), .B2(new_n218), .C1(new_n219), .C2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT9), .B(G234), .ZN(new_n223));
  INV_X1    g037(.A(G217), .ZN(new_n224));
  NOR3_X1   g038(.A1(new_n223), .A2(new_n224), .A3(G953), .ZN(new_n225));
  NAND3_X1  g039(.A1(new_n217), .A2(new_n222), .A3(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT94), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT94), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n217), .A2(new_n222), .A3(new_n228), .A4(new_n225), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n217), .A2(new_n222), .ZN(new_n230));
  INV_X1    g044(.A(new_n225), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n227), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(G902), .ZN(new_n234));
  AND3_X1   g048(.A1(new_n233), .A2(KEYINPUT95), .A3(new_n234), .ZN(new_n235));
  AOI21_X1  g049(.A(KEYINPUT95), .B1(new_n233), .B2(new_n234), .ZN(new_n236));
  OAI21_X1  g050(.A(new_n188), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n234), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT95), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n187), .B(G478), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n237), .A2(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(G952), .ZN(new_n242));
  OR2_X1    g056(.A1(new_n242), .A2(KEYINPUT96), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(KEYINPUT96), .ZN(new_n244));
  AOI21_X1  g058(.A(G953), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(G234), .ZN(new_n246));
  INV_X1    g060(.A(G237), .ZN(new_n247));
  OAI21_X1  g061(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(new_n248), .B(KEYINPUT97), .ZN(new_n249));
  OR2_X1    g063(.A1(KEYINPUT70), .A2(G953), .ZN(new_n250));
  NAND2_X1  g064(.A1(KEYINPUT70), .A2(G953), .ZN(new_n251));
  AND2_X1   g065(.A1(new_n250), .A2(new_n251), .ZN(new_n252));
  AOI211_X1 g066(.A(new_n234), .B(new_n252), .C1(G234), .C2(G237), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT21), .B(G898), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(G475), .A2(G902), .ZN(new_n257));
  XNOR2_X1  g071(.A(G113), .B(G122), .ZN(new_n258));
  INV_X1    g072(.A(G104), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n250), .A2(G214), .A3(new_n247), .A4(new_n251), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(new_n195), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g077(.A1(new_n261), .A2(new_n195), .ZN(new_n264));
  OAI211_X1 g078(.A(KEYINPUT18), .B(G131), .C1(new_n263), .C2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(G125), .B(G140), .ZN(new_n266));
  INV_X1    g080(.A(G146), .ZN(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(new_n264), .ZN(new_n269));
  NAND2_X1  g083(.A1(KEYINPUT18), .A2(G131), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n269), .A2(new_n262), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n265), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(G131), .B1(new_n263), .B2(new_n264), .ZN(new_n273));
  INV_X1    g087(.A(G131), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n269), .A2(new_n274), .A3(new_n262), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT17), .ZN(new_n276));
  AND3_X1   g090(.A1(new_n273), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  OAI211_X1 g091(.A(KEYINPUT17), .B(G131), .C1(new_n263), .C2(new_n264), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  NOR3_X1   g093(.A1(new_n279), .A2(KEYINPUT16), .A3(G140), .ZN(new_n280));
  OR2_X1    g094(.A1(new_n280), .A2(KEYINPUT74), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n280), .B1(new_n266), .B2(KEYINPUT16), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT74), .ZN(new_n283));
  OAI21_X1  g097(.A(new_n281), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n284), .A2(new_n267), .ZN(new_n285));
  OAI211_X1 g099(.A(G146), .B(new_n281), .C1(new_n282), .C2(new_n283), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n278), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n260), .B(new_n272), .C1(new_n277), .C2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(KEYINPUT90), .A2(KEYINPUT19), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n266), .A2(new_n290), .ZN(new_n291));
  XOR2_X1   g105(.A(KEYINPUT90), .B(KEYINPUT19), .Z(new_n292));
  OAI211_X1 g106(.A(new_n291), .B(new_n267), .C1(new_n266), .C2(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n286), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT91), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n273), .A2(new_n275), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n286), .A2(KEYINPUT91), .A3(new_n293), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n260), .B1(new_n299), .B2(new_n272), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n257), .B1(new_n289), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(KEYINPUT20), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT20), .ZN(new_n303));
  OAI211_X1 g117(.A(new_n303), .B(new_n257), .C1(new_n289), .C2(new_n300), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n302), .A2(new_n304), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n272), .B1(new_n277), .B2(new_n287), .ZN(new_n306));
  INV_X1    g120(.A(new_n260), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n288), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n309), .A2(new_n234), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(G475), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n305), .A2(new_n311), .ZN(new_n312));
  NOR3_X1   g126(.A1(new_n241), .A2(new_n256), .A3(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(G214), .B1(G237), .B2(G902), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n267), .A2(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n195), .A2(G146), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  NOR3_X1   g131(.A1(new_n317), .A2(KEYINPUT1), .A3(new_n190), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n195), .A2(KEYINPUT1), .A3(G146), .ZN(new_n319));
  XNOR2_X1  g133(.A(G143), .B(G146), .ZN(new_n320));
  OAI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(G128), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT66), .ZN(new_n322));
  NAND2_X1  g136(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n317), .A2(new_n190), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n324), .A2(KEYINPUT66), .A3(new_n319), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n318), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n279), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n320), .A2(KEYINPUT0), .A3(G128), .ZN(new_n328));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G128), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n328), .B1(new_n320), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n330), .A2(G125), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(G224), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(G953), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n332), .B(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT80), .B(G104), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT3), .B1(new_n336), .B2(G107), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n259), .A2(KEYINPUT3), .A3(G107), .ZN(new_n338));
  AOI21_X1  g152(.A(new_n338), .B1(new_n336), .B2(G107), .ZN(new_n339));
  INV_X1    g153(.A(G101), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n337), .A2(new_n339), .A3(new_n340), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT81), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n342), .B1(new_n259), .B2(G107), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n343), .B1(new_n336), .B2(G107), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n259), .A2(KEYINPUT80), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n259), .A2(KEYINPUT80), .ZN(new_n346));
  OAI211_X1 g160(.A(new_n342), .B(new_n213), .C1(new_n345), .C2(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n344), .A2(G101), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n341), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT84), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  XOR2_X1   g165(.A(KEYINPUT2), .B(G113), .Z(new_n352));
  NAND3_X1  g166(.A1(new_n205), .A2(new_n207), .A3(G119), .ZN(new_n353));
  INV_X1    g167(.A(G119), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n354), .A2(G116), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n353), .A3(new_n355), .ZN(new_n356));
  AND3_X1   g170(.A1(new_n353), .A2(KEYINPUT5), .A3(new_n355), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT86), .ZN(new_n358));
  OAI21_X1  g172(.A(new_n358), .B1(new_n355), .B2(KEYINPUT5), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n204), .A2(G119), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT5), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n360), .A2(KEYINPUT86), .A3(new_n361), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n359), .A2(new_n362), .A3(G113), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n356), .B1(new_n357), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(new_n364), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n341), .A2(new_n348), .A3(KEYINPUT84), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n351), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XNOR2_X1  g181(.A(G110), .B(G122), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n340), .B1(new_n337), .B2(new_n339), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT4), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT67), .B(G116), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n360), .B1(new_n372), .B2(G119), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n373), .B(new_n352), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n341), .A2(KEYINPUT4), .ZN(new_n375));
  OAI211_X1 g189(.A(new_n371), .B(new_n374), .C1(new_n375), .C2(new_n369), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n367), .A2(new_n368), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n367), .A2(new_n376), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n368), .A2(KEYINPUT87), .ZN(new_n379));
  AOI22_X1  g193(.A1(new_n377), .A2(KEYINPUT6), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AND3_X1   g194(.A1(new_n378), .A2(KEYINPUT6), .A3(new_n379), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n335), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n368), .B(KEYINPUT8), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n349), .A2(new_n364), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT88), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n349), .A2(new_n364), .A3(KEYINPUT88), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n386), .A2(new_n387), .ZN(new_n388));
  AND3_X1   g202(.A1(new_n341), .A2(new_n348), .A3(KEYINPUT84), .ZN(new_n389));
  AOI21_X1  g203(.A(KEYINPUT84), .B1(new_n341), .B2(new_n348), .ZN(new_n390));
  NOR3_X1   g204(.A1(new_n389), .A2(new_n390), .A3(new_n364), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n383), .B1(new_n388), .B2(new_n391), .ZN(new_n392));
  OAI21_X1  g206(.A(KEYINPUT7), .B1(new_n333), .B2(G953), .ZN(new_n393));
  INV_X1    g207(.A(new_n393), .ZN(new_n394));
  AND3_X1   g208(.A1(new_n327), .A2(new_n331), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n394), .B1(new_n327), .B2(new_n331), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n392), .A2(KEYINPUT89), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(new_n377), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT89), .B1(new_n392), .B2(new_n397), .ZN(new_n400));
  OAI211_X1 g214(.A(new_n382), .B(new_n234), .C1(new_n399), .C2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(G210), .B1(G237), .B2(G902), .ZN(new_n402));
  INV_X1    g216(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(KEYINPUT89), .ZN(new_n405));
  INV_X1    g219(.A(new_n383), .ZN(new_n406));
  AND3_X1   g220(.A1(new_n349), .A2(KEYINPUT88), .A3(new_n364), .ZN(new_n407));
  AOI21_X1  g221(.A(KEYINPUT88), .B1(new_n349), .B2(new_n364), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n406), .B1(new_n409), .B2(new_n367), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n332), .A2(new_n393), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n327), .A2(new_n331), .A3(new_n394), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n405), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(new_n377), .A3(new_n398), .ZN(new_n415));
  NAND4_X1  g229(.A1(new_n415), .A2(new_n234), .A3(new_n402), .A4(new_n382), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n404), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n313), .A2(new_n314), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n252), .A2(G210), .A3(new_n247), .ZN(new_n419));
  XNOR2_X1  g233(.A(KEYINPUT26), .B(G101), .ZN(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  XNOR2_X1  g235(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n421), .B(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(G137), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n424), .A2(G134), .ZN(new_n425));
  OAI21_X1  g239(.A(KEYINPUT11), .B1(new_n189), .B2(G137), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT11), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n427), .A2(new_n424), .A3(G134), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n425), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n429), .A2(new_n274), .ZN(new_n430));
  INV_X1    g244(.A(new_n425), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(G134), .B2(new_n424), .ZN(new_n432));
  NOR3_X1   g246(.A1(new_n189), .A2(KEYINPUT11), .A3(G137), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n274), .B(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT64), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n429), .A2(KEYINPUT64), .A3(new_n274), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n430), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT68), .B1(new_n438), .B2(new_n330), .ZN(new_n439));
  OR2_X1    g253(.A1(new_n429), .A2(new_n274), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n426), .A2(new_n428), .ZN(new_n441));
  AND4_X1   g255(.A1(KEYINPUT64), .A2(new_n441), .A3(new_n274), .A4(new_n431), .ZN(new_n442));
  AOI21_X1  g256(.A(KEYINPUT64), .B1(new_n429), .B2(new_n274), .ZN(new_n443));
  OAI21_X1  g257(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT68), .ZN(new_n445));
  INV_X1    g259(.A(new_n330), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n444), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n439), .A2(new_n447), .ZN(new_n448));
  OAI21_X1  g262(.A(KEYINPUT65), .B1(new_n424), .B2(G134), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT65), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n450), .A2(new_n189), .A3(G137), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n424), .A2(G134), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n449), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G131), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n442), .B2(new_n443), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n455), .A2(KEYINPUT69), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n453), .A2(G131), .ZN(new_n457));
  AOI21_X1  g271(.A(new_n457), .B1(new_n436), .B2(new_n437), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n318), .ZN(new_n461));
  AOI21_X1  g275(.A(KEYINPUT66), .B1(new_n324), .B2(new_n319), .ZN(new_n462));
  AOI21_X1  g276(.A(G128), .B1(new_n315), .B2(new_n316), .ZN(new_n463));
  INV_X1    g277(.A(new_n319), .ZN(new_n464));
  NOR3_X1   g278(.A1(new_n463), .A2(new_n464), .A3(new_n322), .ZN(new_n465));
  OAI21_X1  g279(.A(new_n461), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n456), .A2(new_n460), .A3(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(new_n374), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n448), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n444), .A2(new_n446), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n458), .A2(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n472), .A2(new_n374), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n469), .A2(new_n473), .ZN(new_n474));
  XOR2_X1   g288(.A(KEYINPUT72), .B(KEYINPUT28), .Z(new_n475));
  NAND2_X1  g289(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n374), .B1(new_n444), .B2(new_n446), .ZN(new_n477));
  AOI21_X1  g291(.A(KEYINPUT28), .B1(new_n467), .B2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n478), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n423), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n469), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT30), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n470), .A2(new_n471), .A3(new_n483), .ZN(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n326), .B1(new_n455), .B2(KEYINPUT69), .ZN(new_n486));
  AOI22_X1  g300(.A1(new_n460), .A2(new_n486), .B1(new_n439), .B2(new_n447), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n485), .B1(new_n487), .B2(new_n483), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n482), .B1(new_n488), .B2(new_n374), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT31), .B1(new_n489), .B2(new_n423), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n483), .B1(new_n448), .B2(new_n467), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n374), .B1(new_n491), .B2(new_n484), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n492), .A2(KEYINPUT31), .A3(new_n423), .A4(new_n469), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n481), .B1(new_n490), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(G472), .A2(G902), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n495), .A2(KEYINPUT32), .A3(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT73), .B(KEYINPUT32), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n438), .A2(KEYINPUT68), .A3(new_n330), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n445), .B1(new_n444), .B2(new_n446), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n466), .B1(new_n458), .B2(new_n459), .ZN(new_n501));
  AOI211_X1 g315(.A(KEYINPUT69), .B(new_n457), .C1(new_n436), .C2(new_n437), .ZN(new_n502));
  OAI22_X1  g316(.A1(new_n499), .A2(new_n500), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  AOI21_X1  g317(.A(new_n484), .B1(new_n503), .B2(KEYINPUT30), .ZN(new_n504));
  OAI211_X1 g318(.A(new_n423), .B(new_n469), .C1(new_n504), .C2(new_n468), .ZN(new_n505));
  INV_X1    g319(.A(KEYINPUT31), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n480), .B1(new_n507), .B2(new_n493), .ZN(new_n508));
  INV_X1    g322(.A(new_n496), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n498), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n423), .B1(new_n492), .B2(new_n469), .ZN(new_n511));
  INV_X1    g325(.A(new_n475), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n512), .B1(new_n469), .B2(new_n473), .ZN(new_n513));
  INV_X1    g327(.A(new_n423), .ZN(new_n514));
  NOR3_X1   g328(.A1(new_n513), .A2(new_n514), .A3(new_n478), .ZN(new_n515));
  NOR3_X1   g329(.A1(new_n511), .A2(new_n515), .A3(KEYINPUT29), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n503), .A2(new_n374), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n517), .A2(new_n469), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(KEYINPUT28), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n423), .A2(KEYINPUT29), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(new_n479), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n521), .A2(new_n234), .ZN(new_n522));
  OAI21_X1  g336(.A(G472), .B1(new_n516), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n497), .A2(new_n510), .A3(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n285), .A2(new_n286), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT23), .ZN(new_n526));
  OAI21_X1  g340(.A(new_n526), .B1(new_n354), .B2(G128), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n190), .A2(KEYINPUT23), .A3(G119), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n527), .B(new_n528), .C1(G119), .C2(new_n190), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G110), .ZN(new_n530));
  XOR2_X1   g344(.A(KEYINPUT24), .B(G110), .Z(new_n531));
  XNOR2_X1  g345(.A(G119), .B(G128), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n530), .A2(new_n533), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n525), .A2(new_n534), .ZN(new_n535));
  OAI22_X1  g349(.A1(new_n529), .A2(G110), .B1(new_n532), .B2(new_n531), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT75), .ZN(new_n537));
  XNOR2_X1  g351(.A(new_n536), .B(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n266), .A2(new_n267), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n286), .A2(new_n539), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n252), .A2(G221), .A3(G234), .ZN(new_n543));
  XNOR2_X1  g357(.A(KEYINPUT22), .B(G137), .ZN(new_n544));
  XNOR2_X1  g358(.A(new_n543), .B(new_n544), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n535), .A2(new_n542), .A3(new_n545), .ZN(new_n546));
  INV_X1    g360(.A(new_n545), .ZN(new_n547));
  NOR2_X1   g361(.A1(new_n525), .A2(new_n534), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n547), .B1(new_n548), .B2(new_n541), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n224), .B1(G234), .B2(new_n234), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n551), .A2(new_n234), .ZN(new_n552));
  XNOR2_X1  g366(.A(new_n552), .B(KEYINPUT77), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n546), .A2(new_n549), .A3(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(new_n555), .B(KEYINPUT78), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n546), .A2(new_n549), .A3(new_n234), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT25), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT76), .ZN(new_n559));
  INV_X1    g373(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n546), .A2(new_n549), .A3(new_n234), .A4(new_n559), .ZN(new_n562));
  AOI21_X1  g376(.A(new_n551), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g377(.A1(new_n556), .A2(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(G221), .B1(new_n223), .B2(G902), .ZN(new_n565));
  INV_X1    g379(.A(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G469), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(new_n234), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n466), .B1(new_n351), .B2(new_n366), .ZN(new_n569));
  OR3_X1    g383(.A1(new_n463), .A2(KEYINPUT82), .A3(new_n464), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n321), .A2(KEYINPUT82), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n461), .A3(new_n571), .ZN(new_n572));
  NAND3_X1  g386(.A1(new_n572), .A2(new_n341), .A3(new_n348), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  OAI211_X1 g388(.A(KEYINPUT12), .B(new_n444), .C1(new_n569), .C2(new_n574), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(KEYINPUT85), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n326), .B1(new_n389), .B2(new_n390), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n438), .B1(new_n577), .B2(new_n573), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT85), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(KEYINPUT12), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n444), .B1(new_n569), .B2(new_n574), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT12), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(new_n580), .A3(new_n583), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n351), .A2(KEYINPUT10), .A3(new_n466), .A4(new_n366), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT83), .B(KEYINPUT10), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n573), .A2(new_n586), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n371), .B(new_n446), .C1(new_n375), .C2(new_n369), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n585), .A2(new_n587), .A3(new_n438), .A4(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(new_n252), .ZN(new_n590));
  INV_X1    g404(.A(G227), .ZN(new_n591));
  NOR2_X1   g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g406(.A(G110), .B(G140), .ZN(new_n593));
  XNOR2_X1  g407(.A(new_n593), .B(KEYINPUT79), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n592), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  INV_X1    g410(.A(new_n596), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n584), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n585), .A2(new_n587), .A3(new_n588), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n444), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(new_n589), .ZN(new_n601));
  INV_X1    g415(.A(new_n595), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(G902), .B1(new_n598), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n568), .B1(new_n604), .B2(new_n567), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n584), .A2(new_n589), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n602), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n597), .A2(new_n600), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n607), .A2(G469), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n566), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  NAND4_X1  g424(.A1(new_n418), .A2(new_n524), .A3(new_n564), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(G101), .ZN(G3));
  INV_X1    g426(.A(KEYINPUT98), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n314), .B1(new_n416), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT99), .ZN(new_n616));
  NAND3_X1  g430(.A1(new_n404), .A2(new_n613), .A3(new_n416), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  NOR3_X1   g433(.A1(new_n618), .A2(new_n619), .A3(new_n256), .ZN(new_n620));
  INV_X1    g434(.A(new_n620), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n232), .A2(KEYINPUT33), .A3(new_n226), .ZN(new_n622));
  INV_X1    g436(.A(G478), .ZN(new_n623));
  NOR2_X1   g437(.A1(new_n623), .A2(G902), .ZN(new_n624));
  AND3_X1   g438(.A1(new_n227), .A2(new_n229), .A3(new_n232), .ZN(new_n625));
  OAI211_X1 g439(.A(new_n622), .B(new_n624), .C1(new_n625), .C2(KEYINPUT33), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n238), .A2(new_n623), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n312), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n621), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n604), .A2(new_n567), .ZN(new_n631));
  INV_X1    g445(.A(new_n568), .ZN(new_n632));
  NAND3_X1  g446(.A1(new_n631), .A2(new_n632), .A3(new_n609), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n633), .A2(new_n565), .ZN(new_n634));
  OAI21_X1  g448(.A(G472), .B1(new_n508), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n495), .A2(new_n496), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g451(.A(new_n564), .ZN(new_n638));
  NOR3_X1   g452(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n630), .A2(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT34), .B(G104), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G6));
  AOI21_X1  g456(.A(new_n312), .B1(new_n237), .B2(new_n240), .ZN(new_n643));
  AND2_X1   g457(.A1(new_n620), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n644), .A2(new_n639), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT35), .B(G107), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G9));
  INV_X1    g461(.A(new_n637), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n561), .A2(new_n562), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n550), .ZN(new_n650));
  INV_X1    g464(.A(KEYINPUT36), .ZN(new_n651));
  OR3_X1    g465(.A1(new_n548), .A2(new_n541), .A3(KEYINPUT100), .ZN(new_n652));
  OAI21_X1  g466(.A(KEYINPUT100), .B1(new_n548), .B2(new_n541), .ZN(new_n653));
  AND4_X1   g467(.A1(new_n651), .A2(new_n652), .A3(new_n545), .A4(new_n653), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n652), .A2(new_n653), .B1(new_n651), .B2(new_n545), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n554), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n650), .A2(new_n656), .ZN(new_n657));
  NAND4_X1  g471(.A1(new_n418), .A2(new_n610), .A3(new_n648), .A4(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(KEYINPUT37), .B(G110), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n658), .B(new_n659), .ZN(G12));
  AND3_X1   g474(.A1(new_n524), .A2(new_n610), .A3(new_n657), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n618), .A2(new_n619), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT101), .B(G900), .Z(new_n663));
  NAND2_X1  g477(.A1(new_n253), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g478(.A1(new_n249), .A2(new_n664), .ZN(new_n665));
  INV_X1    g479(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n643), .A2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n661), .A2(new_n662), .A3(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G128), .ZN(G30));
  NAND2_X1  g484(.A1(new_n241), .A2(new_n312), .ZN(new_n671));
  INV_X1    g485(.A(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n314), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n657), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n672), .A2(new_n674), .ZN(new_n675));
  INV_X1    g489(.A(new_n675), .ZN(new_n676));
  OR2_X1    g490(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n417), .B(KEYINPUT38), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n676), .A2(KEYINPUT102), .ZN(new_n679));
  AND3_X1   g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  XOR2_X1   g494(.A(new_n665), .B(KEYINPUT39), .Z(new_n681));
  NAND2_X1  g495(.A1(new_n610), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g496(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n682), .A2(KEYINPUT40), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n518), .A2(new_n514), .ZN(new_n685));
  AND2_X1   g499(.A1(new_n505), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g500(.A(G472), .B1(new_n686), .B2(G902), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n497), .A2(new_n510), .A3(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n680), .A2(new_n683), .A3(new_n684), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  NOR2_X1   g504(.A1(new_n629), .A2(new_n665), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n661), .A2(new_n662), .A3(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G146), .ZN(G48));
  NAND2_X1  g507(.A1(new_n524), .A2(new_n564), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n598), .A2(new_n603), .ZN(new_n695));
  INV_X1    g509(.A(KEYINPUT103), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n695), .A2(new_n696), .A3(new_n234), .ZN(new_n697));
  AOI22_X1  g511(.A1(new_n584), .A2(new_n597), .B1(new_n602), .B2(new_n601), .ZN(new_n698));
  OAI21_X1  g512(.A(KEYINPUT103), .B1(new_n698), .B2(G902), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n697), .A2(new_n699), .A3(G469), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT104), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n566), .B1(new_n604), .B2(new_n567), .ZN(new_n702));
  AND3_X1   g516(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n700), .B2(new_n702), .ZN(new_n704));
  NOR3_X1   g518(.A1(new_n694), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AND2_X1   g519(.A1(new_n630), .A2(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(KEYINPUT41), .B(G113), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT105), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n706), .B(new_n708), .ZN(G15));
  AND2_X1   g523(.A1(new_n644), .A2(new_n705), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(new_n204), .ZN(G18));
  NAND3_X1  g525(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n712));
  OAI21_X1  g526(.A(G469), .B1(new_n604), .B2(new_n696), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n698), .A2(KEYINPUT103), .A3(G902), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n702), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT104), .ZN(new_n716));
  AND3_X1   g530(.A1(new_n404), .A2(new_n613), .A3(new_n416), .ZN(new_n717));
  OAI21_X1  g531(.A(KEYINPUT99), .B1(new_n717), .B2(new_n614), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n719));
  AND4_X1   g533(.A1(new_n712), .A2(new_n716), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  AND3_X1   g534(.A1(new_n524), .A2(new_n313), .A3(new_n657), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  XOR2_X1   g536(.A(KEYINPUT106), .B(G119), .Z(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G21));
  NOR2_X1   g538(.A1(new_n490), .A2(new_n494), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n423), .B1(new_n519), .B2(new_n479), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n496), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n256), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n727), .A2(new_n635), .A3(new_n564), .A4(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n703), .A2(new_n729), .A3(new_n704), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n618), .A2(new_n619), .A3(new_n671), .ZN(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G122), .ZN(G24));
  AND4_X1   g547(.A1(new_n635), .A2(new_n691), .A3(new_n727), .A4(new_n657), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n662), .A2(new_n719), .A3(new_n716), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  NAND3_X1  g550(.A1(new_n597), .A2(KEYINPUT107), .A3(new_n600), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT107), .ZN(new_n738));
  INV_X1    g552(.A(new_n600), .ZN(new_n739));
  OAI21_X1  g553(.A(new_n738), .B1(new_n739), .B2(new_n596), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n737), .A2(new_n740), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n741), .A2(G469), .A3(new_n607), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n605), .A2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(new_n417), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n566), .A2(new_n673), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n743), .A2(new_n744), .A3(new_n745), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n691), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n748), .A2(KEYINPUT42), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n747), .A2(new_n749), .A3(new_n524), .A4(new_n564), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT32), .ZN(new_n751));
  OAI21_X1  g565(.A(new_n751), .B1(new_n508), .B2(new_n509), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n497), .A2(new_n752), .A3(new_n523), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n753), .A2(new_n564), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n743), .A2(new_n744), .A3(new_n691), .A4(new_n745), .ZN(new_n755));
  OAI21_X1  g569(.A(KEYINPUT42), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n750), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(new_n274), .ZN(G33));
  NAND4_X1  g572(.A1(new_n747), .A2(new_n668), .A3(new_n524), .A4(new_n564), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G134), .ZN(G36));
  NAND3_X1  g574(.A1(new_n404), .A2(new_n314), .A3(new_n416), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT43), .ZN(new_n762));
  OAI21_X1  g576(.A(new_n762), .B1(new_n312), .B2(KEYINPUT109), .ZN(new_n763));
  AOI22_X1  g577(.A1(new_n302), .A2(new_n304), .B1(new_n310), .B2(G475), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n628), .A2(new_n764), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n763), .B(new_n765), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n766), .A2(new_n637), .A3(new_n657), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT44), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n761), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  OAI21_X1  g583(.A(new_n769), .B1(new_n768), .B2(new_n767), .ZN(new_n770));
  XOR2_X1   g584(.A(new_n770), .B(KEYINPUT110), .Z(new_n771));
  AND2_X1   g585(.A1(new_n607), .A2(new_n608), .ZN(new_n772));
  OAI21_X1  g586(.A(G469), .B1(new_n772), .B2(KEYINPUT45), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  AND3_X1   g588(.A1(new_n741), .A2(KEYINPUT45), .A3(new_n607), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n775), .B1(new_n773), .B2(KEYINPUT108), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n568), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  AND2_X1   g591(.A1(new_n777), .A2(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n631), .B1(new_n777), .B2(KEYINPUT46), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n565), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n781), .A2(new_n681), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n771), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n424), .ZN(G39));
  OR4_X1    g598(.A1(new_n524), .A2(new_n748), .A3(new_n564), .A4(new_n761), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n785), .B(KEYINPUT111), .Z(new_n786));
  NAND2_X1  g600(.A1(new_n781), .A2(KEYINPUT47), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT47), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n780), .A2(new_n788), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n786), .B1(new_n787), .B2(new_n789), .ZN(new_n790));
  XOR2_X1   g604(.A(new_n790), .B(G140), .Z(G42));
  NAND2_X1  g605(.A1(new_n700), .A2(new_n631), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n792), .A2(KEYINPUT49), .ZN(new_n793));
  NAND4_X1  g607(.A1(new_n793), .A2(new_n564), .A3(new_n745), .A4(new_n765), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(KEYINPUT112), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n678), .A2(new_n688), .ZN(new_n796));
  OAI211_X1 g610(.A(new_n795), .B(new_n796), .C1(KEYINPUT49), .C2(new_n792), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT54), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT52), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n735), .A2(new_n669), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n665), .A2(new_n566), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n650), .A2(new_n656), .A3(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n605), .B2(new_n742), .ZN(new_n803));
  AND2_X1   g617(.A1(new_n688), .A2(new_n803), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n662), .A2(new_n804), .A3(new_n672), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n692), .A2(new_n805), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n799), .B1(new_n800), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n718), .A2(new_n712), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n524), .A2(new_n610), .A3(new_n657), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  AOI22_X1  g624(.A1(new_n810), .A2(new_n691), .B1(new_n731), .B2(new_n804), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n811), .A2(KEYINPUT52), .A3(new_n669), .A4(new_n735), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n807), .A2(new_n812), .A3(KEYINPUT114), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT114), .ZN(new_n814));
  OAI211_X1 g628(.A(new_n814), .B(new_n799), .C1(new_n800), .C2(new_n806), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n720), .A2(new_n721), .B1(new_n730), .B2(new_n731), .ZN(new_n816));
  INV_X1    g630(.A(new_n629), .ZN(new_n817));
  OAI211_X1 g631(.A(new_n705), .B(new_n620), .C1(new_n817), .C2(new_n643), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n643), .A2(new_n817), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n417), .A2(new_n728), .A3(new_n314), .ZN(new_n820));
  NOR2_X1   g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n821), .A2(new_n564), .A3(new_n610), .A4(new_n648), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n611), .A3(new_n658), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n816), .A2(new_n818), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n237), .A2(new_n764), .A3(new_n240), .A4(new_n666), .ZN(new_n825));
  INV_X1    g639(.A(new_n825), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n744), .A2(KEYINPUT113), .A3(new_n826), .A4(new_n314), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT113), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n828), .B1(new_n761), .B2(new_n825), .ZN(new_n829));
  AND2_X1   g643(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  AOI22_X1  g644(.A1(new_n830), .A2(new_n661), .B1(new_n734), .B2(new_n747), .ZN(new_n831));
  NAND4_X1  g645(.A1(new_n831), .A2(new_n756), .A3(new_n750), .A4(new_n759), .ZN(new_n832));
  NOR2_X1   g646(.A1(new_n824), .A2(new_n832), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n813), .A2(new_n815), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(KEYINPUT53), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n807), .A2(new_n812), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n833), .A2(new_n837), .A3(KEYINPUT53), .ZN(new_n838));
  AOI21_X1  g652(.A(new_n798), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  AND2_X1   g653(.A1(new_n807), .A2(new_n812), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n830), .A2(new_n661), .ZN(new_n841));
  INV_X1    g655(.A(new_n734), .ZN(new_n842));
  OAI21_X1  g656(.A(new_n841), .B1(new_n842), .B2(new_n746), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n750), .A2(new_n759), .A3(new_n756), .ZN(new_n844));
  NOR2_X1   g658(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n845), .A2(new_n823), .A3(new_n818), .A4(new_n816), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n835), .B1(new_n840), .B2(new_n846), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n824), .A2(new_n835), .A3(new_n832), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n813), .A3(new_n815), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n847), .A2(new_n798), .A3(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n839), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n716), .A2(new_n719), .ZN(new_n852));
  OR3_X1    g666(.A1(new_n852), .A2(new_n314), .A3(new_n678), .ZN(new_n853));
  OR2_X1    g667(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n854));
  INV_X1    g668(.A(new_n249), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n766), .A2(new_n855), .ZN(new_n856));
  AND2_X1   g670(.A1(new_n727), .A2(new_n635), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n857), .A2(new_n564), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(KEYINPUT115), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n854), .A2(new_n859), .A3(new_n860), .ZN(new_n861));
  XNOR2_X1  g675(.A(new_n861), .B(KEYINPUT50), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n852), .A2(new_n761), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n863), .A2(new_n855), .A3(new_n766), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n857), .A2(new_n657), .ZN(new_n865));
  NOR2_X1   g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  NOR3_X1   g680(.A1(new_n688), .A2(new_n638), .A3(new_n249), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n863), .A2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n868), .A2(new_n312), .A3(new_n628), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n862), .A2(new_n866), .A3(new_n869), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n787), .B(new_n789), .C1(new_n565), .C2(new_n792), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(new_n314), .A3(new_n744), .A4(new_n859), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n870), .A2(KEYINPUT51), .A3(new_n872), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n864), .A2(new_n754), .ZN(new_n877));
  XNOR2_X1  g691(.A(new_n877), .B(KEYINPUT48), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n720), .A2(new_n859), .ZN(new_n879));
  OAI211_X1 g693(.A(new_n879), .B(new_n245), .C1(new_n868), .C2(new_n629), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n878), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT116), .ZN(new_n882));
  AND4_X1   g696(.A1(new_n851), .A2(new_n875), .A3(new_n876), .A4(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(G952), .A2(G953), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n797), .B1(new_n883), .B2(new_n884), .ZN(G75));
  NOR2_X1   g699(.A1(new_n252), .A2(G952), .ZN(new_n886));
  INV_X1    g700(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n234), .B1(new_n847), .B2(new_n849), .ZN(new_n888));
  AOI21_X1  g702(.A(KEYINPUT56), .B1(new_n888), .B2(G210), .ZN(new_n889));
  NOR2_X1   g703(.A1(new_n380), .A2(new_n381), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n890), .B(KEYINPUT117), .Z(new_n891));
  XNOR2_X1  g705(.A(new_n335), .B(KEYINPUT55), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n891), .B(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n887), .B1(new_n889), .B2(new_n893), .ZN(new_n894));
  AOI21_X1  g708(.A(new_n894), .B1(new_n889), .B2(new_n893), .ZN(G51));
  AND3_X1   g709(.A1(new_n848), .A2(new_n815), .A3(new_n813), .ZN(new_n896));
  AOI21_X1  g710(.A(KEYINPUT53), .B1(new_n833), .B2(new_n837), .ZN(new_n897));
  OAI21_X1  g711(.A(KEYINPUT54), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n847), .A2(new_n798), .A3(new_n849), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n568), .B(KEYINPUT57), .ZN(new_n901));
  AOI21_X1  g715(.A(new_n698), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  OR2_X1    g716(.A1(new_n902), .A2(KEYINPUT118), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n888), .A2(new_n774), .A3(new_n776), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n904), .B1(new_n902), .B2(KEYINPUT118), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n886), .B1(new_n903), .B2(new_n905), .ZN(G54));
  NAND3_X1  g720(.A1(new_n888), .A2(KEYINPUT58), .A3(G475), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n289), .A2(new_n300), .ZN(new_n908));
  AND2_X1   g722(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n907), .A2(new_n908), .ZN(new_n910));
  NOR3_X1   g724(.A1(new_n909), .A2(new_n910), .A3(new_n886), .ZN(G60));
  OR2_X1    g725(.A1(new_n625), .A2(KEYINPUT33), .ZN(new_n912));
  AND2_X1   g726(.A1(new_n912), .A2(new_n622), .ZN(new_n913));
  INV_X1    g727(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(G478), .A2(G902), .ZN(new_n915));
  XOR2_X1   g729(.A(new_n915), .B(KEYINPUT59), .Z(new_n916));
  NOR2_X1   g730(.A1(new_n914), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n918), .B1(new_n898), .B2(new_n899), .ZN(new_n919));
  OAI21_X1  g733(.A(KEYINPUT119), .B1(new_n919), .B2(new_n886), .ZN(new_n920));
  AOI21_X1  g734(.A(new_n798), .B1(new_n847), .B2(new_n849), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n917), .B1(new_n850), .B2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(KEYINPUT119), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n922), .A2(new_n923), .A3(new_n887), .ZN(new_n924));
  INV_X1    g738(.A(new_n916), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n925), .B1(new_n839), .B2(new_n850), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n926), .A2(new_n914), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n920), .A2(new_n924), .A3(new_n927), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT120), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n920), .A2(new_n924), .A3(new_n927), .A4(KEYINPUT120), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n930), .A2(new_n931), .ZN(G63));
  NAND2_X1  g746(.A1(G217), .A2(G902), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT60), .Z(new_n934));
  OAI21_X1  g748(.A(new_n934), .B1(new_n896), .B2(new_n897), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n546), .A2(new_n549), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n886), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n654), .A2(new_n655), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT121), .Z(new_n939));
  OAI21_X1  g753(.A(new_n937), .B1(new_n935), .B2(new_n939), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT61), .Z(G66));
  OAI21_X1  g755(.A(G953), .B1(new_n254), .B2(new_n333), .ZN(new_n942));
  INV_X1    g756(.A(new_n824), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n942), .B1(new_n943), .B2(new_n590), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT122), .Z(new_n945));
  OAI21_X1  g759(.A(new_n891), .B1(G898), .B2(new_n252), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(G69));
  OAI21_X1  g761(.A(new_n291), .B1(new_n266), .B2(new_n292), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n488), .B(new_n948), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AND2_X1   g764(.A1(new_n950), .A2(KEYINPUT125), .ZN(new_n951));
  INV_X1    g765(.A(G900), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n590), .B1(new_n591), .B2(new_n952), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n800), .B1(new_n810), .B2(new_n691), .ZN(new_n956));
  INV_X1    g770(.A(new_n956), .ZN(new_n957));
  NOR3_X1   g771(.A1(new_n783), .A2(new_n844), .A3(new_n957), .ZN(new_n958));
  INV_X1    g772(.A(new_n754), .ZN(new_n959));
  NAND4_X1  g773(.A1(new_n781), .A2(new_n681), .A3(new_n731), .A4(new_n959), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT124), .ZN(new_n961));
  INV_X1    g775(.A(new_n790), .ZN(new_n962));
  NAND4_X1  g776(.A1(new_n958), .A2(new_n961), .A3(new_n252), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n949), .B1(G900), .B2(new_n590), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n956), .A2(new_n689), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n967));
  XOR2_X1   g781(.A(new_n967), .B(KEYINPUT123), .Z(new_n968));
  NOR4_X1   g782(.A1(new_n694), .A2(new_n682), .A3(new_n761), .A4(new_n819), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n783), .A2(new_n790), .A3(new_n969), .ZN(new_n970));
  OR2_X1    g784(.A1(new_n966), .A2(KEYINPUT62), .ZN(new_n971));
  NAND3_X1  g785(.A1(new_n968), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n972), .A2(new_n252), .ZN(new_n973));
  OAI211_X1 g787(.A(new_n955), .B(new_n965), .C1(new_n973), .C2(new_n950), .ZN(new_n974));
  INV_X1    g788(.A(new_n965), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n950), .B1(new_n972), .B2(new_n252), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n954), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n974), .A2(new_n977), .ZN(G72));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT63), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT126), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n958), .A2(new_n962), .A3(new_n961), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(new_n824), .ZN(new_n983));
  XNOR2_X1  g797(.A(new_n489), .B(KEYINPUT127), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n984), .A2(new_n423), .ZN(new_n985));
  AOI21_X1  g799(.A(new_n886), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n981), .B1(new_n972), .B2(new_n824), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n984), .A2(new_n423), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n836), .A2(new_n838), .ZN(new_n990));
  INV_X1    g804(.A(new_n511), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n980), .B1(new_n991), .B2(new_n505), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n990), .A2(new_n992), .ZN(new_n993));
  AND3_X1   g807(.A1(new_n986), .A2(new_n989), .A3(new_n993), .ZN(G57));
endmodule


