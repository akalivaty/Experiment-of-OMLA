//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 1 1 1 1 0 1 0 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 0 1 1 1 1 1 0 0 0 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:53 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1092, new_n1093,
    new_n1094, new_n1095, new_n1096, new_n1097, new_n1098, new_n1099,
    new_n1100, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1126, new_n1127, new_n1128, new_n1129, new_n1130,
    new_n1131, new_n1132, new_n1133, new_n1134, new_n1135, new_n1136,
    new_n1137, new_n1138, new_n1139, new_n1140, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1288, new_n1289,
    new_n1290, new_n1291, new_n1292, new_n1293, new_n1294, new_n1295,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1316, new_n1317, new_n1318, new_n1319, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1327,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1405, new_n1406, new_n1407,
    new_n1408, new_n1409;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AOI211_X1 g0005(.A(G50), .B(G77), .C1(new_n204), .C2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n204), .A2(new_n205), .ZN(new_n215));
  INV_X1    g0015(.A(G50), .ZN(new_n216));
  NOR2_X1   g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND2_X1  g0017(.A1(G1), .A2(G13), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n218), .A2(new_n209), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  AND2_X1   g0020(.A1(KEYINPUT65), .A2(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(KEYINPUT65), .A2(G238), .ZN(new_n222));
  OR2_X1    g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  AND2_X1   g0023(.A1(new_n223), .A2(G68), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n225));
  AOI22_X1  g0025(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G107), .A2(G264), .ZN(new_n228));
  NAND4_X1  g0028(.A1(new_n225), .A2(new_n226), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n211), .B1(new_n224), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n214), .B(new_n220), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(KEYINPUT2), .B(G226), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XOR2_X1   g0036(.A(G264), .B(G270), .Z(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G358));
  XOR2_X1   g0040(.A(G50), .B(G58), .Z(new_n241));
  XNOR2_X1  g0041(.A(new_n241), .B(KEYINPUT66), .ZN(new_n242));
  XNOR2_X1  g0042(.A(G68), .B(G77), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  AND2_X1   g0048(.A1(KEYINPUT3), .A2(G33), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT3), .A2(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G77), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT67), .B(G1698), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n253), .A2(G222), .B1(G223), .B2(G1698), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n252), .B1(new_n254), .B2(new_n251), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT68), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g0057(.A1(G33), .A2(G41), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(new_n218), .ZN(new_n259));
  OAI211_X1 g0059(.A(KEYINPUT68), .B(new_n252), .C1(new_n254), .C2(new_n251), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G41), .ZN(new_n262));
  INV_X1    g0062(.A(G45), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  AND2_X1   g0064(.A1(G1), .A2(G13), .ZN(new_n265));
  NAND2_X1  g0065(.A1(G33), .A2(G41), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n208), .A2(new_n264), .B1(new_n265), .B2(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(G274), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n268), .B1(new_n265), .B2(new_n266), .ZN(new_n269));
  AOI21_X1  g0069(.A(G1), .B1(new_n262), .B2(new_n263), .ZN(new_n270));
  AOI22_X1  g0070(.A1(new_n267), .A2(G226), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n261), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(G200), .ZN(new_n273));
  NAND3_X1  g0073(.A1(new_n261), .A2(G190), .A3(new_n271), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g0075(.A(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(new_n218), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n209), .B1(new_n215), .B2(new_n216), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT8), .B(G58), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n209), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G150), .ZN(new_n282));
  NOR2_X1   g0082(.A1(G20), .A2(G33), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  OAI22_X1  g0084(.A1(new_n280), .A2(new_n281), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n278), .B1(new_n279), .B2(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT69), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  OAI211_X1 g0088(.A(KEYINPUT69), .B(new_n278), .C1(new_n279), .C2(new_n285), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n290));
  INV_X1    g0090(.A(new_n290), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(new_n278), .ZN(new_n292));
  AOI21_X1  g0092(.A(new_n216), .B1(new_n208), .B2(G20), .ZN(new_n293));
  AOI22_X1  g0093(.A1(new_n292), .A2(new_n293), .B1(new_n216), .B2(new_n291), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n288), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT9), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n276), .A2(KEYINPUT75), .A3(KEYINPUT10), .A4(new_n296), .ZN(new_n297));
  NAND2_X1  g0097(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n298));
  OR2_X1    g0098(.A1(KEYINPUT75), .A2(KEYINPUT10), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT9), .ZN(new_n300));
  XNOR2_X1  g0100(.A(new_n295), .B(new_n300), .ZN(new_n301));
  OAI211_X1 g0101(.A(new_n298), .B(new_n299), .C1(new_n275), .C2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n272), .A2(G179), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT70), .ZN(new_n306));
  INV_X1    g0106(.A(G169), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n306), .B1(new_n272), .B2(new_n307), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n305), .B(new_n295), .C1(new_n304), .C2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n303), .A2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n292), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n313));
  INV_X1    g0113(.A(KEYINPUT8), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n314), .A2(G58), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n313), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n208), .A2(G20), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI22_X1  g0118(.A1(new_n312), .A2(new_n318), .B1(new_n290), .B2(new_n316), .ZN(new_n319));
  AND2_X1   g0119(.A1(new_n277), .A2(new_n218), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n202), .A2(new_n203), .ZN(new_n321));
  OAI21_X1  g0121(.A(G20), .B1(new_n215), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G159), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n322), .B1(new_n323), .B2(new_n284), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT79), .ZN(new_n325));
  NOR3_X1   g0125(.A1(new_n249), .A2(new_n250), .A3(G20), .ZN(new_n326));
  OAI21_X1  g0126(.A(new_n325), .B1(new_n326), .B2(KEYINPUT7), .ZN(new_n327));
  INV_X1    g0127(.A(KEYINPUT3), .ZN(new_n328));
  INV_X1    g0128(.A(G33), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(KEYINPUT3), .A2(G33), .ZN(new_n331));
  NAND4_X1  g0131(.A1(new_n330), .A2(KEYINPUT7), .A3(new_n209), .A4(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n332), .A2(KEYINPUT80), .ZN(new_n333));
  INV_X1    g0133(.A(KEYINPUT80), .ZN(new_n334));
  NAND4_X1  g0134(.A1(new_n251), .A2(new_n334), .A3(KEYINPUT7), .A4(new_n209), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n330), .A2(new_n209), .A3(new_n331), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT7), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n336), .A2(KEYINPUT79), .A3(new_n337), .ZN(new_n338));
  NAND4_X1  g0138(.A1(new_n327), .A2(new_n333), .A3(new_n335), .A4(new_n338), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n324), .B1(new_n339), .B2(G68), .ZN(new_n340));
  AOI21_X1  g0140(.A(new_n320), .B1(new_n340), .B2(KEYINPUT16), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT7), .B1(new_n251), .B2(new_n209), .ZN(new_n342));
  INV_X1    g0142(.A(new_n332), .ZN(new_n343));
  OAI21_X1  g0143(.A(G68), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI211_X1 g0144(.A(new_n204), .B(new_n205), .C1(new_n202), .C2(new_n203), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n345), .A2(G20), .B1(G159), .B2(new_n283), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT16), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n319), .B1(new_n341), .B2(new_n348), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n269), .A2(new_n270), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n264), .A2(new_n208), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n265), .A2(new_n266), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(G232), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n350), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n330), .A2(new_n331), .ZN(new_n356));
  NAND3_X1  g0156(.A1(new_n356), .A2(G226), .A3(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G87), .ZN(new_n358));
  INV_X1    g0158(.A(G223), .ZN(new_n359));
  INV_X1    g0159(.A(G1698), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(KEYINPUT67), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT67), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(G1698), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n361), .B(new_n363), .C1(new_n249), .C2(new_n250), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n357), .B(new_n358), .C1(new_n359), .C2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n355), .B1(new_n365), .B2(new_n259), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n366), .A2(G179), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n307), .B2(new_n366), .ZN(new_n368));
  INV_X1    g0168(.A(new_n368), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT18), .B1(new_n349), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n339), .A2(G68), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(KEYINPUT16), .A3(new_n346), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n372), .A2(new_n348), .A3(new_n278), .ZN(new_n373));
  INV_X1    g0173(.A(new_n319), .ZN(new_n374));
  INV_X1    g0174(.A(G190), .ZN(new_n375));
  AOI211_X1 g0175(.A(new_n375), .B(new_n355), .C1(new_n365), .C2(new_n259), .ZN(new_n376));
  INV_X1    g0176(.A(G200), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n365), .A2(new_n259), .ZN(new_n378));
  INV_X1    g0178(.A(new_n355), .ZN(new_n379));
  AOI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n374), .A3(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(KEYINPUT17), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  INV_X1    g0184(.A(KEYINPUT18), .ZN(new_n385));
  AOI211_X1 g0185(.A(new_n320), .B(new_n347), .C1(new_n340), .C2(KEYINPUT16), .ZN(new_n386));
  OAI211_X1 g0186(.A(new_n385), .B(new_n368), .C1(new_n386), .C2(new_n319), .ZN(new_n387));
  NAND4_X1  g0187(.A1(new_n373), .A2(new_n381), .A3(KEYINPUT17), .A4(new_n374), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n370), .A2(new_n384), .A3(new_n387), .A4(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(G179), .ZN(new_n391));
  OAI21_X1  g0191(.A(G1698), .B1(new_n221), .B2(new_n222), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n361), .A2(new_n363), .A3(G232), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(new_n356), .ZN(new_n394));
  INV_X1    g0194(.A(G107), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n352), .B1(new_n251), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT71), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n267), .A2(G244), .B1(new_n269), .B2(new_n270), .ZN(new_n399));
  AND3_X1   g0199(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n398), .B1(new_n397), .B2(new_n399), .ZN(new_n401));
  OAI21_X1  g0201(.A(new_n391), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n402), .A2(KEYINPUT73), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n397), .A2(new_n399), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n404), .A2(KEYINPUT71), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT73), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n407), .A2(new_n408), .A3(new_n391), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n403), .A2(new_n409), .ZN(new_n410));
  NAND3_X1  g0210(.A1(new_n405), .A2(new_n307), .A3(new_n406), .ZN(new_n411));
  INV_X1    g0211(.A(G77), .ZN(new_n412));
  OAI22_X1  g0212(.A1(new_n280), .A2(new_n284), .B1(new_n209), .B2(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT72), .ZN(new_n414));
  XNOR2_X1  g0214(.A(KEYINPUT15), .B(G87), .ZN(new_n415));
  OAI22_X1  g0215(.A1(new_n413), .A2(new_n414), .B1(new_n281), .B2(new_n415), .ZN(new_n416));
  AND2_X1   g0216(.A1(new_n413), .A2(new_n414), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n278), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n412), .B1(new_n208), .B2(G20), .ZN(new_n419));
  AOI22_X1  g0219(.A1(new_n292), .A2(new_n419), .B1(new_n412), .B2(new_n291), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n411), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT74), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT74), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n411), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n410), .A2(new_n423), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n407), .A2(G190), .ZN(new_n427));
  INV_X1    g0227(.A(new_n421), .ZN(new_n428));
  OAI211_X1 g0228(.A(new_n427), .B(new_n428), .C1(new_n377), .C2(new_n407), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n283), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n431), .B1(new_n412), .B2(new_n281), .ZN(new_n432));
  AOI21_X1  g0232(.A(KEYINPUT11), .B1(new_n432), .B2(new_n278), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT76), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n432), .A2(KEYINPUT11), .A3(new_n278), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n436), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT76), .B1(new_n438), .B2(new_n433), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n292), .A2(G68), .A3(new_n317), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT12), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n441), .B1(new_n291), .B2(new_n203), .ZN(new_n442));
  NOR3_X1   g0242(.A1(new_n290), .A2(KEYINPUT12), .A3(G68), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n440), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT77), .ZN(new_n446));
  OAI211_X1 g0246(.A(new_n440), .B(new_n446), .C1(new_n442), .C2(new_n443), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n437), .A2(new_n439), .A3(new_n445), .A4(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n361), .A2(new_n363), .A3(G226), .ZN(new_n449));
  NAND2_X1  g0249(.A1(G232), .A2(G1698), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n251), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(G97), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n329), .A2(new_n452), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n259), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(KEYINPUT13), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n267), .A2(G238), .B1(new_n269), .B2(new_n270), .ZN(new_n456));
  AND3_X1   g0256(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI21_X1  g0257(.A(new_n455), .B1(new_n454), .B2(new_n456), .ZN(new_n458));
  OAI21_X1  g0258(.A(G169), .B1(new_n457), .B2(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT78), .B1(new_n459), .B2(KEYINPUT14), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT14), .ZN(new_n461));
  OAI211_X1 g0261(.A(new_n461), .B(G169), .C1(new_n457), .C2(new_n458), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n454), .A2(new_n456), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(KEYINPUT13), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n464), .A2(G179), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n462), .A2(new_n466), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n460), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n459), .A2(KEYINPUT78), .A3(KEYINPUT14), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n448), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(G200), .B1(new_n457), .B2(new_n458), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n464), .A2(G190), .A3(new_n465), .ZN(new_n472));
  AND3_X1   g0272(.A1(new_n448), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n311), .A2(new_n390), .A3(new_n430), .A4(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n208), .A2(G45), .ZN(new_n477));
  OR2_X1    g0277(.A1(KEYINPUT5), .A2(G41), .ZN(new_n478));
  NAND2_X1  g0278(.A1(KEYINPUT5), .A2(G41), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n269), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n479), .ZN(new_n482));
  NOR2_X1   g0282(.A1(new_n263), .A2(G1), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n352), .ZN(new_n485));
  INV_X1    g0285(.A(G257), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n481), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  INV_X1    g0287(.A(new_n487), .ZN(new_n488));
  INV_X1    g0288(.A(KEYINPUT83), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n356), .A2(new_n253), .A3(G244), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(KEYINPUT82), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT4), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT82), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n356), .A2(new_n253), .A3(new_n493), .A4(G244), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n491), .A2(new_n492), .A3(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(G250), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n496));
  NAND2_X1  g0296(.A1(G33), .A2(G283), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(G244), .ZN(new_n499));
  NOR2_X1   g0299(.A1(new_n364), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n498), .B1(new_n500), .B2(KEYINPUT4), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n489), .B1(new_n502), .B2(new_n259), .ZN(new_n503));
  AOI211_X1 g0303(.A(KEYINPUT83), .B(new_n352), .C1(new_n495), .C2(new_n501), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n488), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G200), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n208), .A2(G33), .ZN(new_n507));
  NAND4_X1  g0307(.A1(new_n290), .A2(new_n507), .A3(new_n218), .A4(new_n277), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(G97), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n509), .B1(G97), .B2(new_n291), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(KEYINPUT81), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT81), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n509), .B(new_n512), .C1(G97), .C2(new_n291), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n511), .A2(new_n513), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT6), .ZN(new_n515));
  NOR3_X1   g0315(.A1(new_n515), .A2(new_n452), .A3(G107), .ZN(new_n516));
  XNOR2_X1  g0316(.A(G97), .B(G107), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n516), .B1(new_n515), .B2(new_n517), .ZN(new_n518));
  OAI22_X1  g0318(.A1(new_n518), .A2(new_n209), .B1(new_n412), .B2(new_n284), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n336), .A2(new_n337), .ZN(new_n520));
  AOI21_X1  g0320(.A(new_n395), .B1(new_n520), .B2(new_n332), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n278), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n514), .A2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n487), .B1(new_n502), .B2(new_n259), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n523), .B1(new_n524), .B2(G190), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n391), .B(new_n488), .C1(new_n503), .C2(new_n504), .ZN(new_n526));
  NAND4_X1  g0326(.A1(new_n356), .A2(new_n253), .A3(KEYINPUT4), .A4(G244), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n527), .A2(new_n497), .A3(new_n496), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT4), .B1(new_n490), .B2(KEYINPUT82), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n528), .B1(new_n494), .B2(new_n529), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n488), .B1(new_n530), .B2(new_n352), .ZN(new_n531));
  AOI22_X1  g0331(.A1(new_n531), .A2(new_n307), .B1(new_n522), .B2(new_n514), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n506), .A2(new_n525), .B1(new_n526), .B2(new_n532), .ZN(new_n533));
  OAI211_X1 g0333(.A(G257), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n534));
  NAND2_X1  g0334(.A1(G33), .A2(G294), .ZN(new_n535));
  INV_X1    g0335(.A(G250), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n534), .B(new_n535), .C1(new_n364), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n480), .A2(new_n259), .ZN(new_n538));
  AOI22_X1  g0338(.A1(new_n537), .A2(new_n259), .B1(new_n538), .B2(G264), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n539), .A2(new_n391), .A3(new_n481), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n539), .A2(new_n481), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(new_n307), .ZN(new_n542));
  INV_X1    g0342(.A(G116), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n543), .A2(KEYINPUT85), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT85), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G116), .ZN(new_n546));
  AOI21_X1  g0346(.A(new_n329), .B1(new_n544), .B2(new_n546), .ZN(new_n547));
  INV_X1    g0347(.A(KEYINPUT23), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(new_n209), .B2(G107), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n395), .A2(KEYINPUT23), .A3(G20), .ZN(new_n550));
  AOI22_X1  g0350(.A1(new_n547), .A2(new_n209), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g0351(.A(KEYINPUT22), .ZN(new_n552));
  AOI21_X1  g0352(.A(G20), .B1(new_n330), .B2(new_n331), .ZN(new_n553));
  AOI21_X1  g0353(.A(new_n552), .B1(new_n553), .B2(G87), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n209), .B(G87), .C1(new_n249), .C2(new_n250), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n556));
  OAI21_X1  g0356(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(KEYINPUT24), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n555), .A2(KEYINPUT22), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n356), .A2(new_n552), .A3(new_n209), .A4(G87), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT24), .ZN(new_n562));
  NAND3_X1  g0362(.A1(new_n561), .A2(new_n562), .A3(new_n551), .ZN(new_n563));
  AOI21_X1  g0363(.A(new_n320), .B1(new_n558), .B2(new_n563), .ZN(new_n564));
  INV_X1    g0364(.A(new_n508), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n291), .A2(KEYINPUT25), .A3(new_n395), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT25), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(new_n290), .B2(G107), .ZN(new_n568));
  AOI22_X1  g0368(.A1(G107), .A2(new_n565), .B1(new_n566), .B2(new_n568), .ZN(new_n569));
  INV_X1    g0369(.A(new_n569), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n540), .B(new_n542), .C1(new_n564), .C2(new_n570), .ZN(new_n571));
  AND3_X1   g0371(.A1(new_n561), .A2(new_n562), .A3(new_n551), .ZN(new_n572));
  AOI21_X1  g0372(.A(new_n562), .B1(new_n561), .B2(new_n551), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n278), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  AND3_X1   g0374(.A1(new_n539), .A2(new_n375), .A3(new_n481), .ZN(new_n575));
  AOI21_X1  g0375(.A(G200), .B1(new_n539), .B2(new_n481), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n574), .B(new_n569), .C1(new_n575), .C2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n578), .A2(KEYINPUT93), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT93), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n571), .A2(new_n577), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n544), .A2(new_n546), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n583), .A2(G33), .ZN(new_n584));
  OAI211_X1 g0384(.A(G244), .B(G1698), .C1(new_n249), .C2(new_n250), .ZN(new_n585));
  INV_X1    g0385(.A(G238), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n584), .B(new_n585), .C1(new_n586), .C2(new_n364), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n259), .ZN(new_n588));
  NOR3_X1   g0388(.A1(new_n259), .A2(new_n536), .A3(new_n483), .ZN(new_n589));
  OAI21_X1  g0389(.A(G274), .B1(new_n258), .B2(new_n218), .ZN(new_n590));
  OAI21_X1  g0390(.A(KEYINPUT84), .B1(new_n590), .B2(new_n477), .ZN(new_n591));
  INV_X1    g0391(.A(KEYINPUT84), .ZN(new_n592));
  NAND3_X1  g0392(.A1(new_n269), .A2(new_n592), .A3(new_n483), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n589), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n588), .A2(new_n391), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n588), .A2(new_n594), .A3(KEYINPUT86), .A4(new_n391), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT89), .ZN(new_n600));
  NAND3_X1  g0400(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n209), .ZN(new_n602));
  INV_X1    g0402(.A(G87), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n603), .A2(new_n452), .A3(new_n395), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n602), .A2(KEYINPUT87), .A3(new_n604), .ZN(new_n605));
  AOI21_X1  g0405(.A(KEYINPUT87), .B1(new_n602), .B2(new_n604), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n209), .B(G68), .C1(new_n249), .C2(new_n250), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n209), .A2(G33), .A3(G97), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT19), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n609), .A2(KEYINPUT88), .A3(new_n610), .ZN(new_n611));
  AOI21_X1  g0411(.A(KEYINPUT88), .B1(new_n609), .B2(new_n610), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n608), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n600), .B1(new_n607), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n602), .A2(new_n604), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT87), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g0417(.A1(new_n602), .A2(KEYINPUT87), .A3(new_n604), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n609), .A2(new_n610), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT88), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n609), .A2(KEYINPUT88), .A3(new_n610), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND4_X1  g0424(.A1(new_n619), .A2(KEYINPUT89), .A3(new_n608), .A4(new_n624), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n614), .A2(new_n625), .A3(new_n278), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n415), .A2(new_n291), .ZN(new_n627));
  OR2_X1    g0427(.A1(new_n508), .A2(new_n415), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(G169), .B1(new_n588), .B2(new_n594), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n599), .A2(new_n629), .A3(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n588), .A2(new_n594), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n377), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n588), .A2(new_n375), .A3(new_n594), .ZN(new_n635));
  NAND2_X1  g0435(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n565), .A2(G87), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(new_n637), .A3(new_n627), .A4(new_n626), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n632), .A2(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n486), .B1(new_n330), .B2(new_n331), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n253), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n356), .A2(G264), .A3(G1698), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n251), .A2(G303), .ZN(new_n643));
  NAND3_X1  g0443(.A1(new_n641), .A2(new_n642), .A3(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n644), .A2(new_n259), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n538), .A2(G270), .B1(new_n269), .B2(new_n480), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n307), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n544), .A2(new_n546), .A3(G20), .ZN(new_n648));
  OAI211_X1 g0448(.A(new_n497), .B(new_n209), .C1(G33), .C2(new_n452), .ZN(new_n649));
  NOR2_X1   g0449(.A1(KEYINPUT90), .A2(KEYINPUT20), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n648), .A2(new_n278), .A3(new_n649), .A4(new_n650), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n320), .A2(G116), .A3(new_n290), .A4(new_n507), .ZN(new_n652));
  AND2_X1   g0452(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n648), .A2(new_n278), .A3(new_n649), .ZN(new_n654));
  XOR2_X1   g0454(.A(KEYINPUT90), .B(KEYINPUT20), .Z(new_n655));
  INV_X1    g0455(.A(new_n583), .ZN(new_n656));
  AOI22_X1  g0456(.A1(new_n654), .A2(new_n655), .B1(new_n291), .B2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT91), .ZN(new_n658));
  AND3_X1   g0458(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n658), .B1(new_n653), .B2(new_n657), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n647), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  XOR2_X1   g0461(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n662));
  NAND2_X1  g0462(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  AOI22_X1  g0463(.A1(new_n640), .A2(new_n253), .B1(new_n251), .B2(G303), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n352), .B1(new_n664), .B2(new_n642), .ZN(new_n665));
  INV_X1    g0465(.A(G270), .ZN(new_n666));
  OAI21_X1  g0466(.A(new_n481), .B1(new_n485), .B2(new_n666), .ZN(new_n667));
  OAI211_X1 g0467(.A(KEYINPUT21), .B(G169), .C1(new_n665), .C2(new_n667), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n645), .A2(new_n646), .A3(G179), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n653), .A2(new_n657), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(KEYINPUT91), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n653), .A2(new_n657), .A3(new_n658), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n670), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n645), .A2(new_n646), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G200), .ZN(new_n677));
  NAND3_X1  g0477(.A1(new_n645), .A2(new_n646), .A3(G190), .ZN(new_n678));
  NAND4_X1  g0478(.A1(new_n677), .A2(new_n673), .A3(new_n672), .A4(new_n678), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n663), .A2(new_n675), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n639), .A2(new_n680), .ZN(new_n681));
  AND4_X1   g0481(.A1(new_n476), .A2(new_n533), .A3(new_n582), .A4(new_n681), .ZN(G372));
  INV_X1    g0482(.A(KEYINPUT97), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT96), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n426), .A2(new_n473), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n684), .B1(new_n470), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n384), .A2(new_n388), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  AOI22_X1  g0488(.A1(new_n403), .A2(new_n409), .B1(new_n422), .B2(KEYINPUT74), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n448), .A2(new_n472), .A3(new_n471), .ZN(new_n690));
  NAND3_X1  g0490(.A1(new_n689), .A2(new_n425), .A3(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(new_n469), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n692), .A2(new_n460), .A3(new_n467), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n691), .B(KEYINPUT96), .C1(new_n693), .C2(new_n448), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n686), .A2(new_n688), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n370), .A2(new_n387), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n303), .B1(new_n695), .B2(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n683), .B1(new_n698), .B2(new_n310), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n691), .B1(new_n693), .B2(new_n448), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n687), .B1(new_n700), .B2(new_n684), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n696), .B1(new_n701), .B2(new_n694), .ZN(new_n702));
  OAI211_X1 g0502(.A(KEYINPUT97), .B(new_n309), .C1(new_n702), .C2(new_n303), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n699), .A2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n571), .A2(new_n663), .A3(new_n675), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n588), .A2(new_n391), .A3(new_n594), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n706), .A2(new_n630), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n629), .A2(new_n707), .ZN(new_n708));
  AND3_X1   g0508(.A1(new_n638), .A2(new_n577), .A3(new_n708), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n533), .A2(new_n705), .A3(new_n709), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  XNOR2_X1  g0511(.A(new_n708), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g0512(.A1(new_n638), .A2(new_n526), .A3(new_n708), .A4(new_n532), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  AND2_X1   g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  NAND4_X1  g0515(.A1(new_n632), .A2(new_n638), .A3(new_n526), .A4(new_n532), .ZN(new_n716));
  XNOR2_X1  g0516(.A(KEYINPUT95), .B(KEYINPUT26), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  OAI211_X1 g0518(.A(new_n710), .B(new_n712), .C1(new_n715), .C2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n704), .B1(new_n475), .B2(new_n720), .ZN(G369));
  NAND3_X1  g0521(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n722));
  OR2_X1    g0522(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(KEYINPUT27), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n723), .A2(G213), .A3(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(G343), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n674), .A2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT98), .ZN(new_n729));
  AND2_X1   g0529(.A1(new_n729), .A2(new_n680), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n663), .A2(new_n675), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n729), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g0532(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(G330), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n727), .B1(new_n564), .B2(new_n570), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n582), .A2(new_n735), .ZN(new_n736));
  INV_X1    g0536(.A(new_n571), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(new_n727), .ZN(new_n738));
  AND2_X1   g0538(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n734), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n727), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n582), .A2(new_n731), .A3(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n737), .A2(new_n742), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n745), .ZN(G399));
  INV_X1    g0546(.A(new_n212), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(G41), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n604), .A2(G116), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n749), .A2(G1), .A3(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n217), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n751), .B1(new_n752), .B2(new_n749), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT28), .ZN(new_n754));
  INV_X1    g0554(.A(new_n713), .ZN(new_n755));
  AOI22_X1  g0555(.A1(new_n755), .A2(KEYINPUT26), .B1(new_n716), .B2(new_n717), .ZN(new_n756));
  AND3_X1   g0556(.A1(new_n626), .A2(new_n637), .A3(new_n627), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(new_n636), .B1(new_n629), .B2(new_n707), .ZN(new_n758));
  NAND3_X1  g0558(.A1(new_n705), .A2(new_n758), .A3(new_n577), .ZN(new_n759));
  OAI21_X1  g0559(.A(KEYINPUT83), .B1(new_n530), .B2(new_n352), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n502), .A2(new_n489), .A3(new_n259), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n487), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n525), .B1(new_n762), .B2(new_n377), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n526), .A2(new_n532), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g0565(.A(new_n712), .B1(new_n759), .B2(new_n765), .ZN(new_n766));
  OAI21_X1  g0566(.A(new_n742), .B1(new_n756), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT29), .ZN(new_n768));
  NAND4_X1  g0568(.A1(new_n582), .A2(new_n681), .A3(new_n533), .A4(new_n742), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT99), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n539), .A2(new_n588), .A3(new_n594), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n771), .A2(new_n669), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n770), .B1(new_n772), .B2(new_n524), .ZN(new_n773));
  INV_X1    g0573(.A(KEYINPUT30), .ZN(new_n774));
  NAND4_X1  g0574(.A1(new_n541), .A2(new_n676), .A3(new_n633), .A4(new_n391), .ZN(new_n775));
  OAI22_X1  g0575(.A1(new_n773), .A2(new_n774), .B1(new_n762), .B2(new_n775), .ZN(new_n776));
  AOI211_X1 g0576(.A(new_n770), .B(KEYINPUT30), .C1(new_n772), .C2(new_n524), .ZN(new_n777));
  OAI21_X1  g0577(.A(new_n727), .B1(new_n776), .B2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(KEYINPUT31), .ZN(new_n779));
  NAND2_X1  g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  OAI211_X1 g0580(.A(KEYINPUT31), .B(new_n727), .C1(new_n776), .C2(new_n777), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n769), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G330), .ZN(new_n783));
  INV_X1    g0583(.A(KEYINPUT29), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n719), .A2(new_n784), .A3(new_n742), .ZN(new_n785));
  NAND3_X1  g0585(.A1(new_n768), .A2(new_n783), .A3(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n754), .B1(new_n787), .B2(G1), .ZN(G364));
  NOR2_X1   g0588(.A1(G13), .A2(G33), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n733), .A2(G20), .A3(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n218), .B1(G20), .B2(new_n307), .ZN(new_n792));
  NAND2_X1  g0592(.A1(G20), .A2(G179), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND3_X1  g0594(.A1(new_n794), .A2(G190), .A3(new_n377), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(G322), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n793), .A2(new_n377), .ZN(new_n798));
  AND3_X1   g0598(.A1(new_n798), .A2(KEYINPUT101), .A3(new_n375), .ZN(new_n799));
  AOI21_X1  g0599(.A(KEYINPUT101), .B1(new_n798), .B2(new_n375), .ZN(new_n800));
  NOR2_X1   g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(KEYINPUT33), .B(G317), .Z(new_n802));
  OAI21_X1  g0602(.A(new_n797), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT103), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n798), .A2(G190), .ZN(new_n805));
  INV_X1    g0605(.A(G326), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n209), .A2(G179), .ZN(new_n807));
  NAND3_X1  g0607(.A1(new_n807), .A2(G190), .A3(G200), .ZN(new_n808));
  INV_X1    g0608(.A(G303), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n805), .A2(new_n806), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NAND3_X1  g0610(.A1(new_n807), .A2(new_n375), .A3(G200), .ZN(new_n811));
  INV_X1    g0611(.A(new_n811), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(G283), .B2(new_n812), .ZN(new_n813));
  NOR2_X1   g0613(.A1(G190), .A2(G200), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n807), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n815), .ZN(new_n816));
  OR2_X1    g0616(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n816), .A2(KEYINPUT102), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(G329), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n794), .A2(new_n814), .ZN(new_n822));
  INV_X1    g0622(.A(G311), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n251), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  NOR3_X1   g0624(.A1(new_n375), .A2(G179), .A3(G200), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n825), .A2(new_n209), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n824), .B1(G294), .B2(new_n827), .ZN(new_n828));
  AND4_X1   g0628(.A1(new_n804), .A2(new_n813), .A3(new_n821), .A4(new_n828), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n812), .A2(G107), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n816), .A2(G159), .ZN(new_n831));
  OAI221_X1 g0631(.A(new_n830), .B1(new_n216), .B2(new_n805), .C1(new_n831), .C2(KEYINPUT32), .ZN(new_n832));
  NOR2_X1   g0632(.A1(new_n826), .A2(new_n452), .ZN(new_n833));
  INV_X1    g0633(.A(new_n808), .ZN(new_n834));
  AOI21_X1  g0634(.A(new_n833), .B1(G87), .B2(new_n834), .ZN(new_n835));
  OAI21_X1  g0635(.A(new_n356), .B1(new_n822), .B2(new_n412), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(new_n831), .B2(KEYINPUT32), .ZN(new_n837));
  XOR2_X1   g0637(.A(new_n795), .B(KEYINPUT100), .Z(new_n838));
  OAI211_X1 g0638(.A(new_n835), .B(new_n837), .C1(new_n202), .C2(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(new_n801), .ZN(new_n840));
  AOI211_X1 g0640(.A(new_n832), .B(new_n839), .C1(G68), .C2(new_n840), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n792), .B1(new_n829), .B2(new_n841), .ZN(new_n842));
  INV_X1    g0642(.A(G13), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n843), .A2(G20), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n208), .B1(new_n844), .B2(G45), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NOR2_X1   g0646(.A1(new_n748), .A2(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n790), .A2(G20), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n848), .A2(new_n792), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n747), .A2(new_n251), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G355), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n852), .B1(G116), .B2(new_n212), .ZN(new_n853));
  OR2_X1    g0653(.A1(new_n244), .A2(new_n263), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n747), .A2(new_n356), .ZN(new_n855));
  INV_X1    g0655(.A(new_n855), .ZN(new_n856));
  AOI21_X1  g0656(.A(new_n856), .B1(new_n217), .B2(new_n263), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n853), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n842), .B(new_n847), .C1(new_n850), .C2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n791), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g0660(.A(new_n860), .B(KEYINPUT104), .ZN(new_n861));
  INV_X1    g0661(.A(new_n734), .ZN(new_n862));
  NOR2_X1   g0662(.A1(new_n862), .A2(new_n847), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n863), .B1(G330), .B2(new_n733), .ZN(new_n864));
  INV_X1    g0664(.A(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n861), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G396));
  NOR2_X1   g0667(.A1(new_n428), .A2(new_n742), .ZN(new_n868));
  AOI21_X1  g0668(.A(new_n868), .B1(new_n426), .B2(new_n429), .ZN(new_n869));
  INV_X1    g0669(.A(new_n868), .ZN(new_n870));
  AOI21_X1  g0670(.A(new_n870), .B1(new_n689), .B2(new_n425), .ZN(new_n871));
  NOR2_X1   g0671(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n639), .A2(new_n764), .ZN(new_n873));
  INV_X1    g0673(.A(new_n717), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n873), .A2(new_n874), .B1(new_n714), .B2(new_n713), .ZN(new_n875));
  OAI211_X1 g0675(.A(new_n742), .B(new_n872), .C1(new_n875), .C2(new_n766), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n876), .A2(KEYINPUT106), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT106), .ZN(new_n878));
  NAND4_X1  g0678(.A1(new_n719), .A2(new_n878), .A3(new_n742), .A4(new_n872), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g0680(.A(new_n708), .B(KEYINPUT94), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n705), .A2(new_n758), .A3(new_n577), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n882), .B2(new_n533), .ZN(new_n883));
  OAI22_X1  g0683(.A1(new_n755), .A2(KEYINPUT26), .B1(new_n716), .B2(new_n717), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n727), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n880), .B1(new_n885), .B2(new_n872), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n847), .B1(new_n886), .B2(new_n783), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n887), .B1(new_n783), .B2(new_n886), .ZN(new_n888));
  INV_X1    g0688(.A(new_n847), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n792), .A2(new_n789), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n889), .B1(new_n412), .B2(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(new_n792), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n811), .A2(new_n603), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n833), .A2(new_n893), .ZN(new_n894));
  OAI221_X1 g0694(.A(new_n894), .B1(new_n395), .B2(new_n808), .C1(new_n809), .C2(new_n805), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n356), .B1(new_n796), .B2(G294), .ZN(new_n896));
  OAI221_X1 g0696(.A(new_n896), .B1(new_n656), .B2(new_n822), .C1(new_n819), .C2(new_n823), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n895), .B(new_n897), .C1(G283), .C2(new_n840), .ZN(new_n898));
  OAI22_X1  g0698(.A1(new_n216), .A2(new_n808), .B1(new_n811), .B2(new_n203), .ZN(new_n899));
  INV_X1    g0699(.A(KEYINPUT105), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n251), .B1(new_n827), .B2(G58), .ZN(new_n903));
  INV_X1    g0703(.A(G132), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n902), .B(new_n903), .C1(new_n819), .C2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n805), .ZN(new_n906));
  INV_X1    g0706(.A(new_n822), .ZN(new_n907));
  AOI22_X1  g0707(.A1(new_n906), .A2(G137), .B1(new_n907), .B2(G159), .ZN(new_n908));
  INV_X1    g0708(.A(G143), .ZN(new_n909));
  OAI221_X1 g0709(.A(new_n908), .B1(new_n282), .B2(new_n801), .C1(new_n838), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  AOI211_X1 g0711(.A(new_n901), .B(new_n905), .C1(new_n911), .C2(KEYINPUT34), .ZN(new_n912));
  OR2_X1    g0712(.A1(new_n911), .A2(KEYINPUT34), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n898), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  OAI221_X1 g0714(.A(new_n891), .B1(new_n892), .B2(new_n914), .C1(new_n872), .C2(new_n790), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n888), .A2(new_n915), .ZN(G384));
  NOR2_X1   g0716(.A1(new_n844), .A2(new_n208), .ZN(new_n917));
  INV_X1    g0717(.A(G330), .ZN(new_n918));
  INV_X1    g0718(.A(new_n448), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n468), .A2(new_n469), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n919), .B(new_n727), .C1(new_n920), .C2(new_n473), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n919), .A2(new_n727), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n690), .B(new_n922), .C1(new_n693), .C2(new_n448), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n782), .A2(new_n872), .A3(new_n924), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT107), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(KEYINPUT107), .A2(KEYINPUT40), .ZN(new_n928));
  NAND4_X1  g0728(.A1(new_n782), .A2(new_n872), .A3(new_n924), .A4(new_n928), .ZN(new_n929));
  INV_X1    g0729(.A(KEYINPUT16), .ZN(new_n930));
  INV_X1    g0730(.A(new_n338), .ZN(new_n931));
  AOI21_X1  g0731(.A(KEYINPUT79), .B1(new_n336), .B2(new_n337), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AND2_X1   g0733(.A1(new_n333), .A2(new_n335), .ZN(new_n934));
  AOI21_X1  g0734(.A(new_n203), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n930), .B1(new_n935), .B2(new_n324), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n319), .B1(new_n341), .B2(new_n936), .ZN(new_n937));
  OAI21_X1  g0737(.A(new_n382), .B1(new_n937), .B2(new_n725), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n369), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT37), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n373), .A2(new_n374), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n941), .A2(new_n368), .ZN(new_n942));
  INV_X1    g0742(.A(new_n725), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(KEYINPUT37), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n942), .A2(new_n944), .A3(new_n945), .A4(new_n382), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n940), .A2(new_n946), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n937), .A2(new_n725), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n389), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT38), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n947), .A2(new_n949), .A3(KEYINPUT38), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n927), .A2(new_n929), .A3(new_n954), .ZN(new_n955));
  AND3_X1   g0755(.A1(new_n947), .A2(new_n949), .A3(KEYINPUT38), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n382), .B1(new_n349), .B2(new_n369), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n349), .A2(new_n725), .ZN(new_n958));
  OAI21_X1  g0758(.A(KEYINPUT37), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(new_n946), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n389), .A2(new_n958), .ZN(new_n961));
  AOI21_X1  g0761(.A(KEYINPUT38), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n956), .A2(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(KEYINPUT40), .B1(new_n963), .B2(new_n925), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n955), .A2(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n476), .A2(new_n782), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n918), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n967), .B1(new_n966), .B2(new_n965), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n968), .B(KEYINPUT108), .Z(new_n969));
  INV_X1    g0769(.A(new_n969), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n426), .A2(new_n727), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(new_n877), .B2(new_n879), .ZN(new_n972));
  AND2_X1   g0772(.A1(new_n921), .A2(new_n923), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n952), .A2(new_n953), .ZN(new_n974));
  NOR3_X1   g0774(.A1(new_n972), .A2(new_n973), .A3(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(KEYINPUT39), .ZN(new_n976));
  OAI21_X1  g0776(.A(new_n976), .B1(new_n956), .B2(new_n962), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n952), .A2(KEYINPUT39), .A3(new_n953), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n470), .A2(new_n742), .ZN(new_n979));
  INV_X1    g0779(.A(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n977), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n696), .A2(new_n725), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n975), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n475), .B1(new_n768), .B2(new_n785), .ZN(new_n985));
  AOI21_X1  g0785(.A(new_n985), .B1(new_n699), .B2(new_n703), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n984), .B(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n917), .B1(new_n970), .B2(new_n987), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n988), .B1(new_n970), .B2(new_n987), .ZN(new_n989));
  INV_X1    g0789(.A(new_n518), .ZN(new_n990));
  OR2_X1    g0790(.A1(new_n990), .A2(KEYINPUT35), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n990), .A2(KEYINPUT35), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n991), .A2(G116), .A3(new_n219), .A4(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n993), .B(KEYINPUT36), .ZN(new_n994));
  NOR3_X1   g0794(.A1(new_n752), .A2(new_n412), .A3(new_n321), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n203), .A2(G50), .ZN(new_n996));
  OAI211_X1 g0796(.A(G1), .B(new_n843), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NAND3_X1  g0797(.A1(new_n989), .A2(new_n994), .A3(new_n997), .ZN(G367));
  OAI221_X1 g0798(.A(new_n849), .B1(new_n212), .B2(new_n415), .C1(new_n856), .C2(new_n239), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n999), .A2(new_n847), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G150), .A2(new_n796), .B1(new_n816), .B2(G137), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n216), .B2(new_n822), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n826), .A2(new_n203), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n805), .A2(new_n909), .B1(new_n808), .B2(new_n202), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n251), .B1(new_n812), .B2(G77), .ZN(new_n1006));
  AOI22_X1  g0806(.A1(new_n840), .A2(G159), .B1(KEYINPUT111), .B2(new_n1006), .ZN(new_n1007));
  OAI211_X1 g0807(.A(new_n1005), .B(new_n1007), .C1(KEYINPUT111), .C2(new_n1006), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT46), .ZN(new_n1009));
  NOR3_X1   g0809(.A1(new_n808), .A2(new_n1009), .A3(new_n543), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n251), .B1(new_n815), .B2(new_n1011), .C1(new_n452), .C2(new_n811), .ZN(new_n1012));
  AOI211_X1 g0812(.A(new_n1010), .B(new_n1012), .C1(G311), .C2(new_n906), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1009), .B1(new_n656), .B2(new_n808), .ZN(new_n1014));
  OAI211_X1 g0814(.A(new_n1013), .B(new_n1014), .C1(new_n809), .C2(new_n838), .ZN(new_n1015));
  INV_X1    g0815(.A(KEYINPUT110), .ZN(new_n1016));
  INV_X1    g0816(.A(G283), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n826), .A2(new_n395), .B1(new_n822), .B2(new_n1017), .ZN(new_n1018));
  AOI22_X1  g0818(.A1(new_n840), .A2(G294), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1019), .B1(new_n1016), .B2(new_n1018), .ZN(new_n1020));
  OAI21_X1  g0820(.A(new_n1008), .B1(new_n1015), .B2(new_n1020), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(KEYINPUT47), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1000), .B1(new_n1022), .B2(new_n792), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n757), .A2(new_n742), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n881), .A2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g0825(.A(new_n758), .B1(new_n757), .B2(new_n742), .ZN(new_n1026));
  NAND3_X1  g0826(.A1(new_n1025), .A2(new_n848), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n1023), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g0828(.A(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(KEYINPUT44), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n523), .A2(new_n727), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n533), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n526), .A2(new_n532), .A3(new_n727), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1030), .B1(new_n745), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1034), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n743), .A2(new_n744), .ZN(new_n1037));
  NAND3_X1  g0837(.A1(new_n1036), .A2(new_n1037), .A3(KEYINPUT44), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1035), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n745), .A2(KEYINPUT45), .A3(new_n1034), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT45), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1042));
  NAND2_X1  g0842(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1039), .A2(new_n1043), .A3(new_n741), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n741), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n731), .A2(new_n742), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n736), .A2(new_n738), .A3(new_n1047), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1048), .A2(new_n743), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(new_n734), .ZN(new_n1050));
  NOR2_X1   g0850(.A1(new_n1050), .A2(new_n786), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n786), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g0852(.A(new_n748), .B(KEYINPUT41), .Z(new_n1053));
  OAI21_X1  g0853(.A(new_n845), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(KEYINPUT43), .ZN(new_n1056));
  XNOR2_X1  g0856(.A(new_n1056), .B(KEYINPUT109), .ZN(new_n1057));
  OR3_X1    g0857(.A1(new_n1036), .A2(KEYINPUT42), .A3(new_n743), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n764), .B1(new_n1032), .B2(new_n571), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n742), .ZN(new_n1060));
  OAI21_X1  g0860(.A(KEYINPUT42), .B1(new_n1036), .B2(new_n743), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n1058), .A2(new_n1060), .A3(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1055), .A2(KEYINPUT43), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1057), .A2(new_n1062), .A3(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1057), .B1(new_n1063), .B2(new_n1062), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n1065), .A2(new_n1066), .B1(new_n741), .B2(new_n1036), .ZN(new_n1067));
  NAND2_X1  g0867(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1068));
  INV_X1    g0868(.A(new_n1057), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NOR2_X1   g0870(.A1(new_n741), .A2(new_n1036), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1070), .A2(new_n1071), .A3(new_n1064), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1029), .B1(new_n1054), .B2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(KEYINPUT112), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1039), .A2(new_n1043), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n740), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1039), .A2(new_n1043), .A3(new_n741), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n787), .B1(new_n1079), .B2(new_n1050), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1053), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n846), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1067), .A2(new_n1072), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1028), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT112), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AND2_X1   g0886(.A1(new_n1075), .A2(new_n1086), .ZN(G387));
  XNOR2_X1  g0887(.A(KEYINPUT113), .B(G150), .ZN(new_n1088));
  OAI22_X1  g0888(.A1(new_n795), .A2(new_n216), .B1(new_n815), .B2(new_n1088), .ZN(new_n1089));
  AOI211_X1 g0889(.A(new_n251), .B(new_n1089), .C1(G68), .C2(new_n907), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n840), .A2(new_n316), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(G159), .A2(new_n906), .B1(new_n812), .B2(G97), .ZN(new_n1092));
  NOR2_X1   g0892(.A1(new_n826), .A2(new_n415), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n1093), .B1(G77), .B2(new_n834), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n356), .B1(new_n816), .B2(G326), .ZN(new_n1096));
  INV_X1    g0896(.A(G294), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n826), .A2(new_n1017), .B1(new_n808), .B2(new_n1097), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(new_n906), .A2(G322), .B1(new_n907), .B2(G303), .ZN(new_n1099));
  OAI221_X1 g0899(.A(new_n1099), .B1(new_n823), .B2(new_n801), .C1(new_n838), .C2(new_n1011), .ZN(new_n1100));
  INV_X1    g0900(.A(KEYINPUT48), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1098), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n1101), .B2(new_n1100), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT49), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n1096), .B1(new_n656), .B2(new_n811), .C1(new_n1103), .C2(new_n1104), .ZN(new_n1105));
  AND2_X1   g0905(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1095), .B1(new_n1105), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1107), .A2(new_n792), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n750), .ZN(new_n1109));
  AOI22_X1  g0909(.A1(new_n851), .A2(new_n1109), .B1(new_n395), .B2(new_n747), .ZN(new_n1110));
  NOR2_X1   g0910(.A1(new_n236), .A2(new_n263), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n316), .A2(new_n216), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1112), .B(KEYINPUT50), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n750), .B(new_n263), .C1(new_n203), .C2(new_n412), .ZN(new_n1114));
  OAI21_X1  g0914(.A(new_n855), .B1(new_n1113), .B2(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1110), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n889), .B1(new_n1116), .B2(new_n849), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1108), .A2(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1118), .B1(new_n739), .B2(new_n848), .ZN(new_n1119));
  INV_X1    g0919(.A(new_n1050), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n1119), .B1(new_n1120), .B2(new_n846), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1120), .A2(new_n787), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n748), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n1120), .A2(new_n787), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1121), .B1(new_n1123), .B2(new_n1124), .ZN(G393));
  INV_X1    g0925(.A(KEYINPUT114), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1077), .A2(new_n1126), .A3(new_n1078), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1044), .B1(new_n1045), .B2(KEYINPUT114), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n1128), .A3(new_n1122), .ZN(new_n1129));
  AOI21_X1  g0929(.A(new_n749), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1036), .A2(new_n848), .ZN(new_n1131));
  OAI221_X1 g0931(.A(new_n849), .B1(new_n452), .B2(new_n212), .C1(new_n856), .C2(new_n247), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n847), .ZN(new_n1133));
  OAI221_X1 g0933(.A(new_n830), .B1(new_n1017), .B2(new_n808), .C1(new_n656), .C2(new_n826), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n356), .B1(new_n816), .B2(G322), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1097), .B2(new_n822), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n805), .A2(new_n1011), .B1(new_n795), .B2(new_n823), .ZN(new_n1138));
  XNOR2_X1  g0938(.A(new_n1138), .B(KEYINPUT52), .ZN(new_n1139));
  OAI211_X1 g0939(.A(new_n1137), .B(new_n1139), .C1(new_n809), .C2(new_n801), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n805), .A2(new_n282), .B1(new_n795), .B2(new_n323), .ZN(new_n1141));
  XOR2_X1   g0941(.A(new_n1141), .B(KEYINPUT51), .Z(new_n1142));
  NOR2_X1   g0942(.A1(new_n808), .A2(new_n203), .ZN(new_n1143));
  AOI211_X1 g0943(.A(new_n893), .B(new_n1143), .C1(G77), .C2(new_n827), .ZN(new_n1144));
  OAI221_X1 g0944(.A(new_n356), .B1(new_n815), .B2(new_n909), .C1(new_n280), .C2(new_n822), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1145), .ZN(new_n1146));
  OAI211_X1 g0946(.A(new_n1144), .B(new_n1146), .C1(new_n216), .C2(new_n801), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1140), .B1(new_n1142), .B2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1133), .B1(new_n1148), .B2(new_n792), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(new_n1129), .A2(new_n1130), .B1(new_n1131), .B2(new_n1149), .ZN(new_n1150));
  NOR3_X1   g0950(.A1(new_n1044), .A2(new_n1045), .A3(KEYINPUT114), .ZN(new_n1151));
  NOR3_X1   g0951(.A1(new_n1076), .A2(new_n1126), .A3(new_n740), .ZN(new_n1152));
  OAI21_X1  g0952(.A(KEYINPUT115), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(KEYINPUT115), .ZN(new_n1154));
  NAND3_X1  g0954(.A1(new_n1127), .A2(new_n1128), .A3(new_n1154), .ZN(new_n1155));
  NAND3_X1  g0955(.A1(new_n1153), .A2(new_n846), .A3(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1150), .A2(new_n1156), .ZN(G390));
  OAI211_X1 g0957(.A(new_n742), .B(new_n872), .C1(new_n756), .C2(new_n766), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n971), .ZN(new_n1159));
  AOI21_X1  g0959(.A(new_n973), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  NOR3_X1   g0960(.A1(new_n1160), .A2(new_n963), .A3(new_n980), .ZN(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n878), .B1(new_n885), .B2(new_n872), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n876), .A2(KEYINPUT106), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n1159), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n980), .B1(new_n1165), .B2(new_n924), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n977), .A2(new_n978), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n1167), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1169));
  NAND4_X1  g0969(.A1(new_n782), .A2(G330), .A3(new_n924), .A4(new_n872), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1170), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1169), .A2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n979), .B1(new_n972), .B2(new_n973), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(new_n1167), .ZN(new_n1174));
  NAND3_X1  g0974(.A1(new_n1174), .A2(new_n1170), .A3(new_n1162), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n782), .A2(G330), .A3(new_n872), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1176), .A2(new_n973), .ZN(new_n1177));
  AOI22_X1  g0977(.A1(new_n880), .A2(new_n1159), .B1(new_n1177), .B2(new_n1170), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1179));
  AND3_X1   g0979(.A1(new_n1177), .A2(new_n1170), .A3(new_n1179), .ZN(new_n1180));
  NOR2_X1   g0980(.A1(new_n1178), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n985), .ZN(new_n1182));
  NOR2_X1   g0982(.A1(new_n783), .A2(new_n475), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  NAND3_X1  g0984(.A1(new_n704), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  NOR2_X1   g0985(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1172), .A2(new_n1175), .A3(new_n1186), .ZN(new_n1187));
  OAI211_X1 g0987(.A(new_n986), .B(new_n1184), .C1(new_n1178), .C2(new_n1180), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1170), .B1(new_n1174), .B2(new_n1162), .ZN(new_n1189));
  AOI211_X1 g0989(.A(new_n1171), .B(new_n1161), .C1(new_n1173), .C2(new_n1167), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1187), .A2(new_n1191), .A3(new_n748), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n834), .A2(G87), .B1(new_n812), .B2(G68), .ZN(new_n1193));
  OAI221_X1 g0993(.A(new_n1193), .B1(new_n412), .B2(new_n826), .C1(new_n1017), .C2(new_n805), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n356), .B1(new_n907), .B2(G97), .ZN(new_n1195));
  OAI221_X1 g0995(.A(new_n1195), .B1(new_n543), .B2(new_n795), .C1(new_n819), .C2(new_n1097), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G107), .C2(new_n840), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(KEYINPUT54), .B(G143), .ZN(new_n1198));
  INV_X1    g0998(.A(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n251), .B1(new_n907), .B2(new_n1199), .ZN(new_n1200));
  INV_X1    g1000(.A(G125), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1200), .B1(new_n904), .B2(new_n795), .C1(new_n819), .C2(new_n1201), .ZN(new_n1202));
  NOR2_X1   g1002(.A1(new_n808), .A2(new_n1088), .ZN(new_n1203));
  XOR2_X1   g1003(.A(new_n1203), .B(KEYINPUT53), .Z(new_n1204));
  AOI22_X1  g1004(.A1(new_n827), .A2(G159), .B1(new_n812), .B2(G50), .ZN(new_n1205));
  INV_X1    g1005(.A(G128), .ZN(new_n1206));
  INV_X1    g1006(.A(G137), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1205), .B1(new_n1206), .B2(new_n805), .C1(new_n801), .C2(new_n1207), .ZN(new_n1208));
  NOR3_X1   g1008(.A1(new_n1202), .A2(new_n1204), .A3(new_n1208), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n792), .B1(new_n1197), .B2(new_n1209), .ZN(new_n1210));
  AOI21_X1  g1010(.A(new_n889), .B1(new_n280), .B2(new_n890), .ZN(new_n1211));
  OAI211_X1 g1011(.A(new_n1210), .B(new_n1211), .C1(new_n1168), .C2(new_n790), .ZN(new_n1212));
  INV_X1    g1012(.A(KEYINPUT116), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1189), .A2(new_n1190), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1213), .B1(new_n1214), .B2(new_n846), .ZN(new_n1215));
  NOR4_X1   g1015(.A1(new_n1189), .A2(new_n1190), .A3(KEYINPUT116), .A4(new_n845), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1192), .B(new_n1212), .C1(new_n1215), .C2(new_n1216), .ZN(G378));
  NOR3_X1   g1017(.A1(new_n1189), .A2(new_n1190), .A3(new_n1188), .ZN(new_n1218));
  AND2_X1   g1018(.A1(new_n981), .A2(new_n982), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1165), .A2(new_n924), .A3(new_n954), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(new_n925), .A2(new_n926), .B1(new_n953), .B2(new_n952), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(new_n946), .A2(new_n959), .B1(new_n389), .B2(new_n958), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n953), .B1(new_n1222), .B2(KEYINPUT38), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1223), .A2(new_n782), .A3(new_n872), .A4(new_n924), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n929), .A2(new_n1221), .B1(new_n1224), .B2(KEYINPUT40), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1219), .B(new_n1220), .C1(new_n1225), .C2(new_n918), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n295), .A2(new_n943), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n311), .B(new_n1227), .Z(new_n1228));
  XNOR2_X1  g1028(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1229));
  AND2_X1   g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT118), .ZN(new_n1232));
  NOR3_X1   g1032(.A1(new_n1230), .A2(new_n1231), .A3(new_n1232), .ZN(new_n1233));
  AOI21_X1  g1033(.A(new_n918), .B1(new_n955), .B2(new_n964), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1234), .B1(new_n975), .B2(new_n983), .ZN(new_n1235));
  AND3_X1   g1035(.A1(new_n1226), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1233), .B1(new_n1226), .B2(new_n1235), .ZN(new_n1237));
  OAI22_X1  g1037(.A1(new_n1218), .A2(new_n1185), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(KEYINPUT57), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  AOI211_X1 g1040(.A(new_n1183), .B(new_n985), .C1(new_n699), .C2(new_n703), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1187), .A2(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(new_n1233), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n965), .A2(G330), .ZN(new_n1244));
  NOR2_X1   g1044(.A1(new_n984), .A2(new_n1244), .ZN(new_n1245));
  NOR3_X1   g1045(.A1(new_n1234), .A2(new_n975), .A3(new_n983), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1243), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(new_n1226), .A2(new_n1233), .A3(new_n1235), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1242), .A2(new_n1249), .A3(KEYINPUT57), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1240), .A2(new_n748), .A3(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT119), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n845), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1253));
  NOR3_X1   g1053(.A1(new_n1230), .A2(new_n1231), .A3(new_n790), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n889), .B1(new_n216), .B2(new_n890), .ZN(new_n1255));
  NOR2_X1   g1055(.A1(G33), .A2(G41), .ZN(new_n1256));
  AOI211_X1 g1056(.A(G50), .B(new_n1256), .C1(new_n251), .C2(new_n262), .ZN(new_n1257));
  AOI211_X1 g1057(.A(G41), .B(new_n356), .C1(new_n796), .C2(G107), .ZN(new_n1258));
  OAI21_X1  g1058(.A(new_n1258), .B1(new_n415), .B2(new_n822), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1259), .B1(G283), .B2(new_n820), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n805), .A2(new_n543), .B1(new_n811), .B2(new_n202), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n1003), .B(new_n1261), .C1(G77), .C2(new_n834), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n1260), .B(new_n1262), .C1(new_n452), .C2(new_n801), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT58), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1257), .B1(new_n1263), .B2(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1265), .B1(new_n1264), .B2(new_n1263), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n795), .A2(new_n1206), .ZN(new_n1267));
  OAI22_X1  g1067(.A1(new_n805), .A2(new_n1201), .B1(new_n808), .B2(new_n1198), .ZN(new_n1268));
  AOI211_X1 g1068(.A(new_n1267), .B(new_n1268), .C1(G150), .C2(new_n827), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n840), .A2(G132), .B1(G137), .B2(new_n907), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1270), .A2(KEYINPUT117), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1270), .A2(KEYINPUT117), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1269), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  OR2_X1    g1074(.A1(new_n1274), .A2(KEYINPUT59), .ZN(new_n1275));
  INV_X1    g1075(.A(G124), .ZN(new_n1276));
  OAI221_X1 g1076(.A(new_n1256), .B1(new_n815), .B2(new_n1276), .C1(new_n323), .C2(new_n811), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(new_n1274), .B2(KEYINPUT59), .ZN(new_n1278));
  AOI21_X1  g1078(.A(new_n1266), .B1(new_n1275), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1255), .B1(new_n1279), .B2(new_n892), .ZN(new_n1280));
  NOR2_X1   g1080(.A1(new_n1254), .A2(new_n1280), .ZN(new_n1281));
  OAI21_X1  g1081(.A(new_n1252), .B1(new_n1253), .B2(new_n1281), .ZN(new_n1282));
  OAI21_X1  g1082(.A(new_n846), .B1(new_n1236), .B2(new_n1237), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1281), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1283), .A2(KEYINPUT119), .A3(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1282), .A2(new_n1285), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1251), .A2(new_n1286), .ZN(G375));
  NAND2_X1  g1087(.A1(new_n1181), .A2(new_n1185), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1288), .A2(new_n1188), .A3(new_n1081), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1177), .A2(new_n1170), .A3(new_n1179), .ZN(new_n1290));
  AND2_X1   g1090(.A1(new_n1177), .A2(new_n1170), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1290), .B1(new_n1291), .B2(new_n972), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n973), .A2(new_n789), .ZN(new_n1293));
  NOR3_X1   g1093(.A1(new_n792), .A2(G68), .A3(new_n789), .ZN(new_n1294));
  OAI221_X1 g1094(.A(new_n251), .B1(new_n822), .B2(new_n395), .C1(new_n1017), .C2(new_n795), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1295), .B1(new_n820), .B2(G303), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n840), .A2(new_n583), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1093), .B1(G77), .B2(new_n812), .ZN(new_n1298));
  AOI22_X1  g1098(.A1(G294), .A2(new_n906), .B1(new_n834), .B2(G97), .ZN(new_n1299));
  NAND4_X1  g1099(.A1(new_n1296), .A2(new_n1297), .A3(new_n1298), .A4(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(KEYINPUT120), .ZN(new_n1301));
  OR2_X1    g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1303));
  OAI221_X1 g1103(.A(new_n356), .B1(new_n822), .B2(new_n282), .C1(new_n811), .C2(new_n202), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n838), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1304), .B1(new_n1305), .B2(G137), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n820), .A2(G128), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n840), .A2(new_n1199), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n826), .A2(new_n216), .B1(new_n808), .B2(new_n323), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(G132), .B2(new_n906), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  NAND3_X1  g1111(.A1(new_n1302), .A2(new_n1303), .A3(new_n1311), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n889), .B(new_n1294), .C1(new_n1312), .C2(new_n792), .ZN(new_n1313));
  AOI22_X1  g1113(.A1(new_n1292), .A2(new_n846), .B1(new_n1293), .B2(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1289), .A2(new_n1314), .ZN(G381));
  AND2_X1   g1115(.A1(new_n1150), .A2(new_n1156), .ZN(new_n1316));
  INV_X1    g1116(.A(G384), .ZN(new_n1317));
  OAI211_X1 g1117(.A(new_n866), .B(new_n1121), .C1(new_n1123), .C2(new_n1124), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1318), .ZN(new_n1319));
  NAND3_X1  g1119(.A1(new_n1316), .A2(new_n1317), .A3(new_n1319), .ZN(new_n1320));
  NOR3_X1   g1120(.A1(G387), .A2(G381), .A3(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(G378), .ZN(new_n1322));
  AOI21_X1  g1122(.A(new_n749), .B1(new_n1238), .B2(new_n1239), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n1323), .A2(new_n1250), .B1(new_n1282), .B2(new_n1285), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1321), .A2(new_n1322), .A3(new_n1324), .ZN(new_n1325));
  XOR2_X1   g1125(.A(new_n1325), .B(KEYINPUT121), .Z(G407));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n726), .A3(new_n1322), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(G407), .A2(G213), .A3(new_n1327), .ZN(G409));
  NAND3_X1  g1128(.A1(new_n1075), .A2(new_n1086), .A3(new_n1316), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(G393), .A2(G396), .ZN(new_n1330));
  AOI22_X1  g1130(.A1(new_n1074), .A2(G390), .B1(new_n1318), .B2(new_n1330), .ZN(new_n1331));
  NAND2_X1  g1131(.A1(new_n1329), .A2(new_n1331), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1330), .A2(new_n1318), .ZN(new_n1333));
  INV_X1    g1133(.A(KEYINPUT125), .ZN(new_n1334));
  XNOR2_X1  g1134(.A(new_n1333), .B(new_n1334), .ZN(new_n1335));
  NOR2_X1   g1135(.A1(new_n1316), .A2(new_n1084), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1074), .A2(G390), .ZN(new_n1337));
  OAI21_X1  g1137(.A(new_n1335), .B1(new_n1336), .B2(new_n1337), .ZN(new_n1338));
  NAND2_X1  g1138(.A1(new_n1332), .A2(new_n1338), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1339), .ZN(new_n1340));
  INV_X1    g1140(.A(G213), .ZN(new_n1341));
  NOR2_X1   g1141(.A1(new_n1341), .A2(G343), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1342), .A2(G2897), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  NOR2_X1   g1144(.A1(new_n1241), .A2(new_n1292), .ZN(new_n1345));
  OAI21_X1  g1145(.A(KEYINPUT60), .B1(new_n1186), .B2(new_n1345), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT60), .ZN(new_n1347));
  AOI21_X1  g1147(.A(new_n749), .B1(new_n1288), .B2(new_n1347), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1346), .A2(new_n1348), .ZN(new_n1349));
  AOI21_X1  g1149(.A(G384), .B1(new_n1349), .B2(new_n1314), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n748), .B1(new_n1345), .B2(KEYINPUT60), .ZN(new_n1351));
  AOI21_X1  g1151(.A(new_n1347), .B1(new_n1288), .B2(new_n1188), .ZN(new_n1352));
  OAI211_X1 g1152(.A(G384), .B(new_n1314), .C1(new_n1351), .C2(new_n1352), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1353), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1344), .B1(new_n1350), .B2(new_n1354), .ZN(new_n1355));
  INV_X1    g1155(.A(KEYINPUT123), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1355), .A2(new_n1356), .ZN(new_n1357));
  OAI21_X1  g1157(.A(new_n1314), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1358), .A2(new_n1317), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1353), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(KEYINPUT123), .A3(new_n1344), .ZN(new_n1361));
  NAND3_X1  g1161(.A1(new_n1359), .A2(new_n1353), .A3(new_n1343), .ZN(new_n1362));
  INV_X1    g1162(.A(KEYINPUT122), .ZN(new_n1363));
  NAND2_X1  g1163(.A1(new_n1362), .A2(new_n1363), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1359), .A2(KEYINPUT122), .A3(new_n1353), .A4(new_n1343), .ZN(new_n1365));
  AOI22_X1  g1165(.A1(new_n1357), .A2(new_n1361), .B1(new_n1364), .B2(new_n1365), .ZN(new_n1366));
  NOR2_X1   g1166(.A1(new_n1253), .A2(new_n1281), .ZN(new_n1367));
  NAND3_X1  g1167(.A1(new_n1242), .A2(new_n1249), .A3(new_n1081), .ZN(new_n1368));
  AOI21_X1  g1168(.A(G378), .B1(new_n1367), .B2(new_n1368), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1369), .B1(new_n1324), .B2(G378), .ZN(new_n1370));
  OAI21_X1  g1170(.A(new_n1366), .B1(new_n1370), .B2(new_n1342), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1251), .A2(new_n1286), .A3(G378), .ZN(new_n1372));
  NAND2_X1  g1172(.A1(new_n1367), .A2(new_n1368), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1322), .A2(new_n1373), .ZN(new_n1374));
  NAND2_X1  g1174(.A1(new_n1372), .A2(new_n1374), .ZN(new_n1375));
  INV_X1    g1175(.A(new_n1342), .ZN(new_n1376));
  INV_X1    g1176(.A(new_n1360), .ZN(new_n1377));
  XOR2_X1   g1177(.A(KEYINPUT127), .B(KEYINPUT62), .Z(new_n1378));
  NAND4_X1  g1178(.A1(new_n1375), .A2(new_n1376), .A3(new_n1377), .A4(new_n1378), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT61), .ZN(new_n1380));
  NAND3_X1  g1180(.A1(new_n1371), .A2(new_n1379), .A3(new_n1380), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(KEYINPUT127), .A2(KEYINPUT62), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1342), .B1(new_n1372), .B2(new_n1374), .ZN(new_n1383));
  AOI21_X1  g1183(.A(new_n1382), .B1(new_n1383), .B2(new_n1377), .ZN(new_n1384));
  OAI21_X1  g1184(.A(new_n1340), .B1(new_n1381), .B2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(new_n1364), .A2(new_n1365), .ZN(new_n1386));
  AOI21_X1  g1186(.A(KEYINPUT123), .B1(new_n1360), .B2(new_n1344), .ZN(new_n1387));
  AOI211_X1 g1187(.A(new_n1356), .B(new_n1343), .C1(new_n1359), .C2(new_n1353), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1386), .B1(new_n1387), .B2(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1389), .A2(KEYINPUT124), .ZN(new_n1390));
  INV_X1    g1190(.A(new_n1383), .ZN(new_n1391));
  INV_X1    g1191(.A(KEYINPUT124), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1366), .A2(new_n1392), .ZN(new_n1393));
  NAND3_X1  g1193(.A1(new_n1390), .A2(new_n1391), .A3(new_n1393), .ZN(new_n1394));
  NAND2_X1  g1194(.A1(new_n1383), .A2(new_n1377), .ZN(new_n1395));
  INV_X1    g1195(.A(KEYINPUT63), .ZN(new_n1396));
  NAND2_X1  g1196(.A1(new_n1395), .A2(new_n1396), .ZN(new_n1397));
  NAND3_X1  g1197(.A1(new_n1383), .A2(KEYINPUT63), .A3(new_n1377), .ZN(new_n1398));
  INV_X1    g1198(.A(KEYINPUT126), .ZN(new_n1399));
  AOI21_X1  g1199(.A(new_n1399), .B1(new_n1339), .B2(new_n1380), .ZN(new_n1400));
  AOI211_X1 g1200(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1332), .C2(new_n1338), .ZN(new_n1401));
  NOR2_X1   g1201(.A1(new_n1400), .A2(new_n1401), .ZN(new_n1402));
  NAND4_X1  g1202(.A1(new_n1394), .A2(new_n1397), .A3(new_n1398), .A4(new_n1402), .ZN(new_n1403));
  NAND2_X1  g1203(.A1(new_n1385), .A2(new_n1403), .ZN(G405));
  NAND2_X1  g1204(.A1(G375), .A2(new_n1322), .ZN(new_n1405));
  NAND2_X1  g1205(.A1(new_n1405), .A2(new_n1372), .ZN(new_n1406));
  NAND2_X1  g1206(.A1(new_n1406), .A2(new_n1377), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1405), .A2(new_n1372), .A3(new_n1360), .ZN(new_n1408));
  NAND2_X1  g1208(.A1(new_n1407), .A2(new_n1408), .ZN(new_n1409));
  XNOR2_X1  g1209(.A(new_n1409), .B(new_n1340), .ZN(G402));
endmodule


