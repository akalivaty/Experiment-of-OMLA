//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 0 0 0 0 1 1 1 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n725, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n984, new_n985,
    new_n986, new_n987, new_n988, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  XNOR2_X1  g001(.A(new_n187), .B(KEYINPUT80), .ZN(new_n188));
  OAI21_X1  g002(.A(G210), .B1(G237), .B2(G902), .ZN(new_n189));
  INV_X1    g003(.A(new_n189), .ZN(new_n190));
  INV_X1    g004(.A(G224), .ZN(new_n191));
  NOR2_X1   g005(.A1(new_n191), .A2(G953), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n193), .A2(KEYINPUT7), .ZN(new_n194));
  INV_X1    g008(.A(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G146), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G143), .ZN(new_n197));
  INV_X1    g011(.A(G143), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G146), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(KEYINPUT66), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(KEYINPUT66), .A2(G128), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(G143), .B2(new_n196), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(KEYINPUT67), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(G128), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(KEYINPUT1), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n210), .A2(new_n197), .A3(new_n199), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT65), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  XNOR2_X1  g027(.A(G143), .B(G146), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n214), .A2(KEYINPUT65), .A3(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  OAI211_X1 g031(.A(KEYINPUT67), .B(new_n200), .C1(new_n203), .C2(new_n205), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n208), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT83), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT0), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n214), .B1(new_n223), .B2(new_n209), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT0), .B(G128), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n200), .A2(new_n225), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n224), .A2(new_n226), .A3(G125), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n227), .B1(new_n219), .B2(new_n220), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n195), .B1(new_n222), .B2(new_n228), .ZN(new_n229));
  AOI21_X1  g043(.A(KEYINPUT65), .B1(new_n214), .B2(new_n210), .ZN(new_n230));
  AND4_X1   g044(.A1(KEYINPUT65), .A2(new_n210), .A3(new_n197), .A4(new_n199), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n218), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n197), .A2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n233), .B1(new_n202), .B2(new_n201), .ZN(new_n234));
  AOI21_X1  g048(.A(KEYINPUT67), .B1(new_n234), .B2(new_n200), .ZN(new_n235));
  NOR2_X1   g049(.A1(new_n232), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n236), .A2(KEYINPUT83), .A3(new_n217), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n237), .A2(new_n221), .A3(new_n227), .A4(new_n194), .ZN(new_n238));
  NAND2_X1  g052(.A1(new_n229), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(G119), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G116), .ZN(new_n241));
  INV_X1    g055(.A(G116), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G119), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT2), .B(G113), .ZN(new_n245));
  OAI21_X1  g059(.A(KEYINPUT68), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g060(.A(G116), .B(G119), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT68), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT2), .ZN(new_n249));
  NOR2_X1   g063(.A1(new_n249), .A2(G113), .ZN(new_n250));
  INV_X1    g064(.A(G113), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n251), .A2(KEYINPUT2), .ZN(new_n252));
  OAI211_X1 g066(.A(new_n247), .B(new_n248), .C1(new_n250), .C2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n246), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n244), .A2(new_n255), .ZN(new_n256));
  OAI21_X1  g070(.A(G113), .B1(new_n241), .B2(KEYINPUT5), .ZN(new_n257));
  OAI21_X1  g071(.A(KEYINPUT81), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  INV_X1    g072(.A(G107), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n259), .A2(KEYINPUT76), .A3(G104), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n260), .A2(KEYINPUT3), .ZN(new_n261));
  INV_X1    g075(.A(G101), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT3), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n263), .A2(new_n259), .A3(KEYINPUT76), .A4(G104), .ZN(new_n264));
  INV_X1    g078(.A(G104), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G107), .ZN(new_n266));
  NAND4_X1  g080(.A1(new_n261), .A2(new_n262), .A3(new_n264), .A4(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n265), .A2(G107), .ZN(new_n268));
  NOR2_X1   g082(.A1(new_n259), .A2(G104), .ZN(new_n269));
  OAI21_X1  g083(.A(G101), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n267), .A2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(new_n257), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n247), .A2(KEYINPUT5), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT81), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n272), .A2(new_n273), .A3(new_n274), .ZN(new_n275));
  AND4_X1   g089(.A1(new_n254), .A2(new_n258), .A3(new_n271), .A4(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(G122), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(G110), .ZN(new_n280));
  INV_X1    g094(.A(G110), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G122), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT82), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n283), .B1(new_n280), .B2(new_n282), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n278), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n280), .A2(new_n282), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT82), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(new_n284), .A3(new_n277), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n287), .A2(new_n290), .ZN(new_n291));
  AOI22_X1  g105(.A1(new_n246), .A2(new_n253), .B1(new_n273), .B2(new_n272), .ZN(new_n292));
  OAI21_X1  g106(.A(new_n291), .B1(new_n292), .B2(new_n271), .ZN(new_n293));
  NOR2_X1   g107(.A1(new_n276), .A2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n261), .A2(new_n264), .A3(new_n266), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G101), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT77), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(KEYINPUT77), .A3(G101), .ZN(new_n299));
  NAND4_X1  g113(.A1(new_n298), .A2(KEYINPUT4), .A3(new_n267), .A4(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n244), .A2(new_n245), .ZN(new_n301));
  AOI21_X1  g115(.A(new_n269), .B1(KEYINPUT3), .B2(new_n260), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n262), .B1(new_n302), .B2(new_n264), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT4), .ZN(new_n304));
  AOI22_X1  g118(.A1(new_n254), .A2(new_n301), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  AND3_X1   g119(.A1(new_n258), .A2(new_n254), .A3(new_n275), .ZN(new_n306));
  INV_X1    g120(.A(new_n271), .ZN(new_n307));
  AOI22_X1  g121(.A1(new_n300), .A2(new_n305), .B1(new_n306), .B2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n285), .A2(new_n286), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n294), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n239), .A2(new_n311), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n312), .A2(KEYINPUT85), .A3(new_n313), .ZN(new_n314));
  NAND4_X1  g128(.A1(new_n307), .A2(new_n254), .A3(new_n258), .A4(new_n275), .ZN(new_n315));
  INV_X1    g129(.A(new_n305), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n299), .A2(KEYINPUT4), .A3(new_n267), .ZN(new_n317));
  NOR2_X1   g131(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI21_X1  g133(.A(new_n315), .B1(new_n316), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(new_n309), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n308), .A2(new_n310), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(new_n322), .A3(KEYINPUT6), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n308), .A2(KEYINPUT6), .A3(new_n310), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n192), .B1(new_n222), .B2(new_n228), .ZN(new_n325));
  NAND4_X1  g139(.A1(new_n237), .A2(new_n221), .A3(new_n227), .A4(new_n193), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n314), .A2(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(KEYINPUT85), .B1(new_n312), .B2(new_n313), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n190), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n312), .A2(new_n313), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT85), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  NAND4_X1  g148(.A1(new_n334), .A2(new_n189), .A3(new_n328), .A4(new_n314), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n188), .B1(new_n331), .B2(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(G469), .ZN(new_n337));
  OAI21_X1  g151(.A(new_n200), .B1(new_n205), .B2(new_n209), .ZN(new_n338));
  OAI21_X1  g152(.A(new_n338), .B1(new_n230), .B2(new_n231), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n307), .A2(new_n339), .ZN(new_n340));
  NAND4_X1  g154(.A1(new_n271), .A2(new_n208), .A3(new_n216), .A4(new_n218), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(KEYINPUT11), .ZN(new_n343));
  INV_X1    g157(.A(G134), .ZN(new_n344));
  OAI21_X1  g158(.A(new_n343), .B1(new_n344), .B2(G137), .ZN(new_n345));
  INV_X1    g159(.A(G137), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n346), .A2(KEYINPUT11), .A3(G134), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n344), .A2(G137), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n347), .A3(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(G131), .ZN(new_n350));
  INV_X1    g164(.A(G131), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n345), .A2(new_n347), .A3(new_n351), .A4(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g167(.A(KEYINPUT12), .B1(new_n342), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT12), .ZN(new_n355));
  INV_X1    g169(.A(new_n353), .ZN(new_n356));
  AOI211_X1 g170(.A(new_n355), .B(new_n356), .C1(new_n340), .C2(new_n341), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  AOI22_X1  g172(.A1(new_n303), .A2(new_n304), .B1(new_n226), .B2(new_n224), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n359), .B1(new_n317), .B2(new_n318), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT78), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n353), .B(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n214), .B1(G128), .B2(new_n233), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n364), .B1(new_n213), .B2(new_n215), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n365), .B2(new_n271), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n208), .A2(new_n216), .A3(new_n218), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n367), .A2(KEYINPUT10), .A3(new_n307), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n360), .A2(new_n362), .A3(new_n366), .A4(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(G110), .B(G140), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n370), .B(KEYINPUT75), .ZN(new_n371));
  INV_X1    g185(.A(G953), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n372), .A2(G227), .ZN(new_n373));
  XNOR2_X1  g187(.A(new_n371), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n358), .A2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n360), .A2(new_n366), .A3(new_n368), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n353), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n374), .B1(new_n378), .B2(new_n369), .ZN(new_n379));
  OAI211_X1 g193(.A(new_n337), .B(new_n313), .C1(new_n376), .C2(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G469), .A2(G902), .ZN(new_n381));
  OAI21_X1  g195(.A(new_n369), .B1(new_n354), .B2(new_n357), .ZN(new_n382));
  INV_X1    g196(.A(new_n374), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n378), .A2(new_n369), .A3(new_n374), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n384), .A2(G469), .A3(new_n385), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n380), .A2(new_n381), .A3(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT9), .B(G234), .ZN(new_n388));
  OAI21_X1  g202(.A(G221), .B1(new_n388), .B2(G902), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT79), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n387), .A2(KEYINPUT79), .A3(new_n389), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n336), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(G140), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G125), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n217), .A2(G140), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n396), .A2(new_n397), .A3(KEYINPUT16), .ZN(new_n398));
  OR3_X1    g212(.A1(new_n217), .A2(KEYINPUT16), .A3(G140), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n398), .A2(new_n399), .A3(G146), .ZN(new_n400));
  XNOR2_X1  g214(.A(G125), .B(G140), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n196), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT66), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n209), .ZN(new_n404));
  NAND2_X1  g218(.A1(KEYINPUT66), .A2(G128), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n404), .A2(KEYINPUT23), .A3(G119), .A4(new_n405), .ZN(new_n406));
  OAI21_X1  g220(.A(KEYINPUT23), .B1(new_n209), .B2(G119), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n209), .A2(G119), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND3_X1   g223(.A1(new_n406), .A2(new_n409), .A3(new_n281), .ZN(new_n410));
  XOR2_X1   g224(.A(KEYINPUT24), .B(G110), .Z(new_n411));
  NAND3_X1  g225(.A1(new_n404), .A2(G119), .A3(new_n405), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n240), .A2(G128), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n411), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  OAI211_X1 g228(.A(new_n400), .B(new_n402), .C1(new_n410), .C2(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(KEYINPUT72), .ZN(new_n416));
  AND3_X1   g230(.A1(new_n406), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n416), .B1(new_n406), .B2(new_n409), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n417), .A2(new_n418), .A3(new_n281), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n412), .A3(new_n413), .ZN(new_n420));
  AND3_X1   g234(.A1(new_n398), .A2(G146), .A3(new_n399), .ZN(new_n421));
  AOI21_X1  g235(.A(G146), .B1(new_n398), .B2(new_n399), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n420), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n415), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(KEYINPUT22), .B(G137), .ZN(new_n425));
  NAND3_X1  g239(.A1(new_n372), .A2(G221), .A3(G234), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n425), .B(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g243(.A(new_n415), .B(new_n427), .C1(new_n419), .C2(new_n423), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n429), .A2(new_n313), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT25), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT25), .ZN(new_n433));
  NAND4_X1  g247(.A1(new_n429), .A2(new_n433), .A3(new_n313), .A4(new_n430), .ZN(new_n434));
  XOR2_X1   g248(.A(KEYINPUT71), .B(G217), .Z(new_n435));
  AOI21_X1  g249(.A(new_n435), .B1(G234), .B2(new_n313), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n432), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT73), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n432), .A2(KEYINPUT73), .A3(new_n434), .A4(new_n436), .ZN(new_n440));
  NOR2_X1   g254(.A1(new_n436), .A2(G902), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n429), .A2(new_n430), .A3(new_n441), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(KEYINPUT74), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n439), .A2(new_n440), .A3(new_n443), .ZN(new_n444));
  NOR2_X1   g258(.A1(G237), .A2(G953), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G210), .ZN(new_n446));
  XNOR2_X1  g260(.A(new_n446), .B(KEYINPUT27), .ZN(new_n447));
  XNOR2_X1  g261(.A(KEYINPUT26), .B(G101), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  NOR2_X1   g263(.A1(new_n344), .A2(G137), .ZN(new_n450));
  NOR2_X1   g264(.A1(new_n346), .A2(G134), .ZN(new_n451));
  OAI21_X1  g265(.A(G131), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n352), .A2(new_n452), .ZN(new_n453));
  INV_X1    g267(.A(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n454), .B1(new_n232), .B2(new_n235), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n254), .A2(new_n301), .ZN(new_n456));
  INV_X1    g270(.A(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n224), .A2(new_n226), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n353), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n455), .A2(new_n457), .A3(new_n459), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n460), .B(KEYINPUT28), .ZN(new_n461));
  OR2_X1    g275(.A1(new_n453), .A2(KEYINPUT64), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n453), .A2(KEYINPUT64), .ZN(new_n463));
  NAND3_X1  g277(.A1(new_n367), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n459), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(new_n456), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n449), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT31), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n460), .A2(new_n449), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(KEYINPUT69), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT69), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n460), .A2(new_n471), .A3(new_n449), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n455), .A2(new_n459), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(KEYINPUT30), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT30), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n464), .A2(new_n476), .A3(new_n459), .ZN(new_n477));
  AOI21_X1  g291(.A(new_n457), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g292(.A(new_n468), .B1(new_n473), .B2(new_n478), .ZN(new_n479));
  AND3_X1   g293(.A1(new_n460), .A2(new_n471), .A3(new_n449), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n471), .B1(new_n460), .B2(new_n449), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n475), .A2(new_n477), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n456), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n482), .A2(KEYINPUT31), .A3(new_n484), .ZN(new_n485));
  AOI21_X1  g299(.A(new_n467), .B1(new_n479), .B2(new_n485), .ZN(new_n486));
  NOR2_X1   g300(.A1(G472), .A2(G902), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n487), .B(KEYINPUT70), .ZN(new_n488));
  OAI21_X1  g302(.A(KEYINPUT32), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  INV_X1    g303(.A(new_n467), .ZN(new_n490));
  AOI21_X1  g304(.A(KEYINPUT31), .B1(new_n482), .B2(new_n484), .ZN(new_n491));
  NOR4_X1   g305(.A1(new_n478), .A2(new_n480), .A3(new_n481), .A4(new_n468), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n490), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT32), .ZN(new_n494));
  INV_X1    g308(.A(new_n488), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n489), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n474), .A2(new_n456), .ZN(new_n498));
  AND2_X1   g312(.A1(new_n461), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(new_n449), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT29), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G902), .B1(new_n499), .B2(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n461), .A2(new_n466), .A3(new_n449), .ZN(new_n504));
  INV_X1    g318(.A(new_n460), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n478), .A2(new_n505), .ZN(new_n506));
  OAI211_X1 g320(.A(new_n504), .B(new_n501), .C1(new_n506), .C2(new_n449), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n503), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G472), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n444), .B1(new_n497), .B2(new_n509), .ZN(new_n510));
  NOR3_X1   g324(.A1(new_n201), .A2(new_n202), .A3(new_n198), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n209), .A2(G143), .ZN(new_n512));
  OAI21_X1  g326(.A(KEYINPUT90), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n404), .A2(G143), .A3(new_n405), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT90), .ZN(new_n515));
  INV_X1    g329(.A(new_n512), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n513), .A2(new_n344), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n279), .A2(G116), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n242), .A2(G122), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  XNOR2_X1  g335(.A(new_n521), .B(G107), .ZN(new_n522));
  AND2_X1   g336(.A1(new_n512), .A2(KEYINPUT13), .ZN(new_n523));
  NOR2_X1   g337(.A1(new_n512), .A2(KEYINPUT13), .ZN(new_n524));
  NOR3_X1   g338(.A1(new_n523), .A2(new_n511), .A3(new_n524), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n518), .B(new_n522), .C1(new_n344), .C2(new_n525), .ZN(new_n526));
  NOR3_X1   g340(.A1(new_n435), .A2(G953), .A3(new_n388), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT91), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n515), .B1(new_n514), .B2(new_n516), .ZN(new_n530));
  OAI21_X1  g344(.A(G134), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n518), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n259), .B1(new_n519), .B2(KEYINPUT14), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n533), .B(new_n521), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n528), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  AOI211_X1 g350(.A(KEYINPUT91), .B(new_n534), .C1(new_n531), .C2(new_n518), .ZN(new_n537));
  OAI211_X1 g351(.A(new_n526), .B(new_n527), .C1(new_n536), .C2(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT92), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n529), .A2(new_n530), .A3(G134), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n344), .B1(new_n513), .B2(new_n517), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n535), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(KEYINPUT91), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n532), .A2(new_n528), .A3(new_n535), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT92), .ZN(new_n546));
  NAND4_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n526), .A4(new_n527), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n526), .B1(new_n536), .B2(new_n537), .ZN(new_n548));
  INV_X1    g362(.A(new_n527), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n539), .A2(new_n547), .A3(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(G478), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(KEYINPUT15), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n555));
  OAI21_X1  g369(.A(new_n313), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n556), .B1(new_n555), .B2(new_n554), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n551), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(KEYINPUT94), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n313), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n553), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT94), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n551), .A2(new_n562), .A3(new_n557), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n559), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(G234), .A2(G237), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n565), .A2(G952), .A3(new_n372), .ZN(new_n566));
  INV_X1    g380(.A(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n565), .A2(G902), .A3(G953), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT21), .B(G898), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n569), .B2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(new_n571), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n445), .A2(G214), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n573), .A2(new_n198), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n445), .A2(G143), .A3(G214), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT87), .B1(new_n576), .B2(G131), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT17), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n576), .A2(G131), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT87), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n574), .A2(new_n580), .A3(new_n351), .A4(new_n575), .ZN(new_n581));
  NAND4_X1  g395(.A1(new_n577), .A2(new_n578), .A3(new_n579), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n421), .A2(new_n422), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n576), .A2(KEYINPUT17), .A3(G131), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n582), .A2(new_n583), .A3(new_n584), .ZN(new_n585));
  XNOR2_X1  g399(.A(G113), .B(G122), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(new_n265), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT86), .ZN(new_n588));
  NAND2_X1  g402(.A1(KEYINPUT18), .A2(G131), .ZN(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n588), .B1(new_n576), .B2(new_n590), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n574), .A2(KEYINPUT86), .A3(new_n575), .A4(new_n589), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  OR2_X1    g407(.A1(new_n401), .A2(new_n196), .ZN(new_n594));
  AOI22_X1  g408(.A1(new_n594), .A2(new_n402), .B1(new_n576), .B2(new_n590), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n585), .A2(new_n587), .A3(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n587), .B1(new_n585), .B2(new_n596), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n313), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G475), .ZN(new_n601));
  INV_X1    g415(.A(new_n587), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n577), .A2(new_n579), .A3(new_n581), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n401), .B(KEYINPUT19), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n421), .B1(new_n604), .B2(new_n196), .ZN(new_n605));
  AND2_X1   g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  AND2_X1   g420(.A1(new_n593), .A2(new_n595), .ZN(new_n607));
  OAI211_X1 g421(.A(KEYINPUT88), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT88), .ZN(new_n609));
  AOI22_X1  g423(.A1(new_n603), .A2(new_n605), .B1(new_n593), .B2(new_n595), .ZN(new_n610));
  OAI21_X1  g424(.A(new_n609), .B1(new_n610), .B2(new_n587), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n611), .A3(new_n597), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT20), .ZN(new_n613));
  NOR2_X1   g427(.A1(G475), .A2(G902), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT89), .ZN(new_n615));
  AND3_X1   g429(.A1(new_n612), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n613), .B1(new_n612), .B2(new_n615), .ZN(new_n617));
  OAI211_X1 g431(.A(new_n572), .B(new_n601), .C1(new_n616), .C2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT95), .B1(new_n564), .B2(new_n618), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n551), .A2(new_n557), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n620), .A2(new_n562), .B1(new_n560), .B2(new_n553), .ZN(new_n621));
  INV_X1    g435(.A(new_n618), .ZN(new_n622));
  INV_X1    g436(.A(KEYINPUT95), .ZN(new_n623));
  NAND4_X1  g437(.A1(new_n621), .A2(new_n622), .A3(new_n623), .A4(new_n559), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n619), .A2(new_n624), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n394), .A2(new_n510), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(G101), .ZN(G3));
  NAND2_X1  g441(.A1(new_n392), .A2(new_n393), .ZN(new_n628));
  OAI21_X1  g442(.A(G472), .B1(new_n486), .B2(G902), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n493), .A2(new_n495), .ZN(new_n630));
  INV_X1    g444(.A(new_n444), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n628), .A2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT33), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n548), .B2(new_n549), .ZN(new_n635));
  AOI22_X1  g449(.A1(new_n551), .A2(new_n634), .B1(new_n538), .B2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n552), .B1(new_n636), .B2(new_n313), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n551), .A2(new_n552), .A3(new_n313), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  OAI21_X1  g453(.A(KEYINPUT96), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g454(.A1(new_n616), .A2(new_n617), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n601), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT96), .ZN(new_n643));
  AOI221_X4 g457(.A(G902), .B1(new_n538), .B2(new_n635), .C1(new_n551), .C2(new_n634), .ZN(new_n644));
  OAI211_X1 g458(.A(new_n638), .B(new_n643), .C1(new_n644), .C2(new_n552), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n640), .A2(new_n642), .A3(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n187), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n331), .B2(new_n335), .ZN(new_n648));
  AND2_X1   g462(.A1(new_n648), .A2(new_n572), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n633), .A2(new_n646), .A3(new_n649), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT34), .B(G104), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G6));
  INV_X1    g466(.A(KEYINPUT97), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n601), .A2(new_n653), .ZN(new_n654));
  NAND3_X1  g468(.A1(new_n600), .A2(KEYINPUT97), .A3(G475), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n654), .B(new_n655), .C1(new_n616), .C2(new_n617), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n571), .B(KEYINPUT98), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n656), .A2(new_n658), .ZN(new_n659));
  AND3_X1   g473(.A1(new_n648), .A2(new_n564), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n633), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(new_n259), .ZN(new_n662));
  XNOR2_X1  g476(.A(KEYINPUT99), .B(KEYINPUT35), .ZN(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  NAND2_X1  g478(.A1(new_n629), .A2(new_n630), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n428), .A2(KEYINPUT36), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT100), .ZN(new_n667));
  INV_X1    g481(.A(new_n424), .ZN(new_n668));
  OR2_X1    g482(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n667), .A2(new_n668), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n669), .A2(new_n441), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g485(.A1(new_n439), .A2(new_n440), .A3(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT101), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n439), .A2(KEYINPUT101), .A3(new_n440), .A4(new_n671), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n665), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n394), .A2(new_n625), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n678), .B(new_n679), .ZN(G12));
  AOI21_X1  g494(.A(new_n676), .B1(new_n497), .B2(new_n509), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n387), .A2(KEYINPUT79), .A3(new_n389), .ZN(new_n682));
  AOI21_X1  g496(.A(KEYINPUT79), .B1(new_n387), .B2(new_n389), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g498(.A(new_n564), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n566), .B1(new_n568), .B2(G900), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n641), .A2(new_n654), .A3(new_n655), .A4(new_n686), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n681), .A2(new_n684), .A3(new_n648), .A4(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XNOR2_X1  g504(.A(new_n686), .B(KEYINPUT39), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n684), .A2(new_n691), .ZN(new_n692));
  XOR2_X1   g506(.A(new_n692), .B(KEYINPUT40), .Z(new_n693));
  NAND2_X1  g507(.A1(new_n331), .A2(new_n335), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(KEYINPUT38), .ZN(new_n695));
  INV_X1    g509(.A(G472), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n482), .A2(new_n484), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n498), .A2(new_n460), .ZN(new_n698));
  OAI21_X1  g512(.A(new_n697), .B1(new_n449), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g513(.A(new_n696), .B1(new_n699), .B2(new_n313), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n672), .B1(new_n497), .B2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(new_n642), .ZN(new_n703));
  NOR3_X1   g517(.A1(new_n685), .A2(new_n703), .A3(new_n647), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n693), .A2(new_n695), .A3(new_n702), .A4(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G143), .ZN(G45));
  AOI21_X1  g520(.A(new_n494), .B1(new_n493), .B2(new_n495), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n486), .A2(KEYINPUT32), .A3(new_n488), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n509), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n676), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n684), .A2(new_n709), .A3(new_n648), .A4(new_n710), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n640), .A2(new_n645), .A3(new_n642), .A4(new_n686), .ZN(new_n712));
  NOR2_X1   g526(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(new_n196), .ZN(G48));
  INV_X1    g528(.A(new_n389), .ZN(new_n715));
  OAI21_X1  g529(.A(new_n313), .B1(new_n376), .B2(new_n379), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n716), .A2(G469), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n717), .A2(KEYINPUT102), .A3(new_n380), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT102), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n716), .A2(new_n719), .A3(G469), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n715), .B1(new_n718), .B2(new_n720), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n646), .A2(new_n510), .A3(new_n649), .A4(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(KEYINPUT41), .B(G113), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n722), .B(new_n723), .ZN(G15));
  NAND3_X1  g538(.A1(new_n660), .A2(new_n510), .A3(new_n721), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G116), .ZN(G18));
  AND2_X1   g540(.A1(new_n721), .A2(new_n648), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n727), .A2(new_n625), .A3(new_n681), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  AND3_X1   g543(.A1(new_n694), .A2(new_n564), .A3(new_n187), .ZN(new_n730));
  AOI211_X1 g544(.A(new_n715), .B(new_n658), .C1(new_n718), .C2(new_n720), .ZN(new_n731));
  OAI22_X1  g545(.A1(new_n491), .A2(new_n492), .B1(new_n449), .B2(new_n499), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n732), .A2(new_n495), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n629), .A2(new_n733), .A3(new_n631), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n730), .A2(new_n642), .A3(new_n731), .A4(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AND4_X1   g550(.A1(new_n642), .A2(new_n640), .A3(new_n645), .A4(new_n686), .ZN(new_n737));
  AND3_X1   g551(.A1(new_n629), .A2(new_n733), .A3(new_n672), .ZN(new_n738));
  AND3_X1   g552(.A1(new_n738), .A2(new_n648), .A3(new_n721), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n740), .B(G125), .ZN(G27));
  NAND3_X1  g555(.A1(new_n331), .A2(new_n335), .A3(new_n187), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT103), .ZN(new_n743));
  AND3_X1   g557(.A1(new_n387), .A2(new_n743), .A3(new_n389), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n743), .B1(new_n387), .B2(new_n389), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT42), .ZN(new_n746));
  NOR4_X1   g560(.A1(new_n742), .A2(new_n744), .A3(new_n745), .A4(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT104), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n497), .A2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n489), .A2(new_n496), .A3(KEYINPUT104), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n509), .A3(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n737), .A2(new_n747), .A3(new_n751), .A4(new_n631), .ZN(new_n752));
  NOR2_X1   g566(.A1(new_n744), .A2(new_n745), .ZN(new_n753));
  AND3_X1   g567(.A1(new_n331), .A2(new_n335), .A3(new_n187), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n753), .A2(new_n709), .A3(new_n631), .A4(new_n754), .ZN(new_n755));
  OAI21_X1  g569(.A(new_n746), .B1(new_n755), .B2(new_n712), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n752), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  INV_X1    g572(.A(new_n755), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n688), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NAND2_X1  g575(.A1(new_n640), .A2(new_n645), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n762), .A2(new_n642), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT43), .ZN(new_n764));
  OAI21_X1  g578(.A(new_n764), .B1(new_n642), .B2(KEYINPUT106), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n763), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n665), .A2(new_n672), .ZN(new_n769));
  INV_X1    g583(.A(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n768), .A2(KEYINPUT44), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n742), .B(KEYINPUT107), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(KEYINPUT108), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT108), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n771), .A2(new_n775), .A3(new_n772), .ZN(new_n776));
  AOI21_X1  g590(.A(KEYINPUT44), .B1(new_n768), .B2(new_n770), .ZN(new_n777));
  AOI21_X1  g591(.A(KEYINPUT45), .B1(new_n384), .B2(new_n385), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n778), .A2(new_n337), .ZN(new_n779));
  NAND3_X1  g593(.A1(new_n384), .A2(KEYINPUT45), .A3(new_n385), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n381), .ZN(new_n782));
  INV_X1    g596(.A(new_n380), .ZN(new_n783));
  NOR2_X1   g597(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n381), .ZN(new_n785));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n786));
  AND2_X1   g600(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g601(.A1(new_n785), .A2(new_n786), .ZN(new_n788));
  OAI21_X1  g602(.A(new_n784), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  AND3_X1   g603(.A1(new_n789), .A2(new_n389), .A3(new_n691), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  NOR2_X1   g605(.A1(new_n777), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n774), .A2(new_n776), .A3(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G137), .ZN(G39));
  NAND2_X1  g608(.A1(new_n789), .A2(new_n389), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT47), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n795), .B(new_n796), .ZN(new_n797));
  NOR4_X1   g611(.A1(new_n712), .A2(new_n709), .A3(new_n631), .A4(new_n742), .ZN(new_n798));
  OR2_X1    g612(.A1(new_n798), .A2(KEYINPUT109), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n798), .A2(KEYINPUT109), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n797), .A2(new_n799), .A3(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT110), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n797), .A2(KEYINPUT110), .A3(new_n799), .A4(new_n800), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(G140), .ZN(G42));
  AND3_X1   g620(.A1(new_n768), .A2(new_n567), .A3(new_n734), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n727), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n372), .A2(G952), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n754), .A2(new_n721), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n497), .A2(new_n701), .ZN(new_n812));
  NOR4_X1   g626(.A1(new_n811), .A2(new_n812), .A3(new_n444), .A4(new_n566), .ZN(new_n813));
  AOI21_X1  g627(.A(new_n810), .B1(new_n813), .B2(new_n646), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n808), .A2(new_n809), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n809), .B1(new_n808), .B2(new_n814), .ZN(new_n816));
  AOI211_X1 g630(.A(new_n566), .B(new_n811), .C1(new_n766), .C2(new_n767), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n751), .A2(new_n631), .ZN(new_n818));
  AOI21_X1  g632(.A(KEYINPUT48), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n817), .A2(KEYINPUT48), .A3(new_n818), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n815), .A2(new_n816), .A3(new_n819), .A4(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT51), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n718), .A2(new_n720), .ZN(new_n823));
  NOR4_X1   g637(.A1(new_n695), .A2(new_n187), .A3(new_n715), .A4(new_n823), .ZN(new_n824));
  NAND2_X1  g638(.A1(new_n807), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT50), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n823), .A2(new_n389), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n807), .B(new_n772), .C1(new_n797), .C2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n817), .A2(new_n738), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n813), .A2(new_n703), .A3(new_n762), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n822), .B1(new_n826), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n821), .A2(new_n832), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n489), .A2(new_n496), .B1(G472), .B2(new_n508), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n628), .A2(new_n834), .A3(new_n676), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n835), .A2(new_n737), .A3(new_n648), .ZN(new_n836));
  AND3_X1   g650(.A1(new_n648), .A2(new_n564), .A3(new_n642), .ZN(new_n837));
  INV_X1    g651(.A(new_n390), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n837), .A2(new_n702), .A3(new_n838), .A4(new_n686), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n836), .A2(new_n689), .A3(new_n740), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n840), .A2(KEYINPUT52), .ZN(new_n841));
  INV_X1    g655(.A(new_n688), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n738), .A2(new_n648), .A3(new_n721), .ZN(new_n843));
  OAI22_X1  g657(.A1(new_n711), .A2(new_n842), .B1(new_n843), .B2(new_n712), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT52), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n845), .A2(new_n846), .A3(new_n836), .A4(new_n839), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n841), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n188), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n694), .A2(new_n849), .A3(new_n657), .ZN(new_n850));
  NOR3_X1   g664(.A1(new_n628), .A2(new_n850), .A3(new_n632), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT112), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n852), .B1(new_n762), .B2(new_n703), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n640), .A2(new_n645), .A3(KEYINPUT112), .A4(new_n642), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n850), .ZN(new_n856));
  INV_X1    g670(.A(new_n632), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n685), .A2(new_n642), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n856), .A2(new_n857), .A3(new_n684), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n626), .A2(new_n678), .A3(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n855), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n745), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n387), .A2(new_n743), .A3(new_n389), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n738), .A2(new_n754), .A3(new_n862), .A4(new_n863), .ZN(new_n864));
  OAI22_X1  g678(.A1(new_n755), .A2(new_n842), .B1(new_n864), .B2(new_n712), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n684), .A2(new_n709), .A3(new_n710), .ZN(new_n867));
  OR3_X1    g681(.A1(new_n742), .A2(new_n687), .A3(new_n564), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n742), .A2(new_n687), .A3(new_n564), .ZN(new_n870));
  NAND4_X1  g684(.A1(new_n681), .A2(new_n870), .A3(KEYINPUT113), .A4(new_n684), .ZN(new_n871));
  AOI21_X1  g685(.A(new_n865), .B1(new_n869), .B2(new_n871), .ZN(new_n872));
  AND4_X1   g686(.A1(new_n722), .A2(new_n725), .A3(new_n728), .A4(new_n735), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n861), .A2(new_n872), .A3(new_n873), .A4(new_n757), .ZN(new_n874));
  AOI21_X1  g688(.A(new_n848), .B1(KEYINPUT114), .B2(new_n874), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n752), .A2(new_n756), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n722), .A2(new_n725), .A3(new_n728), .A4(new_n735), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT114), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n879), .A3(new_n861), .A4(new_n872), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT53), .B1(new_n875), .B2(new_n880), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n626), .A2(new_n678), .A3(new_n859), .ZN(new_n882));
  INV_X1    g696(.A(new_n865), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n869), .A2(new_n871), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n851), .A2(new_n853), .A3(new_n854), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n882), .A2(new_n883), .A3(new_n884), .A4(new_n885), .ZN(new_n886));
  AND3_X1   g700(.A1(new_n725), .A2(new_n728), .A3(new_n735), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n757), .A2(new_n887), .A3(new_n722), .ZN(new_n888));
  OAI21_X1  g702(.A(KEYINPUT114), .B1(new_n886), .B2(new_n888), .ZN(new_n889));
  AND2_X1   g703(.A1(new_n841), .A2(new_n847), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n844), .A2(KEYINPUT52), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT53), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AND4_X1   g707(.A1(new_n880), .A2(new_n889), .A3(new_n890), .A4(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT54), .B1(new_n881), .B2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n880), .A2(new_n889), .A3(new_n890), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n896), .A2(new_n892), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT54), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n861), .A2(new_n872), .A3(KEYINPUT115), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT115), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n886), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n891), .A2(KEYINPUT53), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n888), .A2(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n890), .A2(new_n899), .A3(new_n901), .A4(new_n903), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n897), .A2(new_n898), .A3(new_n904), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n895), .A2(new_n905), .ZN(new_n906));
  NOR3_X1   g720(.A1(new_n826), .A2(new_n822), .A3(new_n831), .ZN(new_n907));
  NOR3_X1   g721(.A1(new_n833), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NOR2_X1   g722(.A1(G952), .A2(G953), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n763), .A2(new_n631), .A3(new_n849), .A4(new_n389), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT111), .ZN(new_n911));
  NOR2_X1   g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n910), .A2(new_n911), .ZN(new_n913));
  AND2_X1   g727(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n823), .A2(KEYINPUT49), .ZN(new_n915));
  NOR4_X1   g729(.A1(new_n695), .A2(new_n914), .A3(new_n915), .A4(new_n812), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n913), .A2(new_n916), .ZN(new_n917));
  OAI22_X1  g731(.A1(new_n908), .A2(new_n909), .B1(new_n912), .B2(new_n917), .ZN(G75));
  NOR2_X1   g732(.A1(new_n372), .A2(G952), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n919), .B(KEYINPUT118), .ZN(new_n920));
  INV_X1    g734(.A(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(KEYINPUT56), .ZN(new_n922));
  AND4_X1   g736(.A1(new_n890), .A2(new_n899), .A3(new_n901), .A4(new_n903), .ZN(new_n923));
  OAI21_X1  g737(.A(G902), .B1(new_n881), .B2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(G210), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n922), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n323), .A2(new_n324), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT117), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n327), .B(KEYINPUT55), .ZN(new_n929));
  XOR2_X1   g743(.A(new_n928), .B(new_n929), .Z(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n926), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n926), .A2(new_n931), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n921), .B1(new_n932), .B2(new_n933), .ZN(G51));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n881), .B2(new_n923), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n905), .ZN(new_n936));
  INV_X1    g750(.A(new_n936), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n381), .B(KEYINPUT57), .ZN(new_n938));
  OAI22_X1  g752(.A1(new_n937), .A2(new_n938), .B1(new_n379), .B2(new_n376), .ZN(new_n939));
  INV_X1    g753(.A(new_n924), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n781), .B(KEYINPUT119), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n919), .B1(new_n939), .B2(new_n942), .ZN(G54));
  INV_X1    g757(.A(new_n612), .ZN(new_n944));
  NAND2_X1  g758(.A1(KEYINPUT58), .A2(G475), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n924), .B2(new_n945), .ZN(new_n946));
  INV_X1    g760(.A(new_n919), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n924), .A2(new_n944), .A3(new_n945), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n949), .ZN(G60));
  INV_X1    g764(.A(KEYINPUT121), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n636), .B(KEYINPUT120), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT59), .Z(new_n955));
  NOR2_X1   g769(.A1(new_n953), .A2(new_n955), .ZN(new_n956));
  NOR3_X1   g770(.A1(new_n881), .A2(KEYINPUT54), .A3(new_n923), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n898), .B1(new_n897), .B2(new_n904), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n959), .A2(new_n920), .ZN(new_n960));
  INV_X1    g774(.A(new_n955), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n952), .B1(new_n906), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n951), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n875), .A2(new_n880), .A3(new_n893), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n898), .B1(new_n897), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n961), .B1(new_n957), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n953), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n921), .B1(new_n936), .B2(new_n956), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n967), .A2(new_n968), .A3(KEYINPUT121), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n963), .A2(new_n969), .ZN(G63));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n429), .A2(new_n430), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n881), .A2(new_n923), .ZN(new_n973));
  NAND2_X1  g787(.A1(G217), .A2(G902), .ZN(new_n974));
  XNOR2_X1  g788(.A(new_n974), .B(KEYINPUT60), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n972), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n976), .A2(new_n920), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n669), .A2(new_n670), .ZN(new_n978));
  NOR3_X1   g792(.A1(new_n973), .A2(new_n978), .A3(new_n975), .ZN(new_n979));
  OAI21_X1  g793(.A(new_n971), .B1(new_n977), .B2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n979), .ZN(new_n981));
  NAND4_X1  g795(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n920), .A4(new_n976), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(G66));
  OAI21_X1  g797(.A(G953), .B1(new_n570), .B2(new_n191), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n861), .A2(new_n873), .ZN(new_n985));
  INV_X1    g799(.A(new_n985), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n984), .B1(new_n986), .B2(G953), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n928), .B1(G898), .B2(new_n372), .ZN(new_n988));
  XNOR2_X1  g802(.A(new_n987), .B(new_n988), .ZN(G69));
  NOR2_X1   g803(.A1(new_n844), .A2(new_n713), .ZN(new_n990));
  INV_X1    g804(.A(KEYINPUT124), .ZN(new_n991));
  XNOR2_X1  g805(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n992), .A2(new_n705), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n993), .B(KEYINPUT62), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n853), .A2(new_n854), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n995), .B1(new_n685), .B2(new_n642), .ZN(new_n996));
  OR2_X1    g810(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n997));
  INV_X1    g811(.A(new_n692), .ZN(new_n998));
  NOR3_X1   g812(.A1(new_n834), .A2(new_n444), .A3(new_n742), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n996), .A2(KEYINPUT125), .ZN(new_n1000));
  NAND4_X1  g814(.A1(new_n997), .A2(new_n998), .A3(new_n999), .A4(new_n1000), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n805), .A2(new_n793), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g816(.A(new_n372), .B1(new_n994), .B2(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n483), .B(KEYINPUT122), .Z(new_n1004));
  XNOR2_X1  g818(.A(new_n1004), .B(new_n604), .ZN(new_n1005));
  XNOR2_X1  g819(.A(new_n1005), .B(KEYINPUT123), .ZN(new_n1006));
  AND2_X1   g820(.A1(new_n805), .A2(new_n793), .ZN(new_n1007));
  NAND2_X1  g821(.A1(new_n757), .A2(new_n760), .ZN(new_n1008));
  INV_X1    g822(.A(KEYINPUT127), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n818), .A2(new_n837), .ZN(new_n1010));
  OAI21_X1  g824(.A(new_n1009), .B1(new_n791), .B2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n790), .A2(KEYINPUT127), .A3(new_n837), .A4(new_n818), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n1008), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AND2_X1   g827(.A1(new_n1013), .A2(new_n992), .ZN(new_n1014));
  NAND3_X1  g828(.A1(new_n1007), .A2(new_n372), .A3(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1005), .B1(G900), .B2(G953), .ZN(new_n1016));
  AOI22_X1  g830(.A1(new_n1003), .A2(new_n1006), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n372), .B1(G227), .B2(G900), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1014), .A2(new_n793), .A3(new_n805), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1016), .B1(new_n1019), .B2(G953), .ZN(new_n1020));
  INV_X1    g834(.A(KEYINPUT126), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1018), .B1(new_n1020), .B2(new_n1021), .ZN(new_n1022));
  XNOR2_X1  g836(.A(new_n1017), .B(new_n1022), .ZN(G72));
  XOR2_X1   g837(.A(new_n993), .B(KEYINPUT62), .Z(new_n1024));
  NAND4_X1  g838(.A1(new_n1024), .A2(new_n1007), .A3(new_n986), .A4(new_n1001), .ZN(new_n1025));
  NAND2_X1  g839(.A1(G472), .A2(G902), .ZN(new_n1026));
  XOR2_X1   g840(.A(new_n1026), .B(KEYINPUT63), .Z(new_n1027));
  AOI211_X1 g841(.A(new_n500), .B(new_n506), .C1(new_n1025), .C2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n1027), .B1(new_n1019), .B2(new_n985), .ZN(new_n1029));
  NAND3_X1  g843(.A1(new_n1029), .A2(new_n500), .A3(new_n506), .ZN(new_n1030));
  OAI21_X1  g844(.A(new_n697), .B1(new_n449), .B2(new_n506), .ZN(new_n1031));
  OAI211_X1 g845(.A(new_n1027), .B(new_n1031), .C1(new_n881), .C2(new_n894), .ZN(new_n1032));
  NAND3_X1  g846(.A1(new_n1030), .A2(new_n947), .A3(new_n1032), .ZN(new_n1033));
  NOR2_X1   g847(.A1(new_n1028), .A2(new_n1033), .ZN(G57));
endmodule


