//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 1 1 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 1 1 0 0 1 1 1 1 0 0 1 1 1 0 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:10 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1317,
    new_n1318, new_n1319, new_n1320, new_n1321, new_n1322, new_n1323;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  XOR2_X1   g0007(.A(KEYINPUT65), .B(G238), .Z(new_n208));
  INV_X1    g0008(.A(G68), .ZN(new_n209));
  OR2_X1    g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G97), .A2(G257), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G58), .A2(G232), .ZN(new_n212));
  INV_X1    g0012(.A(G87), .ZN(new_n213));
  INV_X1    g0013(.A(G250), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n212), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  AOI21_X1  g0015(.A(new_n215), .B1(G107), .B2(G264), .ZN(new_n216));
  INV_X1    g0016(.A(G226), .ZN(new_n217));
  INV_X1    g0017(.A(G244), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n202), .A2(new_n217), .B1(new_n205), .B2(new_n218), .ZN(new_n219));
  AOI21_X1  g0019(.A(new_n219), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND4_X1  g0020(.A1(new_n210), .A2(new_n211), .A3(new_n216), .A4(new_n220), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G20), .ZN(new_n222));
  NAND2_X1  g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XOR2_X1   g0023(.A(new_n223), .B(KEYINPUT1), .Z(new_n224));
  NOR2_X1   g0024(.A1(new_n222), .A2(G13), .ZN(new_n225));
  OAI211_X1 g0025(.A(new_n225), .B(G250), .C1(G257), .C2(G264), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT0), .ZN(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NOR2_X1   g0029(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g0030(.A(new_n230), .ZN(new_n231));
  INV_X1    g0031(.A(new_n201), .ZN(new_n232));
  NAND2_X1  g0032(.A1(new_n232), .A2(G50), .ZN(new_n233));
  OAI211_X1 g0033(.A(new_n224), .B(new_n227), .C1(new_n231), .C2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n236), .B(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G250), .B(G257), .Z(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G107), .B(G116), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT66), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G87), .B(G97), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G58), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n247), .B(new_n250), .ZN(G351));
  INV_X1    g0051(.A(G1), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G13), .A3(G20), .ZN(new_n253));
  INV_X1    g0053(.A(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G116), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g0056(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n257), .A2(new_n228), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n252), .A2(G33), .ZN(new_n260));
  NAND4_X1  g0060(.A1(new_n259), .A2(G116), .A3(new_n253), .A4(new_n260), .ZN(new_n261));
  AOI22_X1  g0061(.A1(new_n257), .A2(new_n228), .B1(G20), .B2(new_n255), .ZN(new_n262));
  NAND2_X1  g0062(.A1(G33), .A2(G283), .ZN(new_n263));
  INV_X1    g0063(.A(G97), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n263), .B(new_n229), .C1(G33), .C2(new_n264), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n262), .A2(KEYINPUT20), .A3(new_n265), .ZN(new_n266));
  AOI21_X1  g0066(.A(KEYINPUT20), .B1(new_n262), .B2(new_n265), .ZN(new_n267));
  OAI211_X1 g0067(.A(new_n256), .B(new_n261), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT84), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n262), .A2(new_n265), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT20), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n262), .A2(KEYINPUT20), .A3(new_n265), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT84), .ZN(new_n275));
  NAND4_X1  g0075(.A1(new_n274), .A2(new_n275), .A3(new_n256), .A4(new_n261), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n269), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT3), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n280), .A2(G33), .ZN(new_n281));
  INV_X1    g0081(.A(G1698), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n282), .A2(G257), .ZN(new_n283));
  NAND2_X1  g0083(.A1(G264), .A2(G1698), .ZN(new_n284));
  NAND4_X1  g0084(.A1(new_n279), .A2(new_n281), .A3(new_n283), .A4(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G41), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n286), .A2(G1), .A3(G13), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  XNOR2_X1  g0088(.A(KEYINPUT3), .B(G33), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n285), .B(new_n288), .C1(G303), .C2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G45), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n291), .A2(G1), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT5), .A2(G41), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT5), .A2(G41), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n295), .A2(G270), .A3(new_n287), .ZN(new_n296));
  OAI211_X1 g0096(.A(new_n292), .B(G274), .C1(new_n294), .C2(new_n293), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n290), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  NAND3_X1  g0099(.A1(new_n277), .A2(new_n299), .A3(G179), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n269), .A2(new_n276), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(G200), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n299), .A2(G190), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n301), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT21), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n299), .A2(new_n306), .ZN(new_n307));
  AND3_X1   g0107(.A1(new_n277), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n305), .B1(new_n277), .B2(new_n307), .ZN(new_n309));
  OAI211_X1 g0109(.A(new_n300), .B(new_n304), .C1(new_n308), .C2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n279), .A2(new_n281), .ZN(new_n312));
  AOI21_X1  g0112(.A(new_n312), .B1(G222), .B2(new_n282), .ZN(new_n313));
  INV_X1    g0113(.A(G223), .ZN(new_n314));
  OAI21_X1  g0114(.A(new_n313), .B1(new_n314), .B2(new_n282), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n288), .C1(G77), .C2(new_n289), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n252), .B1(G41), .B2(G45), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT67), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n252), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n320));
  AND3_X1   g0120(.A1(new_n319), .A2(new_n287), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(G226), .ZN(new_n322));
  INV_X1    g0122(.A(G274), .ZN(new_n323));
  OR2_X1    g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n316), .A2(new_n322), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  NOR2_X1   g0126(.A1(new_n326), .A2(G169), .ZN(new_n327));
  NOR2_X1   g0127(.A1(G20), .A2(G33), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G150), .ZN(new_n329));
  XNOR2_X1  g0129(.A(KEYINPUT8), .B(G58), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(KEYINPUT68), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT68), .ZN(new_n332));
  INV_X1    g0132(.A(G58), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n333), .A3(KEYINPUT8), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n229), .A2(G33), .ZN(new_n336));
  OAI221_X1 g0136(.A(new_n329), .B1(new_n335), .B2(new_n336), .C1(new_n229), .C2(new_n204), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n337), .A2(new_n258), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n254), .A2(new_n202), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n258), .B1(new_n252), .B2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n340), .A2(G50), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NOR2_X1   g0143(.A1(new_n325), .A2(G179), .ZN(new_n344));
  NOR3_X1   g0144(.A1(new_n327), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n326), .A2(G190), .ZN(new_n346));
  NAND4_X1  g0146(.A1(new_n338), .A2(KEYINPUT9), .A3(new_n339), .A4(new_n341), .ZN(new_n347));
  AND2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT10), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n325), .A2(G200), .ZN(new_n350));
  INV_X1    g0150(.A(KEYINPUT9), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n342), .A2(new_n351), .ZN(new_n352));
  NAND4_X1  g0152(.A1(new_n348), .A2(new_n349), .A3(new_n350), .A4(new_n352), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n352), .A2(new_n346), .A3(new_n350), .A4(new_n347), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n354), .A2(KEYINPUT10), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n345), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT75), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT16), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT74), .B1(new_n280), .B2(G33), .ZN(new_n360));
  INV_X1    g0160(.A(KEYINPUT74), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n361), .A2(new_n278), .A3(KEYINPUT3), .ZN(new_n362));
  NAND3_X1  g0162(.A1(new_n360), .A2(new_n362), .A3(new_n281), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G20), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n363), .A2(new_n365), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n364), .B1(new_n289), .B2(G20), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n209), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(G58), .A2(G68), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n370), .B2(new_n201), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  INV_X1    g0172(.A(new_n328), .ZN(new_n373));
  OAI21_X1  g0173(.A(new_n371), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n359), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT73), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n229), .B1(new_n232), .B2(new_n369), .ZN(new_n377));
  NOR2_X1   g0177(.A1(new_n373), .A2(new_n372), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI211_X1 g0179(.A(new_n371), .B(KEYINPUT73), .C1(new_n372), .C2(new_n373), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g0181(.A(KEYINPUT7), .B1(new_n312), .B2(new_n229), .ZN(new_n382));
  INV_X1    g0182(.A(new_n365), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n289), .A2(new_n383), .ZN(new_n384));
  OAI21_X1  g0184(.A(G68), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n381), .A2(new_n385), .A3(KEYINPUT16), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n375), .A2(new_n386), .A3(new_n258), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n335), .A2(new_n254), .ZN(new_n388));
  INV_X1    g0188(.A(new_n340), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n388), .B1(new_n335), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n387), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n217), .A2(G1698), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n314), .A2(new_n282), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n289), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(G33), .A2(G87), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n395), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n397), .A2(new_n288), .ZN(new_n398));
  NAND4_X1  g0198(.A1(new_n319), .A2(G232), .A3(new_n287), .A4(new_n320), .ZN(new_n399));
  NAND4_X1  g0199(.A1(new_n398), .A2(G179), .A3(new_n324), .A4(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n399), .A2(new_n324), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n287), .B1(new_n395), .B2(new_n396), .ZN(new_n402));
  OAI21_X1  g0202(.A(G169), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n400), .A2(new_n403), .ZN(new_n404));
  AND3_X1   g0204(.A1(new_n392), .A2(KEYINPUT18), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(KEYINPUT18), .B1(new_n392), .B2(new_n404), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n358), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(KEYINPUT18), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n367), .B1(new_n289), .B2(new_n383), .ZN(new_n409));
  AOI22_X1  g0209(.A1(new_n409), .A2(G68), .B1(new_n379), .B2(new_n380), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n259), .B1(new_n410), .B2(KEYINPUT16), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n390), .B1(new_n411), .B2(new_n375), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n400), .A2(new_n403), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n408), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n392), .A2(KEYINPUT18), .A3(new_n404), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n414), .A2(KEYINPUT75), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g0216(.A(G200), .B1(new_n401), .B2(new_n402), .ZN(new_n417));
  NAND4_X1  g0217(.A1(new_n398), .A2(G190), .A3(new_n324), .A4(new_n399), .ZN(new_n418));
  NAND4_X1  g0218(.A1(new_n387), .A2(new_n417), .A3(new_n418), .A4(new_n391), .ZN(new_n419));
  XNOR2_X1  g0219(.A(new_n419), .B(KEYINPUT17), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n407), .A2(new_n416), .A3(new_n420), .ZN(new_n421));
  NOR2_X1   g0221(.A1(new_n357), .A2(new_n421), .ZN(new_n422));
  NAND4_X1  g0222(.A1(new_n279), .A2(new_n281), .A3(G226), .A4(new_n282), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(KEYINPUT69), .ZN(new_n424));
  INV_X1    g0224(.A(KEYINPUT69), .ZN(new_n425));
  NAND4_X1  g0225(.A1(new_n289), .A2(new_n425), .A3(G226), .A4(new_n282), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(G33), .A2(G97), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n289), .A2(G232), .A3(G1698), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n427), .A2(new_n428), .A3(new_n429), .ZN(new_n430));
  INV_X1    g0230(.A(KEYINPUT70), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n427), .A2(KEYINPUT70), .A3(new_n428), .A4(new_n429), .ZN(new_n433));
  NAND3_X1  g0233(.A1(new_n432), .A2(new_n288), .A3(new_n433), .ZN(new_n434));
  INV_X1    g0234(.A(KEYINPUT13), .ZN(new_n435));
  INV_X1    g0235(.A(new_n324), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n321), .B2(G238), .ZN(new_n437));
  AND3_X1   g0237(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n435), .B1(new_n434), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g0239(.A(G169), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(KEYINPUT14), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n438), .A2(new_n439), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G179), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(G169), .C1(new_n438), .C2(new_n439), .ZN(new_n445));
  NAND3_X1  g0245(.A1(new_n441), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n373), .A2(new_n202), .B1(new_n336), .B2(new_n205), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n229), .A2(G68), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n258), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT11), .ZN(new_n450));
  AOI211_X1 g0250(.A(G68), .B(new_n253), .C1(KEYINPUT72), .C2(KEYINPUT12), .ZN(new_n451));
  NOR2_X1   g0251(.A1(KEYINPUT72), .A2(KEYINPUT12), .ZN(new_n452));
  XNOR2_X1  g0252(.A(new_n451), .B(new_n452), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n450), .B(new_n453), .C1(new_n209), .C2(new_n389), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(new_n454), .ZN(new_n456));
  INV_X1    g0256(.A(G190), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n438), .A2(new_n439), .A3(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(KEYINPUT71), .ZN(new_n460));
  INV_X1    g0260(.A(new_n439), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n434), .A2(new_n435), .A3(new_n437), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n460), .B1(new_n463), .B2(G200), .ZN(new_n464));
  OAI211_X1 g0264(.A(new_n460), .B(G200), .C1(new_n438), .C2(new_n439), .ZN(new_n465));
  INV_X1    g0265(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n456), .B(new_n459), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  AOI21_X1  g0267(.A(new_n436), .B1(new_n321), .B2(G244), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n282), .A2(G232), .ZN(new_n469));
  OAI211_X1 g0269(.A(new_n289), .B(new_n469), .C1(new_n208), .C2(new_n282), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n470), .B1(G107), .B2(new_n289), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n471), .B2(new_n287), .ZN(new_n472));
  OR2_X1    g0272(.A1(new_n472), .A2(G179), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n253), .A2(G77), .ZN(new_n474));
  INV_X1    g0274(.A(new_n330), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT15), .B(G87), .Z(new_n476));
  INV_X1    g0276(.A(new_n336), .ZN(new_n477));
  AOI22_X1  g0277(.A1(new_n475), .A2(new_n328), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(new_n229), .B2(new_n205), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n474), .B1(new_n479), .B2(new_n258), .ZN(new_n480));
  OAI21_X1  g0280(.A(new_n480), .B1(new_n205), .B2(new_n389), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n472), .A2(new_n306), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n473), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NOR2_X1   g0283(.A1(new_n389), .A2(new_n205), .ZN(new_n484));
  AOI211_X1 g0284(.A(new_n474), .B(new_n484), .C1(new_n479), .C2(new_n258), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n472), .A2(G200), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n485), .B(new_n486), .C1(new_n457), .C2(new_n472), .ZN(new_n487));
  AND2_X1   g0287(.A1(new_n483), .A2(new_n487), .ZN(new_n488));
  AND4_X1   g0288(.A1(new_n422), .A2(new_n455), .A3(new_n467), .A4(new_n488), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n295), .A2(G257), .A3(new_n287), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(new_n297), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n218), .A2(G1698), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(new_n279), .A3(new_n281), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT4), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(KEYINPUT77), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT77), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(KEYINPUT4), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n289), .A2(new_n492), .A3(new_n495), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n279), .A2(new_n281), .A3(G250), .A4(G1698), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n499), .A2(new_n500), .A3(new_n263), .A4(new_n501), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n491), .B1(new_n502), .B2(new_n288), .ZN(new_n503));
  NOR2_X1   g0303(.A1(new_n503), .A2(G169), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n502), .A2(new_n288), .ZN(new_n505));
  INV_X1    g0305(.A(G179), .ZN(new_n506));
  INV_X1    g0306(.A(new_n491), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n505), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT79), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT79), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n510), .A3(new_n506), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n504), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g0312(.A1(new_n280), .A2(G33), .ZN(new_n513));
  NOR2_X1   g0313(.A1(new_n278), .A2(KEYINPUT3), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n229), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n364), .A2(new_n515), .B1(new_n363), .B2(new_n365), .ZN(new_n516));
  INV_X1    g0316(.A(G107), .ZN(new_n517));
  OAI21_X1  g0317(.A(KEYINPUT76), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n517), .A2(KEYINPUT6), .A3(G97), .ZN(new_n519));
  XOR2_X1   g0319(.A(G97), .B(G107), .Z(new_n520));
  OAI21_X1  g0320(.A(new_n519), .B1(new_n520), .B2(KEYINPUT6), .ZN(new_n521));
  AOI22_X1  g0321(.A1(new_n521), .A2(G20), .B1(G77), .B2(new_n328), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n366), .A2(new_n367), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT76), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n523), .A2(new_n524), .A3(G107), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n518), .A2(new_n522), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(new_n258), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n254), .A2(new_n264), .ZN(new_n528));
  NAND4_X1  g0328(.A1(new_n253), .A2(new_n260), .A3(new_n228), .A4(new_n257), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n528), .B1(new_n529), .B2(new_n264), .ZN(new_n530));
  INV_X1    g0330(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n512), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT78), .ZN(new_n534));
  INV_X1    g0334(.A(G200), .ZN(new_n535));
  OAI21_X1  g0335(.A(new_n534), .B1(new_n503), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n503), .A2(G190), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n503), .A2(new_n534), .A3(G190), .ZN(new_n539));
  NAND4_X1  g0339(.A1(new_n538), .A2(new_n527), .A3(new_n531), .A4(new_n539), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n252), .A2(new_n517), .A3(G13), .A4(G20), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n541), .A2(KEYINPUT25), .ZN(new_n542));
  NOR2_X1   g0342(.A1(new_n229), .A2(G107), .ZN(new_n543));
  INV_X1    g0343(.A(KEYINPUT25), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(new_n252), .A4(G13), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n542), .B(new_n545), .C1(new_n529), .C2(new_n517), .ZN(new_n546));
  XNOR2_X1  g0346(.A(new_n546), .B(KEYINPUT86), .ZN(new_n547));
  AND2_X1   g0347(.A1(KEYINPUT85), .A2(G87), .ZN(new_n548));
  NAND4_X1  g0348(.A1(new_n279), .A2(new_n281), .A3(new_n548), .A4(new_n229), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(KEYINPUT22), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT22), .ZN(new_n551));
  NAND4_X1  g0351(.A1(new_n289), .A2(new_n551), .A3(new_n229), .A4(new_n548), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n550), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n543), .A2(KEYINPUT23), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT23), .ZN(new_n555));
  OAI21_X1  g0355(.A(new_n555), .B1(new_n229), .B2(G107), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n554), .A2(new_n556), .B1(new_n477), .B2(G116), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n553), .A2(KEYINPUT24), .A3(new_n557), .ZN(new_n558));
  AOI21_X1  g0358(.A(KEYINPUT24), .B1(new_n553), .B2(new_n557), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AOI21_X1  g0360(.A(new_n547), .B1(new_n560), .B2(new_n258), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n295), .A2(G264), .A3(new_n287), .ZN(new_n562));
  NAND2_X1  g0362(.A1(G257), .A2(G1698), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n563), .B1(new_n214), .B2(G1698), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n289), .A2(new_n564), .B1(G33), .B2(G294), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n562), .B(new_n297), .C1(new_n565), .C2(new_n287), .ZN(new_n566));
  OR2_X1    g0366(.A1(new_n566), .A2(new_n457), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(G200), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n561), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  AND3_X1   g0369(.A1(new_n533), .A2(new_n540), .A3(new_n569), .ZN(new_n570));
  OR2_X1    g0370(.A1(G238), .A2(G1698), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n218), .A2(G1698), .ZN(new_n572));
  NAND4_X1  g0372(.A1(new_n279), .A2(new_n571), .A3(new_n281), .A4(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(G33), .A2(G116), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n288), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n252), .A2(G45), .A3(G274), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n577), .A2(KEYINPUT80), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT80), .ZN(new_n579));
  NAND4_X1  g0379(.A1(new_n579), .A2(new_n252), .A3(G45), .A4(G274), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n291), .B2(G1), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n252), .A2(KEYINPUT81), .A3(G45), .ZN(new_n584));
  NAND4_X1  g0384(.A1(new_n287), .A2(new_n583), .A3(G250), .A4(new_n584), .ZN(new_n585));
  AND2_X1   g0385(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n576), .A2(new_n586), .A3(G179), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n287), .B1(new_n573), .B2(new_n574), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n581), .A2(new_n585), .ZN(new_n589));
  OAI21_X1  g0389(.A(G169), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT82), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT82), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n587), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n595), .A2(KEYINPUT83), .A3(new_n229), .ZN(new_n596));
  INV_X1    g0396(.A(new_n596), .ZN(new_n597));
  AOI21_X1  g0397(.A(KEYINPUT83), .B1(new_n595), .B2(new_n229), .ZN(new_n598));
  NOR3_X1   g0398(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n279), .A2(new_n281), .A3(new_n229), .A4(G68), .ZN(new_n601));
  INV_X1    g0401(.A(KEYINPUT19), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n602), .B1(new_n336), .B2(new_n264), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n258), .B1(new_n600), .B2(new_n604), .ZN(new_n605));
  INV_X1    g0405(.A(new_n476), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n254), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n605), .B(new_n607), .C1(new_n529), .C2(new_n606), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n592), .A2(new_n594), .A3(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n595), .A2(new_n229), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT83), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(new_n599), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n596), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n614), .A2(new_n601), .A3(new_n603), .ZN(new_n615));
  AOI22_X1  g0415(.A1(new_n615), .A2(new_n258), .B1(new_n254), .B2(new_n606), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n588), .A2(new_n589), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n617), .A2(G190), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n588), .B2(new_n589), .ZN(new_n619));
  OR2_X1    g0419(.A1(new_n529), .A2(new_n213), .ZN(new_n620));
  NAND4_X1  g0420(.A1(new_n616), .A2(new_n618), .A3(new_n619), .A4(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n609), .A2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT87), .ZN(new_n623));
  AND3_X1   g0423(.A1(new_n566), .A2(new_n623), .A3(G169), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n623), .B1(new_n566), .B2(G169), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n566), .A2(new_n506), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n624), .A2(new_n625), .A3(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(KEYINPUT88), .B1(new_n561), .B2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n566), .A2(G169), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT87), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n566), .A2(new_n623), .A3(G169), .ZN(new_n631));
  OAI211_X1 g0431(.A(new_n630), .B(new_n631), .C1(new_n506), .C2(new_n566), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n553), .A2(new_n557), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT24), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n553), .A2(KEYINPUT24), .A3(new_n557), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n258), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n547), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT88), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n632), .A2(new_n639), .A3(new_n640), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n622), .B1(new_n628), .B2(new_n641), .ZN(new_n642));
  AND4_X1   g0442(.A1(new_n311), .A2(new_n489), .A3(new_n570), .A4(new_n642), .ZN(G372));
  NAND2_X1  g0443(.A1(new_n353), .A2(new_n355), .ZN(new_n644));
  INV_X1    g0444(.A(new_n420), .ZN(new_n645));
  INV_X1    g0445(.A(new_n483), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n467), .A2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n645), .B1(new_n647), .B2(new_n455), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n405), .A2(new_n406), .ZN(new_n649));
  OAI21_X1  g0449(.A(new_n644), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  INV_X1    g0450(.A(new_n345), .ZN(new_n651));
  AND2_X1   g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n512), .A2(new_n532), .A3(new_n609), .A4(new_n621), .ZN(new_n653));
  INV_X1    g0453(.A(KEYINPUT26), .ZN(new_n654));
  OAI21_X1  g0454(.A(KEYINPUT90), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND2_X1   g0455(.A1(new_n512), .A2(new_n532), .ZN(new_n656));
  AND2_X1   g0456(.A1(new_n609), .A2(new_n621), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT90), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n656), .A2(new_n657), .A3(new_n658), .A4(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT89), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n605), .A2(new_n620), .A3(new_n607), .ZN(new_n661));
  INV_X1    g0461(.A(new_n619), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n660), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n616), .A2(KEYINPUT89), .A3(new_n619), .A4(new_n620), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n663), .A2(new_n618), .A3(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n608), .A2(new_n591), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n654), .B1(new_n667), .B2(new_n533), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n655), .A2(new_n659), .A3(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n632), .A2(new_n639), .ZN(new_n670));
  OAI211_X1 g0470(.A(new_n670), .B(new_n300), .C1(new_n308), .C2(new_n309), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n665), .A2(new_n666), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n570), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n666), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n489), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n652), .A2(new_n675), .ZN(G369));
  NAND2_X1  g0476(.A1(new_n628), .A2(new_n641), .ZN(new_n677));
  INV_X1    g0477(.A(G13), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G20), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n252), .ZN(new_n680));
  OR2_X1    g0480(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n680), .A2(KEYINPUT27), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n681), .A2(G213), .A3(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(G343), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n677), .B(new_n569), .C1(new_n561), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT91), .ZN(new_n688));
  OR2_X1    g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n687), .A2(new_n688), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n691), .B1(new_n670), .B2(new_n686), .ZN(new_n692));
  OAI21_X1  g0492(.A(new_n300), .B1(new_n308), .B2(new_n309), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n301), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  OAI21_X1  g0495(.A(new_n695), .B1(new_n310), .B2(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G330), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n632), .A2(new_n639), .A3(new_n686), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n693), .A2(new_n686), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n689), .A2(new_n690), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n699), .A2(new_n700), .A3(new_n703), .ZN(G399));
  INV_X1    g0504(.A(new_n225), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G41), .ZN(new_n706));
  INV_X1    g0506(.A(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n613), .A2(G116), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n707), .A2(G1), .A3(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n709), .B1(new_n233), .B2(new_n707), .ZN(new_n710));
  XNOR2_X1  g0510(.A(new_n710), .B(KEYINPUT28), .ZN(new_n711));
  NAND3_X1  g0511(.A1(new_n533), .A2(new_n540), .A3(new_n569), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n712), .A2(new_n667), .ZN(new_n713));
  AOI22_X1  g0513(.A1(new_n713), .A2(new_n671), .B1(new_n608), .B2(new_n591), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n685), .B1(new_n714), .B2(new_n669), .ZN(new_n715));
  OR2_X1    g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  INV_X1    g0516(.A(new_n677), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n713), .B1(new_n693), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n608), .A2(new_n591), .A3(KEYINPUT93), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n653), .A2(KEYINPUT26), .ZN(new_n720));
  INV_X1    g0520(.A(KEYINPUT93), .ZN(new_n721));
  AOI21_X1  g0521(.A(new_n720), .B1(new_n721), .B2(new_n666), .ZN(new_n722));
  OAI21_X1  g0522(.A(KEYINPUT26), .B1(new_n667), .B2(new_n533), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n718), .A2(new_n719), .A3(new_n722), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT29), .A3(new_n686), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n716), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g0526(.A1(new_n570), .A2(new_n311), .A3(new_n642), .A4(new_n686), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n505), .A2(new_n507), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n562), .B1(new_n565), .B2(new_n287), .ZN(new_n729));
  NOR4_X1   g0529(.A1(new_n728), .A2(new_n587), .A3(new_n298), .A4(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT30), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n728), .A2(new_n566), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(KEYINPUT92), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(new_n298), .ZN(new_n734));
  OAI21_X1  g0534(.A(new_n506), .B1(new_n732), .B2(KEYINPUT92), .ZN(new_n735));
  NOR3_X1   g0535(.A1(new_n734), .A2(new_n735), .A3(new_n617), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n685), .B1(new_n731), .B2(new_n736), .ZN(new_n737));
  NAND3_X1  g0537(.A1(new_n727), .A2(KEYINPUT31), .A3(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n737), .A2(KEYINPUT31), .ZN(new_n739));
  AND2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(G330), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n726), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n711), .B1(new_n743), .B2(G1), .ZN(G364));
  NOR2_X1   g0544(.A1(new_n705), .A2(new_n289), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n745), .B1(G45), .B2(new_n233), .ZN(new_n746));
  XNOR2_X1  g0546(.A(new_n746), .B(KEYINPUT94), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n291), .B2(new_n250), .ZN(new_n748));
  INV_X1    g0548(.A(G355), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n289), .A2(new_n225), .ZN(new_n750));
  OAI221_X1 g0550(.A(new_n748), .B1(G116), .B2(new_n225), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(G1), .B(G13), .C1(new_n229), .C2(G169), .ZN(new_n752));
  OR2_X1    g0552(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(KEYINPUT95), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  NOR2_X1   g0555(.A1(G13), .A2(G33), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(G20), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n758), .ZN(new_n759));
  XNOR2_X1  g0559(.A(new_n759), .B(KEYINPUT96), .ZN(new_n760));
  NAND2_X1  g0560(.A1(new_n751), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n252), .B1(new_n679), .B2(G45), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n706), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n229), .A2(new_n457), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n506), .A2(G200), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n289), .B1(new_n768), .B2(G322), .ZN(new_n769));
  INV_X1    g0569(.A(G294), .ZN(new_n770));
  NOR2_X1   g0570(.A1(G179), .A2(G200), .ZN(new_n771));
  AOI21_X1  g0571(.A(new_n229), .B1(new_n771), .B2(G190), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n506), .A2(new_n535), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n229), .A2(G190), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g0575(.A(KEYINPUT33), .B(G317), .Z(new_n776));
  OAI221_X1 g0576(.A(new_n769), .B1(new_n770), .B2(new_n772), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n535), .A2(G179), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n774), .A2(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n774), .A2(new_n771), .ZN(new_n781));
  INV_X1    g0581(.A(new_n781), .ZN(new_n782));
  AOI22_X1  g0582(.A1(G283), .A2(new_n780), .B1(new_n782), .B2(G329), .ZN(new_n783));
  INV_X1    g0583(.A(G303), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n765), .A2(new_n778), .ZN(new_n785));
  INV_X1    g0585(.A(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n774), .A2(new_n766), .ZN(new_n787));
  OAI221_X1 g0587(.A(new_n783), .B1(new_n784), .B2(new_n785), .C1(new_n786), .C2(new_n787), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n765), .A2(new_n773), .ZN(new_n789));
  INV_X1    g0589(.A(new_n789), .ZN(new_n790));
  AOI211_X1 g0590(.A(new_n777), .B(new_n788), .C1(G326), .C2(new_n790), .ZN(new_n791));
  NOR2_X1   g0591(.A1(new_n785), .A2(new_n213), .ZN(new_n792));
  INV_X1    g0592(.A(new_n792), .ZN(new_n793));
  OAI221_X1 g0593(.A(new_n793), .B1(new_n787), .B2(new_n205), .C1(new_n333), .C2(new_n767), .ZN(new_n794));
  OR3_X1    g0594(.A1(new_n781), .A2(KEYINPUT32), .A3(new_n372), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT32), .B1(new_n781), .B2(new_n372), .ZN(new_n796));
  OAI211_X1 g0596(.A(new_n795), .B(new_n796), .C1(new_n264), .C2(new_n772), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n779), .A2(new_n517), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n289), .B1(new_n775), .B2(new_n209), .C1(new_n202), .C2(new_n789), .ZN(new_n799));
  NOR4_X1   g0599(.A1(new_n794), .A2(new_n797), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n755), .B1(new_n791), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n761), .A2(new_n764), .A3(new_n801), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n802), .A2(KEYINPUT97), .ZN(new_n804));
  INV_X1    g0604(.A(new_n758), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n803), .B(new_n804), .C1(new_n696), .C2(new_n805), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n696), .A2(G330), .ZN(new_n807));
  INV_X1    g0607(.A(new_n764), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n697), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n806), .B1(new_n807), .B2(new_n809), .ZN(G396));
  INV_X1    g0610(.A(KEYINPUT99), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n481), .A2(new_n685), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n483), .A2(new_n487), .A3(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n813), .A2(KEYINPUT98), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(KEYINPUT98), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n811), .B1(new_n715), .B2(new_n816), .ZN(new_n817));
  AND4_X1   g0617(.A1(new_n811), .A2(new_n674), .A3(new_n686), .A4(new_n816), .ZN(new_n818));
  OAI22_X1  g0618(.A1(new_n814), .A2(new_n815), .B1(new_n483), .B2(new_n686), .ZN(new_n819));
  OAI22_X1  g0619(.A1(new_n817), .A2(new_n818), .B1(new_n715), .B2(new_n819), .ZN(new_n820));
  XOR2_X1   g0620(.A(new_n820), .B(new_n741), .Z(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n808), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n779), .A2(new_n213), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n823), .B1(G294), .B2(new_n768), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n824), .B1(new_n517), .B2(new_n785), .ZN(new_n825));
  INV_X1    g0625(.A(new_n787), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n825), .B1(G116), .B2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(G283), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n312), .B1(new_n775), .B2(new_n828), .C1(new_n784), .C2(new_n789), .ZN(new_n829));
  INV_X1    g0629(.A(new_n772), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n829), .B1(G97), .B2(new_n830), .ZN(new_n831));
  OAI211_X1 g0631(.A(new_n827), .B(new_n831), .C1(new_n786), .C2(new_n781), .ZN(new_n832));
  INV_X1    g0632(.A(new_n775), .ZN(new_n833));
  AOI22_X1  g0633(.A1(G143), .A2(new_n768), .B1(new_n833), .B2(G150), .ZN(new_n834));
  NAND2_X1  g0634(.A1(new_n790), .A2(G137), .ZN(new_n835));
  OAI211_X1 g0635(.A(new_n834), .B(new_n835), .C1(new_n372), .C2(new_n787), .ZN(new_n836));
  INV_X1    g0636(.A(KEYINPUT34), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n836), .A2(new_n837), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n779), .A2(new_n209), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n289), .B1(new_n785), .B2(new_n202), .ZN(new_n841));
  AOI211_X1 g0641(.A(new_n840), .B(new_n841), .C1(G58), .C2(new_n830), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n838), .A2(new_n839), .A3(new_n842), .ZN(new_n843));
  INV_X1    g0643(.A(G132), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n781), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n832), .B1(new_n843), .B2(new_n845), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n808), .B1(new_n846), .B2(new_n755), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n755), .A2(new_n756), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI221_X1 g0649(.A(new_n847), .B1(G77), .B2(new_n849), .C1(new_n819), .C2(new_n757), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n822), .A2(new_n850), .ZN(G384));
  OAI21_X1  g0651(.A(new_n411), .B1(KEYINPUT16), .B2(new_n410), .ZN(new_n852));
  AOI21_X1  g0652(.A(new_n683), .B1(new_n852), .B2(new_n391), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n421), .A2(new_n853), .ZN(new_n854));
  OR2_X1    g0654(.A1(new_n412), .A2(new_n683), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  AND2_X1   g0656(.A1(new_n419), .A2(new_n856), .ZN(new_n857));
  AND3_X1   g0657(.A1(new_n392), .A2(KEYINPUT100), .A3(new_n404), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT100), .B1(new_n392), .B2(new_n404), .ZN(new_n859));
  OAI211_X1 g0659(.A(new_n855), .B(new_n857), .C1(new_n858), .C2(new_n859), .ZN(new_n860));
  AOI22_X1  g0660(.A1(new_n852), .A2(new_n391), .B1(new_n413), .B2(new_n683), .ZN(new_n861));
  INV_X1    g0661(.A(new_n419), .ZN(new_n862));
  OAI21_X1  g0662(.A(KEYINPUT37), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n854), .A2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n854), .A2(KEYINPUT38), .A3(new_n864), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g0669(.A(G200), .B1(new_n438), .B2(new_n439), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(KEYINPUT71), .ZN(new_n871));
  AOI211_X1 g0671(.A(new_n454), .B(new_n458), .C1(new_n871), .C2(new_n465), .ZN(new_n872));
  OAI211_X1 g0672(.A(new_n454), .B(new_n685), .C1(new_n872), .C2(new_n446), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n454), .A2(new_n685), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n455), .A2(new_n467), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n873), .A2(new_n875), .ZN(new_n876));
  AND3_X1   g0676(.A1(new_n738), .A2(new_n739), .A3(new_n819), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n869), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT40), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n738), .A2(new_n739), .A3(new_n819), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n881), .B1(new_n875), .B2(new_n873), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n412), .A2(new_n683), .ZN(new_n883));
  INV_X1    g0683(.A(new_n858), .ZN(new_n884));
  INV_X1    g0684(.A(new_n859), .ZN(new_n885));
  AOI21_X1  g0685(.A(new_n883), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(KEYINPUT101), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n413), .B1(new_n387), .B2(new_n391), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n887), .B1(new_n862), .B2(new_n888), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n419), .B(KEYINPUT101), .C1(new_n412), .C2(new_n413), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n889), .A2(new_n855), .A3(new_n890), .ZN(new_n891));
  AOI22_X1  g0691(.A1(new_n857), .A2(new_n886), .B1(new_n891), .B2(KEYINPUT37), .ZN(new_n892));
  INV_X1    g0692(.A(new_n649), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n855), .B1(new_n893), .B2(new_n420), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n866), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n868), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n882), .A2(KEYINPUT40), .A3(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n880), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n489), .A2(new_n740), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n898), .B(new_n899), .Z(new_n900));
  NAND2_X1  g0700(.A1(new_n900), .A2(G330), .ZN(new_n901));
  XNOR2_X1  g0701(.A(new_n901), .B(KEYINPUT102), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n489), .A2(new_n716), .A3(new_n725), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n652), .A2(new_n903), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n902), .B(new_n904), .Z(new_n905));
  NOR2_X1   g0705(.A1(new_n483), .A2(new_n685), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n907), .B1(new_n817), .B2(new_n818), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n869), .A3(new_n876), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n649), .A2(new_n683), .ZN(new_n910));
  INV_X1    g0710(.A(KEYINPUT39), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n896), .A2(new_n911), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n446), .A2(new_n454), .A3(new_n686), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  OAI211_X1 g0714(.A(new_n912), .B(new_n914), .C1(new_n911), .C2(new_n869), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n909), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n905), .B(new_n916), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n252), .B2(new_n679), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n255), .B1(new_n521), .B2(KEYINPUT35), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n230), .C1(KEYINPUT35), .C2(new_n521), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT36), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n369), .A2(G77), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n233), .A2(new_n922), .B1(G50), .B2(new_n209), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n923), .A2(G1), .A3(new_n678), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n918), .A2(new_n921), .A3(new_n924), .ZN(G367));
  INV_X1    g0725(.A(new_n745), .ZN(new_n926));
  OAI221_X1 g0726(.A(new_n759), .B1(new_n225), .B2(new_n606), .C1(new_n242), .C2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n772), .A2(new_n209), .ZN(new_n928));
  INV_X1    g0728(.A(new_n785), .ZN(new_n929));
  AOI22_X1  g0729(.A1(G58), .A2(new_n929), .B1(new_n782), .B2(G137), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n790), .A2(G143), .ZN(new_n931));
  OAI211_X1 g0731(.A(new_n930), .B(new_n931), .C1(new_n372), .C2(new_n775), .ZN(new_n932));
  AOI211_X1 g0732(.A(new_n928), .B(new_n932), .C1(G150), .C2(new_n768), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n289), .B1(new_n779), .B2(new_n205), .ZN(new_n934));
  XOR2_X1   g0734(.A(new_n934), .B(KEYINPUT107), .Z(new_n935));
  OAI211_X1 g0735(.A(new_n933), .B(new_n935), .C1(new_n202), .C2(new_n787), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n767), .A2(new_n784), .ZN(new_n937));
  NOR2_X1   g0737(.A1(new_n779), .A2(new_n264), .ZN(new_n938));
  XNOR2_X1  g0738(.A(KEYINPUT106), .B(G317), .ZN(new_n939));
  OAI22_X1  g0739(.A1(new_n789), .A2(new_n786), .B1(new_n781), .B2(new_n939), .ZN(new_n940));
  AOI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(G294), .C2(new_n833), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n787), .A2(new_n828), .B1(new_n772), .B2(new_n517), .ZN(new_n942));
  XNOR2_X1  g0742(.A(new_n942), .B(KEYINPUT105), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n929), .A2(KEYINPUT46), .A3(G116), .ZN(new_n944));
  AOI21_X1  g0744(.A(KEYINPUT46), .B1(new_n929), .B2(G116), .ZN(new_n945));
  NOR2_X1   g0745(.A1(new_n945), .A2(new_n289), .ZN(new_n946));
  NAND4_X1  g0746(.A1(new_n941), .A2(new_n943), .A3(new_n944), .A4(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n936), .B1(new_n937), .B2(new_n947), .ZN(new_n948));
  XOR2_X1   g0748(.A(new_n948), .B(KEYINPUT47), .Z(new_n949));
  INV_X1    g0749(.A(new_n755), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n764), .B(new_n927), .C1(new_n949), .C2(new_n950), .ZN(new_n951));
  XOR2_X1   g0751(.A(new_n951), .B(KEYINPUT108), .Z(new_n952));
  NAND2_X1  g0752(.A1(new_n661), .A2(new_n685), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n672), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n954), .B1(new_n666), .B2(new_n953), .ZN(new_n955));
  OR2_X1    g0755(.A1(new_n955), .A2(new_n805), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n952), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n656), .A2(new_n685), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n532), .A2(new_n685), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n533), .A2(new_n959), .A3(new_n540), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n958), .A2(new_n960), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n703), .A2(new_n700), .A3(new_n961), .ZN(new_n962));
  XOR2_X1   g0762(.A(KEYINPUT104), .B(KEYINPUT45), .Z(new_n963));
  XNOR2_X1  g0763(.A(new_n962), .B(new_n963), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT44), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n703), .A2(new_n700), .ZN(new_n966));
  INV_X1    g0766(.A(new_n961), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  AOI211_X1 g0768(.A(KEYINPUT44), .B(new_n961), .C1(new_n703), .C2(new_n700), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n699), .B1(new_n964), .B2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n971), .ZN(new_n972));
  OAI21_X1  g0772(.A(new_n703), .B1(new_n692), .B2(new_n702), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n973), .A2(new_n698), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n697), .B(new_n703), .C1(new_n692), .C2(new_n702), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n742), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n964), .A2(new_n970), .A3(new_n699), .ZN(new_n977));
  NAND3_X1  g0777(.A1(new_n972), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n743), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n706), .B(KEYINPUT41), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n763), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT103), .ZN(new_n982));
  OR2_X1    g0782(.A1(new_n703), .A2(new_n960), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n982), .B1(new_n983), .B2(KEYINPUT42), .ZN(new_n984));
  OR4_X1    g0784(.A1(new_n982), .A2(new_n703), .A3(KEYINPUT42), .A4(new_n960), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n983), .A2(KEYINPUT42), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n533), .B1(new_n960), .B2(new_n677), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n686), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n984), .A2(new_n985), .A3(new_n986), .A4(new_n988), .ZN(new_n989));
  NOR2_X1   g0789(.A1(new_n699), .A2(new_n967), .ZN(new_n990));
  INV_X1    g0790(.A(new_n990), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n992));
  NAND3_X1  g0792(.A1(new_n989), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n993), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n991), .B1(new_n989), .B2(new_n992), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n994), .A2(new_n995), .B1(KEYINPUT43), .B2(new_n955), .ZN(new_n996));
  INV_X1    g0796(.A(new_n995), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n955), .A2(KEYINPUT43), .ZN(new_n998));
  NAND3_X1  g0798(.A1(new_n997), .A2(new_n998), .A3(new_n993), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n957), .B1(new_n981), .B2(new_n1000), .ZN(G387));
  NAND2_X1  g0801(.A1(new_n974), .A2(new_n975), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n763), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n782), .A2(G326), .ZN(new_n1004));
  XNOR2_X1  g0804(.A(KEYINPUT109), .B(G322), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n790), .A2(new_n1005), .B1(new_n826), .B2(G303), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n1006), .B1(new_n786), .B2(new_n775), .C1(new_n767), .C2(new_n939), .ZN(new_n1007));
  XNOR2_X1  g0807(.A(new_n1007), .B(KEYINPUT48), .ZN(new_n1008));
  OAI221_X1 g0808(.A(new_n1008), .B1(new_n828), .B2(new_n772), .C1(new_n770), .C2(new_n785), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  AOI211_X1 g0810(.A(new_n289), .B(new_n1004), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n1011), .B1(new_n1010), .B2(new_n1009), .C1(new_n255), .C2(new_n779), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n606), .A2(new_n772), .ZN(new_n1013));
  INV_X1    g0813(.A(G150), .ZN(new_n1014));
  OAI221_X1 g0814(.A(new_n289), .B1(new_n781), .B2(new_n1014), .C1(new_n264), .C2(new_n779), .ZN(new_n1015));
  AOI211_X1 g0815(.A(new_n1013), .B(new_n1015), .C1(G77), .C2(new_n929), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n789), .A2(new_n372), .B1(new_n767), .B2(new_n202), .ZN(new_n1017));
  INV_X1    g0817(.A(new_n335), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1017), .B1(new_n1018), .B2(new_n833), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n1016), .B(new_n1019), .C1(new_n209), .C2(new_n787), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n950), .B1(new_n1012), .B2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n760), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n745), .B1(new_n239), .B2(new_n291), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1023), .B1(new_n708), .B2(new_n750), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n475), .A2(new_n202), .ZN(new_n1025));
  AOI211_X1 g0825(.A(G116), .B(new_n613), .C1(new_n1025), .C2(KEYINPUT50), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(G68), .A2(G77), .ZN(new_n1027));
  OR2_X1    g0827(.A1(new_n1025), .A2(KEYINPUT50), .ZN(new_n1028));
  NAND4_X1  g0828(.A1(new_n1026), .A2(new_n291), .A3(new_n1027), .A4(new_n1028), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n1024), .A2(new_n1029), .B1(new_n517), .B2(new_n705), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n764), .B1(new_n1022), .B2(new_n1030), .C1(new_n692), .C2(new_n805), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n706), .B1(new_n1002), .B2(new_n743), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1003), .B1(new_n1021), .B2(new_n1031), .C1(new_n1032), .C2(new_n976), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n967), .A2(new_n758), .ZN(new_n1034));
  OAI221_X1 g0834(.A(new_n759), .B1(new_n264), .B2(new_n225), .C1(new_n247), .C2(new_n926), .ZN(new_n1035));
  OAI22_X1  g0835(.A1(new_n787), .A2(new_n770), .B1(new_n772), .B2(new_n255), .ZN(new_n1036));
  AOI21_X1  g0836(.A(new_n1036), .B1(G303), .B2(new_n833), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT110), .Z(new_n1038));
  NAND2_X1  g0838(.A1(new_n782), .A2(new_n1005), .ZN(new_n1039));
  AOI22_X1  g0839(.A1(G317), .A2(new_n790), .B1(new_n768), .B2(G311), .ZN(new_n1040));
  XOR2_X1   g0840(.A(new_n1040), .B(KEYINPUT52), .Z(new_n1041));
  AOI211_X1 g0841(.A(new_n289), .B(new_n798), .C1(G283), .C2(new_n929), .ZN(new_n1042));
  NAND4_X1  g0842(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .A4(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n782), .A2(G143), .ZN(new_n1044));
  OAI221_X1 g0844(.A(new_n1044), .B1(new_n202), .B2(new_n775), .C1(new_n330), .C2(new_n787), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n823), .B(new_n1045), .C1(G68), .C2(new_n929), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n830), .A2(G77), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n789), .A2(new_n1014), .B1(new_n767), .B2(new_n372), .ZN(new_n1048));
  XNOR2_X1  g0848(.A(new_n1048), .B(KEYINPUT51), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1043), .B1(new_n1050), .B2(new_n312), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n808), .B1(new_n1051), .B2(new_n755), .ZN(new_n1052));
  AND3_X1   g0852(.A1(new_n1034), .A2(new_n1035), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n976), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n977), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1054), .B1(new_n1055), .B2(new_n971), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1056), .A2(new_n978), .A3(new_n706), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(KEYINPUT111), .ZN(new_n1058));
  INV_X1    g0858(.A(KEYINPUT111), .ZN(new_n1059));
  NAND4_X1  g0859(.A1(new_n1056), .A2(new_n978), .A3(new_n1059), .A4(new_n706), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1053), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n972), .A2(new_n763), .A3(new_n977), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1061), .A2(new_n1062), .ZN(G390));
  NOR2_X1   g0863(.A1(new_n772), .A2(new_n372), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT54), .B(G143), .Z(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n289), .B1(new_n844), .B2(new_n767), .C1(new_n1066), .C2(new_n787), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n1064), .B(new_n1067), .C1(G137), .C2(new_n833), .ZN(new_n1068));
  INV_X1    g0868(.A(G125), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n779), .A2(new_n202), .B1(new_n781), .B2(new_n1069), .ZN(new_n1070));
  NAND3_X1  g0870(.A1(new_n929), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1071));
  INV_X1    g0871(.A(KEYINPUT53), .ZN(new_n1072));
  OAI21_X1  g0872(.A(new_n1072), .B1(new_n785), .B2(new_n1014), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n1070), .B1(new_n1071), .B2(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(G128), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1068), .B(new_n1074), .C1(new_n1075), .C2(new_n789), .ZN(new_n1076));
  XNOR2_X1  g0876(.A(new_n1076), .B(KEYINPUT116), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n767), .A2(new_n255), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n775), .A2(new_n517), .B1(new_n781), .B2(new_n770), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1078), .B(new_n1079), .C1(G283), .C2(new_n790), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n840), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n289), .B(new_n792), .C1(G97), .C2(new_n826), .ZN(new_n1082));
  NAND4_X1  g0882(.A1(new_n1080), .A2(new_n1081), .A3(new_n1047), .A4(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1077), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n808), .B1(new_n1084), .B2(new_n755), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n869), .A2(new_n911), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1086), .B1(new_n911), .B2(new_n896), .ZN(new_n1087));
  OAI221_X1 g0887(.A(new_n1085), .B1(new_n1018), .B2(new_n849), .C1(new_n1087), .C2(new_n757), .ZN(new_n1088));
  XOR2_X1   g0888(.A(new_n1088), .B(KEYINPUT117), .Z(new_n1089));
  AND3_X1   g0889(.A1(new_n455), .A2(new_n467), .A3(new_n874), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n874), .B1(new_n455), .B2(new_n467), .ZN(new_n1091));
  OAI211_X1 g0891(.A(new_n877), .B(G330), .C1(new_n1090), .C2(new_n1091), .ZN(new_n1092));
  AND3_X1   g0892(.A1(new_n655), .A2(new_n659), .A3(new_n668), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n672), .A2(new_n533), .A3(new_n540), .A4(new_n569), .ZN(new_n1094));
  INV_X1    g0894(.A(new_n671), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n666), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n686), .B(new_n816), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT99), .ZN(new_n1098));
  NAND4_X1  g0898(.A1(new_n674), .A2(new_n811), .A3(new_n686), .A4(new_n816), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n906), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NOR2_X1   g0900(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n913), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n912), .B1(new_n911), .B2(new_n869), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n891), .A2(KEYINPUT37), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1105), .A2(new_n860), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n883), .B1(new_n645), .B2(new_n649), .ZN(new_n1107));
  AOI21_X1  g0907(.A(KEYINPUT38), .B1(new_n1106), .B2(new_n1107), .ZN(new_n1108));
  AOI221_X4 g0908(.A(new_n866), .B1(new_n860), .B2(new_n863), .C1(new_n421), .C2(new_n853), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n913), .B1(new_n1108), .B2(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n724), .A2(new_n686), .A3(new_n816), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(new_n907), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n1110), .B1(new_n1112), .B2(new_n876), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1092), .B1(new_n1104), .B2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1092), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1116), .B(new_n1113), .C1(new_n1102), .C2(new_n1103), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1115), .A2(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(KEYINPUT115), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1118), .A2(new_n1119), .A3(new_n763), .ZN(new_n1120));
  AOI21_X1  g0920(.A(new_n914), .B1(new_n908), .B2(new_n876), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1114), .B1(new_n1121), .B2(new_n1087), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n1116), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1104), .A2(new_n1114), .A3(new_n1092), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g0925(.A(KEYINPUT115), .B1(new_n1125), .B2(new_n762), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1089), .A2(new_n1120), .A3(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n738), .A2(new_n739), .A3(G330), .A4(new_n819), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n882), .A2(G330), .B1(new_n1101), .B2(new_n1128), .ZN(new_n1129));
  OAI21_X1  g0929(.A(KEYINPUT112), .B1(new_n1129), .B2(new_n1100), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n1129), .A2(new_n907), .A3(new_n1111), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1128), .A2(new_n873), .A3(new_n875), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1092), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(KEYINPUT112), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n908), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n1130), .A2(new_n1131), .A3(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n489), .A2(G330), .A3(new_n740), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n652), .A2(new_n903), .A3(new_n1137), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1136), .A2(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n1140), .A2(KEYINPUT113), .ZN(new_n1141));
  INV_X1    g0941(.A(KEYINPUT113), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1142), .A3(new_n1139), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n1125), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1123), .A2(new_n1124), .A3(new_n1139), .A4(new_n1136), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1146), .A2(new_n706), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1147), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1145), .A2(new_n1148), .A3(KEYINPUT114), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT114), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1118), .B1(new_n1141), .B2(new_n1143), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n1150), .B1(new_n1151), .B2(new_n1147), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1127), .B1(new_n1149), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g0953(.A(new_n1153), .ZN(G378));
  INV_X1    g0954(.A(KEYINPUT57), .ZN(new_n1155));
  AND3_X1   g0955(.A1(new_n880), .A2(G330), .A3(new_n897), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n916), .A2(new_n1156), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n880), .A2(G330), .A3(new_n897), .ZN(new_n1158));
  NAND4_X1  g0958(.A1(new_n1158), .A2(new_n910), .A3(new_n909), .A4(new_n915), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n357), .A2(KEYINPUT55), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT55), .ZN(new_n1162));
  NOR2_X1   g0962(.A1(new_n356), .A2(new_n1162), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n343), .A2(new_n683), .ZN(new_n1164));
  NOR3_X1   g0964(.A1(new_n1161), .A2(new_n1163), .A3(new_n1164), .ZN(new_n1165));
  INV_X1    g0965(.A(new_n1165), .ZN(new_n1166));
  XNOR2_X1  g0966(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1164), .B1(new_n1161), .B2(new_n1163), .ZN(new_n1168));
  AND3_X1   g0968(.A1(new_n1166), .A2(new_n1167), .A3(new_n1168), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1167), .B1(new_n1166), .B2(new_n1168), .ZN(new_n1170));
  NOR2_X1   g0970(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  NAND2_X1  g0972(.A1(new_n1160), .A2(new_n1172), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(new_n1157), .A2(new_n1159), .A3(new_n1171), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1138), .B1(new_n1118), .B2(new_n1136), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1155), .B1(new_n1175), .B2(new_n1176), .ZN(new_n1177));
  AND3_X1   g0977(.A1(new_n1157), .A2(new_n1171), .A3(new_n1159), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1171), .B1(new_n1157), .B2(new_n1159), .ZN(new_n1179));
  NOR2_X1   g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1146), .A2(new_n1139), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(KEYINPUT57), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1177), .A2(new_n1182), .A3(new_n706), .ZN(new_n1183));
  AOI22_X1  g0983(.A1(new_n790), .A2(G116), .B1(new_n826), .B2(new_n476), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1184), .B1(new_n264), .B2(new_n775), .C1(new_n517), .C2(new_n767), .ZN(new_n1185));
  AOI211_X1 g0985(.A(new_n928), .B(new_n1185), .C1(G283), .C2(new_n782), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n780), .A2(G58), .ZN(new_n1187));
  AOI211_X1 g0987(.A(G41), .B(new_n289), .C1(new_n929), .C2(G77), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT118), .ZN(new_n1189));
  OR2_X1    g0989(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1189), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1186), .A2(new_n1187), .A3(new_n1190), .A4(new_n1191), .ZN(new_n1192));
  XOR2_X1   g0992(.A(new_n1192), .B(KEYINPUT58), .Z(new_n1193));
  OAI22_X1  g0993(.A1(new_n767), .A2(new_n1075), .B1(new_n772), .B2(new_n1014), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n929), .A2(new_n1065), .B1(new_n826), .B2(G137), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1195), .B1(new_n844), .B2(new_n775), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1194), .B(new_n1196), .C1(G125), .C2(new_n790), .ZN(new_n1197));
  XNOR2_X1  g0997(.A(new_n1197), .B(KEYINPUT59), .ZN(new_n1198));
  AOI21_X1  g0998(.A(G41), .B1(new_n782), .B2(G124), .ZN(new_n1199));
  AOI21_X1  g0999(.A(G33), .B1(new_n780), .B2(G159), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1198), .A2(new_n1199), .A3(new_n1200), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G41), .B1(KEYINPUT3), .B2(G33), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1201), .B1(G50), .B2(new_n1202), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n755), .B1(new_n1193), .B2(new_n1203), .ZN(new_n1204));
  AND2_X1   g1004(.A1(new_n1204), .A2(new_n764), .ZN(new_n1205));
  OAI221_X1 g1005(.A(new_n1205), .B1(G50), .B2(new_n849), .C1(new_n1171), .C2(new_n757), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT120), .ZN(new_n1207));
  OR2_X1    g1007(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1209));
  AOI22_X1  g1009(.A1(new_n763), .A2(new_n1180), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1183), .A2(new_n1210), .ZN(G375));
  AND3_X1   g1011(.A1(new_n1133), .A2(new_n1134), .A3(new_n908), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1134), .B1(new_n1133), .B2(new_n908), .ZN(new_n1213));
  NOR2_X1   g1013(.A1(new_n1212), .A2(new_n1213), .ZN(new_n1214));
  INV_X1    g1014(.A(KEYINPUT121), .ZN(new_n1215));
  NAND4_X1  g1015(.A1(new_n1214), .A2(new_n1215), .A3(new_n1138), .A4(new_n1131), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1138), .A2(new_n1130), .A3(new_n1131), .A4(new_n1135), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1217), .A2(KEYINPUT121), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(new_n1216), .A2(new_n1218), .ZN(new_n1219));
  NAND3_X1  g1019(.A1(new_n1144), .A2(new_n980), .A3(new_n1219), .ZN(new_n1220));
  XOR2_X1   g1020(.A(new_n1220), .B(KEYINPUT122), .Z(new_n1221));
  NAND2_X1  g1021(.A1(new_n1136), .A2(new_n763), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n312), .B1(new_n779), .B2(new_n205), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n1223), .B(new_n1013), .C1(G303), .C2(new_n782), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n785), .A2(new_n264), .ZN(new_n1225));
  OAI22_X1  g1025(.A1(new_n767), .A2(new_n828), .B1(new_n787), .B2(new_n517), .ZN(new_n1226));
  AOI211_X1 g1026(.A(new_n1225), .B(new_n1226), .C1(G294), .C2(new_n790), .ZN(new_n1227));
  OAI211_X1 g1027(.A(new_n1224), .B(new_n1227), .C1(new_n255), .C2(new_n775), .ZN(new_n1228));
  OAI22_X1  g1028(.A1(new_n785), .A2(new_n372), .B1(new_n781), .B2(new_n1075), .ZN(new_n1229));
  XOR2_X1   g1029(.A(new_n1229), .B(KEYINPUT123), .Z(new_n1230));
  OAI211_X1 g1030(.A(new_n1230), .B(new_n289), .C1(new_n202), .C2(new_n772), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(G132), .A2(new_n790), .B1(new_n833), .B2(new_n1065), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n826), .A2(G150), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n768), .A2(G137), .ZN(new_n1234));
  NAND4_X1  g1034(.A1(new_n1232), .A2(new_n1187), .A3(new_n1233), .A4(new_n1234), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1228), .B1(new_n1231), .B2(new_n1235), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n808), .B1(new_n1236), .B2(new_n755), .ZN(new_n1237));
  OAI221_X1 g1037(.A(new_n1237), .B1(G68), .B2(new_n849), .C1(new_n876), .C2(new_n757), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1222), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1221), .A2(new_n1240), .ZN(G381));
  OR4_X1    g1041(.A1(G396), .A2(G390), .A3(G384), .A4(G393), .ZN(new_n1242));
  AOI21_X1  g1042(.A(new_n1127), .B1(new_n1145), .B2(new_n1148), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(new_n1183), .A3(new_n1210), .ZN(new_n1244));
  OR4_X1    g1044(.A1(G387), .A2(new_n1242), .A3(G381), .A4(new_n1244), .ZN(G407));
  OAI211_X1 g1045(.A(G407), .B(G213), .C1(G343), .C2(new_n1244), .ZN(G409));
  XNOR2_X1  g1046(.A(G393), .B(G396), .ZN(new_n1247));
  NAND3_X1  g1047(.A1(G387), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1248), .ZN(new_n1249));
  AOI21_X1  g1049(.A(G387), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n1247), .B1(new_n1249), .B2(new_n1250), .ZN(new_n1251));
  INV_X1    g1051(.A(G387), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(G390), .A2(new_n1252), .ZN(new_n1253));
  NOR2_X1   g1053(.A1(new_n1247), .A2(KEYINPUT126), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1253), .A2(new_n1254), .A3(new_n1248), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1249), .A2(KEYINPUT126), .ZN(new_n1256));
  AND3_X1   g1056(.A1(new_n1251), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1251), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT127), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1259), .A2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1127), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1145), .A2(new_n1148), .ZN(new_n1264));
  AND3_X1   g1064(.A1(new_n1180), .A2(new_n1181), .A3(new_n980), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1206), .B1(new_n1175), .B2(new_n762), .ZN(new_n1266));
  OAI211_X1 g1066(.A(new_n1263), .B(new_n1264), .C1(new_n1265), .C2(new_n1266), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1267), .B1(G375), .B2(new_n1153), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n684), .A2(G213), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1268), .A2(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT60), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1271), .A2(KEYINPUT124), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1272), .B1(new_n1136), .B2(new_n1139), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT124), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(KEYINPUT60), .ZN(new_n1275));
  INV_X1    g1075(.A(new_n1275), .ZN(new_n1276));
  AOI22_X1  g1076(.A1(new_n1218), .A2(new_n1216), .B1(new_n1273), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(new_n706), .B1(new_n1217), .B2(new_n1271), .ZN(new_n1278));
  OAI21_X1  g1078(.A(KEYINPUT125), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1278), .ZN(new_n1281));
  XNOR2_X1  g1081(.A(new_n1217), .B(new_n1215), .ZN(new_n1282));
  AOI211_X1 g1082(.A(new_n1275), .B(new_n1272), .C1(new_n1136), .C2(new_n1139), .ZN(new_n1283));
  OAI211_X1 g1083(.A(new_n1280), .B(new_n1281), .C1(new_n1282), .C2(new_n1283), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(new_n1279), .A2(new_n1284), .ZN(new_n1285));
  AOI21_X1  g1085(.A(G384), .B1(new_n1285), .B2(new_n1240), .ZN(new_n1286));
  INV_X1    g1086(.A(G384), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1287), .B(new_n1239), .C1(new_n1279), .C2(new_n1284), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n684), .A2(G213), .A3(G2897), .ZN(new_n1289));
  NOR3_X1   g1089(.A1(new_n1286), .A2(new_n1288), .A3(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1272), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1140), .A2(new_n1276), .A3(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(new_n1219), .A2(new_n1293), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1280), .B1(new_n1294), .B2(new_n1281), .ZN(new_n1295));
  AOI211_X1 g1095(.A(KEYINPUT125), .B(new_n1278), .C1(new_n1219), .C2(new_n1293), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1240), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1287), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1285), .A2(G384), .A3(new_n1240), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1291), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1270), .B1(new_n1290), .B2(new_n1300), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1286), .A2(new_n1288), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1302), .A2(new_n1269), .A3(new_n1268), .ZN(new_n1303));
  AOI21_X1  g1103(.A(KEYINPUT62), .B1(new_n1301), .B2(new_n1303), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1303), .A2(KEYINPUT62), .ZN(new_n1305));
  INV_X1    g1105(.A(KEYINPUT61), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1305), .A2(new_n1306), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1262), .B1(new_n1304), .B2(new_n1307), .ZN(new_n1308));
  OAI21_X1  g1108(.A(new_n1289), .B1(new_n1286), .B2(new_n1288), .ZN(new_n1309));
  NAND3_X1  g1109(.A1(new_n1298), .A2(new_n1299), .A3(new_n1291), .ZN(new_n1310));
  AOI22_X1  g1110(.A1(new_n1309), .A2(new_n1310), .B1(new_n1268), .B2(new_n1269), .ZN(new_n1311));
  INV_X1    g1111(.A(KEYINPUT63), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1303), .B1(new_n1311), .B2(new_n1312), .ZN(new_n1313));
  OR2_X1    g1113(.A1(new_n1303), .A2(new_n1312), .ZN(new_n1314));
  NAND4_X1  g1114(.A1(new_n1313), .A2(new_n1306), .A3(new_n1257), .A4(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1308), .A2(new_n1315), .ZN(G405));
  AND2_X1   g1116(.A1(G375), .A2(new_n1243), .ZN(new_n1317));
  NOR2_X1   g1117(.A1(G375), .A2(new_n1153), .ZN(new_n1318));
  OR3_X1    g1118(.A1(new_n1302), .A2(new_n1317), .A3(new_n1318), .ZN(new_n1319));
  OAI21_X1  g1119(.A(new_n1302), .B1(new_n1317), .B2(new_n1318), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1319), .A2(new_n1320), .ZN(new_n1321));
  NAND2_X1  g1121(.A1(new_n1262), .A2(new_n1321), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1259), .A2(new_n1319), .A3(new_n1261), .A4(new_n1320), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1322), .A2(new_n1323), .ZN(G402));
endmodule


