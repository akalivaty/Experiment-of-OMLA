

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738;

  XNOR2_X1 U371 ( .A(n475), .B(n474), .ZN(n672) );
  NOR2_X2 U372 ( .A1(n539), .A2(n538), .ZN(n540) );
  XNOR2_X2 U373 ( .A(n459), .B(G469), .ZN(n552) );
  NOR2_X1 U374 ( .A1(n546), .A2(n561), .ZN(n375) );
  XNOR2_X1 U375 ( .A(n532), .B(KEYINPUT33), .ZN(n667) );
  XNOR2_X1 U376 ( .A(n517), .B(n516), .ZN(n531) );
  AND2_X1 U377 ( .A1(n669), .A2(n670), .ZN(n550) );
  XOR2_X1 U378 ( .A(KEYINPUT71), .B(G131), .Z(n438) );
  BUF_X1 U379 ( .A(n552), .Z(n350) );
  BUF_X2 U380 ( .A(n545), .Z(n622) );
  NOR2_X1 U381 ( .A1(n529), .A2(n669), .ZN(n548) );
  NOR2_X1 U382 ( .A1(G902), .A2(G237), .ZN(n426) );
  XNOR2_X1 U383 ( .A(n522), .B(n521), .ZN(n529) );
  NOR2_X1 U384 ( .A1(n531), .A2(n520), .ZN(n522) );
  NOR2_X1 U385 ( .A1(n570), .A2(n358), .ZN(n576) );
  XNOR2_X1 U386 ( .A(n360), .B(n359), .ZN(n358) );
  INV_X1 U387 ( .A(KEYINPUT82), .ZN(n359) );
  XNOR2_X1 U388 ( .A(G113), .B(G143), .ZN(n387) );
  AND2_X1 U389 ( .A1(n380), .A2(n381), .ZN(n379) );
  INV_X1 U390 ( .A(KEYINPUT44), .ZN(n381) );
  INV_X1 U391 ( .A(n561), .ZN(n380) );
  OR2_X1 U392 ( .A1(n735), .A2(n543), .ZN(n544) );
  XNOR2_X1 U393 ( .A(n362), .B(n352), .ZN(n536) );
  OR2_X1 U394 ( .A1(n616), .A2(G902), .ZN(n362) );
  XNOR2_X1 U395 ( .A(n511), .B(n510), .ZN(n563) );
  XNOR2_X1 U396 ( .A(n382), .B(n363), .ZN(n720) );
  XNOR2_X1 U397 ( .A(n364), .B(KEYINPUT10), .ZN(n363) );
  INV_X1 U398 ( .A(G140), .ZN(n364) );
  XNOR2_X1 U399 ( .A(n366), .B(n592), .ZN(n365) );
  XNOR2_X1 U400 ( .A(n548), .B(n523), .ZN(n525) );
  NAND2_X1 U401 ( .A1(n658), .A2(KEYINPUT47), .ZN(n360) );
  XNOR2_X1 U402 ( .A(n557), .B(n361), .ZN(n658) );
  INV_X1 U403 ( .A(KEYINPUT104), .ZN(n361) );
  NAND2_X1 U404 ( .A1(n656), .A2(n653), .ZN(n557) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n431) );
  XNOR2_X1 U406 ( .A(n409), .B(n408), .ZN(n719) );
  XNOR2_X1 U407 ( .A(n412), .B(n371), .ZN(n370) );
  XNOR2_X1 U408 ( .A(n411), .B(KEYINPUT18), .ZN(n371) );
  INV_X1 U409 ( .A(n382), .ZN(n412) );
  XNOR2_X1 U410 ( .A(n719), .B(n368), .ZN(n440) );
  XNOR2_X1 U411 ( .A(n410), .B(KEYINPUT68), .ZN(n368) );
  XNOR2_X1 U412 ( .A(KEYINPUT69), .B(G101), .ZN(n410) );
  AND2_X1 U413 ( .A1(n591), .A2(n367), .ZN(n366) );
  NOR2_X1 U414 ( .A1(n586), .A2(n732), .ZN(n367) );
  XNOR2_X1 U415 ( .A(n428), .B(n427), .ZN(n509) );
  XNOR2_X1 U416 ( .A(n418), .B(n455), .ZN(n424) );
  XNOR2_X1 U417 ( .A(n416), .B(KEYINPUT76), .ZN(n418) );
  XNOR2_X1 U418 ( .A(G119), .B(G128), .ZN(n464) );
  XNOR2_X1 U419 ( .A(n392), .B(n391), .ZN(n616) );
  XNOR2_X1 U420 ( .A(n390), .B(n389), .ZN(n391) );
  XNOR2_X1 U421 ( .A(n386), .B(n720), .ZN(n392) );
  NAND2_X1 U422 ( .A1(n377), .A2(n376), .ZN(n378) );
  XNOR2_X1 U423 ( .A(n406), .B(n405), .ZN(n498) );
  XNOR2_X1 U424 ( .A(n536), .B(KEYINPUT100), .ZN(n495) );
  NOR2_X1 U425 ( .A1(n563), .A2(n515), .ZN(n517) );
  BUF_X1 U426 ( .A(n623), .Z(n633) );
  OR2_X1 U427 ( .A1(n723), .A2(G952), .ZN(n627) );
  XNOR2_X1 U428 ( .A(n372), .B(KEYINPUT32), .ZN(n735) );
  NAND2_X1 U429 ( .A1(n530), .A2(n374), .ZN(n373) );
  AND2_X1 U430 ( .A1(n495), .A2(n498), .ZN(n650) );
  XNOR2_X1 U431 ( .A(n527), .B(n526), .ZN(n734) );
  NOR2_X1 U432 ( .A1(n525), .A2(n524), .ZN(n527) );
  NOR2_X1 U433 ( .A1(n705), .A2(n704), .ZN(n706) );
  AND2_X1 U434 ( .A1(n365), .A2(n354), .ZN(n351) );
  XOR2_X1 U435 ( .A(KEYINPUT13), .B(G475), .Z(n352) );
  AND2_X1 U436 ( .A1(G214), .A2(n431), .ZN(n353) );
  AND2_X1 U437 ( .A1(n736), .A2(n598), .ZN(n354) );
  NOR2_X1 U438 ( .A1(n734), .A2(n544), .ZN(n355) );
  NAND2_X1 U439 ( .A1(n542), .A2(n541), .ZN(n356) );
  XOR2_X1 U440 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n357) );
  XNOR2_X1 U441 ( .A(n369), .B(n440), .ZN(n425) );
  XNOR2_X1 U442 ( .A(n415), .B(n370), .ZN(n369) );
  NOR2_X1 U443 ( .A1(n529), .A2(n373), .ZN(n372) );
  INV_X1 U444 ( .A(n580), .ZN(n374) );
  NAND2_X1 U445 ( .A1(n375), .A2(n355), .ZN(n376) );
  NAND2_X1 U446 ( .A1(n356), .A2(n379), .ZN(n377) );
  XNOR2_X2 U447 ( .A(n378), .B(n357), .ZN(n695) );
  XNOR2_X1 U448 ( .A(n404), .B(n403), .ZN(n629) );
  XNOR2_X1 U449 ( .A(n402), .B(n401), .ZN(n403) );
  INV_X1 U450 ( .A(KEYINPUT17), .ZN(n411) );
  XNOR2_X1 U451 ( .A(G125), .B(G146), .ZN(n382) );
  XNOR2_X1 U452 ( .A(n385), .B(n353), .ZN(n386) );
  INV_X1 U453 ( .A(KEYINPUT19), .ZN(n510) );
  INV_X1 U454 ( .A(n599), .ZN(n600) );
  INV_X1 U455 ( .A(KEYINPUT108), .ZN(n523) );
  XNOR2_X1 U456 ( .A(n540), .B(KEYINPUT35), .ZN(n545) );
  INV_X1 U457 ( .A(n624), .ZN(n625) );
  INV_X1 U458 ( .A(KEYINPUT109), .ZN(n526) );
  XNOR2_X1 U459 ( .A(n626), .B(n625), .ZN(n628) );
  XOR2_X1 U460 ( .A(KEYINPUT98), .B(KEYINPUT12), .Z(n384) );
  XNOR2_X1 U461 ( .A(KEYINPUT97), .B(KEYINPUT99), .ZN(n383) );
  XNOR2_X1 U462 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U463 ( .A(n438), .B(KEYINPUT11), .Z(n390) );
  XOR2_X1 U464 ( .A(G122), .B(G104), .Z(n388) );
  XNOR2_X1 U465 ( .A(n388), .B(n387), .ZN(n389) );
  INV_X1 U466 ( .A(n495), .ZN(n407) );
  XOR2_X1 U467 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n395) );
  INV_X1 U468 ( .A(KEYINPUT64), .ZN(n393) );
  XNOR2_X2 U469 ( .A(n393), .B(G953), .ZN(n723) );
  NAND2_X1 U470 ( .A1(G234), .A2(n723), .ZN(n394) );
  XNOR2_X1 U471 ( .A(n395), .B(n394), .ZN(n463) );
  NAND2_X1 U472 ( .A1(G217), .A2(n463), .ZN(n404) );
  XNOR2_X2 U473 ( .A(G143), .B(G128), .ZN(n409) );
  XOR2_X1 U474 ( .A(G122), .B(G116), .Z(n396) );
  XNOR2_X1 U475 ( .A(n409), .B(n396), .ZN(n400) );
  XOR2_X1 U476 ( .A(KEYINPUT101), .B(KEYINPUT9), .Z(n398) );
  XNOR2_X1 U477 ( .A(G107), .B(KEYINPUT102), .ZN(n397) );
  XNOR2_X1 U478 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U479 ( .A(n400), .B(n399), .Z(n402) );
  XOR2_X1 U480 ( .A(G134), .B(KEYINPUT7), .Z(n401) );
  INV_X1 U481 ( .A(G902), .ZN(n470) );
  NAND2_X1 U482 ( .A1(n629), .A2(n470), .ZN(n406) );
  XNOR2_X1 U483 ( .A(KEYINPUT103), .B(G478), .ZN(n405) );
  INV_X1 U484 ( .A(n498), .ZN(n535) );
  NAND2_X1 U485 ( .A1(n407), .A2(n535), .ZN(n656) );
  INV_X1 U486 ( .A(n656), .ZN(n646) );
  INV_X1 U487 ( .A(KEYINPUT4), .ZN(n408) );
  XOR2_X1 U488 ( .A(KEYINPUT80), .B(KEYINPUT88), .Z(n414) );
  NAND2_X1 U489 ( .A1(G224), .A2(n723), .ZN(n413) );
  XNOR2_X1 U490 ( .A(n414), .B(n413), .ZN(n415) );
  XOR2_X1 U491 ( .A(KEYINPUT16), .B(G122), .Z(n416) );
  XNOR2_X1 U492 ( .A(G104), .B(G110), .ZN(n417) );
  XNOR2_X1 U493 ( .A(n417), .B(G107), .ZN(n455) );
  XNOR2_X1 U494 ( .A(G119), .B(G116), .ZN(n421) );
  INV_X1 U495 ( .A(KEYINPUT72), .ZN(n419) );
  XNOR2_X1 U496 ( .A(n419), .B(KEYINPUT73), .ZN(n420) );
  XNOR2_X1 U497 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U498 ( .A(G113), .B(KEYINPUT3), .Z(n422) );
  XNOR2_X1 U499 ( .A(n423), .B(n422), .ZN(n436) );
  XNOR2_X1 U500 ( .A(n424), .B(n436), .ZN(n713) );
  XNOR2_X1 U501 ( .A(n425), .B(n713), .ZN(n608) );
  XNOR2_X1 U502 ( .A(KEYINPUT15), .B(G902), .ZN(n599) );
  NAND2_X1 U503 ( .A1(n608), .A2(n599), .ZN(n428) );
  XNOR2_X1 U504 ( .A(KEYINPUT77), .B(n426), .ZN(n446) );
  AND2_X1 U505 ( .A1(n446), .A2(G210), .ZN(n427) );
  BUF_X1 U506 ( .A(n509), .Z(n429) );
  INV_X1 U507 ( .A(KEYINPUT38), .ZN(n430) );
  XNOR2_X1 U508 ( .A(n429), .B(n430), .ZN(n662) );
  NAND2_X1 U509 ( .A1(n431), .A2(G210), .ZN(n432) );
  XNOR2_X1 U510 ( .A(n432), .B(KEYINPUT78), .ZN(n434) );
  XNOR2_X1 U511 ( .A(KEYINPUT95), .B(KEYINPUT5), .ZN(n433) );
  XNOR2_X1 U512 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U513 ( .A(n436), .B(n435), .ZN(n439) );
  XNOR2_X1 U514 ( .A(G137), .B(G134), .ZN(n437) );
  XNOR2_X1 U515 ( .A(n438), .B(n437), .ZN(n456) );
  XNOR2_X1 U516 ( .A(n439), .B(n456), .ZN(n442) );
  XNOR2_X1 U517 ( .A(n440), .B(G146), .ZN(n454) );
  INV_X1 U518 ( .A(n454), .ZN(n441) );
  XNOR2_X1 U519 ( .A(n442), .B(n441), .ZN(n603) );
  NAND2_X1 U520 ( .A1(n603), .A2(n470), .ZN(n445) );
  XNOR2_X1 U521 ( .A(KEYINPUT96), .B(G472), .ZN(n443) );
  XNOR2_X1 U522 ( .A(n443), .B(KEYINPUT75), .ZN(n444) );
  XNOR2_X1 U523 ( .A(n445), .B(n444), .ZN(n555) );
  NAND2_X1 U524 ( .A1(n446), .A2(G214), .ZN(n661) );
  INV_X1 U525 ( .A(n661), .ZN(n447) );
  OR2_X1 U526 ( .A1(n555), .A2(n447), .ZN(n450) );
  INV_X1 U527 ( .A(KEYINPUT112), .ZN(n448) );
  XNOR2_X1 U528 ( .A(n448), .B(KEYINPUT30), .ZN(n449) );
  XNOR2_X1 U529 ( .A(n450), .B(n449), .ZN(n491) );
  XOR2_X1 U530 ( .A(G140), .B(KEYINPUT79), .Z(n452) );
  NAND2_X1 U531 ( .A1(G227), .A2(n723), .ZN(n451) );
  XNOR2_X1 U532 ( .A(n452), .B(n451), .ZN(n453) );
  XNOR2_X1 U533 ( .A(n454), .B(n453), .ZN(n458) );
  XOR2_X1 U534 ( .A(KEYINPUT91), .B(n456), .Z(n721) );
  XNOR2_X1 U535 ( .A(n455), .B(n721), .ZN(n457) );
  XNOR2_X1 U536 ( .A(n458), .B(n457), .ZN(n635) );
  NAND2_X1 U537 ( .A1(n635), .A2(n470), .ZN(n459) );
  XOR2_X1 U538 ( .A(KEYINPUT92), .B(KEYINPUT83), .Z(n461) );
  XNOR2_X1 U539 ( .A(KEYINPUT24), .B(KEYINPUT23), .ZN(n460) );
  XNOR2_X1 U540 ( .A(n461), .B(n460), .ZN(n462) );
  XOR2_X1 U541 ( .A(n720), .B(n462), .Z(n469) );
  NAND2_X1 U542 ( .A1(n463), .A2(G221), .ZN(n467) );
  XOR2_X1 U543 ( .A(G110), .B(G137), .Z(n465) );
  XNOR2_X1 U544 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U545 ( .A(n467), .B(n466), .ZN(n468) );
  XNOR2_X1 U546 ( .A(n469), .B(n468), .ZN(n624) );
  NAND2_X1 U547 ( .A1(n624), .A2(n470), .ZN(n475) );
  XOR2_X1 U548 ( .A(KEYINPUT20), .B(KEYINPUT93), .Z(n472) );
  NAND2_X1 U549 ( .A1(G234), .A2(n599), .ZN(n471) );
  XNOR2_X1 U550 ( .A(n472), .B(n471), .ZN(n484) );
  NAND2_X1 U551 ( .A1(n484), .A2(G217), .ZN(n473) );
  XNOR2_X1 U552 ( .A(n473), .B(KEYINPUT25), .ZN(n474) );
  NAND2_X1 U553 ( .A1(G234), .A2(G237), .ZN(n476) );
  XNOR2_X1 U554 ( .A(n476), .B(KEYINPUT14), .ZN(n481) );
  NAND2_X1 U555 ( .A1(n481), .A2(G902), .ZN(n477) );
  XNOR2_X1 U556 ( .A(n477), .B(KEYINPUT90), .ZN(n512) );
  OR2_X1 U557 ( .A1(n723), .A2(n512), .ZN(n478) );
  NOR2_X1 U558 ( .A1(G900), .A2(n478), .ZN(n480) );
  INV_X1 U559 ( .A(KEYINPUT110), .ZN(n479) );
  XNOR2_X1 U560 ( .A(n480), .B(n479), .ZN(n483) );
  NAND2_X1 U561 ( .A1(G952), .A2(n481), .ZN(n688) );
  NOR2_X1 U562 ( .A1(n688), .A2(G953), .ZN(n514) );
  INV_X1 U563 ( .A(n514), .ZN(n482) );
  NAND2_X1 U564 ( .A1(n483), .A2(n482), .ZN(n487) );
  NAND2_X1 U565 ( .A1(n484), .A2(G221), .ZN(n485) );
  XNOR2_X1 U566 ( .A(n485), .B(KEYINPUT21), .ZN(n673) );
  INV_X1 U567 ( .A(n673), .ZN(n486) );
  AND2_X1 U568 ( .A1(n487), .A2(n486), .ZN(n577) );
  INV_X1 U569 ( .A(n577), .ZN(n488) );
  NOR2_X1 U570 ( .A1(n672), .A2(n488), .ZN(n489) );
  AND2_X1 U571 ( .A1(n350), .A2(n489), .ZN(n490) );
  NAND2_X1 U572 ( .A1(n491), .A2(n490), .ZN(n572) );
  INV_X1 U573 ( .A(n572), .ZN(n492) );
  NAND2_X1 U574 ( .A1(n662), .A2(n492), .ZN(n494) );
  XNOR2_X1 U575 ( .A(KEYINPUT74), .B(KEYINPUT39), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n494), .B(n493), .ZN(n496) );
  NAND2_X1 U577 ( .A1(n646), .A2(n496), .ZN(n598) );
  XNOR2_X1 U578 ( .A(n598), .B(G134), .ZN(G36) );
  NAND2_X1 U579 ( .A1(n650), .A2(n496), .ZN(n497) );
  XNOR2_X1 U580 ( .A(n497), .B(KEYINPUT40), .ZN(n587) );
  XNOR2_X1 U581 ( .A(n587), .B(G131), .ZN(G33) );
  INV_X1 U582 ( .A(n536), .ZN(n499) );
  NAND2_X1 U583 ( .A1(n499), .A2(n498), .ZN(n664) );
  NAND2_X1 U584 ( .A1(n662), .A2(n661), .ZN(n659) );
  NOR2_X1 U585 ( .A1(n664), .A2(n659), .ZN(n500) );
  XNOR2_X1 U586 ( .A(n500), .B(KEYINPUT41), .ZN(n691) );
  NAND2_X1 U587 ( .A1(n672), .A2(n577), .ZN(n501) );
  OR2_X1 U588 ( .A1(n555), .A2(n501), .ZN(n503) );
  XNOR2_X1 U589 ( .A(KEYINPUT115), .B(KEYINPUT28), .ZN(n502) );
  XNOR2_X1 U590 ( .A(n503), .B(n502), .ZN(n564) );
  INV_X1 U591 ( .A(KEYINPUT114), .ZN(n504) );
  XNOR2_X1 U592 ( .A(n350), .B(n504), .ZN(n562) );
  INV_X1 U593 ( .A(n562), .ZN(n505) );
  NAND2_X1 U594 ( .A1(n564), .A2(n505), .ZN(n506) );
  NOR2_X1 U595 ( .A1(n691), .A2(n506), .ZN(n508) );
  XOR2_X1 U596 ( .A(KEYINPUT116), .B(KEYINPUT42), .Z(n507) );
  XNOR2_X1 U597 ( .A(n508), .B(n507), .ZN(n588) );
  XNOR2_X1 U598 ( .A(n588), .B(G137), .ZN(G39) );
  NAND2_X1 U599 ( .A1(n509), .A2(n661), .ZN(n511) );
  XNOR2_X1 U600 ( .A(G898), .B(KEYINPUT89), .ZN(n710) );
  NAND2_X1 U601 ( .A1(G953), .A2(n710), .ZN(n715) );
  NOR2_X1 U602 ( .A1(n715), .A2(n512), .ZN(n513) );
  NOR2_X1 U603 ( .A1(n514), .A2(n513), .ZN(n515) );
  XNOR2_X1 U604 ( .A(KEYINPUT67), .B(KEYINPUT0), .ZN(n516) );
  INV_X1 U605 ( .A(n664), .ZN(n518) );
  NAND2_X1 U606 ( .A1(n518), .A2(n486), .ZN(n519) );
  XOR2_X1 U607 ( .A(KEYINPUT105), .B(n519), .Z(n520) );
  INV_X1 U608 ( .A(KEYINPUT22), .ZN(n521) );
  XNOR2_X2 U609 ( .A(n552), .B(KEYINPUT1), .ZN(n669) );
  NAND2_X1 U610 ( .A1(n555), .A2(n672), .ZN(n524) );
  NAND2_X1 U611 ( .A1(n672), .A2(n669), .ZN(n528) );
  XNOR2_X1 U612 ( .A(n528), .B(KEYINPUT107), .ZN(n530) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT6), .ZN(n580) );
  NOR2_X1 U614 ( .A1(n734), .A2(n735), .ZN(n542) );
  INV_X1 U615 ( .A(n531), .ZN(n533) );
  NOR2_X1 U616 ( .A1(n672), .A2(n673), .ZN(n670) );
  NAND2_X1 U617 ( .A1(n550), .A2(n580), .ZN(n532) );
  NAND2_X1 U618 ( .A1(n533), .A2(n667), .ZN(n534) );
  XNOR2_X1 U619 ( .A(n534), .B(KEYINPUT34), .ZN(n539) );
  AND2_X1 U620 ( .A1(n536), .A2(n535), .ZN(n571) );
  INV_X1 U621 ( .A(n571), .ZN(n537) );
  XOR2_X1 U622 ( .A(KEYINPUT81), .B(n537), .Z(n538) );
  XNOR2_X1 U623 ( .A(n545), .B(KEYINPUT70), .ZN(n541) );
  NAND2_X1 U624 ( .A1(KEYINPUT44), .A2(KEYINPUT70), .ZN(n543) );
  INV_X1 U625 ( .A(n622), .ZN(n546) );
  NOR2_X1 U626 ( .A1(n580), .A2(n672), .ZN(n547) );
  NAND2_X1 U627 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U628 ( .A(n549), .B(KEYINPUT106), .ZN(n738) );
  INV_X1 U629 ( .A(n555), .ZN(n676) );
  NAND2_X1 U630 ( .A1(n550), .A2(n676), .ZN(n680) );
  NOR2_X1 U631 ( .A1(n531), .A2(n680), .ZN(n551) );
  XNOR2_X1 U632 ( .A(n551), .B(KEYINPUT31), .ZN(n655) );
  NAND2_X1 U633 ( .A1(n350), .A2(n670), .ZN(n553) );
  NOR2_X1 U634 ( .A1(n531), .A2(n553), .ZN(n554) );
  XNOR2_X1 U635 ( .A(KEYINPUT94), .B(n554), .ZN(n556) );
  NAND2_X1 U636 ( .A1(n556), .A2(n555), .ZN(n643) );
  NAND2_X1 U637 ( .A1(n655), .A2(n643), .ZN(n559) );
  INV_X1 U638 ( .A(n650), .ZN(n653) );
  INV_X1 U639 ( .A(n658), .ZN(n558) );
  NAND2_X1 U640 ( .A1(n559), .A2(n558), .ZN(n560) );
  NAND2_X1 U641 ( .A1(n738), .A2(n560), .ZN(n561) );
  NOR2_X1 U642 ( .A1(n658), .A2(KEYINPUT47), .ZN(n566) );
  NOR2_X1 U643 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n567) );
  NOR2_X1 U645 ( .A1(n566), .A2(n567), .ZN(n569) );
  INV_X1 U646 ( .A(n567), .ZN(n651) );
  NOR2_X1 U647 ( .A1(n651), .A2(KEYINPUT47), .ZN(n568) );
  NOR2_X1 U648 ( .A1(n569), .A2(n568), .ZN(n570) );
  NAND2_X1 U649 ( .A1(n571), .A2(n429), .ZN(n573) );
  NOR2_X1 U650 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U651 ( .A(n574), .B(KEYINPUT113), .Z(n731) );
  INV_X1 U652 ( .A(n731), .ZN(n575) );
  NAND2_X1 U653 ( .A1(n576), .A2(n575), .ZN(n586) );
  NAND2_X1 U654 ( .A1(n577), .A2(n661), .ZN(n579) );
  NAND2_X1 U655 ( .A1(n672), .A2(n650), .ZN(n578) );
  NOR2_X1 U656 ( .A1(n579), .A2(n578), .ZN(n581) );
  AND2_X1 U657 ( .A1(n581), .A2(n580), .ZN(n594) );
  NAND2_X1 U658 ( .A1(n594), .A2(n429), .ZN(n583) );
  INV_X1 U659 ( .A(KEYINPUT36), .ZN(n582) );
  XNOR2_X1 U660 ( .A(n583), .B(n582), .ZN(n584) );
  NAND2_X1 U661 ( .A1(n584), .A2(n669), .ZN(n585) );
  XNOR2_X1 U662 ( .A(n585), .B(KEYINPUT117), .ZN(n732) );
  NAND2_X1 U663 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U664 ( .A(KEYINPUT65), .B(KEYINPUT46), .ZN(n589) );
  XNOR2_X1 U665 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U666 ( .A(KEYINPUT86), .B(KEYINPUT48), .ZN(n592) );
  INV_X1 U667 ( .A(n669), .ZN(n593) );
  NAND2_X1 U668 ( .A1(n594), .A2(n593), .ZN(n595) );
  XOR2_X1 U669 ( .A(n595), .B(KEYINPUT43), .Z(n596) );
  NOR2_X1 U670 ( .A1(n596), .A2(n429), .ZN(n597) );
  XNOR2_X1 U671 ( .A(n597), .B(KEYINPUT111), .ZN(n736) );
  NAND2_X1 U672 ( .A1(n695), .A2(n351), .ZN(n699) );
  INV_X1 U673 ( .A(KEYINPUT2), .ZN(n697) );
  XNOR2_X1 U674 ( .A(n699), .B(KEYINPUT2), .ZN(n601) );
  AND2_X2 U675 ( .A1(n601), .A2(n600), .ZN(n623) );
  NAND2_X1 U676 ( .A1(n623), .A2(G472), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT87), .B(KEYINPUT62), .Z(n602) );
  XNOR2_X1 U678 ( .A(n603), .B(n602), .ZN(n604) );
  XNOR2_X1 U679 ( .A(n605), .B(n604), .ZN(n606) );
  NAND2_X1 U680 ( .A1(n606), .A2(n627), .ZN(n607) );
  XNOR2_X1 U681 ( .A(n607), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U682 ( .A1(n623), .A2(G210), .ZN(n612) );
  XNOR2_X1 U683 ( .A(KEYINPUT124), .B(KEYINPUT54), .ZN(n609) );
  XOR2_X1 U684 ( .A(n609), .B(KEYINPUT55), .Z(n610) );
  XNOR2_X1 U685 ( .A(n608), .B(n610), .ZN(n611) );
  XNOR2_X1 U686 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U687 ( .A1(n613), .A2(n627), .ZN(n615) );
  INV_X1 U688 ( .A(KEYINPUT56), .ZN(n614) );
  XNOR2_X1 U689 ( .A(n615), .B(n614), .ZN(G51) );
  NAND2_X1 U690 ( .A1(n623), .A2(G475), .ZN(n618) );
  XNOR2_X1 U691 ( .A(n616), .B(KEYINPUT59), .ZN(n617) );
  XNOR2_X1 U692 ( .A(n618), .B(n617), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n619), .A2(n627), .ZN(n621) );
  INV_X1 U694 ( .A(KEYINPUT60), .ZN(n620) );
  XNOR2_X1 U695 ( .A(n621), .B(n620), .ZN(G60) );
  XNOR2_X1 U696 ( .A(n622), .B(G122), .ZN(G24) );
  NAND2_X1 U697 ( .A1(n633), .A2(G217), .ZN(n626) );
  INV_X1 U698 ( .A(n627), .ZN(n638) );
  NOR2_X1 U699 ( .A1(n628), .A2(n638), .ZN(G66) );
  NAND2_X1 U700 ( .A1(n633), .A2(G478), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n629), .B(KEYINPUT125), .ZN(n630) );
  XNOR2_X1 U702 ( .A(n631), .B(n630), .ZN(n632) );
  NOR2_X1 U703 ( .A1(n632), .A2(n638), .ZN(G63) );
  NAND2_X1 U704 ( .A1(n633), .A2(G469), .ZN(n637) );
  XNOR2_X1 U705 ( .A(KEYINPUT57), .B(KEYINPUT58), .ZN(n634) );
  XNOR2_X1 U706 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U707 ( .A(n637), .B(n636), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n639), .A2(n638), .ZN(G54) );
  NOR2_X1 U709 ( .A1(n643), .A2(n653), .ZN(n640) );
  XOR2_X1 U710 ( .A(G104), .B(n640), .Z(G6) );
  XOR2_X1 U711 ( .A(KEYINPUT26), .B(KEYINPUT118), .Z(n642) );
  XNOR2_X1 U712 ( .A(G107), .B(KEYINPUT27), .ZN(n641) );
  XNOR2_X1 U713 ( .A(n642), .B(n641), .ZN(n645) );
  NOR2_X1 U714 ( .A1(n643), .A2(n656), .ZN(n644) );
  XOR2_X1 U715 ( .A(n645), .B(n644), .Z(G9) );
  XOR2_X1 U716 ( .A(KEYINPUT29), .B(KEYINPUT119), .Z(n648) );
  NAND2_X1 U717 ( .A1(n651), .A2(n646), .ZN(n647) );
  XNOR2_X1 U718 ( .A(n648), .B(n647), .ZN(n649) );
  XOR2_X1 U719 ( .A(G128), .B(n649), .Z(G30) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(n652), .B(G146), .ZN(G48) );
  NOR2_X1 U722 ( .A1(n653), .A2(n655), .ZN(n654) );
  XOR2_X1 U723 ( .A(G113), .B(n654), .Z(G15) );
  NOR2_X1 U724 ( .A1(n656), .A2(n655), .ZN(n657) );
  XOR2_X1 U725 ( .A(G116), .B(n657), .Z(G18) );
  NOR2_X1 U726 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U727 ( .A(KEYINPUT122), .B(n660), .ZN(n666) );
  NOR2_X1 U728 ( .A1(n662), .A2(n661), .ZN(n663) );
  NOR2_X1 U729 ( .A1(n664), .A2(n663), .ZN(n665) );
  NOR2_X1 U730 ( .A1(n666), .A2(n665), .ZN(n668) );
  INV_X1 U731 ( .A(n667), .ZN(n690) );
  NOR2_X1 U732 ( .A1(n668), .A2(n690), .ZN(n685) );
  NOR2_X1 U733 ( .A1(n670), .A2(n669), .ZN(n671) );
  XOR2_X1 U734 ( .A(KEYINPUT50), .B(n671), .Z(n679) );
  XOR2_X1 U735 ( .A(KEYINPUT121), .B(KEYINPUT49), .Z(n675) );
  NAND2_X1 U736 ( .A1(n673), .A2(n672), .ZN(n674) );
  XNOR2_X1 U737 ( .A(n675), .B(n674), .ZN(n677) );
  NOR2_X1 U738 ( .A1(n677), .A2(n676), .ZN(n678) );
  NAND2_X1 U739 ( .A1(n679), .A2(n678), .ZN(n681) );
  NAND2_X1 U740 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U741 ( .A(KEYINPUT51), .B(n682), .ZN(n683) );
  NOR2_X1 U742 ( .A1(n683), .A2(n691), .ZN(n684) );
  NOR2_X1 U743 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U744 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  NOR2_X1 U745 ( .A1(n688), .A2(n687), .ZN(n689) );
  XNOR2_X1 U746 ( .A(KEYINPUT123), .B(n689), .ZN(n694) );
  NOR2_X1 U747 ( .A1(n691), .A2(n690), .ZN(n692) );
  NOR2_X1 U748 ( .A1(n692), .A2(G953), .ZN(n693) );
  NAND2_X1 U749 ( .A1(n694), .A2(n693), .ZN(n705) );
  XNOR2_X1 U750 ( .A(n695), .B(KEYINPUT85), .ZN(n696) );
  NOR2_X1 U751 ( .A1(n696), .A2(KEYINPUT2), .ZN(n701) );
  NOR2_X1 U752 ( .A1(n697), .A2(KEYINPUT85), .ZN(n698) );
  AND2_X1 U753 ( .A1(n699), .A2(n698), .ZN(n700) );
  NOR2_X1 U754 ( .A1(n701), .A2(n700), .ZN(n703) );
  NOR2_X1 U755 ( .A1(n351), .A2(KEYINPUT2), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n703), .A2(n702), .ZN(n704) );
  XNOR2_X1 U757 ( .A(KEYINPUT53), .B(n706), .ZN(G75) );
  INV_X1 U758 ( .A(n695), .ZN(n707) );
  NOR2_X1 U759 ( .A1(n707), .A2(G953), .ZN(n712) );
  NAND2_X1 U760 ( .A1(G953), .A2(G224), .ZN(n708) );
  XOR2_X1 U761 ( .A(KEYINPUT61), .B(n708), .Z(n709) );
  NOR2_X1 U762 ( .A1(n710), .A2(n709), .ZN(n711) );
  NOR2_X1 U763 ( .A1(n712), .A2(n711), .ZN(n718) );
  XOR2_X1 U764 ( .A(G101), .B(n713), .Z(n714) );
  NAND2_X1 U765 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U766 ( .A(n716), .B(KEYINPUT126), .ZN(n717) );
  XNOR2_X1 U767 ( .A(n718), .B(n717), .ZN(G69) );
  XOR2_X1 U768 ( .A(n720), .B(n719), .Z(n722) );
  XNOR2_X1 U769 ( .A(n722), .B(n721), .ZN(n725) );
  XOR2_X1 U770 ( .A(n725), .B(n351), .Z(n724) );
  NAND2_X1 U771 ( .A1(n724), .A2(n723), .ZN(n730) );
  XNOR2_X1 U772 ( .A(G227), .B(n725), .ZN(n726) );
  NAND2_X1 U773 ( .A1(n726), .A2(G900), .ZN(n727) );
  XOR2_X1 U774 ( .A(KEYINPUT127), .B(n727), .Z(n728) );
  NAND2_X1 U775 ( .A1(G953), .A2(n728), .ZN(n729) );
  NAND2_X1 U776 ( .A1(n730), .A2(n729), .ZN(G72) );
  XOR2_X1 U777 ( .A(G143), .B(n731), .Z(G45) );
  XNOR2_X1 U778 ( .A(G125), .B(n732), .ZN(n733) );
  XNOR2_X1 U779 ( .A(n733), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U780 ( .A(n734), .B(G110), .Z(G12) );
  XOR2_X1 U781 ( .A(G119), .B(n735), .Z(G21) );
  XNOR2_X1 U782 ( .A(G140), .B(KEYINPUT120), .ZN(n737) );
  XNOR2_X1 U783 ( .A(n737), .B(n736), .ZN(G42) );
  XNOR2_X1 U784 ( .A(G101), .B(n738), .ZN(G3) );
endmodule

