//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 0 1 0 0 0 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:21 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1231,
    new_n1232, new_n1233, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1301, new_n1302;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(new_n206));
  XNOR2_X1  g0006(.A(new_n206), .B(KEYINPUT64), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT0), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G238), .ZN(new_n216));
  INV_X1    g0016(.A(G87), .ZN(new_n217));
  INV_X1    g0017(.A(G250), .ZN(new_n218));
  OAI221_X1 g0018(.A(new_n215), .B1(new_n203), .B2(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n211), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OR2_X1    g0023(.A1(new_n223), .A2(KEYINPUT1), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(new_n203), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n225), .A2(G50), .ZN(new_n226));
  XOR2_X1   g0026(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  NAND2_X1  g0027(.A1(G1), .A2(G13), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n228), .A2(new_n209), .ZN(new_n229));
  INV_X1    g0029(.A(new_n229), .ZN(new_n230));
  OR2_X1    g0030(.A1(new_n227), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n214), .A2(new_n224), .A3(new_n231), .ZN(new_n232));
  AOI21_X1  g0032(.A(new_n232), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n234), .B(KEYINPUT66), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G238), .B(G244), .ZN(new_n238));
  INV_X1    g0038(.A(G232), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n238), .B(new_n239), .ZN(new_n240));
  XNOR2_X1  g0040(.A(KEYINPUT2), .B(G226), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n237), .B(new_n242), .ZN(G358));
  NAND2_X1  g0043(.A1(new_n201), .A2(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n203), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XOR2_X1   g0049(.A(G87), .B(G97), .Z(new_n250));
  XOR2_X1   g0050(.A(G107), .B(G116), .Z(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XNOR2_X1  g0052(.A(new_n249), .B(new_n252), .ZN(G351));
  INV_X1    g0053(.A(KEYINPUT81), .ZN(new_n254));
  XNOR2_X1  g0054(.A(KEYINPUT5), .B(G41), .ZN(new_n255));
  INV_X1    g0055(.A(G45), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(G1), .ZN(new_n257));
  INV_X1    g0057(.A(new_n228), .ZN(new_n258));
  NAND2_X1  g0058(.A1(G33), .A2(G41), .ZN(new_n259));
  AOI22_X1  g0059(.A1(new_n255), .A2(new_n257), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n261));
  AOI21_X1  g0061(.A(new_n261), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  AOI22_X1  g0062(.A1(new_n260), .A2(G270), .B1(new_n255), .B2(new_n262), .ZN(new_n263));
  AND2_X1   g0063(.A1(KEYINPUT3), .A2(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(KEYINPUT3), .A2(G33), .ZN(new_n265));
  OAI211_X1 g0065(.A(G264), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G1698), .ZN(new_n267));
  OAI211_X1 g0067(.A(G257), .B(new_n267), .C1(new_n264), .C2(new_n265), .ZN(new_n268));
  OR2_X1    g0068(.A1(KEYINPUT3), .A2(G33), .ZN(new_n269));
  NAND2_X1  g0069(.A1(KEYINPUT3), .A2(G33), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n269), .A2(G303), .A3(new_n270), .ZN(new_n271));
  NAND3_X1  g0071(.A1(new_n266), .A2(new_n268), .A3(new_n271), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n259), .A2(G1), .A3(G13), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(new_n263), .A2(new_n275), .A3(G190), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n208), .A2(G13), .A3(G20), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G116), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n208), .A2(G33), .ZN(new_n281));
  NAND3_X1  g0081(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n282));
  NAND4_X1  g0082(.A1(new_n277), .A2(new_n281), .A3(new_n228), .A4(new_n282), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n283), .B2(new_n279), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n282), .A2(new_n228), .B1(G20), .B2(new_n279), .ZN(new_n285));
  NAND2_X1  g0085(.A1(G33), .A2(G283), .ZN(new_n286));
  INV_X1    g0086(.A(G97), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n286), .B(new_n209), .C1(G33), .C2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(KEYINPUT20), .B1(new_n285), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  NAND3_X1  g0090(.A1(new_n285), .A2(KEYINPUT20), .A3(new_n288), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n284), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n276), .A2(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G200), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n294), .B1(new_n263), .B2(new_n275), .ZN(new_n295));
  OAI21_X1  g0095(.A(new_n254), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n263), .A2(new_n275), .ZN(new_n297));
  NAND2_X1  g0097(.A1(new_n297), .A2(G200), .ZN(new_n298));
  NAND4_X1  g0098(.A1(new_n298), .A2(KEYINPUT81), .A3(new_n292), .A4(new_n276), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n296), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(G33), .A2(G116), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n301), .A2(G20), .ZN(new_n302));
  INV_X1    g0102(.A(KEYINPUT23), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n303), .B1(new_n209), .B2(G107), .ZN(new_n304));
  INV_X1    g0104(.A(G107), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n305), .A2(KEYINPUT23), .A3(G20), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n302), .B1(new_n304), .B2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT22), .ZN(new_n308));
  AOI21_X1  g0108(.A(G20), .B1(new_n269), .B2(new_n270), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n308), .B1(new_n309), .B2(G87), .ZN(new_n310));
  OAI211_X1 g0110(.A(new_n209), .B(G87), .C1(new_n264), .C2(new_n265), .ZN(new_n311));
  NOR2_X1   g0111(.A1(new_n311), .A2(KEYINPUT22), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n307), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(KEYINPUT24), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT24), .ZN(new_n315));
  OAI211_X1 g0115(.A(new_n315), .B(new_n307), .C1(new_n310), .C2(new_n312), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n282), .A2(new_n228), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n208), .A2(new_n305), .A3(G13), .A4(G20), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT25), .ZN(new_n321));
  OAI21_X1  g0121(.A(KEYINPUT82), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n320), .A2(new_n321), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(KEYINPUT82), .A3(new_n321), .ZN(new_n325));
  INV_X1    g0125(.A(new_n283), .ZN(new_n326));
  AOI22_X1  g0126(.A1(new_n324), .A2(new_n325), .B1(G107), .B2(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n262), .A2(new_n255), .ZN(new_n328));
  AND2_X1   g0128(.A1(KEYINPUT5), .A2(G41), .ZN(new_n329));
  NOR2_X1   g0129(.A1(KEYINPUT5), .A2(G41), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(new_n257), .ZN(new_n332));
  OAI211_X1 g0132(.A(G264), .B(new_n273), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n328), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g0134(.A(G250), .B(new_n267), .C1(new_n264), .C2(new_n265), .ZN(new_n335));
  OAI211_X1 g0135(.A(G257), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n336));
  INV_X1    g0136(.A(G33), .ZN(new_n337));
  INV_X1    g0137(.A(G294), .ZN(new_n338));
  OAI211_X1 g0138(.A(new_n335), .B(new_n336), .C1(new_n337), .C2(new_n338), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(new_n274), .ZN(new_n340));
  INV_X1    g0140(.A(G190), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n334), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n328), .A2(new_n333), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n343), .B1(new_n274), .B2(new_n339), .ZN(new_n344));
  OAI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(G200), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n319), .A2(new_n327), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n300), .A2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n318), .ZN(new_n348));
  NAND4_X1  g0148(.A1(new_n348), .A2(G116), .A3(new_n277), .A4(new_n281), .ZN(new_n349));
  AND3_X1   g0149(.A1(new_n285), .A2(KEYINPUT20), .A3(new_n288), .ZN(new_n350));
  OAI211_X1 g0150(.A(new_n280), .B(new_n349), .C1(new_n350), .C2(new_n289), .ZN(new_n351));
  NAND4_X1  g0151(.A1(new_n297), .A2(new_n351), .A3(KEYINPUT21), .A4(G169), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n297), .A2(G169), .A3(new_n351), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT21), .ZN(new_n354));
  AND3_X1   g0154(.A1(new_n263), .A2(G179), .A3(new_n275), .ZN(new_n355));
  AOI22_X1  g0155(.A1(new_n353), .A2(new_n354), .B1(new_n355), .B2(new_n351), .ZN(new_n356));
  INV_X1    g0156(.A(new_n327), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n357), .B1(new_n317), .B2(new_n318), .ZN(new_n358));
  INV_X1    g0158(.A(G179), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n334), .A2(new_n340), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n360), .B1(new_n344), .B2(G169), .ZN(new_n361));
  OAI211_X1 g0161(.A(new_n352), .B(new_n356), .C1(new_n358), .C2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n347), .A2(new_n362), .ZN(new_n363));
  XNOR2_X1  g0163(.A(KEYINPUT15), .B(G87), .ZN(new_n364));
  INV_X1    g0164(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n326), .A2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT79), .ZN(new_n367));
  NOR2_X1   g0167(.A1(new_n365), .A2(new_n277), .ZN(new_n368));
  NAND3_X1  g0168(.A1(KEYINPUT19), .A2(G33), .A3(G97), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(new_n209), .ZN(new_n370));
  NOR2_X1   g0170(.A1(G97), .A2(G107), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n371), .A2(new_n217), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n372), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(KEYINPUT78), .ZN(new_n374));
  INV_X1    g0174(.A(KEYINPUT78), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n370), .A2(new_n372), .A3(new_n375), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n209), .B(G68), .C1(new_n264), .C2(new_n265), .ZN(new_n377));
  INV_X1    g0177(.A(KEYINPUT19), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n209), .A2(G33), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n378), .B1(new_n379), .B2(new_n287), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n374), .A2(new_n376), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  AOI211_X1 g0181(.A(new_n367), .B(new_n368), .C1(new_n381), .C2(new_n318), .ZN(new_n382));
  AOI22_X1  g0182(.A1(new_n209), .A2(new_n369), .B1(new_n371), .B2(new_n217), .ZN(new_n383));
  OAI211_X1 g0183(.A(new_n377), .B(new_n380), .C1(new_n383), .C2(new_n375), .ZN(new_n384));
  INV_X1    g0184(.A(new_n376), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n318), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  INV_X1    g0186(.A(new_n368), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT79), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n366), .B1(new_n382), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT80), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n267), .B1(new_n269), .B2(new_n270), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(G244), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n269), .A2(new_n270), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n394), .A2(G238), .A3(new_n267), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n393), .A2(new_n395), .A3(new_n301), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n396), .A2(new_n274), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n257), .A2(new_n218), .ZN(new_n398));
  AOI22_X1  g0198(.A1(new_n398), .A2(new_n273), .B1(G274), .B2(new_n257), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  INV_X1    g0200(.A(G169), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT80), .B(new_n366), .C1(new_n382), .C2(new_n388), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n397), .A2(new_n359), .A3(new_n399), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n391), .A2(new_n402), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n269), .A2(new_n209), .A3(new_n270), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(KEYINPUT7), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n264), .A2(new_n265), .ZN(new_n408));
  INV_X1    g0208(.A(KEYINPUT7), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(new_n409), .A3(new_n209), .ZN(new_n410));
  AND3_X1   g0210(.A1(new_n407), .A2(new_n410), .A3(G107), .ZN(new_n411));
  NOR2_X1   g0211(.A1(G20), .A2(G33), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(G77), .ZN(new_n413));
  XNOR2_X1  g0213(.A(G97), .B(G107), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT6), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n415), .A2(new_n287), .ZN(new_n416));
  AOI22_X1  g0216(.A1(new_n414), .A2(new_n415), .B1(new_n305), .B2(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n413), .B1(new_n417), .B2(new_n209), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n318), .B1(new_n411), .B2(new_n418), .ZN(new_n419));
  OR3_X1    g0219(.A1(new_n277), .A2(KEYINPUT75), .A3(G97), .ZN(new_n420));
  OAI21_X1  g0220(.A(KEYINPUT75), .B1(new_n277), .B2(G97), .ZN(new_n421));
  AOI22_X1  g0221(.A1(G97), .A2(new_n326), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT76), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n419), .A2(new_n422), .A3(new_n423), .ZN(new_n424));
  AND2_X1   g0224(.A1(G97), .A2(G107), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n415), .B1(new_n425), .B2(new_n371), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n305), .A2(KEYINPUT6), .A3(G97), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI22_X1  g0228(.A1(new_n428), .A2(G20), .B1(G77), .B2(new_n412), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n407), .A2(new_n410), .A3(G107), .ZN(new_n430));
  AOI21_X1  g0230(.A(new_n348), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(new_n422), .ZN(new_n432));
  OAI21_X1  g0232(.A(KEYINPUT76), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  AND2_X1   g0234(.A1(new_n260), .A2(G257), .ZN(new_n435));
  NAND4_X1  g0235(.A1(new_n394), .A2(KEYINPUT4), .A3(G244), .A4(new_n267), .ZN(new_n436));
  INV_X1    g0236(.A(new_n286), .ZN(new_n437));
  OAI211_X1 g0237(.A(G244), .B(new_n267), .C1(new_n264), .C2(new_n265), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT4), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n437), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT77), .B1(new_n392), .B2(G250), .ZN(new_n441));
  OAI211_X1 g0241(.A(G250), .B(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT77), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n436), .B(new_n440), .C1(new_n441), .C2(new_n444), .ZN(new_n445));
  AOI21_X1  g0245(.A(new_n435), .B1(new_n445), .B2(new_n274), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n294), .B1(new_n446), .B2(new_n328), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n434), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n446), .A2(G190), .A3(new_n328), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n419), .A2(new_n422), .ZN(new_n450));
  XNOR2_X1  g0250(.A(new_n442), .B(KEYINPUT77), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n438), .A2(new_n439), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n452), .A2(new_n436), .A3(new_n286), .ZN(new_n453));
  OAI21_X1  g0253(.A(new_n274), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(new_n435), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n454), .A2(G179), .A3(new_n328), .A4(new_n455), .ZN(new_n456));
  INV_X1    g0256(.A(new_n328), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n457), .B(new_n435), .C1(new_n445), .C2(new_n274), .ZN(new_n458));
  OAI21_X1  g0258(.A(new_n456), .B1(new_n458), .B2(new_n401), .ZN(new_n459));
  AOI22_X1  g0259(.A1(new_n448), .A2(new_n449), .B1(new_n450), .B2(new_n459), .ZN(new_n460));
  OR2_X1    g0260(.A1(new_n382), .A2(new_n388), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n400), .A2(G200), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n397), .A2(G190), .A3(new_n399), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n326), .A2(G87), .ZN(new_n464));
  NAND4_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n463), .A4(new_n464), .ZN(new_n465));
  NAND4_X1  g0265(.A1(new_n363), .A2(new_n405), .A3(new_n460), .A4(new_n465), .ZN(new_n466));
  AOI22_X1  g0266(.A1(new_n204), .A2(G20), .B1(G150), .B2(new_n412), .ZN(new_n467));
  NAND2_X1  g0267(.A1(KEYINPUT68), .A2(G58), .ZN(new_n468));
  XNOR2_X1  g0268(.A(new_n468), .B(KEYINPUT8), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n470), .B2(new_n379), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(new_n318), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n277), .A2(G50), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n318), .B1(new_n208), .B2(G20), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(G50), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n476), .A2(KEYINPUT9), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT9), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n478), .B1(new_n472), .B2(new_n475), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n480));
  INV_X1    g0280(.A(G274), .ZN(new_n481));
  OR2_X1    g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n273), .A2(new_n480), .ZN(new_n483));
  INV_X1    g0283(.A(G226), .ZN(new_n484));
  OAI21_X1  g0284(.A(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n392), .A2(G223), .B1(new_n408), .B2(G77), .ZN(new_n486));
  INV_X1    g0286(.A(G222), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n394), .A2(new_n267), .ZN(new_n488));
  OAI21_X1  g0288(.A(new_n486), .B1(new_n487), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(new_n485), .B1(new_n489), .B2(new_n274), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI22_X1  g0291(.A1(new_n477), .A2(new_n479), .B1(new_n341), .B2(new_n491), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT10), .ZN(new_n493));
  OAI22_X1  g0293(.A1(new_n490), .A2(new_n294), .B1(KEYINPUT69), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n493), .A2(KEYINPUT69), .ZN(new_n495));
  INV_X1    g0295(.A(new_n495), .ZN(new_n496));
  OR3_X1    g0296(.A1(new_n492), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n490), .A2(new_n294), .ZN(new_n498));
  OAI211_X1 g0298(.A(KEYINPUT69), .B(new_n493), .C1(new_n492), .C2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NOR2_X1   g0300(.A1(new_n491), .A2(G179), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n476), .B1(new_n490), .B2(G169), .ZN(new_n502));
  OR2_X1    g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n278), .A2(new_n203), .ZN(new_n505));
  OAI21_X1  g0305(.A(KEYINPUT12), .B1(new_n505), .B2(KEYINPUT71), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(KEYINPUT71), .ZN(new_n507));
  XNOR2_X1  g0307(.A(new_n506), .B(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n209), .A2(new_n337), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n509), .A2(new_n201), .B1(new_n209), .B2(G68), .ZN(new_n510));
  INV_X1    g0310(.A(G77), .ZN(new_n511));
  NOR2_X1   g0311(.A1(new_n379), .A2(new_n511), .ZN(new_n512));
  OAI21_X1  g0312(.A(new_n318), .B1(new_n510), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n513), .B(KEYINPUT11), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n474), .A2(G68), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n508), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n239), .A2(G1698), .ZN(new_n517));
  OAI221_X1 g0317(.A(new_n517), .B1(G226), .B2(G1698), .C1(new_n264), .C2(new_n265), .ZN(new_n518));
  NAND2_X1  g0318(.A1(G33), .A2(G97), .ZN(new_n519));
  AOI21_X1  g0319(.A(new_n273), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n482), .B1(new_n483), .B2(new_n216), .ZN(new_n521));
  OAI21_X1  g0321(.A(KEYINPUT13), .B1(new_n520), .B2(new_n521), .ZN(new_n522));
  NOR2_X1   g0322(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT13), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n341), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n516), .B1(new_n522), .B2(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n523), .A2(new_n524), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT70), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n527), .A2(new_n528), .A3(new_n522), .ZN(new_n529));
  OAI211_X1 g0329(.A(KEYINPUT70), .B(KEYINPUT13), .C1(new_n520), .C2(new_n521), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(G200), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g0332(.A1(new_n392), .A2(G238), .B1(new_n408), .B2(G107), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n533), .B1(new_n239), .B2(new_n488), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(new_n274), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n480), .A2(new_n481), .ZN(new_n536));
  AND2_X1   g0336(.A1(new_n273), .A2(new_n480), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n536), .B1(new_n537), .B2(G244), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n535), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(new_n401), .ZN(new_n540));
  INV_X1    g0340(.A(new_n538), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n534), .B2(new_n274), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n359), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n277), .A2(G77), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n474), .B2(G77), .ZN(new_n545));
  XOR2_X1   g0345(.A(KEYINPUT8), .B(G58), .Z(new_n546));
  AOI22_X1  g0346(.A1(new_n546), .A2(new_n412), .B1(G20), .B2(G77), .ZN(new_n547));
  OR2_X1    g0347(.A1(new_n364), .A2(new_n379), .ZN(new_n548));
  AND2_X1   g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n545), .B1(new_n549), .B2(new_n348), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n540), .A2(new_n543), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n550), .B1(G190), .B2(new_n542), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n552), .B1(new_n294), .B2(new_n542), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n532), .A2(new_n551), .A3(new_n553), .ZN(new_n554));
  NOR3_X1   g0354(.A1(new_n500), .A2(new_n504), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n529), .A2(G169), .A3(new_n530), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT14), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT14), .A4(G169), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n527), .A2(G179), .A3(new_n522), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(new_n516), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT16), .ZN(new_n564));
  NAND2_X1  g0364(.A1(G58), .A2(G68), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n225), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n566), .A2(G20), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT72), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n412), .A2(G159), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  AOI21_X1  g0370(.A(new_n209), .B1(new_n225), .B2(new_n565), .ZN(new_n571));
  INV_X1    g0371(.A(new_n569), .ZN(new_n572));
  OAI21_X1  g0372(.A(KEYINPUT72), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND2_X1   g0373(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n407), .A2(new_n410), .A3(G68), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n564), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n575), .A2(new_n564), .A3(new_n570), .A4(new_n573), .ZN(new_n577));
  INV_X1    g0377(.A(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n318), .B1(new_n576), .B2(new_n578), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n536), .B1(new_n537), .B2(G232), .ZN(new_n580));
  NOR2_X1   g0380(.A1(G223), .A2(G1698), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n581), .B1(new_n484), .B2(G1698), .ZN(new_n582));
  AOI22_X1  g0382(.A1(new_n582), .A2(new_n394), .B1(G33), .B2(G87), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n580), .B1(new_n273), .B2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n294), .ZN(new_n585));
  XNOR2_X1  g0385(.A(new_n580), .B(KEYINPUT73), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n341), .B1(new_n583), .B2(new_n273), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n585), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n470), .B1(new_n208), .B2(G20), .ZN(new_n589));
  NOR2_X1   g0389(.A1(new_n278), .A2(new_n318), .ZN(new_n590));
  AOI22_X1  g0390(.A1(new_n589), .A2(new_n590), .B1(new_n278), .B2(new_n470), .ZN(new_n591));
  NAND3_X1  g0391(.A1(new_n579), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT17), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n482), .B1(new_n483), .B2(new_n239), .ZN(new_n595));
  XNOR2_X1  g0395(.A(new_n595), .B(KEYINPUT73), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n583), .A2(new_n273), .ZN(new_n597));
  NOR2_X1   g0397(.A1(new_n597), .A2(G179), .ZN(new_n598));
  AOI22_X1  g0398(.A1(new_n596), .A2(new_n598), .B1(new_n401), .B2(new_n584), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n570), .A2(new_n573), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n407), .A2(new_n410), .A3(G68), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT16), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n348), .B1(new_n602), .B2(new_n577), .ZN(new_n603));
  INV_X1    g0403(.A(new_n591), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n599), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n605), .A2(KEYINPUT18), .ZN(new_n606));
  INV_X1    g0406(.A(KEYINPUT18), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n599), .B(new_n607), .C1(new_n603), .C2(new_n604), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n579), .A2(new_n588), .A3(KEYINPUT17), .A4(new_n591), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n594), .A2(new_n606), .A3(new_n608), .A4(new_n609), .ZN(new_n610));
  INV_X1    g0410(.A(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n555), .A2(new_n563), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT74), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g0414(.A1(new_n555), .A2(KEYINPUT74), .A3(new_n563), .A4(new_n611), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n466), .B1(new_n614), .B2(new_n615), .ZN(G372));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n615), .ZN(new_n617));
  NAND4_X1  g0417(.A1(new_n405), .A2(new_n465), .A3(new_n450), .A4(new_n459), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n618), .A2(KEYINPUT26), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n353), .A2(new_n354), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n355), .A2(new_n351), .ZN(new_n621));
  AND3_X1   g0421(.A1(new_n620), .A2(new_n352), .A3(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n334), .A2(new_n340), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n623), .A2(new_n401), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n348), .B1(new_n314), .B2(new_n316), .ZN(new_n625));
  OAI211_X1 g0425(.A(new_n360), .B(new_n624), .C1(new_n625), .C2(new_n357), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n622), .A2(new_n626), .B1(new_n358), .B2(new_n345), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n396), .A2(KEYINPUT83), .A3(new_n274), .ZN(new_n628));
  AOI21_X1  g0428(.A(KEYINPUT83), .B1(new_n396), .B2(new_n274), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n399), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n630), .A2(new_n401), .ZN(new_n631));
  NAND4_X1  g0431(.A1(new_n391), .A2(new_n403), .A3(new_n404), .A4(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n630), .A2(G200), .ZN(new_n633));
  NAND4_X1  g0433(.A1(new_n461), .A2(new_n633), .A3(new_n463), .A4(new_n464), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n460), .A2(new_n627), .A3(new_n632), .A4(new_n634), .ZN(new_n635));
  AND2_X1   g0435(.A1(new_n459), .A2(new_n434), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT26), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n632), .A2(new_n634), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n619), .A2(new_n635), .A3(new_n632), .A4(new_n638), .ZN(new_n639));
  AND2_X1   g0439(.A1(new_n617), .A2(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n606), .A2(new_n608), .ZN(new_n641));
  INV_X1    g0441(.A(new_n561), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n642), .B1(new_n558), .B2(new_n559), .ZN(new_n643));
  INV_X1    g0443(.A(new_n516), .ZN(new_n644));
  INV_X1    g0444(.A(new_n532), .ZN(new_n645));
  OAI22_X1  g0445(.A1(new_n643), .A2(new_n644), .B1(new_n645), .B2(new_n551), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT84), .ZN(new_n647));
  OR2_X1    g0447(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n594), .A2(new_n609), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n649), .B1(new_n646), .B2(new_n647), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n641), .B1(new_n648), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n503), .B1(new_n651), .B2(new_n500), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n640), .A2(new_n652), .ZN(G369));
  NAND3_X1  g0453(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n654));
  OR2_X1    g0454(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(KEYINPUT27), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n655), .A2(G213), .A3(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(G343), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n659), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n622), .B(new_n300), .C1(new_n292), .C2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n620), .A2(new_n352), .A3(new_n621), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(new_n351), .A3(new_n659), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  INV_X1    g0465(.A(G330), .ZN(new_n666));
  NOR2_X1   g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n346), .B1(new_n358), .B2(new_n660), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n668), .A2(new_n626), .ZN(new_n669));
  INV_X1    g0469(.A(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n626), .A2(new_n659), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n622), .A2(new_n659), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n671), .B1(new_n669), .B2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(G399));
  INV_X1    g0476(.A(new_n212), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n677), .A2(G41), .ZN(new_n678));
  INV_X1    g0478(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n372), .A2(G116), .ZN(new_n680));
  NAND3_X1  g0480(.A1(new_n679), .A2(G1), .A3(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n226), .B2(new_n679), .ZN(new_n682));
  XNOR2_X1  g0482(.A(new_n682), .B(KEYINPUT28), .ZN(new_n683));
  OAI211_X1 g0483(.A(new_n635), .B(new_n632), .C1(KEYINPUT26), .C2(new_n618), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n632), .A2(new_n634), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n637), .B1(new_n685), .B2(new_n636), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n660), .B1(new_n684), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n687), .A2(KEYINPUT29), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n639), .A2(new_n689), .A3(new_n660), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT85), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n355), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g0493(.A(KEYINPUT85), .B1(new_n297), .B2(new_n359), .ZN(new_n694));
  AND2_X1   g0494(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n400), .A2(new_n623), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n695), .A2(KEYINPUT30), .A3(new_n446), .A4(new_n696), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n696), .A2(new_n693), .A3(new_n446), .A4(new_n694), .ZN(new_n698));
  INV_X1    g0498(.A(KEYINPUT30), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n623), .A2(new_n359), .A3(new_n297), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n454), .A2(new_n328), .A3(new_n455), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n630), .A3(new_n702), .ZN(new_n703));
  INV_X1    g0503(.A(KEYINPUT86), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND4_X1  g0505(.A1(new_n701), .A2(new_n630), .A3(new_n702), .A4(KEYINPUT86), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n697), .A2(new_n700), .A3(new_n705), .A4(new_n706), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n707), .A2(new_n659), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n405), .A2(new_n465), .ZN(new_n709));
  NAND4_X1  g0509(.A1(new_n622), .A2(new_n626), .A3(new_n300), .A4(new_n346), .ZN(new_n710));
  INV_X1    g0510(.A(new_n456), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n401), .B1(new_n446), .B2(new_n328), .ZN(new_n712));
  OAI21_X1  g0512(.A(new_n450), .B1(new_n711), .B2(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n702), .A2(G200), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(new_n449), .A3(new_n433), .A4(new_n424), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n710), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n709), .A2(new_n717), .A3(new_n660), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n708), .B1(new_n718), .B2(KEYINPUT31), .ZN(new_n719));
  NAND3_X1  g0519(.A1(new_n697), .A2(new_n700), .A3(new_n703), .ZN(new_n720));
  AND3_X1   g0520(.A1(new_n720), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n721));
  OAI21_X1  g0521(.A(G330), .B1(new_n719), .B2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OR3_X1    g0523(.A1(new_n691), .A2(new_n723), .A3(KEYINPUT87), .ZN(new_n724));
  OAI21_X1  g0524(.A(KEYINPUT87), .B1(new_n691), .B2(new_n723), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n683), .B1(new_n726), .B2(G1), .ZN(G364));
  XNOR2_X1  g0527(.A(new_n667), .B(KEYINPUT88), .ZN(new_n728));
  INV_X1    g0528(.A(G13), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n729), .A2(G20), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT89), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n731), .A2(G45), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G1), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n678), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  OAI211_X1 g0535(.A(new_n728), .B(new_n735), .C1(G330), .C2(new_n664), .ZN(new_n736));
  NOR2_X1   g0536(.A1(G13), .A2(G33), .ZN(new_n737));
  XNOR2_X1  g0537(.A(new_n737), .B(KEYINPUT90), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(new_n209), .ZN(new_n740));
  XOR2_X1   g0540(.A(new_n740), .B(KEYINPUT91), .Z(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n228), .B1(G20), .B2(new_n401), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n677), .A2(new_n408), .ZN(new_n745));
  AOI22_X1  g0545(.A1(new_n745), .A2(G355), .B1(new_n279), .B2(new_n677), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n677), .A2(new_n394), .ZN(new_n747));
  OAI21_X1  g0547(.A(new_n747), .B1(new_n227), .B2(G45), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n248), .A2(new_n256), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n746), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n743), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n209), .A2(new_n341), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n359), .A2(G200), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n209), .A2(G190), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n754), .A2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  AOI22_X1  g0559(.A1(G58), .A2(new_n756), .B1(new_n759), .B2(G77), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n359), .A2(new_n294), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n753), .A2(new_n761), .ZN(new_n762));
  OAI21_X1  g0562(.A(new_n760), .B1(new_n201), .B2(new_n762), .ZN(new_n763));
  XOR2_X1   g0563(.A(new_n763), .B(KEYINPUT92), .Z(new_n764));
  NOR2_X1   g0564(.A1(new_n294), .A2(G179), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n757), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g0566(.A1(new_n753), .A2(new_n765), .ZN(new_n767));
  OAI221_X1 g0567(.A(new_n394), .B1(new_n766), .B2(new_n305), .C1(new_n217), .C2(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(G179), .A2(G200), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n757), .A2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G159), .ZN(new_n771));
  OR3_X1    g0571(.A1(new_n770), .A2(KEYINPUT32), .A3(new_n771), .ZN(new_n772));
  OAI21_X1  g0572(.A(KEYINPUT32), .B1(new_n770), .B2(new_n771), .ZN(new_n773));
  AOI21_X1  g0573(.A(new_n209), .B1(new_n769), .B2(G190), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G97), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n772), .A2(new_n773), .A3(new_n776), .ZN(new_n777));
  AND3_X1   g0577(.A1(new_n761), .A2(KEYINPUT93), .A3(new_n757), .ZN(new_n778));
  AOI21_X1  g0578(.A(KEYINPUT93), .B1(new_n761), .B2(new_n757), .ZN(new_n779));
  NOR2_X1   g0579(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n780), .ZN(new_n781));
  AOI211_X1 g0581(.A(new_n768), .B(new_n777), .C1(G68), .C2(new_n781), .ZN(new_n782));
  INV_X1    g0582(.A(new_n766), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G322), .A2(new_n756), .B1(new_n783), .B2(G283), .ZN(new_n784));
  INV_X1    g0584(.A(new_n762), .ZN(new_n785));
  AOI22_X1  g0585(.A1(G326), .A2(new_n785), .B1(new_n759), .B2(G311), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n775), .A2(G294), .ZN(new_n787));
  INV_X1    g0587(.A(new_n770), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n394), .B1(new_n788), .B2(G329), .ZN(new_n789));
  AND4_X1   g0589(.A1(new_n784), .A2(new_n786), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n767), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n791), .A2(KEYINPUT94), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n791), .A2(KEYINPUT94), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  XNOR2_X1  g0595(.A(KEYINPUT33), .B(G317), .ZN(new_n796));
  AOI22_X1  g0596(.A1(new_n795), .A2(G303), .B1(new_n781), .B2(new_n796), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n764), .A2(new_n782), .B1(new_n790), .B2(new_n797), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n751), .B1(new_n752), .B2(new_n798), .C1(new_n664), .C2(new_n741), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n736), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NOR2_X1   g0601(.A1(new_n539), .A2(G179), .ZN(new_n802));
  OAI21_X1  g0602(.A(new_n550), .B1(new_n542), .B2(G169), .ZN(new_n803));
  OAI21_X1  g0603(.A(KEYINPUT96), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  INV_X1    g0604(.A(KEYINPUT96), .ZN(new_n805));
  NAND4_X1  g0605(.A1(new_n540), .A2(new_n805), .A3(new_n543), .A4(new_n550), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n550), .A2(new_n659), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n804), .A2(new_n553), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(KEYINPUT97), .ZN(new_n809));
  OR2_X1    g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n812), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n639), .A2(new_n813), .A3(new_n660), .ZN(new_n814));
  AND2_X1   g0614(.A1(new_n639), .A2(new_n660), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n551), .A2(new_n660), .ZN(new_n816));
  INV_X1    g0616(.A(new_n816), .ZN(new_n817));
  NAND2_X1  g0617(.A1(new_n812), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n814), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n734), .B1(new_n819), .B2(new_n722), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n820), .B1(new_n722), .B2(new_n819), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n743), .A2(new_n737), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n735), .B1(new_n511), .B2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n794), .A2(new_n201), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n408), .B1(new_n783), .B2(G68), .ZN(new_n825));
  INV_X1    g0625(.A(G132), .ZN(new_n826));
  OAI221_X1 g0626(.A(new_n825), .B1(new_n202), .B2(new_n774), .C1(new_n826), .C2(new_n770), .ZN(new_n827));
  AOI22_X1  g0627(.A1(G137), .A2(new_n785), .B1(new_n756), .B2(G143), .ZN(new_n828));
  INV_X1    g0628(.A(G150), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n828), .B1(new_n771), .B2(new_n758), .C1(new_n829), .C2(new_n780), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT95), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT34), .ZN(new_n832));
  AOI211_X1 g0632(.A(new_n824), .B(new_n827), .C1(new_n831), .C2(new_n832), .ZN(new_n833));
  OR2_X1    g0633(.A1(new_n831), .A2(new_n832), .ZN(new_n834));
  AOI22_X1  g0634(.A1(G303), .A2(new_n785), .B1(new_n759), .B2(G116), .ZN(new_n835));
  AOI22_X1  g0635(.A1(G294), .A2(new_n756), .B1(new_n788), .B2(G311), .ZN(new_n836));
  NOR2_X1   g0636(.A1(new_n766), .A2(new_n217), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n837), .A2(new_n394), .ZN(new_n838));
  AND4_X1   g0638(.A1(new_n776), .A2(new_n835), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI22_X1  g0639(.A1(new_n795), .A2(G107), .B1(G283), .B2(new_n781), .ZN(new_n840));
  AOI22_X1  g0640(.A1(new_n833), .A2(new_n834), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n823), .B1(new_n752), .B2(new_n841), .C1(new_n818), .C2(new_n738), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n821), .A2(new_n842), .ZN(G384));
  NOR2_X1   g0643(.A1(new_n731), .A2(new_n208), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n562), .A2(KEYINPUT100), .A3(new_n516), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n516), .A2(new_n659), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g0647(.A1(new_n645), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT100), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n849), .B1(new_n643), .B2(new_n644), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n845), .A2(new_n848), .A3(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n562), .A2(new_n847), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n818), .ZN(new_n854));
  AND3_X1   g0654(.A1(new_n707), .A2(KEYINPUT31), .A3(new_n659), .ZN(new_n855));
  OAI21_X1  g0655(.A(KEYINPUT102), .B1(new_n719), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT102), .ZN(new_n857));
  INV_X1    g0657(.A(new_n855), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT31), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n361), .B1(new_n319), .B2(new_n327), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n860), .A2(new_n662), .ZN(new_n861));
  AOI22_X1  g0661(.A1(new_n358), .A2(new_n345), .B1(new_n296), .B2(new_n299), .ZN(new_n862));
  NAND4_X1  g0662(.A1(new_n861), .A2(new_n862), .A3(new_n713), .A4(new_n715), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n405), .A2(new_n465), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(new_n859), .B1(new_n865), .B2(new_n660), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n857), .B(new_n858), .C1(new_n866), .C2(new_n708), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n854), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n657), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n603), .B2(new_n604), .ZN(new_n870));
  INV_X1    g0670(.A(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n610), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n592), .A2(new_n605), .A3(new_n870), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n873), .A2(KEYINPUT37), .ZN(new_n874));
  XNOR2_X1  g0674(.A(KEYINPUT101), .B(KEYINPUT37), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n592), .A2(new_n605), .A3(new_n870), .A4(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n872), .A2(new_n877), .A3(KEYINPUT38), .ZN(new_n881));
  AOI21_X1  g0681(.A(KEYINPUT40), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n868), .A2(new_n882), .ZN(new_n883));
  AND3_X1   g0683(.A1(new_n872), .A2(KEYINPUT38), .A3(new_n877), .ZN(new_n884));
  INV_X1    g0684(.A(new_n875), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n873), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n886), .A2(new_n876), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n872), .B2(new_n887), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n884), .A2(new_n888), .ZN(new_n889));
  AOI211_X1 g0689(.A(new_n889), .B(new_n854), .C1(new_n856), .C2(new_n867), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT40), .ZN(new_n891));
  OAI21_X1  g0691(.A(new_n883), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n856), .A2(new_n867), .B1(new_n614), .B2(new_n615), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n666), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n892), .ZN(new_n895));
  XOR2_X1   g0695(.A(new_n895), .B(KEYINPUT103), .Z(new_n896));
  INV_X1    g0696(.A(new_n896), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n641), .A2(new_n657), .ZN(new_n898));
  NAND3_X1  g0698(.A1(new_n880), .A2(KEYINPUT39), .A3(new_n881), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n899), .B1(new_n889), .B2(KEYINPUT39), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n659), .B1(new_n845), .B2(new_n850), .ZN(new_n901));
  INV_X1    g0701(.A(new_n901), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n898), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n880), .A2(new_n881), .ZN(new_n904));
  INV_X1    g0704(.A(new_n853), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n804), .A2(new_n806), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n906), .A2(new_n660), .ZN(new_n907));
  AOI21_X1  g0707(.A(new_n905), .B1(new_n814), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n903), .B1(new_n904), .B2(new_n908), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n652), .B1(new_n691), .B2(new_n617), .ZN(new_n910));
  XNOR2_X1  g0710(.A(new_n909), .B(new_n910), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n844), .B1(new_n897), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n912), .B1(new_n897), .B2(new_n911), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n279), .B(new_n230), .C1(new_n428), .C2(KEYINPUT35), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(KEYINPUT35), .B2(new_n428), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n915), .B(KEYINPUT36), .ZN(new_n916));
  XNOR2_X1  g0716(.A(new_n244), .B(KEYINPUT99), .ZN(new_n917));
  AOI211_X1 g0717(.A(new_n511), .B(new_n226), .C1(G58), .C2(G68), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT98), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n917), .B1(new_n918), .B2(new_n919), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n920), .B1(new_n919), .B2(new_n918), .ZN(new_n921));
  NAND3_X1  g0721(.A1(new_n921), .A2(G1), .A3(new_n729), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n913), .A2(new_n916), .A3(new_n922), .ZN(G367));
  OAI21_X1  g0723(.A(new_n744), .B1(new_n212), .B2(new_n364), .ZN(new_n924));
  AND2_X1   g0724(.A1(new_n237), .A2(new_n747), .ZN(new_n925));
  OAI21_X1  g0725(.A(new_n734), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(G143), .ZN(new_n927));
  OAI22_X1  g0727(.A1(new_n762), .A2(new_n927), .B1(new_n755), .B2(new_n829), .ZN(new_n928));
  AOI211_X1 g0728(.A(new_n408), .B(new_n928), .C1(G58), .C2(new_n791), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n775), .A2(G68), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n781), .A2(G159), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n201), .A2(new_n758), .B1(new_n766), .B2(new_n511), .ZN(new_n932));
  AOI21_X1  g0732(.A(new_n932), .B1(G137), .B2(new_n788), .ZN(new_n933));
  NAND4_X1  g0733(.A1(new_n929), .A2(new_n930), .A3(new_n931), .A4(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n766), .A2(new_n287), .ZN(new_n935));
  AOI211_X1 g0735(.A(new_n394), .B(new_n935), .C1(G317), .C2(new_n788), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n936), .B(KEYINPUT106), .Z(new_n937));
  INV_X1    g0737(.A(G303), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n755), .A2(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(G311), .ZN(new_n940));
  INV_X1    g0740(.A(G283), .ZN(new_n941));
  OAI22_X1  g0741(.A1(new_n762), .A2(new_n940), .B1(new_n758), .B2(new_n941), .ZN(new_n942));
  AOI211_X1 g0742(.A(new_n939), .B(new_n942), .C1(G107), .C2(new_n775), .ZN(new_n943));
  OAI211_X1 g0743(.A(new_n937), .B(new_n943), .C1(new_n338), .C2(new_n780), .ZN(new_n944));
  NOR3_X1   g0744(.A1(new_n767), .A2(KEYINPUT46), .A3(new_n279), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n795), .A2(G116), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n945), .B1(new_n946), .B2(KEYINPUT46), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n934), .B1(new_n944), .B2(new_n947), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n948), .B(KEYINPUT47), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n926), .B1(new_n949), .B2(new_n743), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n461), .A2(new_n464), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n951), .A2(new_n659), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n685), .A2(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n632), .A2(new_n952), .ZN(new_n954));
  NAND3_X1  g0754(.A1(new_n953), .A2(new_n742), .A3(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n950), .A2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n434), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n460), .B1(new_n957), .B2(new_n660), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n636), .A2(new_n659), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  OR3_X1    g0760(.A1(new_n960), .A2(KEYINPUT104), .A3(new_n675), .ZN(new_n961));
  OAI21_X1  g0761(.A(KEYINPUT104), .B1(new_n960), .B2(new_n675), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n961), .A2(KEYINPUT44), .A3(new_n962), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n960), .A2(new_n675), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT45), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n967), .B(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n965), .A2(new_n966), .A3(new_n969), .ZN(new_n970));
  INV_X1    g0770(.A(new_n673), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n965), .A2(new_n673), .A3(new_n966), .A4(new_n969), .ZN(new_n973));
  AND2_X1   g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n672), .B(new_n674), .ZN(new_n975));
  AND2_X1   g0775(.A1(new_n728), .A2(new_n975), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(new_n666), .A3(new_n665), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND3_X1  g0778(.A1(new_n974), .A2(new_n726), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(KEYINPUT105), .ZN(new_n980));
  AOI211_X1 g0780(.A(new_n976), .B(new_n977), .C1(new_n724), .C2(new_n725), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT105), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n981), .A2(new_n982), .A3(new_n974), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n980), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n726), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n678), .B(KEYINPUT41), .Z(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n733), .B1(new_n985), .B2(new_n987), .ZN(new_n988));
  NAND3_X1  g0788(.A1(new_n960), .A2(new_n672), .A3(new_n674), .ZN(new_n989));
  XOR2_X1   g0789(.A(new_n989), .B(KEYINPUT42), .Z(new_n990));
  INV_X1    g0790(.A(new_n960), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n713), .B1(new_n991), .B2(new_n626), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n660), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n953), .A2(new_n954), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n990), .A2(new_n993), .B1(KEYINPUT43), .B2(new_n994), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n994), .A2(KEYINPUT43), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n995), .B(new_n996), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n673), .A2(new_n991), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n997), .B(new_n998), .Z(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n956), .B1(new_n988), .B2(new_n1000), .ZN(G387));
  OAI21_X1  g0801(.A(new_n742), .B1(new_n670), .B2(new_n671), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n745), .ZN(new_n1003));
  OAI22_X1  g0803(.A1(new_n1003), .A2(new_n680), .B1(G107), .B2(new_n212), .ZN(new_n1004));
  AOI211_X1 g0804(.A(new_n677), .B(new_n394), .C1(new_n242), .C2(G45), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n546), .A2(new_n201), .ZN(new_n1006));
  XOR2_X1   g0806(.A(new_n1006), .B(KEYINPUT50), .Z(new_n1007));
  OAI211_X1 g0807(.A(new_n680), .B(new_n256), .C1(new_n203), .C2(new_n511), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT107), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  NAND3_X1  g0811(.A1(new_n1007), .A2(new_n1010), .A3(new_n1011), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1004), .B1(new_n1005), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(new_n744), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n734), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  AOI22_X1  g0815(.A1(G50), .A2(new_n756), .B1(new_n759), .B2(G68), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n771), .B2(new_n762), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n774), .A2(new_n364), .ZN(new_n1018));
  NOR4_X1   g0818(.A1(new_n1017), .A2(new_n408), .A3(new_n935), .A4(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n767), .A2(new_n511), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G150), .B2(new_n788), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1021), .B(KEYINPUT108), .Z(new_n1022));
  OAI211_X1 g0822(.A(new_n1019), .B(new_n1022), .C1(new_n470), .C2(new_n780), .ZN(new_n1023));
  AOI21_X1  g0823(.A(new_n394), .B1(new_n788), .B2(G326), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n767), .A2(new_n338), .B1(new_n774), .B2(new_n941), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n785), .A2(G322), .ZN(new_n1026));
  INV_X1    g0826(.A(G317), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n1026), .B1(new_n938), .B2(new_n758), .C1(new_n1027), .C2(new_n755), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G311), .B2(new_n781), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1025), .B1(new_n1029), .B2(KEYINPUT48), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT48), .B2(new_n1029), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT49), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1024), .B1(new_n279), .B2(new_n766), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  AND2_X1   g0833(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n1023), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n743), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(new_n978), .A2(new_n733), .B1(new_n1002), .B2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n981), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1038), .A2(new_n678), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n726), .A2(new_n978), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1037), .B1(new_n1039), .B2(new_n1040), .ZN(G393));
  NAND2_X1  g0841(.A1(new_n974), .A2(new_n733), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n408), .B1(new_n766), .B2(new_n305), .ZN(new_n1043));
  AOI22_X1  g0843(.A1(G283), .A2(new_n791), .B1(new_n788), .B2(G322), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n338), .B2(new_n758), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1043), .B(new_n1045), .C1(G116), .C2(new_n775), .ZN(new_n1046));
  OAI22_X1  g0846(.A1(new_n762), .A2(new_n1027), .B1(new_n755), .B2(new_n940), .ZN(new_n1047));
  XNOR2_X1  g0847(.A(new_n1047), .B(KEYINPUT52), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1046), .B(new_n1048), .C1(new_n938), .C2(new_n780), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT110), .Z(new_n1050));
  AOI22_X1  g0850(.A1(new_n781), .A2(G50), .B1(new_n546), .B2(new_n759), .ZN(new_n1051));
  OR2_X1    g0851(.A1(new_n1051), .A2(KEYINPUT109), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1051), .A2(KEYINPUT109), .ZN(new_n1053));
  OAI22_X1  g0853(.A1(new_n762), .A2(new_n829), .B1(new_n755), .B2(new_n771), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT51), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n767), .A2(new_n203), .B1(new_n770), .B2(new_n927), .ZN(new_n1056));
  NOR2_X1   g0856(.A1(new_n774), .A2(new_n511), .ZN(new_n1057));
  NOR4_X1   g0857(.A1(new_n1056), .A2(new_n837), .A3(new_n1057), .A4(new_n408), .ZN(new_n1058));
  NAND4_X1  g0858(.A1(new_n1052), .A2(new_n1053), .A3(new_n1055), .A4(new_n1058), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n752), .B1(new_n1050), .B2(new_n1059), .ZN(new_n1060));
  AOI22_X1  g0860(.A1(new_n747), .A2(new_n252), .B1(G97), .B2(new_n677), .ZN(new_n1061));
  AOI211_X1 g0861(.A(new_n735), .B(new_n1060), .C1(new_n744), .C2(new_n1061), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1062), .B1(new_n741), .B2(new_n960), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1042), .A2(new_n1063), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n974), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n679), .B1(new_n1038), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1064), .B1(new_n984), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(G390));
  INV_X1    g0868(.A(new_n854), .ZN(new_n1069));
  OAI21_X1  g0869(.A(KEYINPUT31), .B1(new_n466), .B2(new_n659), .ZN(new_n1070));
  INV_X1    g0870(.A(new_n708), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n857), .B1(new_n1072), .B2(new_n858), .ZN(new_n1073));
  AOI211_X1 g0873(.A(KEYINPUT102), .B(new_n855), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1074));
  OAI211_X1 g0874(.A(G330), .B(new_n1069), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n813), .B(new_n660), .C1(new_n684), .C2(new_n686), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n907), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1077), .A2(new_n853), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n889), .A2(new_n901), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n900), .B1(new_n908), .B2(new_n901), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1075), .B1(new_n1080), .B2(new_n1081), .ZN(new_n1082));
  AND2_X1   g0882(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n723), .A2(new_n1069), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1082), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n900), .A2(new_n739), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n822), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n734), .B1(new_n469), .B2(new_n1087), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n767), .A2(new_n829), .ZN(new_n1089));
  XNOR2_X1  g0889(.A(new_n1089), .B(KEYINPUT112), .ZN(new_n1090));
  OR2_X1    g0890(.A1(new_n1090), .A2(KEYINPUT53), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(KEYINPUT53), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n775), .A2(G159), .ZN(new_n1093));
  INV_X1    g0893(.A(G128), .ZN(new_n1094));
  XNOR2_X1  g0894(.A(KEYINPUT54), .B(G143), .ZN(new_n1095));
  OAI22_X1  g0895(.A1(new_n762), .A2(new_n1094), .B1(new_n758), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g0896(.A(G125), .ZN(new_n1097));
  OAI22_X1  g0897(.A1(new_n755), .A2(new_n826), .B1(new_n770), .B2(new_n1097), .ZN(new_n1098));
  NOR2_X1   g0898(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  NAND4_X1  g0899(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .A4(new_n1099), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n394), .B1(new_n766), .B2(new_n201), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1101), .A2(KEYINPUT111), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1101), .A2(KEYINPUT111), .ZN(new_n1103));
  INV_X1    g0903(.A(G137), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1102), .B(new_n1103), .C1(new_n1104), .C2(new_n780), .ZN(new_n1105));
  AOI211_X1 g0905(.A(new_n394), .B(new_n1057), .C1(G68), .C2(new_n783), .ZN(new_n1106));
  AOI22_X1  g0906(.A1(G283), .A2(new_n785), .B1(new_n759), .B2(G97), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(G116), .A2(new_n756), .B1(new_n788), .B2(G294), .ZN(new_n1108));
  NAND3_X1  g0908(.A1(new_n1106), .A2(new_n1107), .A3(new_n1108), .ZN(new_n1109));
  OAI22_X1  g0909(.A1(new_n794), .A2(new_n217), .B1(new_n305), .B2(new_n780), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n1100), .A2(new_n1105), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n1088), .B1(new_n1111), .B2(new_n743), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(new_n1085), .A2(new_n733), .B1(new_n1086), .B2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n666), .B1(new_n856), .B2(new_n867), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1114), .A2(new_n617), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n910), .A2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g0916(.A(G330), .B(new_n818), .C1(new_n719), .C2(new_n721), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1117), .A2(new_n905), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1075), .A2(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n814), .A2(new_n907), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n907), .B(new_n1076), .C1(new_n722), .C2(new_n854), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n818), .ZN(new_n1124));
  AOI211_X1 g0924(.A(new_n666), .B(new_n1124), .C1(new_n856), .C2(new_n867), .ZN(new_n1125));
  OAI21_X1  g0925(.A(new_n1123), .B1(new_n1125), .B2(new_n853), .ZN(new_n1126));
  AOI21_X1  g0926(.A(new_n1116), .B1(new_n1121), .B2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n678), .B1(new_n1085), .B2(new_n1127), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n1114), .A2(new_n1069), .B1(new_n905), .B2(new_n1117), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1120), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n853), .B1(new_n1114), .B2(new_n818), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n1129), .A2(new_n1130), .B1(new_n1131), .B2(new_n1122), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1116), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1080), .A2(new_n1081), .A3(new_n1084), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n1083), .B2(new_n1075), .ZN(new_n1136));
  NOR2_X1   g0936(.A1(new_n1134), .A2(new_n1136), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1113), .B1(new_n1128), .B2(new_n1137), .ZN(G378));
  INV_X1    g0938(.A(new_n733), .ZN(new_n1139));
  NOR2_X1   g0939(.A1(new_n500), .A2(new_n504), .ZN(new_n1140));
  XOR2_X1   g0940(.A(KEYINPUT117), .B(KEYINPUT56), .Z(new_n1141));
  XNOR2_X1  g0941(.A(new_n1141), .B(KEYINPUT118), .ZN(new_n1142));
  XNOR2_X1  g0942(.A(new_n1140), .B(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n476), .A2(new_n869), .ZN(new_n1144));
  XOR2_X1   g0944(.A(new_n1144), .B(KEYINPUT55), .Z(new_n1145));
  XNOR2_X1  g0945(.A(new_n1145), .B(KEYINPUT116), .ZN(new_n1146));
  XNOR2_X1  g0946(.A(new_n1143), .B(new_n1146), .ZN(new_n1147));
  NOR2_X1   g0947(.A1(new_n1147), .A2(KEYINPUT120), .ZN(new_n1148));
  INV_X1    g0948(.A(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n908), .A2(new_n904), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1150), .B(new_n898), .C1(new_n902), .C2(new_n900), .ZN(new_n1151));
  AND3_X1   g0951(.A1(new_n892), .A2(G330), .A3(new_n1151), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1151), .B1(new_n892), .B2(G330), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n1149), .B1(new_n1152), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(new_n889), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n1155), .B(new_n1069), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n1156), .A2(KEYINPUT40), .B1(new_n868), .B2(new_n882), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n909), .B1(new_n1157), .B2(new_n666), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n892), .A2(G330), .A3(new_n1151), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1148), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n1139), .B1(new_n1154), .B2(new_n1160), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n734), .B1(G50), .B2(new_n1087), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n201), .B1(new_n264), .B2(G41), .ZN(new_n1163));
  XOR2_X1   g0963(.A(new_n1163), .B(KEYINPUT113), .Z(new_n1164));
  AOI22_X1  g0964(.A1(G116), .A2(new_n785), .B1(new_n756), .B2(G107), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n1165), .B1(new_n941), .B2(new_n770), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1166), .B1(G97), .B2(new_n781), .ZN(new_n1167));
  NOR3_X1   g0967(.A1(new_n1020), .A2(G41), .A3(new_n394), .ZN(new_n1168));
  NOR2_X1   g0968(.A1(new_n766), .A2(new_n202), .ZN(new_n1169));
  AOI21_X1  g0969(.A(new_n1169), .B1(new_n365), .B2(new_n759), .ZN(new_n1170));
  NAND4_X1  g0970(.A1(new_n1167), .A2(new_n930), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT58), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1164), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  OR3_X1    g0973(.A1(new_n767), .A2(new_n1095), .A3(KEYINPUT114), .ZN(new_n1174));
  OAI21_X1  g0974(.A(KEYINPUT114), .B1(new_n767), .B2(new_n1095), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1174), .B(new_n1175), .C1(new_n829), .C2(new_n774), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(G125), .A2(new_n785), .B1(new_n756), .B2(G128), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n1104), .B2(new_n758), .ZN(new_n1178));
  AOI211_X1 g0978(.A(new_n1176), .B(new_n1178), .C1(G132), .C2(new_n781), .ZN(new_n1179));
  INV_X1    g0979(.A(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n783), .C2(G159), .ZN(new_n1182));
  XNOR2_X1  g0982(.A(KEYINPUT115), .B(G124), .ZN(new_n1183));
  OAI211_X1 g0983(.A(new_n1181), .B(new_n1182), .C1(new_n770), .C2(new_n1183), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1185));
  OAI221_X1 g0985(.A(new_n1173), .B1(new_n1172), .B2(new_n1171), .C1(new_n1184), .C2(new_n1185), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n1162), .B1(new_n1186), .B2(new_n743), .ZN(new_n1187));
  OAI21_X1  g0987(.A(new_n1187), .B1(new_n1147), .B2(new_n738), .ZN(new_n1188));
  XOR2_X1   g0988(.A(new_n1188), .B(KEYINPUT119), .Z(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  NOR2_X1   g0990(.A1(new_n1161), .A2(new_n1190), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1130), .B1(new_n1075), .B2(new_n1118), .ZN(new_n1192));
  OAI211_X1 g0992(.A(G330), .B(new_n818), .C1(new_n1073), .C2(new_n1074), .ZN(new_n1193));
  AOI21_X1  g0993(.A(new_n1122), .B1(new_n1193), .B2(new_n905), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n1192), .A2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n1133), .B1(new_n1136), .B2(new_n1195), .ZN(new_n1196));
  AND3_X1   g0996(.A1(new_n1158), .A2(new_n1159), .A3(new_n1148), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1148), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1198));
  OAI211_X1 g0998(.A(KEYINPUT57), .B(new_n1196), .C1(new_n1197), .C2(new_n1198), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n678), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1154), .A2(new_n1160), .ZN(new_n1201));
  AOI21_X1  g1001(.A(KEYINPUT57), .B1(new_n1201), .B2(new_n1196), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1191), .B1(new_n1200), .B2(new_n1202), .ZN(G375));
  NAND3_X1  g1003(.A1(new_n1121), .A2(new_n1126), .A3(new_n1116), .ZN(new_n1204));
  NAND3_X1  g1004(.A1(new_n1134), .A2(new_n987), .A3(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(new_n1205), .B(KEYINPUT121), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n905), .A2(new_n737), .ZN(new_n1207));
  OAI22_X1  g1007(.A1(new_n755), .A2(new_n941), .B1(new_n758), .B2(new_n305), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n762), .A2(new_n338), .B1(new_n770), .B2(new_n938), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n408), .B1(new_n766), .B2(new_n511), .ZN(new_n1210));
  NOR4_X1   g1010(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1018), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n287), .B2(new_n794), .C1(new_n279), .C2(new_n780), .ZN(new_n1212));
  OAI221_X1 g1012(.A(new_n394), .B1(new_n774), .B2(new_n201), .C1(new_n202), .C2(new_n766), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n758), .A2(new_n829), .B1(new_n770), .B2(new_n1094), .ZN(new_n1214));
  OAI22_X1  g1014(.A1(new_n762), .A2(new_n826), .B1(new_n755), .B2(new_n1104), .ZN(new_n1215));
  NOR3_X1   g1015(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n780), .B2(new_n1095), .C1(new_n771), .C2(new_n794), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n752), .B1(new_n1212), .B2(new_n1217), .ZN(new_n1218));
  AOI211_X1 g1018(.A(new_n735), .B(new_n1218), .C1(new_n203), .C2(new_n822), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n1132), .A2(new_n733), .B1(new_n1207), .B2(new_n1219), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n1206), .A2(new_n1220), .ZN(G381));
  NOR3_X1   g1021(.A1(G393), .A2(G396), .A3(G384), .ZN(new_n1222));
  XNOR2_X1  g1022(.A(new_n1222), .B(KEYINPUT122), .ZN(new_n1223));
  INV_X1    g1023(.A(G387), .ZN(new_n1224));
  INV_X1    g1024(.A(G381), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1223), .A2(new_n1224), .A3(new_n1067), .A4(new_n1225), .ZN(new_n1226));
  INV_X1    g1026(.A(G375), .ZN(new_n1227));
  INV_X1    g1027(.A(G378), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1227), .A2(new_n1228), .ZN(new_n1229));
  OR2_X1    g1029(.A1(new_n1226), .A2(new_n1229), .ZN(G407));
  NAND2_X1  g1030(.A1(new_n658), .A2(G213), .ZN(new_n1231));
  XOR2_X1   g1031(.A(new_n1231), .B(KEYINPUT123), .Z(new_n1232));
  INV_X1    g1032(.A(new_n1232), .ZN(new_n1233));
  OAI211_X1 g1033(.A(G407), .B(G213), .C1(new_n1229), .C2(new_n1233), .ZN(G409));
  AND2_X1   g1034(.A1(new_n1232), .A2(G2897), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1121), .A2(new_n1126), .A3(new_n1116), .A4(KEYINPUT60), .ZN(new_n1236));
  INV_X1    g1036(.A(KEYINPUT125), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  NAND4_X1  g1038(.A1(new_n1195), .A2(KEYINPUT125), .A3(KEYINPUT60), .A4(new_n1116), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1204), .A2(new_n1240), .ZN(new_n1241));
  AOI21_X1  g1041(.A(new_n679), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1238), .A2(new_n1239), .A3(new_n1241), .A4(new_n1242), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1243), .A2(G384), .A3(new_n1220), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G384), .B1(new_n1243), .B2(new_n1220), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1235), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1243), .A2(new_n1220), .ZN(new_n1247));
  INV_X1    g1047(.A(G384), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1243), .A2(G384), .A3(new_n1220), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n658), .A2(G213), .A3(G2897), .ZN(new_n1251));
  NAND3_X1  g1051(.A1(new_n1249), .A2(new_n1250), .A3(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1246), .A2(new_n1252), .A3(KEYINPUT126), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT126), .ZN(new_n1254));
  OAI211_X1 g1054(.A(new_n1254), .B(new_n1235), .C1(new_n1244), .C2(new_n1245), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1253), .A2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(new_n1258), .A3(new_n1255), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(G375), .A2(G378), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1116), .B1(new_n1085), .B2(new_n1127), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(new_n1160), .B2(new_n1154), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G378), .B1(new_n1262), .B2(new_n987), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1201), .A2(new_n733), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(KEYINPUT124), .A3(new_n1189), .ZN(new_n1265));
  INV_X1    g1065(.A(KEYINPUT124), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n1266), .B1(new_n1161), .B2(new_n1190), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1263), .A2(new_n1265), .A3(new_n1267), .ZN(new_n1268));
  NAND3_X1  g1068(.A1(new_n1260), .A2(new_n1233), .A3(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1257), .A2(new_n1259), .A3(new_n1269), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1244), .A2(new_n1245), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1260), .A2(new_n1231), .A3(new_n1272), .A4(new_n1268), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  NOR3_X1   g1075(.A1(new_n1244), .A2(new_n1245), .A3(new_n1274), .ZN(new_n1276));
  NAND4_X1  g1076(.A1(new_n1260), .A2(new_n1233), .A3(new_n1268), .A4(new_n1276), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1275), .A2(new_n1277), .ZN(new_n1278));
  AND3_X1   g1078(.A1(new_n1270), .A2(new_n1271), .A3(new_n1278), .ZN(new_n1279));
  AOI22_X1  g1079(.A1(new_n980), .A2(new_n983), .B1(new_n724), .B2(new_n725), .ZN(new_n1280));
  OAI21_X1  g1080(.A(new_n1139), .B1(new_n1280), .B2(new_n986), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1281), .A2(new_n999), .ZN(new_n1282));
  AOI21_X1  g1082(.A(G390), .B1(new_n1282), .B2(new_n956), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n956), .ZN(new_n1284));
  AOI211_X1 g1084(.A(new_n1284), .B(new_n1067), .C1(new_n1281), .C2(new_n999), .ZN(new_n1285));
  XNOR2_X1  g1085(.A(G393), .B(new_n800), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1283), .A2(new_n1285), .A3(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(G387), .A2(new_n1067), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1282), .A2(new_n956), .A3(G390), .ZN(new_n1290));
  AOI21_X1  g1090(.A(new_n1286), .B1(new_n1289), .B2(new_n1290), .ZN(new_n1291));
  NOR2_X1   g1091(.A1(new_n1288), .A2(new_n1291), .ZN(new_n1292));
  INV_X1    g1092(.A(new_n1273), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1260), .A2(new_n1231), .A3(new_n1268), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1257), .A2(new_n1294), .A3(new_n1259), .ZN(new_n1295));
  AOI21_X1  g1095(.A(new_n1293), .B1(new_n1295), .B2(KEYINPUT63), .ZN(new_n1296));
  INV_X1    g1096(.A(new_n1269), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1297), .A2(KEYINPUT63), .A3(new_n1272), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1292), .A2(new_n1271), .A3(new_n1298), .ZN(new_n1299));
  OAI22_X1  g1099(.A1(new_n1279), .A2(new_n1292), .B1(new_n1296), .B2(new_n1299), .ZN(G405));
  NAND2_X1  g1100(.A1(new_n1229), .A2(new_n1260), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(new_n1272), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(new_n1292), .ZN(G402));
endmodule


