//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 1 0 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:28 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n511,
    new_n512, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n530, new_n531, new_n532, new_n533, new_n534, new_n535,
    new_n537, new_n539, new_n540, new_n542, new_n543, new_n544, new_n545,
    new_n546, new_n547, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n580, new_n581, new_n582, new_n583, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n596, new_n597, new_n600, new_n602, new_n603, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n812, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XOR2_X1   g012(.A(KEYINPUT66), .B(G69), .Z(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G220), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  OR4_X1    g026(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  NAND2_X1  g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  XNOR2_X1  g035(.A(new_n460), .B(KEYINPUT67), .ZN(new_n461));
  AND2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  NOR2_X1   g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  OAI21_X1  g038(.A(G125), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n459), .B1(new_n461), .B2(new_n464), .ZN(new_n465));
  OAI211_X1 g040(.A(G137), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n466));
  AND2_X1   g041(.A1(new_n459), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G101), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NOR2_X1   g044(.A1(new_n465), .A2(new_n469), .ZN(G160));
  OAI21_X1  g045(.A(KEYINPUT68), .B1(G100), .B2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(new_n471), .ZN(new_n472));
  NOR3_X1   g047(.A1(KEYINPUT68), .A2(G100), .A3(G2105), .ZN(new_n473));
  OAI221_X1 g048(.A(G2104), .B1(G112), .B2(new_n459), .C1(new_n472), .C2(new_n473), .ZN(new_n474));
  XNOR2_X1  g049(.A(new_n474), .B(KEYINPUT69), .ZN(new_n475));
  OR2_X1    g050(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n476));
  NAND2_X1  g051(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n477));
  AOI21_X1  g052(.A(G2105), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n459), .B1(new_n476), .B2(new_n477), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n475), .A2(new_n479), .A3(new_n481), .ZN(G162));
  INV_X1    g057(.A(G114), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n485));
  NAND2_X1  g060(.A1(G126), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n487), .B1(new_n462), .B2(new_n463), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n485), .A2(new_n488), .ZN(new_n489));
  OAI211_X1 g064(.A(G138), .B(new_n459), .C1(new_n462), .C2(new_n463), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n476), .A2(new_n477), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n492), .A2(new_n493), .A3(G138), .A4(new_n459), .ZN(new_n494));
  AOI21_X1  g069(.A(new_n489), .B1(new_n491), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g078(.A(KEYINPUT6), .B(G651), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  XNOR2_X1  g080(.A(KEYINPUT70), .B(G88), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(G543), .ZN(new_n507));
  INV_X1    g082(.A(G50), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n505), .A2(new_n506), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n503), .A2(new_n509), .ZN(G166));
  AND2_X1   g085(.A1(new_n504), .A2(G89), .ZN(new_n511));
  AND2_X1   g086(.A1(G63), .A2(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(new_n500), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NOR2_X1   g088(.A1(KEYINPUT6), .A2(G651), .ZN(new_n514));
  INV_X1    g089(.A(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(KEYINPUT6), .A2(G651), .ZN(new_n516));
  AOI21_X1  g091(.A(new_n497), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n518));
  OR2_X1    g093(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n518), .A2(KEYINPUT7), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n517), .A2(G51), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n513), .A2(new_n521), .ZN(G286));
  INV_X1    g097(.A(G286), .ZN(G168));
  AOI22_X1  g098(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n524));
  NOR2_X1   g099(.A1(new_n524), .A2(new_n502), .ZN(new_n525));
  XNOR2_X1  g100(.A(KEYINPUT71), .B(G90), .ZN(new_n526));
  INV_X1    g101(.A(G52), .ZN(new_n527));
  OAI22_X1  g102(.A1(new_n505), .A2(new_n526), .B1(new_n507), .B2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n525), .A2(new_n528), .ZN(G171));
  AOI22_X1  g104(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n502), .ZN(new_n531));
  INV_X1    g106(.A(G81), .ZN(new_n532));
  INV_X1    g107(.A(G43), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n505), .A2(new_n532), .B1(new_n507), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G860), .ZN(G153));
  NAND4_X1  g111(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT72), .ZN(G176));
  NAND2_X1  g113(.A1(G1), .A2(G3), .ZN(new_n539));
  XNOR2_X1  g114(.A(new_n539), .B(KEYINPUT8), .ZN(new_n540));
  NAND4_X1  g115(.A1(G319), .A2(G483), .A3(G661), .A4(new_n540), .ZN(G188));
  NAND2_X1  g116(.A1(G78), .A2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n500), .ZN(new_n543));
  INV_X1    g118(.A(G65), .ZN(new_n544));
  OAI21_X1  g119(.A(new_n542), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n515), .A2(new_n516), .B1(new_n498), .B2(new_n499), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n545), .A2(G651), .B1(G91), .B2(new_n546), .ZN(new_n547));
  INV_X1    g122(.A(G53), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(KEYINPUT73), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n517), .A2(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(KEYINPUT9), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n517), .A2(new_n552), .A3(new_n549), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n547), .A2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G171), .ZN(G301));
  INV_X1    g131(.A(G166), .ZN(G303));
  INV_X1    g132(.A(KEYINPUT74), .ZN(new_n558));
  OAI21_X1  g133(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n504), .A2(G49), .A3(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  AND3_X1   g136(.A1(new_n500), .A2(new_n504), .A3(G87), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n558), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n546), .A2(G87), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n564), .A2(KEYINPUT74), .A3(new_n559), .A4(new_n560), .ZN(new_n565));
  AND2_X1   g140(.A1(new_n563), .A2(new_n565), .ZN(G288));
  INV_X1    g141(.A(new_n499), .ZN(new_n567));
  NOR2_X1   g142(.A1(KEYINPUT5), .A2(G543), .ZN(new_n568));
  OAI21_X1  g143(.A(G61), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI22_X1  g146(.A1(new_n571), .A2(G651), .B1(new_n546), .B2(G86), .ZN(new_n572));
  AND2_X1   g147(.A1(KEYINPUT6), .A2(G651), .ZN(new_n573));
  OAI211_X1 g148(.A(G48), .B(G543), .C1(new_n573), .C2(new_n514), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT75), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n504), .A2(KEYINPUT75), .A3(G48), .A4(G543), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n572), .A2(new_n578), .ZN(G305));
  AOI22_X1  g154(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n502), .ZN(new_n581));
  INV_X1    g156(.A(G47), .ZN(new_n582));
  INV_X1    g157(.A(G85), .ZN(new_n583));
  OAI221_X1 g158(.A(new_n581), .B1(new_n582), .B2(new_n507), .C1(new_n583), .C2(new_n505), .ZN(G290));
  NAND2_X1  g159(.A1(G301), .A2(G868), .ZN(new_n585));
  AND3_X1   g160(.A1(new_n500), .A2(new_n504), .A3(G92), .ZN(new_n586));
  XNOR2_X1  g161(.A(new_n586), .B(KEYINPUT10), .ZN(new_n587));
  NAND2_X1  g162(.A1(G79), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G66), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n543), .B2(new_n589), .ZN(new_n590));
  AOI22_X1  g165(.A1(new_n590), .A2(G651), .B1(G54), .B2(new_n517), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G284));
  OAI21_X1  g169(.A(new_n585), .B1(new_n593), .B2(G868), .ZN(G321));
  NAND2_X1  g170(.A1(G286), .A2(G868), .ZN(new_n596));
  INV_X1    g171(.A(G299), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G297));
  OAI21_X1  g173(.A(new_n596), .B1(new_n597), .B2(G868), .ZN(G280));
  INV_X1    g174(.A(G559), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n593), .B1(new_n600), .B2(G860), .ZN(G148));
  NAND2_X1  g176(.A1(new_n593), .A2(new_n600), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G868), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n603), .B1(G868), .B2(new_n535), .ZN(G323));
  XNOR2_X1  g179(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g180(.A1(new_n492), .A2(new_n467), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n606), .B(KEYINPUT12), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n607), .B(KEYINPUT13), .ZN(new_n608));
  XNOR2_X1  g183(.A(new_n608), .B(G2100), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n480), .A2(G123), .ZN(new_n610));
  XOR2_X1   g185(.A(new_n610), .B(KEYINPUT77), .Z(new_n611));
  NAND2_X1  g186(.A1(new_n478), .A2(G135), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT76), .ZN(new_n613));
  OR2_X1    g188(.A1(G99), .A2(G2105), .ZN(new_n614));
  OAI211_X1 g189(.A(new_n614), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n615));
  NAND3_X1  g190(.A1(new_n611), .A2(new_n613), .A3(new_n615), .ZN(new_n616));
  OR2_X1    g191(.A1(new_n616), .A2(G2096), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n609), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT78), .ZN(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT15), .B(G2435), .ZN(new_n623));
  OR2_X1    g198(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n622), .A2(new_n623), .ZN(new_n625));
  NAND3_X1  g200(.A1(new_n624), .A2(KEYINPUT14), .A3(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(G1341), .B(G1348), .ZN(new_n627));
  XNOR2_X1  g202(.A(G2443), .B(G2446), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n626), .B(new_n629), .Z(new_n630));
  XOR2_X1   g205(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(G14), .B1(new_n630), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n630), .ZN(G401));
  XNOR2_X1  g211(.A(G2072), .B(G2078), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT17), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2067), .B(G2678), .ZN(new_n639));
  INV_X1    g214(.A(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n638), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(new_n643), .B(KEYINPUT81), .Z(new_n644));
  NAND3_X1  g219(.A1(new_n641), .A2(new_n637), .A3(new_n639), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT80), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT18), .ZN(new_n647));
  NAND2_X1  g222(.A1(new_n638), .A2(new_n639), .ZN(new_n648));
  INV_X1    g223(.A(new_n637), .ZN(new_n649));
  AOI21_X1  g224(.A(new_n641), .B1(new_n649), .B2(new_n640), .ZN(new_n650));
  AOI211_X1 g225(.A(new_n644), .B(new_n647), .C1(new_n648), .C2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(G2096), .B(G2100), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(G227));
  XOR2_X1   g228(.A(G1991), .B(G1996), .Z(new_n654));
  XOR2_X1   g229(.A(G1956), .B(G2474), .Z(new_n655));
  XOR2_X1   g230(.A(G1961), .B(G1966), .Z(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OR2_X1    g232(.A1(new_n657), .A2(KEYINPUT82), .ZN(new_n658));
  XOR2_X1   g233(.A(G1971), .B(G1976), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT19), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n657), .A2(KEYINPUT82), .ZN(new_n661));
  NAND3_X1  g236(.A1(new_n658), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(new_n662), .B(KEYINPUT20), .ZN(new_n663));
  OR2_X1    g238(.A1(new_n655), .A2(new_n656), .ZN(new_n664));
  NAND2_X1  g239(.A1(new_n664), .A2(new_n657), .ZN(new_n665));
  MUX2_X1   g240(.A(new_n665), .B(new_n664), .S(new_n660), .Z(new_n666));
  NAND2_X1  g241(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g242(.A(KEYINPUT83), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(KEYINPUT83), .A3(new_n666), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n672), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n671), .B1(new_n669), .B2(new_n670), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n654), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  INV_X1    g250(.A(new_n674), .ZN(new_n676));
  INV_X1    g251(.A(new_n654), .ZN(new_n677));
  NAND3_X1  g252(.A1(new_n676), .A2(new_n677), .A3(new_n672), .ZN(new_n678));
  XNOR2_X1  g253(.A(G1981), .B(G1986), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n682));
  NOR2_X1   g257(.A1(new_n681), .A2(new_n682), .ZN(G229));
  MUX2_X1   g258(.A(G24), .B(G290), .S(G16), .Z(new_n684));
  XNOR2_X1  g259(.A(new_n684), .B(KEYINPUT87), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G1986), .ZN(new_n686));
  NAND2_X1  g261(.A1(new_n478), .A2(G131), .ZN(new_n687));
  XOR2_X1   g262(.A(new_n687), .B(KEYINPUT84), .Z(new_n688));
  OAI21_X1  g263(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n689));
  INV_X1    g264(.A(G107), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G2105), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT85), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n480), .A2(G119), .ZN(new_n693));
  NAND3_X1  g268(.A1(new_n688), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  MUX2_X1   g269(.A(G25), .B(new_n694), .S(G29), .Z(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT86), .ZN(new_n696));
  XOR2_X1   g271(.A(KEYINPUT35), .B(G1991), .Z(new_n697));
  INV_X1    g272(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  OR2_X1    g274(.A1(new_n696), .A2(new_n698), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n686), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  MUX2_X1   g276(.A(G6), .B(G305), .S(G16), .Z(new_n702));
  XOR2_X1   g277(.A(KEYINPUT32), .B(G1981), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G22), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(G166), .B2(new_n705), .ZN(new_n707));
  INV_X1    g282(.A(G1971), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND3_X1  g284(.A1(new_n564), .A2(new_n559), .A3(new_n560), .ZN(new_n710));
  MUX2_X1   g285(.A(G23), .B(new_n710), .S(G16), .Z(new_n711));
  XNOR2_X1  g286(.A(KEYINPUT33), .B(G1976), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n711), .B(new_n712), .ZN(new_n713));
  NAND3_X1  g288(.A1(new_n704), .A2(new_n709), .A3(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT34), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n701), .A2(KEYINPUT36), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT36), .B1(new_n701), .B2(new_n715), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  INV_X1    g293(.A(G29), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n719), .A2(G26), .ZN(new_n720));
  XOR2_X1   g295(.A(new_n720), .B(KEYINPUT28), .Z(new_n721));
  NAND2_X1  g296(.A1(new_n478), .A2(G140), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n722), .B(KEYINPUT90), .Z(new_n723));
  NAND2_X1  g298(.A1(new_n480), .A2(G128), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n459), .A2(G116), .ZN(new_n725));
  OAI21_X1  g300(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n726));
  OAI211_X1 g301(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n726), .ZN(new_n727));
  AOI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(G29), .ZN(new_n728));
  INV_X1    g303(.A(G2067), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NOR2_X1   g305(.A1(G164), .A2(new_n719), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G27), .B2(new_n719), .ZN(new_n732));
  INV_X1    g307(.A(G2078), .ZN(new_n733));
  OR2_X1    g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  NOR2_X1   g310(.A1(G29), .A2(G32), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n736), .A2(KEYINPUT92), .ZN(new_n737));
  AOI22_X1  g312(.A1(new_n478), .A2(G141), .B1(G105), .B2(new_n467), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n480), .A2(G129), .ZN(new_n739));
  NAND3_X1  g314(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT26), .Z(new_n741));
  NAND3_X1  g316(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n742), .A2(new_n719), .ZN(new_n743));
  MUX2_X1   g318(.A(new_n737), .B(KEYINPUT92), .S(new_n743), .Z(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT27), .B(G1996), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n734), .B(new_n735), .C1(new_n744), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n705), .A2(G5), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(G171), .B2(new_n705), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(G1961), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  INV_X1    g327(.A(G34), .ZN(new_n753));
  AOI21_X1  g328(.A(G29), .B1(new_n753), .B2(KEYINPUT24), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(KEYINPUT24), .B2(new_n753), .ZN(new_n755));
  INV_X1    g330(.A(G160), .ZN(new_n756));
  OAI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(new_n719), .ZN(new_n757));
  OAI22_X1  g332(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n705), .A2(G21), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(G168), .B2(new_n705), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n760), .B(G1966), .ZN(new_n761));
  NOR4_X1   g336(.A1(new_n730), .A2(new_n747), .A3(new_n758), .A4(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(G4), .A2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n593), .B2(G16), .ZN(new_n764));
  XOR2_X1   g339(.A(KEYINPUT88), .B(G1348), .Z(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n719), .A2(G33), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT25), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n478), .A2(G139), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  INV_X1    g347(.A(KEYINPUT91), .ZN(new_n773));
  XNOR2_X1  g348(.A(new_n772), .B(new_n773), .ZN(new_n774));
  AOI22_X1  g349(.A1(new_n492), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n775));
  OR2_X1    g350(.A1(new_n775), .A2(new_n459), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n767), .B1(new_n778), .B2(new_n719), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n766), .B1(G2072), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n705), .A2(G20), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT23), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(new_n597), .B2(new_n705), .ZN(new_n783));
  INV_X1    g358(.A(G1956), .ZN(new_n784));
  XNOR2_X1  g359(.A(new_n783), .B(new_n784), .ZN(new_n785));
  OR2_X1    g360(.A1(new_n779), .A2(G2072), .ZN(new_n786));
  NAND4_X1  g361(.A1(new_n762), .A2(new_n780), .A3(new_n785), .A4(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G29), .A2(G35), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(G162), .B2(G29), .ZN(new_n789));
  XOR2_X1   g364(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  OR2_X1    g366(.A1(new_n791), .A2(G2090), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n791), .A2(G2090), .ZN(new_n793));
  NOR2_X1   g368(.A1(G16), .A2(G19), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n794), .B1(new_n535), .B2(G16), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n795), .B(KEYINPUT89), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(G1341), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT30), .B(G28), .ZN(new_n798));
  OR2_X1    g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  NAND2_X1  g374(.A1(KEYINPUT31), .A2(G11), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n798), .A2(new_n719), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n616), .B2(new_n719), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(KEYINPUT93), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n792), .A2(new_n793), .A3(new_n797), .A4(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n744), .A2(new_n746), .ZN(new_n805));
  AOI22_X1  g380(.A1(new_n750), .A2(new_n751), .B1(new_n752), .B2(new_n757), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT94), .Z(new_n808));
  NOR3_X1   g383(.A1(new_n787), .A2(new_n804), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n718), .A2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n810), .ZN(G311));
  INV_X1    g386(.A(KEYINPUT96), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n810), .B(new_n812), .ZN(G150));
  NOR2_X1   g388(.A1(new_n592), .A2(new_n600), .ZN(new_n814));
  XNOR2_X1  g389(.A(KEYINPUT97), .B(KEYINPUT38), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n814), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n535), .ZN(new_n817));
  AOI22_X1  g392(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n818));
  NOR2_X1   g393(.A1(new_n818), .A2(new_n502), .ZN(new_n819));
  INV_X1    g394(.A(G93), .ZN(new_n820));
  INV_X1    g395(.A(G55), .ZN(new_n821));
  OAI22_X1  g396(.A1(new_n505), .A2(new_n820), .B1(new_n507), .B2(new_n821), .ZN(new_n822));
  OR2_X1    g397(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n817), .A2(new_n823), .ZN(new_n824));
  NOR2_X1   g399(.A1(new_n819), .A2(new_n822), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n535), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  INV_X1    g402(.A(new_n827), .ZN(new_n828));
  XNOR2_X1  g403(.A(new_n816), .B(new_n828), .ZN(new_n829));
  AND2_X1   g404(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n829), .A2(KEYINPUT39), .ZN(new_n831));
  NOR3_X1   g406(.A1(new_n830), .A2(new_n831), .A3(G860), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n823), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  XOR2_X1   g409(.A(new_n834), .B(KEYINPUT37), .Z(new_n835));
  OR2_X1    g410(.A1(new_n832), .A2(new_n835), .ZN(G145));
  XNOR2_X1  g411(.A(new_n616), .B(new_n756), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(G162), .Z(new_n838));
  AOI21_X1  g413(.A(new_n486), .B1(new_n476), .B2(new_n477), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n459), .A2(G114), .ZN(new_n840));
  OAI21_X1  g415(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g417(.A(KEYINPUT99), .B1(new_n839), .B2(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(KEYINPUT99), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n485), .A2(new_n488), .A3(new_n844), .ZN(new_n845));
  AOI21_X1  g420(.A(new_n493), .B1(new_n478), .B2(G138), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n490), .A2(KEYINPUT4), .ZN(new_n847));
  OAI211_X1 g422(.A(new_n843), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(new_n727), .B(new_n848), .Z(new_n849));
  INV_X1    g424(.A(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n742), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n778), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n480), .A2(G130), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n478), .A2(G142), .ZN(new_n854));
  OR2_X1    g429(.A1(G106), .A2(G2105), .ZN(new_n855));
  OAI211_X1 g430(.A(new_n855), .B(G2104), .C1(G118), .C2(new_n459), .ZN(new_n856));
  NAND3_X1  g431(.A1(new_n853), .A2(new_n854), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n777), .A2(new_n742), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n852), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n852), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n850), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(new_n859), .A3(new_n849), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n694), .B(new_n607), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n866), .A2(KEYINPUT100), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n865), .B1(new_n862), .B2(new_n864), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n838), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  INV_X1    g445(.A(new_n838), .ZN(new_n871));
  NAND4_X1  g446(.A1(new_n870), .A2(KEYINPUT100), .A3(new_n871), .A4(new_n866), .ZN(new_n872));
  INV_X1    g447(.A(G37), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n869), .A2(new_n872), .A3(new_n873), .ZN(new_n874));
  XOR2_X1   g449(.A(KEYINPUT101), .B(KEYINPUT40), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(G395));
  XNOR2_X1  g451(.A(new_n597), .B(new_n592), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n877), .B(KEYINPUT41), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n602), .B(new_n827), .ZN(new_n879));
  NOR2_X1   g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT102), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n879), .A2(new_n877), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NOR2_X1   g459(.A1(new_n880), .A2(new_n881), .ZN(new_n885));
  OR3_X1    g460(.A1(new_n884), .A2(new_n885), .A3(KEYINPUT42), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n710), .B(KEYINPUT103), .Z(new_n887));
  XNOR2_X1  g462(.A(new_n887), .B(G305), .ZN(new_n888));
  XNOR2_X1  g463(.A(G290), .B(G166), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(KEYINPUT42), .B1(new_n884), .B2(new_n885), .ZN(new_n892));
  AND3_X1   g467(.A1(new_n886), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n891), .B1(new_n886), .B2(new_n892), .ZN(new_n894));
  OAI21_X1  g469(.A(G868), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n895), .B1(G868), .B2(new_n825), .ZN(G295));
  OAI21_X1  g471(.A(new_n895), .B1(G868), .B2(new_n825), .ZN(G331));
  XNOR2_X1  g472(.A(KEYINPUT104), .B(KEYINPUT44), .ZN(new_n898));
  NAND2_X1  g473(.A1(G171), .A2(KEYINPUT105), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n827), .B(new_n899), .ZN(new_n900));
  OAI21_X1  g475(.A(G286), .B1(G171), .B2(KEYINPUT105), .ZN(new_n901));
  INV_X1    g476(.A(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n828), .A2(new_n899), .ZN(new_n904));
  AOI21_X1  g479(.A(new_n827), .B1(KEYINPUT105), .B2(G171), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n901), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND3_X1  g481(.A1(new_n903), .A2(new_n906), .A3(new_n877), .ZN(new_n907));
  INV_X1    g482(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n878), .B1(new_n903), .B2(new_n906), .ZN(new_n909));
  OAI21_X1  g484(.A(new_n890), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n903), .A2(new_n906), .ZN(new_n911));
  OAI211_X1 g486(.A(new_n891), .B(new_n907), .C1(new_n911), .C2(new_n878), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n873), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT43), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n907), .B1(new_n911), .B2(new_n878), .ZN(new_n916));
  AOI21_X1  g491(.A(G37), .B1(new_n916), .B2(new_n890), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n917), .B2(new_n912), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n898), .B1(new_n914), .B2(new_n918), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT106), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n913), .A2(KEYINPUT43), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n917), .A2(new_n915), .A3(new_n912), .ZN(new_n923));
  NAND3_X1  g498(.A1(new_n922), .A2(new_n923), .A3(KEYINPUT44), .ZN(new_n924));
  OAI211_X1 g499(.A(KEYINPUT106), .B(new_n898), .C1(new_n914), .C2(new_n918), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n924), .A3(new_n925), .ZN(G397));
  INV_X1    g501(.A(G1384), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n848), .A2(new_n927), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT45), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g505(.A1(G160), .A2(G40), .ZN(new_n931));
  NOR2_X1   g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n933), .A2(G1986), .A3(G290), .ZN(new_n934));
  AND2_X1   g509(.A1(G290), .A2(G1986), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n934), .B1(new_n932), .B2(new_n935), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n936), .B(KEYINPUT107), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n727), .B(new_n729), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n742), .A2(G1996), .ZN(new_n939));
  AOI21_X1  g514(.A(new_n933), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(G1996), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n932), .A2(new_n941), .ZN(new_n942));
  OR3_X1    g517(.A1(new_n942), .A2(KEYINPUT108), .A3(new_n742), .ZN(new_n943));
  OAI21_X1  g518(.A(KEYINPUT108), .B1(new_n942), .B2(new_n742), .ZN(new_n944));
  AOI21_X1  g519(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n694), .A2(new_n698), .ZN(new_n946));
  NOR2_X1   g521(.A1(new_n694), .A2(new_n698), .ZN(new_n947));
  OAI21_X1  g522(.A(new_n932), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n945), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n937), .A2(new_n949), .ZN(new_n950));
  XOR2_X1   g525(.A(new_n950), .B(KEYINPUT109), .Z(new_n951));
  INV_X1    g526(.A(KEYINPUT51), .ZN(new_n952));
  INV_X1    g527(.A(G8), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n839), .A2(new_n842), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(new_n846), .B2(new_n847), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n955), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT114), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(G40), .ZN(new_n959));
  NOR3_X1   g534(.A1(new_n465), .A2(new_n959), .A3(new_n469), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n955), .A2(KEYINPUT114), .A3(KEYINPUT45), .A4(new_n927), .ZN(new_n961));
  NAND4_X1  g536(.A1(new_n930), .A2(new_n958), .A3(new_n960), .A4(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1966), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT50), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n848), .A2(new_n964), .A3(new_n927), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n965), .A2(new_n960), .A3(new_n966), .ZN(new_n967));
  AOI22_X1  g542(.A1(new_n962), .A2(new_n963), .B1(new_n752), .B2(new_n967), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n953), .B1(new_n968), .B2(G168), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n962), .A2(new_n963), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n967), .A2(new_n752), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(G286), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n952), .B1(new_n969), .B2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(KEYINPUT51), .B(new_n953), .C1(new_n968), .C2(G168), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n976), .A2(KEYINPUT62), .ZN(new_n978));
  NOR2_X1   g553(.A1(G166), .A2(new_n953), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n979), .B(KEYINPUT55), .ZN(new_n980));
  NOR3_X1   g555(.A1(new_n839), .A2(new_n842), .A3(KEYINPUT99), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n844), .B1(new_n485), .B2(new_n488), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n491), .A2(new_n494), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI211_X1 g560(.A(KEYINPUT113), .B(new_n960), .C1(new_n985), .C2(new_n964), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT113), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n964), .B1(new_n848), .B2(new_n927), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n988), .B2(new_n931), .ZN(new_n989));
  INV_X1    g564(.A(G2090), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n955), .A2(new_n964), .A3(new_n927), .ZN(new_n991));
  NAND4_X1  g566(.A1(new_n986), .A2(new_n989), .A3(new_n990), .A4(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n848), .A2(KEYINPUT45), .A3(new_n927), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n929), .B1(G164), .B2(G1384), .ZN(new_n994));
  NAND3_X1  g569(.A1(new_n993), .A2(new_n960), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n708), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n980), .B1(new_n997), .B2(G8), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n965), .A2(new_n966), .A3(new_n990), .A4(new_n960), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n1000), .A2(G8), .A3(new_n980), .ZN(new_n1001));
  INV_X1    g576(.A(G1981), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n546), .A2(G86), .ZN(new_n1003));
  INV_X1    g578(.A(G61), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n1004), .B1(new_n498), .B2(new_n499), .ZN(new_n1005));
  INV_X1    g580(.A(new_n570), .ZN(new_n1006));
  OAI21_X1  g581(.A(G651), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n578), .A2(new_n1002), .A3(new_n1003), .A4(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT110), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  NAND4_X1  g585(.A1(new_n572), .A2(new_n1010), .A3(new_n1002), .A4(new_n578), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G305), .A2(G1981), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT49), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1012), .A2(KEYINPUT49), .A3(new_n1013), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n960), .A2(new_n848), .A3(new_n927), .ZN(new_n1018));
  INV_X1    g593(.A(new_n1018), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1019), .A2(new_n953), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1016), .A2(new_n1017), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G1976), .ZN(new_n1022));
  OR2_X1    g597(.A1(new_n710), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1023), .A3(G8), .ZN(new_n1024));
  AND2_X1   g599(.A1(new_n1024), .A2(KEYINPUT52), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n563), .A2(new_n1022), .A3(new_n565), .ZN(new_n1026));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1026), .A2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g603(.A1(new_n1024), .A2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g604(.A1(new_n1025), .A2(new_n1029), .ZN(new_n1030));
  NAND3_X1  g605(.A1(new_n1001), .A2(new_n1021), .A3(new_n1030), .ZN(new_n1031));
  AOI21_X1  g606(.A(new_n931), .B1(new_n928), .B2(new_n929), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT53), .ZN(new_n1033));
  NOR2_X1   g608(.A1(new_n1033), .A2(G2078), .ZN(new_n1034));
  NAND4_X1  g609(.A1(new_n1032), .A2(new_n958), .A3(new_n961), .A4(new_n1034), .ZN(new_n1035));
  NAND4_X1  g610(.A1(new_n993), .A2(new_n994), .A3(new_n733), .A4(new_n960), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1033), .ZN(new_n1037));
  NAND3_X1  g612(.A1(new_n965), .A2(new_n960), .A3(new_n966), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1038), .A2(new_n751), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1035), .A2(new_n1037), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(G171), .ZN(new_n1041));
  NOR3_X1   g616(.A1(new_n998), .A2(new_n1031), .A3(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n977), .A2(new_n978), .A3(new_n1042), .ZN(new_n1043));
  NOR2_X1   g618(.A1(G288), .A2(G1976), .ZN(new_n1044));
  AOI22_X1  g619(.A1(new_n1021), .A2(new_n1044), .B1(new_n1009), .B2(new_n1011), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT112), .ZN(new_n1046));
  OR2_X1    g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1048));
  XNOR2_X1  g623(.A(new_n1020), .B(KEYINPUT111), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n1047), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n953), .B1(new_n996), .B2(new_n999), .ZN(new_n1051));
  AND4_X1   g626(.A1(new_n980), .A2(new_n1030), .A3(new_n1021), .A4(new_n1051), .ZN(new_n1052));
  NOR3_X1   g627(.A1(new_n968), .A2(new_n953), .A3(G286), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1051), .A2(new_n980), .ZN(new_n1054));
  NAND4_X1  g629(.A1(new_n1053), .A2(new_n1054), .A3(new_n1021), .A4(new_n1030), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1052), .B1(new_n1055), .B2(KEYINPUT63), .ZN(new_n1056));
  NOR2_X1   g631(.A1(new_n998), .A2(new_n1031), .ZN(new_n1057));
  INV_X1    g632(.A(KEYINPUT63), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1057), .A2(new_n1058), .A3(new_n1053), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1050), .A2(new_n1056), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n931), .B1(new_n985), .B2(KEYINPUT45), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1034), .ZN(new_n1062));
  AOI21_X1  g637(.A(new_n1062), .B1(new_n928), .B2(new_n929), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1061), .A2(new_n1063), .B1(new_n1036), .B2(new_n1033), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT120), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1039), .A2(new_n1065), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n1038), .A2(KEYINPUT120), .A3(new_n751), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(new_n1066), .A3(G301), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(new_n1041), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT54), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  OAI211_X1 g646(.A(new_n1057), .B(new_n1071), .C1(new_n974), .C2(new_n975), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1064), .A2(new_n1066), .A3(new_n1067), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1070), .B1(new_n1073), .B2(G171), .ZN(new_n1074));
  NAND4_X1  g649(.A1(new_n1035), .A2(new_n1037), .A3(G301), .A4(new_n1039), .ZN(new_n1075));
  OR2_X1    g650(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(KEYINPUT121), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1074), .A2(new_n1076), .A3(new_n1077), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1078), .A2(KEYINPUT122), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT122), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1074), .A2(new_n1076), .A3(new_n1080), .A4(new_n1077), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1072), .B1(new_n1079), .B2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT57), .B1(new_n554), .B2(KEYINPUT115), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1083), .A2(G299), .ZN(new_n1084));
  OAI211_X1 g659(.A(new_n547), .B(new_n554), .C1(KEYINPUT115), .C2(KEYINPUT57), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT117), .ZN(new_n1087));
  XNOR2_X1  g662(.A(new_n1086), .B(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g663(.A(KEYINPUT56), .B(G2072), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  NOR2_X1   g665(.A1(new_n995), .A2(new_n1090), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n986), .A2(new_n989), .A3(new_n991), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1091), .B1(new_n1092), .B2(new_n784), .ZN(new_n1093));
  NOR2_X1   g668(.A1(new_n1088), .A2(new_n1093), .ZN(new_n1094));
  INV_X1    g669(.A(G1348), .ZN(new_n1095));
  AOI22_X1  g670(.A1(new_n1038), .A2(new_n1095), .B1(new_n1019), .B2(new_n729), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT116), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(new_n592), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT61), .ZN(new_n1101));
  AND2_X1   g676(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1093), .A2(new_n1086), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1101), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n993), .A2(new_n994), .A3(new_n941), .A4(new_n960), .ZN(new_n1105));
  XOR2_X1   g680(.A(KEYINPUT58), .B(G1341), .Z(new_n1106));
  NAND2_X1  g681(.A1(new_n1018), .A2(new_n1106), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n817), .B1(new_n1105), .B2(new_n1107), .ZN(new_n1108));
  XNOR2_X1  g683(.A(new_n1108), .B(KEYINPUT59), .ZN(new_n1109));
  OR2_X1    g684(.A1(new_n593), .A2(KEYINPUT60), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1096), .A2(KEYINPUT116), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1096), .A2(KEYINPUT116), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n593), .A2(KEYINPUT60), .ZN(new_n1114));
  XNOR2_X1  g689(.A(new_n1114), .B(KEYINPUT119), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1109), .B1(new_n1113), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1115), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1097), .A2(new_n1117), .A3(new_n1110), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1104), .A2(new_n1116), .A3(new_n1118), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1099), .A2(KEYINPUT118), .ZN(new_n1120));
  OAI21_X1  g695(.A(KEYINPUT61), .B1(new_n1088), .B2(new_n1093), .ZN(new_n1121));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n1122));
  AOI21_X1  g697(.A(new_n1122), .B1(new_n1093), .B2(new_n1086), .ZN(new_n1123));
  NOR3_X1   g698(.A1(new_n1120), .A2(new_n1121), .A3(new_n1123), .ZN(new_n1124));
  OAI21_X1  g699(.A(new_n1100), .B1(new_n1119), .B2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1060), .B1(new_n1082), .B2(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT123), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1043), .B1(new_n1126), .B2(new_n1127), .ZN(new_n1128));
  AOI211_X1 g703(.A(KEYINPUT123), .B(new_n1060), .C1(new_n1082), .C2(new_n1125), .ZN(new_n1129));
  OAI21_X1  g704(.A(new_n951), .B1(new_n1128), .B2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n945), .A2(new_n947), .ZN(new_n1131));
  OAI21_X1  g706(.A(new_n1131), .B1(G2067), .B2(new_n727), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1132), .A2(new_n932), .ZN(new_n1133));
  OR2_X1    g708(.A1(new_n1133), .A2(KEYINPUT124), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(KEYINPUT124), .ZN(new_n1135));
  XOR2_X1   g710(.A(new_n942), .B(KEYINPUT46), .Z(new_n1136));
  AOI21_X1  g711(.A(new_n933), .B1(new_n938), .B2(new_n851), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  XOR2_X1   g713(.A(KEYINPUT125), .B(KEYINPUT47), .Z(new_n1139));
  XNOR2_X1  g714(.A(new_n1138), .B(new_n1139), .ZN(new_n1140));
  XOR2_X1   g715(.A(new_n934), .B(KEYINPUT48), .Z(new_n1141));
  AOI21_X1  g716(.A(new_n1140), .B1(new_n949), .B2(new_n1141), .ZN(new_n1142));
  AND3_X1   g717(.A1(new_n1134), .A2(new_n1135), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1130), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g719(.A1(G227), .A2(new_n457), .A3(G401), .ZN(new_n1146));
  INV_X1    g720(.A(new_n682), .ZN(new_n1147));
  AOI21_X1  g721(.A(new_n1146), .B1(new_n680), .B2(new_n1147), .ZN(new_n1148));
  OAI211_X1 g722(.A(new_n1148), .B(new_n874), .C1(new_n914), .C2(new_n918), .ZN(G225));
  INV_X1    g723(.A(KEYINPUT126), .ZN(new_n1150));
  NOR2_X1   g724(.A1(G225), .A2(new_n1150), .ZN(new_n1151));
  NOR3_X1   g725(.A1(G227), .A2(new_n457), .A3(G401), .ZN(new_n1152));
  OAI21_X1  g726(.A(new_n1152), .B1(new_n681), .B2(new_n682), .ZN(new_n1153));
  AOI21_X1  g727(.A(new_n1153), .B1(new_n922), .B2(new_n923), .ZN(new_n1154));
  AOI21_X1  g728(.A(KEYINPUT126), .B1(new_n1154), .B2(new_n874), .ZN(new_n1155));
  NOR2_X1   g729(.A1(new_n1151), .A2(new_n1155), .ZN(G308));
endmodule


