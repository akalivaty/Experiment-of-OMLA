//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 0 1 1 0 0 1 0 1 0 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 0 0 1 0 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:52 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  AND2_X1   g005(.A1(KEYINPUT0), .A2(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n191), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(G143), .B(G146), .ZN(new_n194));
  XNOR2_X1  g008(.A(KEYINPUT0), .B(G128), .ZN(new_n195));
  OAI21_X1  g009(.A(new_n193), .B1(new_n194), .B2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G125), .ZN(new_n197));
  INV_X1    g011(.A(G128), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(KEYINPUT1), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n199), .A2(new_n189), .A3(new_n191), .ZN(new_n200));
  OAI211_X1 g014(.A(new_n190), .B(G146), .C1(new_n198), .C2(KEYINPUT1), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n198), .A2(new_n188), .A3(G143), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n200), .A2(new_n201), .A3(new_n202), .ZN(new_n203));
  OAI21_X1  g017(.A(new_n197), .B1(G125), .B2(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G953), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G224), .ZN(new_n206));
  XOR2_X1   g020(.A(new_n204), .B(new_n206), .Z(new_n207));
  INV_X1    g021(.A(KEYINPUT65), .ZN(new_n208));
  INV_X1    g022(.A(G119), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n208), .B1(new_n209), .B2(G116), .ZN(new_n210));
  INV_X1    g024(.A(G116), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n211), .A2(KEYINPUT65), .A3(G119), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n209), .A2(G116), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n213), .A2(KEYINPUT5), .A3(new_n214), .ZN(new_n215));
  OR2_X1    g029(.A1(new_n214), .A2(KEYINPUT5), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(G113), .A3(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(G104), .ZN(new_n218));
  OAI21_X1  g032(.A(KEYINPUT3), .B1(new_n218), .B2(G107), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n220));
  INV_X1    g034(.A(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(new_n221), .A3(G104), .ZN(new_n222));
  INV_X1    g036(.A(G101), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(G107), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n219), .A2(new_n222), .A3(new_n223), .A4(new_n224), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n221), .A2(G104), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n218), .A2(G107), .ZN(new_n227));
  OAI21_X1  g041(.A(G101), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n225), .A2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(new_n229), .ZN(new_n230));
  AOI22_X1  g044(.A1(new_n210), .A2(new_n212), .B1(G116), .B2(new_n209), .ZN(new_n231));
  AND2_X1   g045(.A1(KEYINPUT2), .A2(G113), .ZN(new_n232));
  INV_X1    g046(.A(KEYINPUT64), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT2), .ZN(new_n234));
  INV_X1    g048(.A(G113), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n233), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  OAI21_X1  g050(.A(KEYINPUT64), .B1(KEYINPUT2), .B2(G113), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n232), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  AND3_X1   g052(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT66), .ZN(new_n239));
  AOI21_X1  g053(.A(KEYINPUT66), .B1(new_n231), .B2(new_n238), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n217), .B(new_n230), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n231), .A2(new_n238), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n231), .A2(new_n238), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n231), .A2(new_n238), .A3(KEYINPUT66), .ZN(new_n246));
  AOI21_X1  g060(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n219), .A2(new_n222), .A3(new_n224), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n248), .A2(G101), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n249), .A2(KEYINPUT4), .A3(new_n225), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT4), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n248), .A2(new_n251), .A3(G101), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  OAI21_X1  g067(.A(new_n241), .B1(new_n247), .B2(new_n253), .ZN(new_n254));
  XOR2_X1   g068(.A(G110), .B(G122), .Z(new_n255));
  NAND2_X1  g069(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n256), .A2(KEYINPUT6), .ZN(new_n257));
  INV_X1    g071(.A(new_n257), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n254), .A2(KEYINPUT82), .A3(new_n255), .ZN(new_n259));
  AOI21_X1  g073(.A(KEYINPUT82), .B1(new_n254), .B2(new_n255), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(new_n255), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n241), .B(new_n262), .C1(new_n247), .C2(new_n253), .ZN(new_n263));
  AND2_X1   g077(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT83), .B1(new_n261), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n263), .A2(KEYINPUT6), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT83), .ZN(new_n267));
  NOR4_X1   g081(.A1(new_n259), .A2(new_n260), .A3(new_n266), .A4(new_n267), .ZN(new_n268));
  OAI211_X1 g082(.A(new_n207), .B(new_n258), .C1(new_n265), .C2(new_n268), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n255), .B(KEYINPUT8), .ZN(new_n270));
  OAI21_X1  g084(.A(new_n217), .B1(new_n239), .B2(new_n240), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(new_n229), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n270), .B1(new_n272), .B2(new_n241), .ZN(new_n273));
  INV_X1    g087(.A(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n206), .A2(KEYINPUT7), .ZN(new_n275));
  XNOR2_X1  g089(.A(new_n204), .B(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n274), .A2(new_n277), .A3(KEYINPUT84), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT84), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n279), .B1(new_n273), .B2(new_n276), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n278), .A2(new_n263), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(G902), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT85), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n281), .A2(new_n285), .A3(new_n282), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n269), .A2(new_n284), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(G210), .B1(G237), .B2(G902), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT86), .ZN(new_n291));
  NAND4_X1  g105(.A1(new_n269), .A2(new_n284), .A3(new_n288), .A4(new_n286), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n290), .A2(new_n291), .A3(new_n292), .ZN(new_n293));
  OR2_X1    g107(.A1(new_n292), .A2(new_n291), .ZN(new_n294));
  INV_X1    g108(.A(KEYINPUT90), .ZN(new_n295));
  NOR2_X1   g109(.A1(G237), .A2(G953), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(G143), .A3(G214), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(G143), .B1(new_n296), .B2(G214), .ZN(new_n299));
  OAI21_X1  g113(.A(G131), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT17), .ZN(new_n301));
  INV_X1    g115(.A(G237), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n302), .A2(new_n205), .A3(G214), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n190), .ZN(new_n304));
  INV_X1    g118(.A(G131), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n305), .A3(new_n297), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n300), .A2(new_n301), .A3(new_n306), .ZN(new_n307));
  XNOR2_X1  g121(.A(G125), .B(G140), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n308), .A2(KEYINPUT16), .ZN(new_n309));
  INV_X1    g123(.A(G125), .ZN(new_n310));
  OR3_X1    g124(.A1(new_n310), .A2(KEYINPUT16), .A3(G140), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(new_n188), .ZN(new_n313));
  OAI211_X1 g127(.A(KEYINPUT17), .B(G131), .C1(new_n298), .C2(new_n299), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n309), .A2(G146), .A3(new_n311), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n307), .A2(new_n313), .A3(new_n314), .A4(new_n315), .ZN(new_n316));
  XOR2_X1   g130(.A(G125), .B(G140), .Z(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G146), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n308), .A2(new_n188), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  AND2_X1   g134(.A1(KEYINPUT18), .A2(G131), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n298), .A2(new_n299), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n321), .B1(new_n322), .B2(KEYINPUT87), .ZN(new_n323));
  AND4_X1   g137(.A1(KEYINPUT87), .A2(new_n304), .A3(new_n321), .A4(new_n297), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n320), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n316), .A2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(G113), .B(G122), .Z(new_n327));
  XNOR2_X1  g141(.A(new_n327), .B(KEYINPUT89), .ZN(new_n328));
  XNOR2_X1  g142(.A(new_n328), .B(new_n218), .ZN(new_n329));
  OAI21_X1  g143(.A(new_n295), .B1(new_n326), .B2(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(new_n328), .B(G104), .ZN(new_n331));
  NAND4_X1  g145(.A1(new_n331), .A2(new_n325), .A3(new_n316), .A4(KEYINPUT90), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT88), .ZN(new_n334));
  NOR3_X1   g148(.A1(new_n317), .A2(new_n334), .A3(KEYINPUT19), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT19), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n308), .A2(new_n336), .ZN(new_n337));
  AOI21_X1  g151(.A(KEYINPUT88), .B1(new_n308), .B2(new_n336), .ZN(new_n338));
  NOR3_X1   g152(.A1(new_n335), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(new_n188), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n300), .A2(new_n306), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n315), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n342), .A2(new_n325), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n329), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n333), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(G475), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n345), .A2(new_n346), .A3(new_n282), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT20), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AOI22_X1  g163(.A1(new_n330), .A2(new_n332), .B1(new_n329), .B2(new_n326), .ZN(new_n350));
  OAI21_X1  g164(.A(G475), .B1(new_n350), .B2(G902), .ZN(new_n351));
  AOI21_X1  g165(.A(G475), .B1(new_n333), .B2(new_n344), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n352), .A2(KEYINPUT20), .A3(new_n282), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(G952), .ZN(new_n355));
  AND2_X1   g169(.A1(new_n355), .A2(KEYINPUT95), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(KEYINPUT95), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n205), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(G237), .ZN(new_n359));
  XNOR2_X1  g173(.A(KEYINPUT73), .B(G902), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  AOI211_X1 g175(.A(new_n205), .B(new_n361), .C1(G234), .C2(G237), .ZN(new_n362));
  XOR2_X1   g176(.A(KEYINPUT21), .B(G898), .Z(new_n363));
  INV_X1    g177(.A(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(new_n359), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n190), .A2(G128), .ZN(new_n366));
  XNOR2_X1  g180(.A(KEYINPUT92), .B(KEYINPUT13), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n198), .A2(G143), .ZN(new_n368));
  INV_X1    g182(.A(new_n368), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT93), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n366), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n372), .B1(new_n371), .B2(new_n370), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n367), .A2(new_n369), .ZN(new_n374));
  OAI21_X1  g188(.A(G134), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n366), .A2(new_n368), .ZN(new_n376));
  OR2_X1    g190(.A1(new_n376), .A2(KEYINPUT94), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(KEYINPUT94), .ZN(new_n378));
  AOI21_X1  g192(.A(G134), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  XNOR2_X1  g194(.A(G116), .B(G122), .ZN(new_n381));
  XNOR2_X1  g195(.A(KEYINPUT91), .B(G107), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n375), .A2(new_n380), .A3(new_n383), .ZN(new_n384));
  OR2_X1    g198(.A1(new_n211), .A2(G122), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n221), .B1(new_n385), .B2(KEYINPUT14), .ZN(new_n386));
  XNOR2_X1  g200(.A(new_n386), .B(new_n381), .ZN(new_n387));
  AND3_X1   g201(.A1(new_n378), .A2(G134), .A3(new_n377), .ZN(new_n388));
  OAI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(new_n379), .ZN(new_n389));
  XOR2_X1   g203(.A(KEYINPUT9), .B(G234), .Z(new_n390));
  INV_X1    g204(.A(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(G217), .ZN(new_n392));
  NOR3_X1   g206(.A1(new_n391), .A2(new_n392), .A3(G953), .ZN(new_n393));
  AND3_X1   g207(.A1(new_n384), .A2(new_n389), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n393), .B1(new_n384), .B2(new_n389), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n361), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(G478), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n397), .A2(KEYINPUT15), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI221_X1 g213(.A(new_n361), .B1(KEYINPUT15), .B2(new_n397), .C1(new_n394), .C2(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NOR3_X1   g215(.A1(new_n354), .A2(new_n365), .A3(new_n401), .ZN(new_n402));
  AND4_X1   g216(.A1(new_n187), .A2(new_n293), .A3(new_n294), .A4(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(KEYINPUT11), .ZN(new_n404));
  INV_X1    g218(.A(G134), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n404), .B1(new_n405), .B2(G137), .ZN(new_n406));
  INV_X1    g220(.A(G137), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n407), .A2(KEYINPUT11), .A3(G134), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n405), .A2(G137), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n406), .A2(new_n408), .A3(new_n305), .A4(new_n409), .ZN(new_n410));
  NOR2_X1   g224(.A1(new_n407), .A2(G134), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n405), .A2(G137), .ZN(new_n412));
  OAI21_X1  g226(.A(G131), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n410), .A2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT67), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n199), .A2(new_n189), .A3(new_n191), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n201), .A2(new_n202), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND4_X1  g232(.A1(new_n200), .A2(KEYINPUT67), .A3(new_n201), .A4(new_n202), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n414), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT30), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n406), .A2(new_n409), .A3(new_n408), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(G131), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n196), .B1(new_n423), .B2(new_n410), .ZN(new_n424));
  NOR3_X1   g238(.A1(new_n420), .A2(new_n421), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n423), .A2(new_n410), .ZN(new_n426));
  INV_X1    g240(.A(new_n196), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND2_X1   g242(.A1(new_n410), .A2(new_n413), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(new_n203), .ZN(new_n430));
  AOI21_X1  g244(.A(KEYINPUT30), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(KEYINPUT68), .B1(new_n425), .B2(new_n431), .ZN(new_n432));
  OAI22_X1  g246(.A1(new_n239), .A2(new_n240), .B1(new_n238), .B2(new_n231), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n418), .A2(new_n419), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n434), .A2(new_n429), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(KEYINPUT30), .A3(new_n428), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT68), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n432), .A2(new_n433), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n247), .A2(new_n435), .A3(new_n428), .ZN(new_n440));
  XNOR2_X1  g254(.A(KEYINPUT26), .B(G101), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n296), .A2(G210), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n441), .B(new_n442), .ZN(new_n443));
  XNOR2_X1  g257(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n444));
  XNOR2_X1  g258(.A(new_n443), .B(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n439), .A2(new_n440), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(KEYINPUT70), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n449));
  NAND4_X1  g263(.A1(new_n439), .A2(new_n449), .A3(new_n440), .A4(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n448), .A2(KEYINPUT31), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT31), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n447), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g268(.A1(new_n420), .A2(new_n424), .ZN(new_n455));
  AOI211_X1 g269(.A(KEYINPUT71), .B(KEYINPUT28), .C1(new_n455), .C2(new_n247), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT71), .ZN(new_n457));
  INV_X1    g271(.A(KEYINPUT28), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n457), .B1(new_n440), .B2(new_n458), .ZN(new_n459));
  NOR2_X1   g273(.A1(new_n456), .A2(new_n459), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n247), .B1(new_n428), .B2(new_n430), .ZN(new_n461));
  NOR3_X1   g275(.A1(new_n433), .A2(new_n420), .A3(new_n424), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT28), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n445), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n454), .A2(new_n465), .ZN(new_n466));
  NOR2_X1   g280(.A1(G472), .A2(G902), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(KEYINPUT32), .A3(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT32), .ZN(new_n469));
  INV_X1    g283(.A(new_n465), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n470), .B1(new_n451), .B2(new_n453), .ZN(new_n471));
  INV_X1    g285(.A(new_n467), .ZN(new_n472));
  OAI21_X1  g286(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT72), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n474), .B1(new_n456), .B2(new_n459), .ZN(new_n475));
  OAI21_X1  g289(.A(KEYINPUT71), .B1(new_n462), .B2(KEYINPUT28), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n440), .A2(new_n457), .A3(new_n458), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n476), .A2(KEYINPUT72), .A3(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n455), .A2(new_n247), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT28), .B1(new_n479), .B2(new_n462), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT29), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n445), .A2(new_n481), .ZN(new_n482));
  NAND4_X1  g296(.A1(new_n475), .A2(new_n478), .A3(new_n480), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(new_n361), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n484), .A2(KEYINPUT74), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n439), .A2(new_n440), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n445), .ZN(new_n487));
  OAI211_X1 g301(.A(new_n487), .B(new_n481), .C1(new_n464), .C2(new_n445), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT74), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n483), .A2(new_n489), .A3(new_n361), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g305(.A1(new_n491), .A2(G472), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n468), .A2(new_n473), .A3(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n392), .B1(new_n361), .B2(G234), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n313), .A2(new_n315), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n209), .A2(G128), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n497), .B1(KEYINPUT75), .B2(KEYINPUT23), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n209), .A2(G128), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n499), .A2(KEYINPUT23), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT75), .ZN(new_n501));
  OAI21_X1  g315(.A(new_n501), .B1(new_n209), .B2(G128), .ZN(new_n502));
  OAI21_X1  g316(.A(new_n498), .B1(new_n500), .B2(new_n502), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n503), .A2(G110), .ZN(new_n504));
  INV_X1    g318(.A(new_n497), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n505), .A2(new_n499), .ZN(new_n506));
  XOR2_X1   g320(.A(KEYINPUT24), .B(G110), .Z(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n496), .A2(new_n504), .A3(new_n508), .ZN(new_n509));
  OAI22_X1  g323(.A1(new_n503), .A2(G110), .B1(new_n506), .B2(new_n507), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(new_n315), .A3(new_n319), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n205), .A2(G221), .A3(G234), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n513), .B(KEYINPUT22), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(G137), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n515), .B1(new_n509), .B2(new_n511), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT25), .ZN(new_n520));
  NOR3_X1   g334(.A1(new_n519), .A2(new_n520), .A3(new_n360), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n520), .B1(new_n519), .B2(new_n360), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n495), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NOR2_X1   g338(.A1(new_n517), .A2(new_n518), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n495), .A2(new_n282), .ZN(new_n526));
  XNOR2_X1  g340(.A(new_n526), .B(KEYINPUT76), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n525), .A2(new_n527), .ZN(new_n528));
  XOR2_X1   g342(.A(new_n528), .B(KEYINPUT77), .Z(new_n529));
  NOR2_X1   g343(.A1(new_n524), .A2(new_n529), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n493), .A2(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G469), .ZN(new_n532));
  OAI211_X1 g346(.A(new_n225), .B(new_n228), .C1(new_n416), .C2(new_n417), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT78), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n203), .A2(KEYINPUT78), .A3(new_n225), .A4(new_n228), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  INV_X1    g351(.A(KEYINPUT10), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(new_n426), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n250), .A2(new_n427), .A3(new_n252), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n434), .A2(KEYINPUT10), .A3(new_n230), .ZN(new_n542));
  NAND4_X1  g356(.A1(new_n539), .A2(new_n540), .A3(new_n541), .A4(new_n542), .ZN(new_n543));
  XNOR2_X1  g357(.A(G110), .B(G140), .ZN(new_n544));
  INV_X1    g358(.A(G227), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n545), .A2(G953), .ZN(new_n546));
  XOR2_X1   g360(.A(new_n544), .B(new_n546), .Z(new_n547));
  AND3_X1   g361(.A1(new_n543), .A2(KEYINPUT81), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g362(.A(KEYINPUT81), .B1(new_n543), .B2(new_n547), .ZN(new_n549));
  AOI21_X1  g363(.A(KEYINPUT12), .B1(new_n426), .B2(KEYINPUT79), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(new_n203), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(new_n229), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n551), .B1(new_n554), .B2(new_n426), .ZN(new_n555));
  AOI22_X1  g369(.A1(new_n535), .A2(new_n536), .B1(new_n552), .B2(new_n229), .ZN(new_n556));
  NOR3_X1   g370(.A1(new_n556), .A2(new_n540), .A3(new_n550), .ZN(new_n557));
  NOR2_X1   g371(.A1(new_n555), .A2(new_n557), .ZN(new_n558));
  NOR3_X1   g372(.A1(new_n548), .A2(new_n549), .A3(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n539), .A2(new_n541), .A3(new_n542), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(new_n426), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n547), .B1(new_n561), .B2(new_n543), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n532), .B(new_n361), .C1(new_n559), .C2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n543), .B1(new_n555), .B2(new_n557), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT80), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n547), .ZN(new_n567));
  OAI211_X1 g381(.A(KEYINPUT80), .B(new_n543), .C1(new_n555), .C2(new_n557), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n561), .A2(new_n547), .A3(new_n543), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n569), .A2(G469), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n532), .A2(new_n282), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n563), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(G221), .B1(new_n391), .B2(G902), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n403), .A2(new_n531), .A3(new_n576), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(G101), .ZN(G3));
  INV_X1    g392(.A(KEYINPUT97), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n290), .A2(new_n292), .ZN(new_n580));
  AOI21_X1  g394(.A(new_n579), .B1(new_n580), .B2(new_n187), .ZN(new_n581));
  INV_X1    g395(.A(new_n187), .ZN(new_n582));
  AOI211_X1 g396(.A(KEYINPUT97), .B(new_n582), .C1(new_n290), .C2(new_n292), .ZN(new_n583));
  NOR3_X1   g397(.A1(new_n581), .A2(new_n583), .A3(new_n365), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n471), .A2(new_n472), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n466), .A2(new_n361), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n586), .B1(new_n587), .B2(G472), .ZN(new_n588));
  NAND4_X1  g402(.A1(new_n588), .A2(KEYINPUT96), .A3(new_n530), .A4(new_n576), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n466), .A2(new_n467), .ZN(new_n590));
  OAI21_X1  g404(.A(G472), .B1(new_n471), .B2(new_n360), .ZN(new_n591));
  NAND4_X1  g405(.A1(new_n576), .A2(new_n590), .A3(new_n530), .A4(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT96), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  NOR2_X1   g409(.A1(new_n396), .A2(G478), .ZN(new_n596));
  INV_X1    g410(.A(KEYINPUT33), .ZN(new_n597));
  INV_X1    g411(.A(new_n393), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(KEYINPUT98), .ZN(new_n599));
  INV_X1    g413(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n600), .B1(new_n394), .B2(new_n395), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n384), .A2(new_n389), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n598), .ZN(new_n603));
  NAND3_X1  g417(.A1(new_n384), .A2(new_n389), .A3(new_n393), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n603), .A2(new_n604), .A3(new_n599), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n601), .A2(new_n605), .A3(new_n361), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n596), .B1(new_n606), .B2(G478), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n354), .A2(new_n607), .ZN(new_n608));
  NOR3_X1   g422(.A1(new_n585), .A2(new_n595), .A3(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT99), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n609), .A2(new_n610), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g428(.A(new_n614), .B(KEYINPUT34), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(new_n218), .ZN(G6));
  INV_X1    g430(.A(new_n401), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n585), .A2(new_n595), .A3(new_n617), .A4(new_n354), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  INV_X1    g434(.A(new_n523), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n494), .B1(new_n621), .B2(new_n521), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n623), .B(new_n512), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(new_n527), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n622), .A2(new_n625), .ZN(new_n626));
  NAND4_X1  g440(.A1(new_n403), .A2(new_n576), .A3(new_n588), .A4(new_n626), .ZN(new_n627));
  XOR2_X1   g441(.A(new_n627), .B(KEYINPUT37), .Z(new_n628));
  XNOR2_X1  g442(.A(new_n628), .B(G110), .ZN(G12));
  NOR2_X1   g443(.A1(new_n581), .A2(new_n583), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n354), .A2(new_n617), .ZN(new_n631));
  INV_X1    g445(.A(G900), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n359), .B1(new_n362), .B2(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n631), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(new_n635), .B(KEYINPUT100), .ZN(new_n636));
  AND2_X1   g450(.A1(new_n493), .A2(new_n626), .ZN(new_n637));
  NAND4_X1  g451(.A1(new_n630), .A2(new_n576), .A3(new_n636), .A4(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(G128), .ZN(G30));
  INV_X1    g453(.A(KEYINPUT38), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT101), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n293), .A2(new_n641), .A3(new_n294), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n641), .B1(new_n293), .B2(new_n294), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n293), .A2(new_n294), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n646), .A2(KEYINPUT101), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n647), .A2(KEYINPUT38), .A3(new_n642), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n645), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n448), .A2(new_n450), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n479), .A2(new_n462), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n652), .A2(new_n446), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n282), .B1(new_n651), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n654), .A2(G472), .ZN(new_n655));
  NAND3_X1  g469(.A1(new_n468), .A2(new_n473), .A3(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(new_n633), .B(KEYINPUT39), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n576), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g473(.A(new_n659), .B(KEYINPUT40), .Z(new_n660));
  AND3_X1   g474(.A1(new_n349), .A2(new_n351), .A3(new_n353), .ZN(new_n661));
  NOR2_X1   g475(.A1(new_n661), .A2(new_n617), .ZN(new_n662));
  INV_X1    g476(.A(new_n626), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n662), .A2(new_n663), .A3(new_n187), .ZN(new_n664));
  XOR2_X1   g478(.A(new_n664), .B(KEYINPUT102), .Z(new_n665));
  NAND4_X1  g479(.A1(new_n649), .A2(new_n656), .A3(new_n660), .A4(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G143), .ZN(G45));
  NOR2_X1   g481(.A1(new_n608), .A2(new_n633), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n630), .A2(new_n576), .A3(new_n637), .A4(new_n668), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n669), .B(G146), .ZN(G48));
  INV_X1    g484(.A(new_n559), .ZN(new_n671));
  INV_X1    g485(.A(new_n562), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n532), .B1(new_n673), .B2(new_n361), .ZN(new_n674));
  INV_X1    g488(.A(new_n563), .ZN(new_n675));
  INV_X1    g489(.A(new_n575), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n493), .A2(new_n530), .A3(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n365), .ZN(new_n679));
  INV_X1    g493(.A(new_n608), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n630), .A2(new_n678), .A3(new_n679), .A4(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(KEYINPUT41), .B(G113), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(KEYINPUT103), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n681), .B(new_n683), .ZN(G15));
  NAND4_X1  g498(.A1(new_n630), .A2(new_n678), .A3(new_n679), .A4(new_n631), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(G116), .ZN(G18));
  NAND4_X1  g500(.A1(new_n630), .A2(new_n402), .A3(new_n637), .A4(new_n677), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G119), .ZN(G21));
  AND3_X1   g502(.A1(new_n475), .A2(new_n480), .A3(new_n478), .ZN(new_n689));
  OAI21_X1  g503(.A(new_n454), .B1(new_n446), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(new_n467), .ZN(new_n691));
  AND4_X1   g505(.A1(new_n530), .A2(new_n677), .A3(new_n591), .A4(new_n691), .ZN(new_n692));
  NAND4_X1  g506(.A1(new_n630), .A2(new_n679), .A3(new_n662), .A4(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G122), .ZN(G24));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n591), .ZN(new_n695));
  NOR2_X1   g509(.A1(new_n695), .A2(new_n663), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT104), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n697), .B1(new_n608), .B2(new_n633), .ZN(new_n698));
  NAND4_X1  g512(.A1(new_n354), .A2(new_n607), .A3(KEYINPUT104), .A4(new_n634), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n630), .A2(new_n677), .A3(new_n696), .A4(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G125), .ZN(G27));
  INV_X1    g516(.A(KEYINPUT42), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n646), .A2(new_n700), .A3(new_n576), .A4(new_n187), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n493), .A2(new_n530), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n574), .A2(new_n575), .ZN(new_n707));
  AOI211_X1 g521(.A(new_n707), .B(new_n582), .C1(new_n293), .C2(new_n294), .ZN(new_n708));
  NAND4_X1  g522(.A1(new_n708), .A2(new_n531), .A3(KEYINPUT42), .A4(new_n700), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(G131), .ZN(G33));
  NAND4_X1  g525(.A1(new_n646), .A2(new_n493), .A3(new_n576), .A4(new_n187), .ZN(new_n712));
  INV_X1    g526(.A(new_n530), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT100), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n635), .B(new_n714), .ZN(new_n715));
  NOR3_X1   g529(.A1(new_n712), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n405), .ZN(G36));
  NAND3_X1  g531(.A1(new_n569), .A2(KEYINPUT45), .A3(new_n570), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT105), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n569), .A2(KEYINPUT105), .A3(KEYINPUT45), .A4(new_n570), .ZN(new_n721));
  AOI21_X1  g535(.A(new_n532), .B1(new_n720), .B2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT45), .B1(new_n569), .B2(new_n570), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n572), .B1(new_n722), .B2(new_n724), .ZN(new_n725));
  OAI21_X1  g539(.A(KEYINPUT106), .B1(new_n725), .B2(KEYINPUT46), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n725), .A2(KEYINPUT46), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT106), .ZN(new_n728));
  INV_X1    g542(.A(KEYINPUT46), .ZN(new_n729));
  AOI211_X1 g543(.A(new_n532), .B(new_n723), .C1(new_n720), .C2(new_n721), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n728), .B(new_n729), .C1(new_n730), .C2(new_n572), .ZN(new_n731));
  NAND4_X1  g545(.A1(new_n726), .A2(new_n563), .A3(new_n727), .A4(new_n731), .ZN(new_n732));
  NAND3_X1  g546(.A1(new_n732), .A2(new_n575), .A3(new_n658), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT107), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g549(.A(new_n588), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n661), .A2(new_n607), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT43), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n737), .B(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n736), .A2(new_n739), .A3(new_n626), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT44), .ZN(new_n741));
  AND2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n582), .B1(new_n293), .B2(new_n294), .ZN(new_n743));
  OAI21_X1  g557(.A(new_n743), .B1(new_n740), .B2(new_n741), .ZN(new_n744));
  NOR2_X1   g558(.A1(new_n742), .A2(new_n744), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n732), .A2(KEYINPUT107), .A3(new_n575), .A4(new_n658), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n735), .A2(new_n745), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G137), .ZN(G39));
  NOR2_X1   g562(.A1(new_n493), .A2(new_n530), .ZN(new_n749));
  AND3_X1   g563(.A1(new_n749), .A2(new_n668), .A3(new_n743), .ZN(new_n750));
  XNOR2_X1  g564(.A(KEYINPUT108), .B(KEYINPUT47), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n732), .A2(new_n575), .A3(new_n751), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n732), .B2(new_n575), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n750), .B1(new_n752), .B2(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  INV_X1    g569(.A(new_n743), .ZN(new_n756));
  INV_X1    g570(.A(new_n677), .ZN(new_n757));
  NOR2_X1   g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g572(.A1(new_n737), .A2(new_n738), .ZN(new_n759));
  AOI21_X1  g573(.A(KEYINPUT43), .B1(new_n661), .B2(new_n607), .ZN(new_n760));
  OAI21_X1  g574(.A(new_n359), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n761), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n531), .A3(new_n762), .ZN(new_n763));
  XNOR2_X1  g577(.A(new_n763), .B(KEYINPUT48), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n530), .A2(new_n359), .ZN(new_n765));
  NOR4_X1   g579(.A1(new_n756), .A2(new_n656), .A3(new_n757), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n358), .B1(new_n766), .B2(new_n680), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n764), .A2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n758), .A2(new_n696), .A3(new_n762), .ZN(new_n769));
  INV_X1    g583(.A(new_n607), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n661), .A3(new_n770), .ZN(new_n771));
  NOR4_X1   g585(.A1(new_n761), .A2(new_n713), .A3(new_n757), .A4(new_n695), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n772), .A2(new_n645), .A3(new_n582), .A4(new_n648), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT50), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  OAI211_X1 g590(.A(new_n769), .B(new_n771), .C1(new_n775), .C2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT115), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NOR2_X1   g593(.A1(new_n752), .A2(new_n753), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n674), .A2(new_n675), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n780), .B1(new_n575), .B2(new_n782), .ZN(new_n783));
  NOR4_X1   g597(.A1(new_n756), .A2(new_n761), .A3(new_n713), .A4(new_n695), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(KEYINPUT114), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n773), .B(new_n774), .ZN(new_n787));
  NAND4_X1  g601(.A1(new_n787), .A2(KEYINPUT115), .A3(new_n769), .A4(new_n771), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n779), .A2(new_n786), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n768), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n681), .A2(new_n685), .A3(new_n687), .ZN(new_n792));
  INV_X1    g606(.A(KEYINPUT109), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n793), .B1(new_n354), .B2(new_n617), .ZN(new_n794));
  AOI21_X1  g608(.A(KEYINPUT20), .B1(new_n352), .B2(new_n282), .ZN(new_n795));
  AOI22_X1  g609(.A1(new_n330), .A2(new_n332), .B1(new_n343), .B2(new_n329), .ZN(new_n796));
  NOR4_X1   g610(.A1(new_n796), .A2(new_n348), .A3(G475), .A4(G902), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT109), .A3(new_n401), .A4(new_n351), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n794), .A2(new_n608), .A3(new_n799), .ZN(new_n800));
  AND4_X1   g614(.A1(new_n187), .A2(new_n293), .A3(new_n800), .A4(new_n294), .ZN(new_n801));
  NAND4_X1  g615(.A1(new_n801), .A2(new_n589), .A3(new_n594), .A4(new_n679), .ZN(new_n802));
  AND3_X1   g616(.A1(new_n802), .A2(new_n627), .A3(new_n577), .ZN(new_n803));
  NAND4_X1  g617(.A1(new_n792), .A2(new_n693), .A3(new_n710), .A4(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(new_n712), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT110), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n354), .A2(new_n401), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n807), .A2(new_n634), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n805), .A2(new_n806), .A3(new_n626), .A4(new_n809), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n743), .A2(new_n493), .A3(new_n576), .A4(new_n626), .ZN(new_n811));
  OAI21_X1  g625(.A(KEYINPUT110), .B1(new_n811), .B2(new_n808), .ZN(new_n812));
  AOI21_X1  g626(.A(new_n716), .B1(new_n810), .B2(new_n812), .ZN(new_n813));
  NOR3_X1   g627(.A1(new_n704), .A2(new_n663), .A3(new_n695), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n804), .A2(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT53), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT111), .ZN(new_n819));
  OAI21_X1  g633(.A(new_n819), .B1(new_n626), .B2(new_n633), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n622), .A2(KEYINPUT111), .A3(new_n625), .A4(new_n634), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AND3_X1   g636(.A1(new_n822), .A2(new_n656), .A3(new_n576), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n630), .A2(new_n823), .A3(new_n662), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n638), .A2(new_n669), .A3(new_n701), .A4(new_n824), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n825), .A2(KEYINPUT52), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n493), .A2(new_n626), .ZN(new_n827));
  NOR3_X1   g641(.A1(new_n827), .A2(new_n581), .A3(new_n583), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n828), .B(new_n576), .C1(new_n636), .C2(new_n668), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT52), .ZN(new_n830));
  NAND4_X1  g644(.A1(new_n829), .A2(new_n830), .A3(new_n701), .A4(new_n824), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT112), .B1(new_n826), .B2(new_n831), .ZN(new_n833));
  OAI211_X1 g647(.A(new_n817), .B(new_n818), .C1(new_n832), .C2(new_n833), .ZN(new_n834));
  AOI211_X1 g648(.A(new_n716), .B(new_n814), .C1(new_n810), .C2(new_n812), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n681), .A2(new_n685), .A3(new_n687), .A4(new_n693), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n802), .A2(new_n627), .A3(new_n577), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(new_n838), .A3(new_n710), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n831), .ZN(new_n840));
  OAI21_X1  g654(.A(KEYINPUT53), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n834), .A2(KEYINPUT54), .A3(new_n841), .ZN(new_n842));
  NAND2_X1  g656(.A1(new_n836), .A2(KEYINPUT113), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n706), .A2(new_n709), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n802), .A2(new_n627), .A3(new_n577), .A4(KEYINPUT53), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n584), .B(new_n678), .C1(new_n680), .C2(new_n631), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT113), .ZN(new_n848));
  NAND4_X1  g662(.A1(new_n847), .A2(new_n848), .A3(new_n687), .A4(new_n693), .ZN(new_n849));
  AND3_X1   g663(.A1(new_n843), .A2(new_n846), .A3(new_n849), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n850), .B(new_n835), .C1(new_n832), .C2(new_n833), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT54), .ZN(new_n852));
  OAI21_X1  g666(.A(new_n818), .B1(new_n839), .B2(new_n840), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n851), .A2(new_n852), .A3(new_n853), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n783), .A2(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n783), .A2(KEYINPUT116), .ZN(new_n856));
  NAND3_X1  g670(.A1(new_n855), .A2(new_n785), .A3(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n777), .A2(new_n790), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n791), .A2(new_n842), .A3(new_n854), .A4(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n772), .A2(new_n630), .ZN(new_n861));
  OAI22_X1  g675(.A1(new_n860), .A2(new_n861), .B1(G952), .B2(G953), .ZN(new_n862));
  OR2_X1    g676(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n782), .A2(KEYINPUT49), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n713), .A2(new_n582), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n863), .A2(new_n864), .A3(new_n575), .A4(new_n865), .ZN(new_n866));
  OR4_X1    g680(.A1(new_n656), .A2(new_n649), .A3(new_n737), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n862), .A2(new_n867), .ZN(G75));
  AOI21_X1  g682(.A(new_n361), .B1(new_n851), .B2(new_n853), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n289), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT56), .ZN(new_n871));
  INV_X1    g685(.A(new_n265), .ZN(new_n872));
  INV_X1    g686(.A(new_n268), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n257), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n874), .B(new_n207), .ZN(new_n875));
  XNOR2_X1  g689(.A(new_n875), .B(KEYINPUT55), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(KEYINPUT117), .B2(new_n871), .ZN(new_n877));
  AND3_X1   g691(.A1(new_n870), .A2(new_n871), .A3(new_n877), .ZN(new_n878));
  AOI21_X1  g692(.A(new_n877), .B1(new_n870), .B2(new_n871), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n205), .A2(G952), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(G51));
  XNOR2_X1  g695(.A(new_n572), .B(KEYINPUT57), .ZN(new_n882));
  INV_X1    g696(.A(new_n854), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n852), .B1(new_n851), .B2(new_n853), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n885), .A2(new_n673), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n869), .A2(new_n730), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n880), .B1(new_n886), .B2(new_n887), .ZN(G54));
  AND2_X1   g702(.A1(KEYINPUT58), .A2(G475), .ZN(new_n889));
  NAND4_X1  g703(.A1(new_n835), .A2(new_n843), .A3(new_n849), .A4(new_n846), .ZN(new_n890));
  NAND3_X1  g704(.A1(new_n826), .A2(KEYINPUT112), .A3(new_n831), .ZN(new_n891));
  INV_X1    g705(.A(KEYINPUT112), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n840), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n890), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(new_n840), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT53), .B1(new_n817), .B2(new_n895), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n360), .B(new_n889), .C1(new_n894), .C2(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n897), .A2(new_n796), .ZN(new_n898));
  INV_X1    g712(.A(new_n880), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n851), .A2(new_n853), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(new_n360), .A3(new_n345), .A4(new_n889), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n898), .A2(new_n899), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT118), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND4_X1  g718(.A1(new_n898), .A2(KEYINPUT118), .A3(new_n901), .A4(new_n899), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(G60));
  NAND2_X1  g720(.A1(new_n601), .A2(new_n605), .ZN(new_n907));
  XNOR2_X1  g721(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n908));
  NAND2_X1  g722(.A1(G478), .A2(G902), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n884), .ZN(new_n911));
  AOI211_X1 g725(.A(new_n907), .B(new_n910), .C1(new_n911), .C2(new_n854), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n910), .B1(new_n854), .B2(new_n842), .ZN(new_n913));
  INV_X1    g727(.A(new_n907), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n899), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  NAND2_X1  g730(.A1(G217), .A2(G902), .ZN(new_n917));
  XOR2_X1   g731(.A(new_n917), .B(KEYINPUT120), .Z(new_n918));
  XOR2_X1   g732(.A(new_n918), .B(KEYINPUT60), .Z(new_n919));
  OAI211_X1 g733(.A(new_n624), .B(new_n919), .C1(new_n894), .C2(new_n896), .ZN(new_n920));
  INV_X1    g734(.A(new_n919), .ZN(new_n921));
  AOI21_X1  g735(.A(new_n921), .B1(new_n851), .B2(new_n853), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n920), .B(new_n899), .C1(new_n922), .C2(new_n525), .ZN(new_n923));
  INV_X1    g737(.A(KEYINPUT61), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT121), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n925), .B(new_n899), .C1(new_n922), .C2(new_n525), .ZN(new_n926));
  NAND3_X1  g740(.A1(new_n923), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n919), .B1(new_n894), .B2(new_n896), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n880), .B1(new_n928), .B2(new_n519), .ZN(new_n929));
  OAI211_X1 g743(.A(new_n929), .B(new_n920), .C1(new_n925), .C2(KEYINPUT61), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n927), .A2(new_n930), .ZN(G66));
  NOR2_X1   g745(.A1(new_n838), .A2(G953), .ZN(new_n932));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n205), .B1(new_n363), .B2(G224), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n935), .B1(new_n933), .B2(new_n934), .ZN(new_n936));
  INV_X1    g750(.A(new_n874), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n937), .B1(G898), .B2(new_n205), .ZN(new_n938));
  XNOR2_X1  g752(.A(new_n936), .B(new_n938), .ZN(G69));
  NAND3_X1  g753(.A1(new_n638), .A2(new_n669), .A3(new_n701), .ZN(new_n940));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n829), .A2(KEYINPUT124), .A3(new_n701), .ZN(new_n943));
  NAND3_X1  g757(.A1(new_n942), .A2(new_n666), .A3(new_n943), .ZN(new_n944));
  INV_X1    g758(.A(KEYINPUT62), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n944), .A2(new_n945), .ZN(new_n946));
  NAND4_X1  g760(.A1(new_n942), .A2(KEYINPUT62), .A3(new_n943), .A4(new_n666), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n747), .A2(new_n754), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n756), .A2(new_n659), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n950), .A2(new_n531), .A3(new_n800), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n948), .A2(new_n949), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n205), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n432), .A2(new_n438), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(new_n339), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n955), .B(KEYINPUT123), .ZN(new_n956));
  NAND2_X1  g770(.A1(G900), .A2(G953), .ZN(new_n957));
  NAND3_X1  g771(.A1(new_n747), .A2(new_n942), .A3(new_n943), .ZN(new_n958));
  AND3_X1   g772(.A1(new_n630), .A2(new_n531), .A3(new_n662), .ZN(new_n959));
  NAND3_X1  g773(.A1(new_n735), .A2(new_n746), .A3(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n716), .B1(new_n706), .B2(new_n709), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(new_n754), .A3(new_n961), .ZN(new_n962));
  NOR2_X1   g776(.A1(new_n958), .A2(new_n962), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n955), .B1(new_n963), .B2(new_n205), .ZN(new_n964));
  AOI22_X1  g778(.A1(new_n953), .A2(new_n956), .B1(new_n957), .B2(new_n964), .ZN(new_n965));
  OAI21_X1  g779(.A(G953), .B1(new_n545), .B2(new_n632), .ZN(new_n966));
  XNOR2_X1  g780(.A(new_n965), .B(new_n966), .ZN(G72));
  NAND2_X1  g781(.A1(G472), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT63), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n650), .B2(new_n487), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n834), .A2(new_n841), .A3(new_n971), .ZN(new_n972));
  NAND3_X1  g786(.A1(new_n439), .A2(new_n440), .A3(new_n445), .ZN(new_n973));
  AND3_X1   g787(.A1(new_n747), .A2(new_n942), .A3(new_n943), .ZN(new_n974));
  AND3_X1   g788(.A1(new_n960), .A2(new_n754), .A3(new_n961), .ZN(new_n975));
  NAND3_X1  g789(.A1(new_n974), .A2(new_n975), .A3(new_n838), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n973), .B1(new_n976), .B2(new_n969), .ZN(new_n977));
  OAI21_X1  g791(.A(KEYINPUT126), .B1(new_n977), .B2(new_n880), .ZN(new_n978));
  INV_X1    g792(.A(KEYINPUT126), .ZN(new_n979));
  AOI21_X1  g793(.A(new_n970), .B1(new_n963), .B2(new_n838), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n979), .B(new_n899), .C1(new_n980), .C2(new_n973), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n972), .B1(new_n978), .B2(new_n981), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n948), .A2(new_n838), .A3(new_n949), .A4(new_n951), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n969), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n984), .A2(new_n446), .A3(new_n486), .ZN(new_n985));
  NAND2_X1  g799(.A1(new_n985), .A2(KEYINPUT125), .ZN(new_n986));
  INV_X1    g800(.A(KEYINPUT125), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n984), .A2(new_n987), .A3(new_n446), .A4(new_n486), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n982), .A2(new_n986), .A3(new_n988), .ZN(G57));
endmodule


