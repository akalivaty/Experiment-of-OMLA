//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  NOR2_X1   g0004(.A1(G97), .A2(G107), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n206), .A2(G87), .ZN(G355));
  NAND2_X1  g0007(.A1(G1), .A2(G20), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT64), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XOR2_X1   g0011(.A(new_n211), .B(KEYINPUT0), .Z(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(G20), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR3_X1   g0015(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT65), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND3_X1  g0021(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n209), .B1(new_n218), .B2(new_n222), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT1), .ZN(new_n224));
  NOR3_X1   g0024(.A1(new_n212), .A2(new_n216), .A3(new_n224), .ZN(G361));
  XNOR2_X1  g0025(.A(G250), .B(G257), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(KEYINPUT66), .ZN(new_n227));
  XOR2_X1   g0027(.A(G264), .B(G270), .Z(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XOR2_X1   g0031(.A(KEYINPUT2), .B(G226), .Z(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n229), .B(new_n233), .ZN(G358));
  XOR2_X1   g0034(.A(G87), .B(G97), .Z(new_n235));
  XNOR2_X1  g0035(.A(G107), .B(G116), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  NAND2_X1  g0037(.A1(new_n202), .A2(G68), .ZN(new_n238));
  INV_X1    g0038(.A(G68), .ZN(new_n239));
  NAND2_X1  g0039(.A1(new_n239), .A2(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n238), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(G58), .B(G77), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n237), .B(new_n243), .ZN(G351));
  INV_X1    g0044(.A(G58), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n245), .A2(KEYINPUT8), .ZN(new_n246));
  INV_X1    g0046(.A(KEYINPUT8), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n247), .A2(G58), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n246), .A2(new_n248), .ZN(new_n249));
  INV_X1    g0049(.A(G33), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(G20), .ZN(new_n251));
  NOR2_X1   g0051(.A1(G20), .A2(G33), .ZN(new_n252));
  AOI22_X1  g0052(.A1(new_n249), .A2(new_n251), .B1(G150), .B2(new_n252), .ZN(new_n253));
  AOI22_X1  g0053(.A1(new_n253), .A2(KEYINPUT68), .B1(G20), .B2(new_n203), .ZN(new_n254));
  OAI21_X1  g0054(.A(new_n254), .B1(KEYINPUT68), .B2(new_n253), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n215), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(new_n256), .A2(new_n215), .ZN(new_n259));
  INV_X1    g0059(.A(G1), .ZN(new_n260));
  NAND3_X1  g0060(.A1(new_n260), .A2(G13), .A3(G20), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n260), .A2(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G50), .ZN(new_n264));
  OAI22_X1  g0064(.A1(new_n262), .A2(new_n264), .B1(G50), .B2(new_n261), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT69), .ZN(new_n266));
  XNOR2_X1  g0066(.A(new_n265), .B(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(new_n258), .A2(new_n267), .ZN(new_n268));
  XNOR2_X1  g0068(.A(new_n268), .B(KEYINPUT72), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT9), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT72), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n268), .B(new_n272), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n273), .A2(KEYINPUT9), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  AND2_X1   g0075(.A1(G1), .A2(G13), .ZN(new_n276));
  NAND2_X1  g0076(.A1(G33), .A2(G41), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(G41), .A2(G45), .ZN(new_n279));
  NOR2_X1   g0079(.A1(new_n279), .A2(G1), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n278), .A2(new_n280), .ZN(new_n281));
  INV_X1    g0081(.A(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT67), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n283), .B1(new_n279), .B2(G1), .ZN(new_n284));
  NAND3_X1  g0084(.A1(new_n277), .A2(G1), .A3(G13), .ZN(new_n285));
  OAI211_X1 g0085(.A(new_n260), .B(KEYINPUT67), .C1(G41), .C2(G45), .ZN(new_n286));
  AND3_X1   g0086(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n282), .B1(new_n287), .B2(G226), .ZN(new_n288));
  INV_X1    g0088(.A(G1698), .ZN(new_n289));
  OR2_X1    g0089(.A1(KEYINPUT3), .A2(G33), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NOR2_X1   g0093(.A1(KEYINPUT3), .A2(G33), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n292), .A2(G223), .B1(new_n295), .B2(G77), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n290), .A2(new_n291), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(G222), .A3(new_n289), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n288), .B1(new_n299), .B2(new_n285), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  INV_X1    g0101(.A(KEYINPUT10), .ZN(new_n302));
  OAI22_X1  g0102(.A1(new_n300), .A2(new_n301), .B1(KEYINPUT73), .B2(new_n302), .ZN(new_n303));
  AOI21_X1  g0103(.A(new_n303), .B1(G200), .B2(new_n300), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n271), .A2(new_n274), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  NAND4_X1  g0108(.A1(new_n271), .A2(new_n274), .A3(new_n306), .A4(new_n304), .ZN(new_n309));
  INV_X1    g0109(.A(G169), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n300), .A2(new_n310), .ZN(new_n311));
  OAI211_X1 g0111(.A(new_n268), .B(new_n311), .C1(G179), .C2(new_n300), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n308), .A2(new_n309), .A3(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n282), .B1(new_n287), .B2(G238), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n297), .A2(G232), .A3(G1698), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n297), .A2(G226), .A3(new_n289), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G33), .A2(G97), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n285), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n314), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n321), .A2(KEYINPUT13), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT13), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n314), .A2(new_n320), .A3(new_n323), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n322), .A2(G190), .A3(new_n324), .ZN(new_n325));
  AOI22_X1  g0125(.A1(new_n252), .A2(G50), .B1(G20), .B2(new_n239), .ZN(new_n326));
  INV_X1    g0126(.A(new_n251), .ZN(new_n327));
  INV_X1    g0127(.A(G77), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AND2_X1   g0129(.A1(new_n329), .A2(new_n257), .ZN(new_n330));
  OR2_X1    g0130(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n331));
  INV_X1    g0131(.A(new_n331), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n330), .A2(KEYINPUT11), .ZN(new_n333));
  INV_X1    g0133(.A(new_n261), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n334), .A2(new_n239), .ZN(new_n335));
  XNOR2_X1  g0135(.A(new_n335), .B(KEYINPUT12), .ZN(new_n336));
  NOR2_X1   g0136(.A1(new_n334), .A2(new_n257), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n337), .A2(G68), .A3(new_n263), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n333), .A2(new_n336), .A3(new_n338), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n332), .A2(new_n339), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n325), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n322), .A2(new_n324), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n342), .A2(G200), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n341), .A2(KEYINPUT74), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(KEYINPUT74), .B1(new_n341), .B2(new_n343), .ZN(new_n345));
  OR2_X1    g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n340), .ZN(new_n347));
  INV_X1    g0147(.A(KEYINPUT14), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n342), .A2(new_n348), .A3(G169), .ZN(new_n349));
  INV_X1    g0149(.A(G179), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n349), .B1(new_n350), .B2(new_n342), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n348), .B1(new_n342), .B2(G169), .ZN(new_n352));
  OAI21_X1  g0152(.A(new_n347), .B1(new_n351), .B2(new_n352), .ZN(new_n353));
  AOI22_X1  g0153(.A1(new_n292), .A2(G238), .B1(new_n295), .B2(G107), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n297), .A2(G232), .A3(new_n289), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n319), .ZN(new_n357));
  AOI21_X1  g0157(.A(new_n282), .B1(new_n287), .B2(G244), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n359), .A2(G179), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n360), .B1(new_n310), .B2(new_n359), .ZN(new_n361));
  XNOR2_X1  g0161(.A(KEYINPUT15), .B(G87), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT70), .ZN(new_n363));
  OR2_X1    g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n363), .ZN(new_n365));
  AND2_X1   g0165(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n366), .A2(KEYINPUT71), .A3(new_n251), .ZN(new_n367));
  AOI22_X1  g0167(.A1(new_n249), .A2(new_n252), .B1(G20), .B2(G77), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(KEYINPUT71), .B1(new_n366), .B2(new_n251), .ZN(new_n370));
  OAI21_X1  g0170(.A(new_n257), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n328), .B1(new_n260), .B2(G20), .ZN(new_n372));
  AOI22_X1  g0172(.A1(new_n337), .A2(new_n372), .B1(new_n328), .B2(new_n334), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n361), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n374), .ZN(new_n376));
  NOR2_X1   g0176(.A1(new_n359), .A2(new_n301), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n377), .B1(G200), .B2(new_n359), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n376), .A2(new_n378), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n346), .A2(new_n353), .A3(new_n375), .A4(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n249), .A2(new_n263), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n262), .A2(new_n381), .B1(new_n249), .B2(new_n261), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NOR2_X1   g0183(.A1(new_n245), .A2(new_n239), .ZN(new_n384));
  OAI21_X1  g0184(.A(G20), .B1(new_n384), .B2(new_n201), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n252), .A2(G159), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(KEYINPUT16), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT75), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n290), .A2(new_n214), .A3(new_n291), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(KEYINPUT7), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n290), .A2(new_n393), .A3(new_n214), .A4(new_n291), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n390), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  NOR2_X1   g0195(.A1(KEYINPUT75), .A2(KEYINPUT7), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n239), .B1(new_n391), .B2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(new_n397), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n389), .B1(new_n395), .B2(new_n398), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n393), .B1(new_n295), .B2(new_n214), .ZN(new_n400));
  NOR4_X1   g0200(.A1(new_n293), .A2(new_n294), .A3(KEYINPUT7), .A4(G20), .ZN(new_n401));
  OAI21_X1  g0201(.A(KEYINPUT75), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NAND3_X1  g0202(.A1(new_n402), .A2(KEYINPUT76), .A3(new_n397), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n388), .B1(new_n399), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n392), .A2(G68), .A3(new_n394), .ZN(new_n405));
  AND2_X1   g0205(.A1(new_n405), .A2(new_n387), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n257), .B1(new_n406), .B2(KEYINPUT16), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n383), .B1(new_n404), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT77), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT77), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n383), .C1(new_n404), .C2(new_n407), .ZN(new_n411));
  NAND4_X1  g0211(.A1(new_n284), .A2(G232), .A3(new_n285), .A4(new_n286), .ZN(new_n412));
  AND2_X1   g0212(.A1(new_n412), .A2(new_n281), .ZN(new_n413));
  OAI211_X1 g0213(.A(G223), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n414));
  OAI211_X1 g0214(.A(G226), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n415));
  NAND2_X1  g0215(.A1(G33), .A2(G87), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(new_n319), .ZN(new_n418));
  AND2_X1   g0218(.A1(new_n413), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(G179), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n420), .B1(new_n310), .B2(new_n419), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n409), .A2(new_n411), .A3(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(KEYINPUT18), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT18), .ZN(new_n424));
  NAND4_X1  g0224(.A1(new_n409), .A2(new_n424), .A3(new_n411), .A4(new_n421), .ZN(new_n425));
  AND3_X1   g0225(.A1(new_n413), .A2(new_n418), .A3(G190), .ZN(new_n426));
  INV_X1    g0226(.A(G200), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n427), .B1(new_n413), .B2(new_n418), .ZN(new_n428));
  NOR2_X1   g0228(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  OAI211_X1 g0229(.A(new_n429), .B(new_n383), .C1(new_n404), .C2(new_n407), .ZN(new_n430));
  XNOR2_X1  g0230(.A(new_n430), .B(KEYINPUT17), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n423), .A2(new_n425), .A3(new_n431), .ZN(new_n432));
  NOR3_X1   g0232(.A1(new_n313), .A2(new_n380), .A3(new_n432), .ZN(new_n433));
  OAI211_X1 g0233(.A(G238), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n434));
  OAI211_X1 g0234(.A(G244), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n435));
  NAND2_X1  g0235(.A1(G33), .A2(G116), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n434), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT80), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n434), .A2(new_n435), .A3(KEYINPUT80), .A4(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n319), .ZN(new_n442));
  INV_X1    g0242(.A(G45), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n443), .A2(G1), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n278), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n260), .A2(G45), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n285), .A2(G250), .A3(new_n446), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n445), .A2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NAND3_X1  g0249(.A1(new_n442), .A2(G190), .A3(new_n449), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n285), .B1(new_n439), .B2(new_n440), .ZN(new_n451));
  OAI21_X1  g0251(.A(G200), .B1(new_n451), .B2(new_n448), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT19), .ZN(new_n453));
  INV_X1    g0253(.A(G97), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n453), .B1(new_n327), .B2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n297), .A2(new_n214), .A3(G68), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n214), .B1(new_n317), .B2(new_n453), .ZN(new_n457));
  OAI21_X1  g0257(.A(new_n457), .B1(G87), .B2(new_n206), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n455), .A2(new_n456), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(new_n257), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n364), .A2(new_n365), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(new_n334), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n260), .A2(G33), .ZN(new_n463));
  AND3_X1   g0263(.A1(new_n259), .A2(new_n261), .A3(new_n463), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n464), .A2(G87), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n460), .A2(new_n462), .A3(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n466), .ZN(new_n467));
  AND3_X1   g0267(.A1(new_n450), .A2(new_n452), .A3(new_n467), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n310), .B1(new_n451), .B2(new_n448), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n337), .A2(new_n463), .ZN(new_n470));
  OAI211_X1 g0270(.A(new_n460), .B(new_n462), .C1(new_n461), .C2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n448), .B1(new_n441), .B2(new_n319), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n473), .B1(new_n474), .B2(new_n350), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n472), .A2(new_n475), .ZN(new_n476));
  NAND3_X1  g0276(.A1(new_n474), .A2(new_n473), .A3(new_n350), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n468), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT6), .ZN(new_n480));
  AND2_X1   g0280(.A1(G97), .A2(G107), .ZN(new_n481));
  OAI21_X1  g0281(.A(new_n480), .B1(new_n481), .B2(new_n205), .ZN(new_n482));
  INV_X1    g0282(.A(G107), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n483), .A2(KEYINPUT6), .A3(G97), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n482), .A2(new_n484), .ZN(new_n485));
  AOI22_X1  g0285(.A1(new_n485), .A2(G20), .B1(G77), .B2(new_n252), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n392), .A2(G107), .A3(new_n394), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n257), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n261), .A2(G97), .ZN(new_n490));
  INV_X1    g0290(.A(new_n490), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(new_n470), .B2(new_n454), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  OAI211_X1 g0294(.A(G244), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n495));
  INV_X1    g0295(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n297), .A2(KEYINPUT4), .A3(G244), .A4(new_n289), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n297), .A2(G250), .A3(G1698), .ZN(new_n500));
  NAND4_X1  g0300(.A1(new_n497), .A2(new_n498), .A3(new_n499), .A4(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(new_n319), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT78), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n285), .A2(G274), .ZN(new_n504));
  NAND2_X1  g0304(.A1(KEYINPUT5), .A2(G41), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g0306(.A1(KEYINPUT5), .A2(G41), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n444), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n504), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT5), .ZN(new_n510));
  INV_X1    g0310(.A(G41), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n446), .B1(new_n512), .B2(new_n505), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n513), .A2(KEYINPUT78), .A3(new_n278), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n513), .A2(new_n319), .ZN(new_n515));
  AOI22_X1  g0315(.A1(new_n509), .A2(new_n514), .B1(new_n515), .B2(G257), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n502), .A2(new_n350), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n494), .A2(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(G169), .B1(new_n502), .B2(new_n516), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n479), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n502), .A2(new_n516), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n521), .A2(new_n310), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n522), .A2(new_n494), .A3(KEYINPUT79), .A4(new_n517), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n521), .A2(G200), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n492), .B1(new_n488), .B2(new_n257), .ZN(new_n525));
  OAI211_X1 g0325(.A(new_n524), .B(new_n525), .C1(new_n301), .C2(new_n521), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n520), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n261), .A2(G116), .ZN(new_n528));
  AOI21_X1  g0328(.A(new_n528), .B1(new_n464), .B2(G116), .ZN(new_n529));
  INV_X1    g0329(.A(G116), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n256), .A2(new_n215), .B1(G20), .B2(new_n530), .ZN(new_n531));
  OAI211_X1 g0331(.A(new_n499), .B(new_n214), .C1(G33), .C2(new_n454), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT20), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n531), .A2(KEYINPUT20), .A3(new_n532), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n529), .A2(new_n537), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n509), .A2(new_n514), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n515), .A2(G270), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n295), .A2(G303), .ZN(new_n541));
  OAI211_X1 g0341(.A(G257), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI211_X1 g0343(.A(G264), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT82), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n292), .A2(KEYINPUT82), .A3(G264), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  OAI211_X1 g0348(.A(new_n539), .B(new_n540), .C1(new_n548), .C2(new_n285), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n538), .B1(new_n549), .B2(G200), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n550), .B1(new_n301), .B2(new_n549), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n310), .B1(new_n529), .B2(new_n537), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(KEYINPUT21), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n547), .A2(new_n546), .ZN(new_n554));
  INV_X1    g0354(.A(new_n543), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n285), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n539), .A2(new_n540), .ZN(new_n558));
  INV_X1    g0358(.A(new_n558), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n557), .A2(new_n559), .A3(G179), .A4(new_n538), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n553), .A2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n556), .A2(new_n558), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n538), .A2(G169), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n562), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n551), .A2(new_n561), .A3(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G257), .B(G1698), .C1(new_n293), .C2(new_n294), .ZN(new_n567));
  OAI211_X1 g0367(.A(G250), .B(new_n289), .C1(new_n293), .C2(new_n294), .ZN(new_n568));
  INV_X1    g0368(.A(G294), .ZN(new_n569));
  OAI211_X1 g0369(.A(new_n567), .B(new_n568), .C1(new_n250), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n319), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n515), .A2(G264), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n571), .A2(new_n539), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g0373(.A1(new_n573), .A2(new_n350), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n570), .A2(KEYINPUT84), .A3(new_n319), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n575), .A2(new_n539), .A3(new_n572), .ZN(new_n576));
  AOI21_X1  g0376(.A(KEYINPUT84), .B1(new_n570), .B2(new_n319), .ZN(new_n577));
  OAI21_X1  g0377(.A(G169), .B1(new_n576), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  XNOR2_X1  g0379(.A(KEYINPUT83), .B(KEYINPUT22), .ZN(new_n580));
  NAND4_X1  g0380(.A1(new_n297), .A2(new_n580), .A3(new_n214), .A4(G87), .ZN(new_n581));
  OAI211_X1 g0381(.A(new_n214), .B(G87), .C1(new_n293), .C2(new_n294), .ZN(new_n582));
  XOR2_X1   g0382(.A(KEYINPUT83), .B(KEYINPUT22), .Z(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n436), .A2(G20), .ZN(new_n585));
  INV_X1    g0385(.A(KEYINPUT23), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n586), .B1(new_n214), .B2(G107), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n483), .A2(KEYINPUT23), .A3(G20), .ZN(new_n588));
  AOI21_X1  g0388(.A(new_n585), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n581), .A2(new_n584), .A3(new_n589), .ZN(new_n590));
  AND2_X1   g0390(.A1(new_n590), .A2(KEYINPUT24), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n590), .A2(KEYINPUT24), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n257), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT25), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n261), .B2(G107), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n334), .A2(KEYINPUT25), .A3(new_n483), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n464), .A2(G107), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n593), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n579), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n573), .A2(new_n427), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT84), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n571), .A2(new_n601), .ZN(new_n602));
  NAND4_X1  g0402(.A1(new_n602), .A2(new_n539), .A3(new_n575), .A4(new_n572), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n600), .B1(new_n603), .B2(G190), .ZN(new_n604));
  INV_X1    g0404(.A(new_n597), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n590), .B(KEYINPUT24), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n605), .B1(new_n606), .B2(new_n257), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n599), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n566), .A2(new_n609), .ZN(new_n610));
  AND4_X1   g0410(.A1(new_n433), .A2(new_n478), .A3(new_n527), .A4(new_n610), .ZN(G372));
  INV_X1    g0411(.A(new_n431), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n375), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n361), .A2(new_n374), .A3(KEYINPUT86), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n346), .A2(new_n614), .A3(new_n615), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n612), .B1(new_n616), .B2(new_n353), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n408), .A2(new_n421), .ZN(new_n618));
  XNOR2_X1  g0418(.A(new_n618), .B(KEYINPUT18), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n308), .B(new_n309), .C1(new_n617), .C2(new_n619), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n312), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n442), .A2(new_n350), .A3(new_n449), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n448), .A2(KEYINPUT85), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT85), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n445), .A2(new_n624), .A3(new_n447), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g0426(.A(new_n310), .B1(new_n451), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g0427(.A1(new_n622), .A2(new_n471), .A3(new_n627), .ZN(new_n628));
  AND3_X1   g0428(.A1(new_n522), .A2(new_n494), .A3(new_n517), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT26), .ZN(new_n630));
  OAI21_X1  g0430(.A(G200), .B1(new_n451), .B2(new_n626), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n450), .A2(new_n467), .A3(new_n631), .ZN(new_n632));
  NAND4_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n628), .A4(new_n632), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n565), .A2(new_n553), .A3(new_n560), .ZN(new_n634));
  AOI22_X1  g0434(.A1(new_n574), .A2(new_n578), .B1(new_n593), .B2(new_n597), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n608), .B(new_n632), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n520), .A2(new_n523), .A3(new_n526), .ZN(new_n637));
  OAI211_X1 g0437(.A(new_n628), .B(new_n633), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n520), .A2(new_n523), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n630), .B1(new_n478), .B2(new_n639), .ZN(new_n640));
  OR2_X1    g0440(.A1(new_n638), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n433), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n621), .A2(new_n642), .ZN(G369));
  NAND3_X1  g0443(.A1(new_n260), .A2(new_n214), .A3(G13), .ZN(new_n644));
  OR2_X1    g0444(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n644), .A2(KEYINPUT27), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n645), .A2(G213), .A3(new_n646), .ZN(new_n647));
  INV_X1    g0447(.A(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT87), .ZN(new_n649));
  OR2_X1    g0449(.A1(new_n649), .A2(G343), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(G343), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n648), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n634), .A2(new_n653), .ZN(new_n654));
  INV_X1    g0454(.A(new_n653), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n635), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g0456(.A(new_n656), .B(KEYINPUT88), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n599), .B(new_n608), .C1(new_n607), .C2(new_n653), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n654), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  NOR2_X1   g0459(.A1(new_n599), .A2(new_n655), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  AOI21_X1  g0461(.A(new_n653), .B1(new_n537), .B2(new_n529), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n634), .A2(new_n662), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n566), .B2(new_n662), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n664), .A2(G330), .ZN(new_n665));
  INV_X1    g0465(.A(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n657), .A2(new_n658), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n661), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g0469(.A(new_n669), .B(KEYINPUT89), .Z(G399));
  INV_X1    g0470(.A(new_n210), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n671), .A2(G41), .ZN(new_n672));
  NOR3_X1   g0472(.A1(new_n206), .A2(G87), .A3(G116), .ZN(new_n673));
  INV_X1    g0473(.A(new_n673), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n672), .A2(new_n260), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n213), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n672), .ZN(new_n677));
  XOR2_X1   g0477(.A(new_n677), .B(KEYINPUT28), .Z(new_n678));
  NAND4_X1  g0478(.A1(new_n610), .A2(new_n478), .A3(new_n527), .A4(new_n653), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n549), .A2(new_n350), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n502), .A2(new_n516), .A3(new_n571), .A4(new_n572), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n680), .A2(new_n681), .A3(new_n474), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT30), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n502), .A2(new_n516), .ZN(new_n685));
  NOR2_X1   g0485(.A1(new_n685), .A2(new_n563), .ZN(new_n686));
  OR2_X1    g0486(.A1(new_n451), .A2(new_n626), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n686), .A2(new_n350), .A3(new_n573), .A4(new_n687), .ZN(new_n688));
  NAND4_X1  g0488(.A1(new_n680), .A2(new_n681), .A3(KEYINPUT30), .A4(new_n474), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n684), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n690), .A2(new_n655), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT31), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n690), .A2(KEYINPUT31), .A3(new_n655), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n679), .A2(new_n693), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n695), .A2(G330), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  AND4_X1   g0497(.A1(KEYINPUT26), .A2(new_n629), .A3(new_n628), .A4(new_n632), .ZN(new_n698));
  INV_X1    g0498(.A(new_n468), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n622), .A2(KEYINPUT81), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n700), .A2(new_n477), .A3(new_n469), .A4(new_n471), .ZN(new_n701));
  AOI21_X1  g0501(.A(new_n525), .B1(new_n685), .B2(new_n350), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT79), .B1(new_n702), .B2(new_n522), .ZN(new_n703));
  INV_X1    g0503(.A(new_n523), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n699), .B(new_n701), .C1(new_n703), .C2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n698), .B1(new_n705), .B2(new_n630), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n628), .B1(new_n636), .B2(new_n637), .ZN(new_n707));
  OAI21_X1  g0507(.A(new_n653), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(KEYINPUT90), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  OAI211_X1 g0510(.A(KEYINPUT90), .B(new_n653), .C1(new_n706), .C2(new_n707), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n712), .A2(KEYINPUT29), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT29), .ZN(new_n714));
  INV_X1    g0514(.A(new_n641), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n655), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n697), .B1(new_n713), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n678), .B1(new_n717), .B2(G1), .ZN(G364));
  INV_X1    g0518(.A(G13), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n719), .A2(G20), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n720), .B(KEYINPUT91), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n721), .A2(G45), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n722), .A2(G1), .ZN(new_n723));
  NOR2_X1   g0523(.A1(new_n672), .A2(new_n723), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n666), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n725), .B1(G330), .B2(new_n664), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n210), .A2(new_n295), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n727), .B1(new_n443), .B2(new_n676), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n728), .B1(new_n443), .B2(new_n243), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n671), .A2(new_n295), .ZN(new_n730));
  INV_X1    g0530(.A(new_n730), .ZN(new_n731));
  XNOR2_X1  g0531(.A(G355), .B(KEYINPUT92), .ZN(new_n732));
  OAI221_X1 g0532(.A(new_n729), .B1(G116), .B2(new_n210), .C1(new_n731), .C2(new_n732), .ZN(new_n733));
  INV_X1    g0533(.A(KEYINPUT93), .ZN(new_n734));
  AND2_X1   g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n215), .B1(G20), .B2(new_n310), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n740), .B1(new_n733), .B2(new_n734), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n724), .B1(new_n735), .B2(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(G20), .A2(G179), .ZN(new_n743));
  XOR2_X1   g0543(.A(new_n743), .B(KEYINPUT94), .Z(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G190), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(new_n427), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n301), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n214), .ZN(new_n748));
  INV_X1    g0548(.A(new_n748), .ZN(new_n749));
  AOI22_X1  g0549(.A1(new_n746), .A2(G326), .B1(G294), .B2(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(new_n750), .B(KEYINPUT95), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n214), .A2(G179), .ZN(new_n752));
  NAND3_X1  g0552(.A1(new_n752), .A2(new_n301), .A3(new_n427), .ZN(new_n753));
  INV_X1    g0553(.A(new_n753), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n297), .B1(new_n754), .B2(G329), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(G190), .A3(G200), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G303), .ZN(new_n758));
  INV_X1    g0558(.A(G283), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n752), .A2(new_n301), .A3(G200), .ZN(new_n760));
  OAI211_X1 g0560(.A(new_n755), .B(new_n758), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n745), .A2(G200), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(G322), .B2(new_n762), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n744), .A2(new_n301), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(G200), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n764), .A2(new_n427), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI22_X1  g0567(.A1(G311), .A2(new_n765), .B1(new_n766), .B2(new_n767), .ZN(new_n768));
  NAND3_X1  g0568(.A1(new_n751), .A2(new_n763), .A3(new_n768), .ZN(new_n769));
  AOI22_X1  g0569(.A1(G50), .A2(new_n746), .B1(new_n762), .B2(G58), .ZN(new_n770));
  AOI22_X1  g0570(.A1(G68), .A2(new_n766), .B1(new_n765), .B2(G77), .ZN(new_n771));
  INV_X1    g0571(.A(new_n760), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n772), .A2(G107), .ZN(new_n773));
  INV_X1    g0573(.A(G159), .ZN(new_n774));
  OAI21_X1  g0574(.A(KEYINPUT32), .B1(new_n753), .B2(new_n774), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n773), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n297), .B1(new_n748), .B2(new_n454), .ZN(new_n777));
  INV_X1    g0577(.A(G87), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n756), .A2(new_n778), .ZN(new_n779));
  NOR3_X1   g0579(.A1(new_n753), .A2(KEYINPUT32), .A3(new_n774), .ZN(new_n780));
  NOR4_X1   g0580(.A1(new_n776), .A2(new_n777), .A3(new_n779), .A4(new_n780), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n770), .A2(new_n771), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n769), .A2(new_n782), .ZN(new_n783));
  AOI21_X1  g0583(.A(new_n742), .B1(new_n739), .B2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(new_n738), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n784), .B1(new_n664), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g0586(.A1(new_n726), .A2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n787), .ZN(G396));
  NAND4_X1  g0588(.A1(new_n614), .A2(new_n374), .A3(new_n615), .A4(new_n655), .ZN(new_n789));
  OAI211_X1 g0589(.A(new_n379), .B(new_n375), .C1(new_n376), .C2(new_n653), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n791), .B1(new_n641), .B2(new_n653), .ZN(new_n792));
  OAI211_X1 g0592(.A(new_n791), .B(new_n653), .C1(new_n638), .C2(new_n640), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NOR3_X1   g0594(.A1(new_n792), .A2(new_n794), .A3(new_n696), .ZN(new_n795));
  XNOR2_X1  g0595(.A(new_n795), .B(KEYINPUT96), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n696), .B1(new_n792), .B2(new_n794), .ZN(new_n797));
  AOI21_X1  g0597(.A(new_n724), .B1(new_n797), .B2(KEYINPUT97), .ZN(new_n798));
  OAI211_X1 g0598(.A(new_n796), .B(new_n798), .C1(KEYINPUT97), .C2(new_n797), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n739), .A2(new_n736), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n724), .B1(G77), .B2(new_n801), .ZN(new_n802));
  AOI22_X1  g0602(.A1(G294), .A2(new_n762), .B1(new_n746), .B2(G303), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n765), .A2(G116), .ZN(new_n804));
  INV_X1    g0604(.A(G311), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n295), .B1(new_n753), .B2(new_n805), .ZN(new_n806));
  OAI22_X1  g0606(.A1(new_n778), .A2(new_n760), .B1(new_n756), .B2(new_n483), .ZN(new_n807));
  AOI211_X1 g0607(.A(new_n806), .B(new_n807), .C1(G97), .C2(new_n749), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n766), .A2(G283), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n803), .A2(new_n804), .A3(new_n808), .A4(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(G143), .A2(new_n762), .B1(new_n765), .B2(G159), .ZN(new_n811));
  INV_X1    g0611(.A(G137), .ZN(new_n812));
  INV_X1    g0612(.A(new_n746), .ZN(new_n813));
  INV_X1    g0613(.A(G150), .ZN(new_n814));
  INV_X1    g0614(.A(new_n766), .ZN(new_n815));
  OAI221_X1 g0615(.A(new_n811), .B1(new_n812), .B2(new_n813), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  XOR2_X1   g0616(.A(new_n816), .B(KEYINPUT34), .Z(new_n817));
  AOI22_X1  g0617(.A1(new_n749), .A2(G58), .B1(new_n757), .B2(G50), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n295), .B1(new_n754), .B2(G132), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(new_n239), .C2(new_n760), .ZN(new_n820));
  OAI21_X1  g0620(.A(new_n810), .B1(new_n817), .B2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n802), .B1(new_n821), .B2(new_n739), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n737), .B2(new_n791), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n799), .A2(new_n823), .ZN(G384));
  NOR2_X1   g0624(.A1(new_n721), .A2(new_n260), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n399), .A2(new_n403), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(new_n387), .ZN(new_n827));
  INV_X1    g0627(.A(KEYINPUT16), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n404), .A2(new_n259), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n382), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NOR2_X1   g0631(.A1(new_n831), .A2(new_n647), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n432), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n833), .A2(KEYINPUT99), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT99), .ZN(new_n835));
  NAND3_X1  g0635(.A1(new_n432), .A2(new_n835), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n834), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n421), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n430), .B1(new_n831), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(KEYINPUT37), .B1(new_n839), .B2(new_n832), .ZN(new_n840));
  NAND3_X1  g0640(.A1(new_n409), .A2(new_n411), .A3(new_n648), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT37), .ZN(new_n842));
  AND2_X1   g0642(.A1(new_n430), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n422), .A2(new_n841), .A3(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT38), .B1(new_n837), .B2(new_n845), .ZN(new_n846));
  AND3_X1   g0646(.A1(new_n432), .A2(new_n835), .A3(new_n832), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n835), .B1(new_n432), .B2(new_n832), .ZN(new_n848));
  OAI211_X1 g0648(.A(KEYINPUT38), .B(new_n845), .C1(new_n847), .C2(new_n848), .ZN(new_n849));
  INV_X1    g0649(.A(new_n849), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n353), .B1(new_n345), .B2(new_n344), .ZN(new_n852));
  NOR2_X1   g0652(.A1(new_n340), .A2(new_n653), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  OAI221_X1 g0654(.A(new_n353), .B1(new_n340), .B2(new_n653), .C1(new_n345), .C2(new_n344), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT40), .ZN(new_n857));
  NAND4_X1  g0657(.A1(new_n856), .A2(new_n695), .A3(new_n857), .A4(new_n791), .ZN(new_n858));
  NAND3_X1  g0658(.A1(new_n856), .A2(new_n695), .A3(new_n791), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n612), .A2(new_n619), .ZN(new_n860));
  INV_X1    g0660(.A(new_n844), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n618), .A2(new_n430), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n842), .B1(new_n863), .B2(new_n841), .ZN(new_n864));
  OAI22_X1  g0664(.A1(new_n860), .A2(new_n841), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT38), .ZN(new_n866));
  NAND2_X1  g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n859), .B1(new_n849), .B2(new_n867), .ZN(new_n868));
  OAI22_X1  g0668(.A1(new_n851), .A2(new_n858), .B1(new_n868), .B2(new_n857), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n869), .A2(new_n433), .A3(new_n695), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(G330), .ZN(new_n871));
  AOI21_X1  g0671(.A(new_n869), .B1(new_n433), .B2(new_n695), .ZN(new_n872));
  OR2_X1    g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n845), .B1(new_n847), .B2(new_n848), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n874), .A2(new_n866), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n849), .A2(new_n867), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT39), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OR2_X1    g0679(.A1(new_n353), .A2(new_n655), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n876), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n875), .A2(new_n849), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n375), .A2(new_n655), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  AND2_X1   g0685(.A1(new_n793), .A2(new_n885), .ZN(new_n886));
  AND2_X1   g0686(.A1(new_n854), .A2(new_n855), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n883), .A2(new_n888), .B1(new_n619), .B2(new_n647), .ZN(new_n889));
  AND2_X1   g0689(.A1(new_n882), .A2(new_n889), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n713), .A2(new_n433), .A3(new_n716), .ZN(new_n891));
  AND3_X1   g0691(.A1(new_n891), .A2(new_n312), .A3(new_n620), .ZN(new_n892));
  XNOR2_X1  g0692(.A(new_n890), .B(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n825), .B1(new_n873), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(new_n893), .B2(new_n873), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n485), .A2(KEYINPUT35), .ZN(new_n896));
  NOR3_X1   g0696(.A1(new_n215), .A2(new_n214), .A3(new_n530), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n485), .B2(KEYINPUT35), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT98), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n896), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n898), .ZN(new_n901));
  XOR2_X1   g0701(.A(new_n901), .B(KEYINPUT36), .Z(new_n902));
  OAI21_X1  g0702(.A(G77), .B1(new_n245), .B2(new_n239), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n238), .B1(new_n903), .B2(new_n213), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n904), .A2(G1), .A3(new_n719), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n895), .A2(new_n902), .A3(new_n905), .ZN(G367));
  NAND2_X1  g0706(.A1(new_n466), .A2(new_n655), .ZN(new_n907));
  OR2_X1    g0707(.A1(new_n628), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n628), .A2(new_n632), .A3(new_n907), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(new_n910), .ZN(new_n911));
  INV_X1    g0711(.A(KEYINPUT43), .ZN(new_n912));
  NOR2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n527), .B1(new_n525), .B2(new_n653), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n629), .A2(new_n655), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n659), .A2(new_n916), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(KEYINPUT42), .ZN(new_n918));
  XOR2_X1   g0718(.A(new_n918), .B(KEYINPUT100), .Z(new_n919));
  INV_X1    g0719(.A(new_n916), .ZN(new_n920));
  OAI211_X1 g0720(.A(new_n520), .B(new_n523), .C1(new_n920), .C2(new_n599), .ZN(new_n921));
  AOI22_X1  g0721(.A1(new_n921), .A2(new_n653), .B1(KEYINPUT42), .B2(new_n917), .ZN(new_n922));
  AOI21_X1  g0722(.A(new_n913), .B1(new_n919), .B2(new_n922), .ZN(new_n923));
  NOR3_X1   g0723(.A1(new_n923), .A2(KEYINPUT43), .A3(new_n910), .ZN(new_n924));
  OAI21_X1  g0724(.A(new_n923), .B1(KEYINPUT43), .B2(new_n910), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  OAI22_X1  g0726(.A1(new_n924), .A2(new_n926), .B1(new_n668), .B2(new_n920), .ZN(new_n927));
  INV_X1    g0727(.A(new_n924), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n668), .A2(new_n920), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n929), .A3(new_n925), .ZN(new_n930));
  XNOR2_X1  g0730(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n672), .B(new_n931), .Z(new_n932));
  NAND3_X1  g0732(.A1(new_n657), .A2(new_n658), .A3(new_n654), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(KEYINPUT106), .ZN(new_n934));
  XNOR2_X1  g0734(.A(new_n934), .B(new_n665), .ZN(new_n935));
  XNOR2_X1  g0735(.A(new_n935), .B(new_n659), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n717), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT103), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n920), .B1(new_n939), .B2(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT104), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n940), .A2(new_n661), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n661), .A2(new_n916), .A3(new_n945), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n661), .A2(new_n916), .ZN(new_n947));
  INV_X1    g0747(.A(new_n945), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n943), .B1(new_n940), .B2(new_n661), .ZN(new_n950));
  NAND4_X1  g0750(.A1(new_n944), .A2(new_n946), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(new_n668), .ZN(new_n952));
  NAND3_X1  g0752(.A1(new_n951), .A2(KEYINPUT105), .A3(new_n952), .ZN(new_n953));
  OR2_X1    g0753(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT105), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND4_X1  g0757(.A1(new_n938), .A2(new_n953), .A3(new_n954), .A4(new_n957), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n932), .B1(new_n958), .B2(new_n717), .ZN(new_n959));
  OAI211_X1 g0759(.A(new_n927), .B(new_n930), .C1(new_n959), .C2(new_n723), .ZN(new_n960));
  AND3_X1   g0760(.A1(new_n229), .A2(new_n210), .A3(new_n295), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n740), .B1(new_n461), .B2(new_n210), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n724), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G303), .A2(new_n762), .B1(new_n746), .B2(G311), .ZN(new_n964));
  INV_X1    g0764(.A(new_n765), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n964), .B1(new_n759), .B2(new_n965), .C1(new_n569), .C2(new_n815), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n760), .A2(new_n454), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n297), .B1(new_n754), .B2(G317), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n968), .B1(new_n483), .B2(new_n748), .ZN(new_n969));
  AND3_X1   g0769(.A1(new_n757), .A2(KEYINPUT46), .A3(G116), .ZN(new_n970));
  AOI21_X1  g0770(.A(KEYINPUT46), .B1(new_n757), .B2(G116), .ZN(new_n971));
  OR4_X1    g0771(.A1(new_n967), .A2(new_n969), .A3(new_n970), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n762), .A2(G150), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT107), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n753), .A2(new_n812), .B1(new_n756), .B2(new_n245), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n973), .B1(new_n974), .B2(new_n975), .C1(new_n965), .C2(new_n202), .ZN(new_n976));
  AOI22_X1  g0776(.A1(new_n746), .A2(G143), .B1(new_n974), .B2(new_n975), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n748), .A2(new_n239), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n295), .B(new_n978), .C1(G77), .C2(new_n772), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n977), .B(new_n979), .C1(new_n774), .C2(new_n815), .ZN(new_n980));
  OAI22_X1  g0780(.A1(new_n966), .A2(new_n972), .B1(new_n976), .B2(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n963), .B1(new_n982), .B2(new_n739), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n785), .B2(new_n910), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n960), .A2(new_n984), .ZN(G387));
  NAND3_X1  g0785(.A1(new_n657), .A2(new_n658), .A3(new_n738), .ZN(new_n986));
  OAI22_X1  g0786(.A1(new_n731), .A2(new_n673), .B1(G107), .B2(new_n210), .ZN(new_n987));
  AOI211_X1 g0787(.A(G45), .B(new_n674), .C1(G68), .C2(G77), .ZN(new_n988));
  INV_X1    g0788(.A(KEYINPUT108), .ZN(new_n989));
  OR2_X1    g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(new_n989), .ZN(new_n991));
  INV_X1    g0791(.A(new_n249), .ZN(new_n992));
  OR3_X1    g0792(.A1(new_n992), .A2(KEYINPUT50), .A3(G50), .ZN(new_n993));
  OAI21_X1  g0793(.A(KEYINPUT50), .B1(new_n992), .B2(G50), .ZN(new_n994));
  NAND4_X1  g0794(.A1(new_n990), .A2(new_n991), .A3(new_n993), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n727), .B1(new_n233), .B2(G45), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n987), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  INV_X1    g0797(.A(new_n740), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n724), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  AOI22_X1  g0799(.A1(G50), .A2(new_n762), .B1(new_n746), .B2(G159), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G68), .A2(new_n765), .B1(new_n766), .B2(new_n249), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n366), .A2(new_n749), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n297), .B1(new_n753), .B2(new_n814), .ZN(new_n1003));
  NOR2_X1   g0803(.A1(new_n756), .A2(new_n328), .ZN(new_n1004));
  NOR3_X1   g0804(.A1(new_n1003), .A2(new_n967), .A3(new_n1004), .ZN(new_n1005));
  NAND4_X1  g0805(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .A4(new_n1005), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n748), .A2(new_n759), .B1(new_n756), .B2(new_n569), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(G303), .A2(new_n765), .B1(new_n762), .B2(G317), .ZN(new_n1008));
  INV_X1    g0808(.A(G322), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1008), .B1(new_n805), .B2(new_n815), .C1(new_n1009), .C2(new_n813), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT48), .ZN(new_n1011));
  AOI21_X1  g0811(.A(new_n1007), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1012), .B1(new_n1011), .B2(new_n1010), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  AND2_X1   g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n297), .B1(new_n754), .B2(G326), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n1016), .B1(new_n530), .B2(new_n760), .ZN(new_n1017));
  XOR2_X1   g0817(.A(new_n1017), .B(KEYINPUT109), .Z(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n1006), .B1(new_n1015), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n999), .B1(new_n1020), .B2(new_n739), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n936), .A2(new_n723), .B1(new_n986), .B2(new_n1021), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n937), .A2(new_n672), .ZN(new_n1023));
  NOR2_X1   g0823(.A1(new_n936), .A2(new_n717), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(G393));
  NOR2_X1   g0825(.A1(new_n727), .A2(new_n237), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n740), .B1(new_n210), .B2(new_n454), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n724), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n916), .A2(new_n785), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(G150), .A2(new_n746), .B1(new_n762), .B2(G159), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT51), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n295), .B1(new_n754), .B2(G143), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n239), .B2(new_n756), .C1(new_n778), .C2(new_n760), .ZN(new_n1033));
  XNOR2_X1  g0833(.A(new_n1033), .B(KEYINPUT111), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1031), .A2(new_n1034), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n765), .A2(new_n249), .B1(G77), .B2(new_n749), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n1036), .B1(new_n202), .B2(new_n815), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT112), .Z(new_n1038));
  AOI22_X1  g0838(.A1(G311), .A2(new_n762), .B1(new_n746), .B2(G317), .ZN(new_n1039));
  XNOR2_X1  g0839(.A(new_n1039), .B(KEYINPUT52), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n748), .A2(new_n530), .B1(new_n756), .B2(new_n759), .ZN(new_n1041));
  OAI211_X1 g0841(.A(new_n773), .B(new_n295), .C1(new_n1009), .C2(new_n753), .ZN(new_n1042));
  AOI211_X1 g0842(.A(new_n1041), .B(new_n1042), .C1(G303), .C2(new_n766), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n569), .B2(new_n965), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1035), .A2(new_n1038), .B1(new_n1040), .B2(new_n1044), .ZN(new_n1045));
  AOI211_X1 g0845(.A(new_n1028), .B(new_n1029), .C1(new_n739), .C2(new_n1045), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n723), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n954), .A2(new_n955), .ZN(new_n1048));
  INV_X1    g0848(.A(KEYINPUT110), .ZN(new_n1049));
  AOI21_X1  g0849(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g0850(.A1(new_n954), .A2(KEYINPUT110), .A3(new_n955), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1046), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1048), .A2(new_n937), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n958), .A2(new_n1053), .A3(new_n672), .ZN(new_n1054));
  AOI21_X1  g0854(.A(KEYINPUT113), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n1052), .A2(KEYINPUT113), .A3(new_n1054), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(G390));
  OAI21_X1  g0858(.A(new_n724), .B1(new_n249), .B2(new_n801), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n737), .B1(new_n876), .B2(new_n879), .ZN(new_n1060));
  XOR2_X1   g0860(.A(KEYINPUT54), .B(G143), .Z(new_n1061));
  XNOR2_X1  g0861(.A(new_n1061), .B(KEYINPUT116), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(G128), .A2(new_n746), .B1(new_n765), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g0863(.A(G132), .ZN(new_n1064));
  INV_X1    g0864(.A(new_n762), .ZN(new_n1065));
  OAI221_X1 g0865(.A(new_n1063), .B1(new_n1064), .B2(new_n1065), .C1(new_n812), .C2(new_n815), .ZN(new_n1066));
  NOR2_X1   g0866(.A1(new_n756), .A2(new_n814), .ZN(new_n1067));
  XOR2_X1   g0867(.A(KEYINPUT117), .B(KEYINPUT53), .Z(new_n1068));
  XNOR2_X1  g0868(.A(new_n1067), .B(new_n1068), .ZN(new_n1069));
  INV_X1    g0869(.A(G125), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n297), .B1(new_n753), .B2(new_n1070), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1071), .B1(G50), .B2(new_n772), .ZN(new_n1072));
  OAI211_X1 g0872(.A(new_n1069), .B(new_n1072), .C1(new_n774), .C2(new_n748), .ZN(new_n1073));
  AOI211_X1 g0873(.A(new_n297), .B(new_n779), .C1(G294), .C2(new_n754), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n749), .A2(G77), .B1(new_n772), .B2(G68), .ZN(new_n1075));
  OAI211_X1 g0875(.A(new_n1074), .B(new_n1075), .C1(new_n965), .C2(new_n454), .ZN(new_n1076));
  AOI22_X1  g0876(.A1(G107), .A2(new_n766), .B1(new_n762), .B2(G116), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n1077), .B1(new_n759), .B2(new_n813), .ZN(new_n1078));
  OAI22_X1  g0878(.A1(new_n1066), .A2(new_n1073), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1079));
  AOI211_X1 g0879(.A(new_n1059), .B(new_n1060), .C1(new_n739), .C2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n793), .A2(new_n885), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n881), .B1(new_n1081), .B2(new_n856), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n1082), .B1(new_n876), .B2(new_n879), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n599), .A2(new_n561), .A3(new_n565), .ZN(new_n1084));
  AND2_X1   g0884(.A1(new_n608), .A2(new_n632), .ZN(new_n1085));
  NAND3_X1  g0885(.A1(new_n527), .A2(new_n1084), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(KEYINPUT26), .B1(new_n478), .B2(new_n639), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1086), .B(new_n628), .C1(new_n1087), .C2(new_n698), .ZN(new_n1088));
  AOI21_X1  g0888(.A(KEYINPUT90), .B1(new_n1088), .B2(new_n653), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n711), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n791), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n887), .B1(new_n1091), .B2(new_n885), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n877), .A2(new_n880), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1083), .A2(new_n1094), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n856), .A2(new_n695), .A3(G330), .A4(new_n791), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n1047), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g0897(.A(new_n1082), .ZN(new_n1098));
  AND3_X1   g0898(.A1(new_n875), .A2(KEYINPUT39), .A3(new_n849), .ZN(new_n1099));
  AOI21_X1  g0899(.A(KEYINPUT39), .B1(new_n849), .B2(new_n867), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1098), .B1(new_n1099), .B2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n884), .B1(new_n712), .B2(new_n791), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n880), .B(new_n877), .C1(new_n1102), .C2(new_n887), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND3_X1  g0904(.A1(new_n695), .A2(G330), .A3(new_n791), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1105), .A2(new_n887), .ZN(new_n1106));
  AOI21_X1  g0906(.A(KEYINPUT114), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(KEYINPUT114), .B(new_n1106), .C1(new_n1083), .C2(new_n1094), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1097), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(KEYINPUT115), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI211_X1 g0912(.A(KEYINPUT115), .B(new_n1097), .C1(new_n1107), .C2(new_n1109), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1080), .B1(new_n1112), .B2(new_n1113), .ZN(new_n1114));
  NOR3_X1   g0914(.A1(new_n1083), .A2(new_n1094), .A3(new_n1106), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1116), .B1(new_n1107), .B2(new_n1109), .ZN(new_n1117));
  AND2_X1   g0917(.A1(new_n1105), .A2(new_n887), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n1106), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1119), .A2(new_n1102), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1105), .A2(new_n887), .ZN(new_n1121));
  AOI21_X1  g0921(.A(new_n886), .B1(new_n1121), .B2(new_n1096), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1120), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n433), .A2(new_n697), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1124), .A2(new_n892), .A3(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1117), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n621), .A2(new_n891), .A3(new_n1125), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1122), .B1(new_n1119), .B2(new_n1102), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g0930(.A(new_n1130), .B(new_n1116), .C1(new_n1107), .C2(new_n1109), .ZN(new_n1131));
  NAND3_X1  g0931(.A1(new_n1127), .A2(new_n672), .A3(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1114), .A2(new_n1132), .ZN(G378));
  INV_X1    g0933(.A(KEYINPUT57), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n882), .A2(new_n889), .ZN(new_n1135));
  NAND3_X1  g0935(.A1(new_n313), .A2(new_n269), .A3(new_n648), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n269), .A2(new_n648), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n308), .A2(new_n309), .A3(new_n312), .A4(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  NAND2_X1  g0941(.A1(new_n1139), .A2(new_n1141), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1136), .A2(new_n1138), .A3(new_n1140), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n869), .B2(G330), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n859), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n857), .B1(new_n877), .B2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n858), .B1(new_n875), .B2(new_n849), .ZN(new_n1148));
  OAI211_X1 g0948(.A(new_n1144), .B(G330), .C1(new_n1147), .C2(new_n1148), .ZN(new_n1149));
  INV_X1    g0949(.A(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1135), .B1(new_n1145), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(G330), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1152), .A2(new_n1143), .A3(new_n1142), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1153), .A2(new_n890), .A3(new_n1149), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1134), .B1(new_n1151), .B2(new_n1154), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1106), .B1(new_n1083), .B2(new_n1094), .ZN(new_n1156));
  INV_X1    g0956(.A(KEYINPUT114), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1156), .A2(new_n1157), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n1115), .B(new_n1126), .C1(new_n1158), .C2(new_n1108), .ZN(new_n1159));
  OAI21_X1  g0959(.A(new_n1155), .B1(new_n1159), .B2(new_n1128), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1128), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n1131), .A2(new_n1161), .B1(new_n1154), .B2(new_n1151), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1160), .B(new_n672), .C1(new_n1162), .C2(KEYINPUT57), .ZN(new_n1163));
  OAI22_X1  g0963(.A1(new_n454), .A2(new_n815), .B1(new_n1065), .B2(new_n483), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1164), .B1(G116), .B2(new_n746), .ZN(new_n1165));
  OAI211_X1 g0965(.A(new_n511), .B(new_n295), .C1(new_n753), .C2(new_n759), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n760), .A2(new_n245), .ZN(new_n1167));
  NOR4_X1   g0967(.A1(new_n1166), .A2(new_n978), .A3(new_n1004), .A4(new_n1167), .ZN(new_n1168));
  OAI211_X1 g0968(.A(new_n1165), .B(new_n1168), .C1(new_n461), .C2(new_n965), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT58), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n295), .A2(new_n511), .ZN(new_n1171));
  AOI21_X1  g0971(.A(G50), .B1(new_n250), .B2(new_n511), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n1169), .A2(new_n1170), .B1(new_n1171), .B2(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G128), .A2(new_n762), .B1(new_n765), .B2(G137), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n1064), .B2(new_n815), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(new_n1062), .A2(new_n757), .B1(G150), .B2(new_n749), .ZN(new_n1176));
  OAI21_X1  g0976(.A(new_n1176), .B1(new_n813), .B2(new_n1070), .ZN(new_n1177));
  NOR2_X1   g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n772), .A2(G159), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n754), .C2(G124), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  NOR2_X1   g0983(.A1(new_n1179), .A2(KEYINPUT59), .ZN(new_n1184));
  OAI221_X1 g0984(.A(new_n1173), .B1(new_n1170), .B2(new_n1169), .C1(new_n1183), .C2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n1185), .A2(new_n739), .ZN(new_n1186));
  OAI211_X1 g0986(.A(new_n1186), .B(new_n724), .C1(G50), .C2(new_n801), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1144), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1187), .B1(new_n1188), .B2(new_n736), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n1151), .A2(new_n1154), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1189), .B1(new_n1190), .B2(new_n723), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1163), .A2(new_n1191), .ZN(G375));
  NAND2_X1  g0992(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n932), .B(KEYINPUT118), .Z(new_n1194));
  INV_X1    g0994(.A(new_n1194), .ZN(new_n1195));
  NAND3_X1  g0995(.A1(new_n1126), .A2(new_n1193), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n887), .A2(new_n736), .ZN(new_n1197));
  OAI21_X1  g0997(.A(new_n724), .B1(G68), .B2(new_n801), .ZN(new_n1198));
  XNOR2_X1  g0998(.A(new_n1198), .B(KEYINPUT119), .ZN(new_n1199));
  AOI22_X1  g0999(.A1(G283), .A2(new_n762), .B1(new_n746), .B2(G294), .ZN(new_n1200));
  OAI221_X1 g1000(.A(new_n1200), .B1(new_n483), .B2(new_n965), .C1(new_n530), .C2(new_n815), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n772), .A2(G77), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n757), .A2(G97), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n297), .B1(new_n754), .B2(G303), .ZN(new_n1204));
  NAND4_X1  g1004(.A1(new_n1002), .A2(new_n1202), .A3(new_n1203), .A4(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n765), .A2(G150), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1167), .ZN(new_n1207));
  AOI21_X1  g1007(.A(new_n295), .B1(new_n754), .B2(G128), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n749), .A2(G50), .B1(new_n757), .B2(G159), .ZN(new_n1209));
  NAND4_X1  g1009(.A1(new_n1206), .A2(new_n1207), .A3(new_n1208), .A4(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n766), .A2(new_n1062), .ZN(new_n1211));
  OAI221_X1 g1011(.A(new_n1211), .B1(new_n1065), .B2(new_n812), .C1(new_n1064), .C2(new_n813), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n1201), .A2(new_n1205), .B1(new_n1210), .B2(new_n1212), .ZN(new_n1213));
  AOI21_X1  g1013(.A(new_n1199), .B1(new_n1213), .B2(new_n739), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n1124), .A2(new_n723), .B1(new_n1197), .B2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1196), .A2(new_n1215), .ZN(G381));
  OR4_X1    g1016(.A1(G396), .A2(G381), .A3(G384), .A4(G393), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(G390), .A2(G387), .A3(new_n1217), .ZN(new_n1218));
  INV_X1    g1018(.A(G378), .ZN(new_n1219));
  NAND4_X1  g1019(.A1(new_n1218), .A2(new_n1219), .A3(new_n1163), .A4(new_n1191), .ZN(G407));
  NAND3_X1  g1020(.A1(new_n650), .A2(new_n651), .A3(G213), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1219), .A2(new_n1222), .ZN(new_n1223));
  OAI211_X1 g1023(.A(G407), .B(G213), .C1(G375), .C2(new_n1223), .ZN(G409));
  INV_X1    g1024(.A(KEYINPUT122), .ZN(new_n1225));
  AND3_X1   g1025(.A1(new_n799), .A2(KEYINPUT121), .A3(new_n823), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1226), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1128), .A2(new_n1129), .A3(KEYINPUT60), .ZN(new_n1228));
  AND2_X1   g1028(.A1(new_n1228), .A2(new_n672), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT60), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1193), .B1(new_n1130), .B2(new_n1230), .ZN(new_n1231));
  NAND2_X1  g1031(.A1(new_n1229), .A2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n1215), .ZN(new_n1233));
  AOI21_X1  g1033(.A(KEYINPUT121), .B1(new_n799), .B2(new_n823), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1227), .B1(new_n1233), .B2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1215), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1237), .B1(new_n1229), .B2(new_n1231), .ZN(new_n1238));
  NOR3_X1   g1038(.A1(new_n1238), .A2(new_n1226), .A3(new_n1234), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1225), .B1(new_n1236), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1222), .A2(G2897), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1233), .A2(new_n1227), .A3(new_n1235), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1238), .A2(KEYINPUT121), .A3(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1242), .A2(KEYINPUT122), .A3(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1240), .A2(new_n1241), .A3(new_n1245), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1247));
  OR2_X1    g1047(.A1(new_n1247), .A2(new_n1241), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1163), .A2(G378), .A3(new_n1191), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1115), .B1(new_n1158), .B2(new_n1108), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1128), .B1(new_n1251), .B2(new_n1130), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1190), .A2(new_n1195), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1191), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1254), .A2(new_n1114), .A3(new_n1132), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(KEYINPUT120), .ZN(new_n1256));
  INV_X1    g1056(.A(KEYINPUT120), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1254), .A2(new_n1114), .A3(new_n1257), .A4(new_n1132), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1250), .A2(new_n1256), .A3(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1249), .B1(new_n1259), .B2(new_n1221), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(G387), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1261));
  INV_X1    g1061(.A(new_n1057), .ZN(new_n1262));
  OAI211_X1 g1062(.A(new_n960), .B(new_n984), .C1(new_n1262), .C2(new_n1055), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n1261), .A2(new_n1263), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(G393), .B(new_n787), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1264), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1261), .A2(new_n1263), .A3(new_n1265), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1267), .A2(new_n1268), .ZN(new_n1269));
  NOR3_X1   g1069(.A1(new_n1260), .A2(new_n1269), .A3(KEYINPUT61), .ZN(new_n1270));
  AND2_X1   g1070(.A1(new_n1240), .A2(new_n1245), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1259), .A2(new_n1221), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(KEYINPUT63), .ZN(new_n1273));
  OR2_X1    g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(KEYINPUT123), .ZN(new_n1275));
  AND3_X1   g1075(.A1(new_n1272), .A2(new_n1275), .A3(new_n1273), .ZN(new_n1276));
  AOI21_X1  g1076(.A(new_n1275), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1277));
  OAI211_X1 g1077(.A(new_n1270), .B(new_n1274), .C1(new_n1276), .C2(new_n1277), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1259), .A2(new_n1221), .ZN(new_n1279));
  INV_X1    g1079(.A(new_n1249), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1279), .A2(new_n1280), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT61), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1281), .A2(new_n1282), .ZN(new_n1283));
  NAND4_X1  g1083(.A1(new_n1259), .A2(KEYINPUT62), .A3(new_n1221), .A4(new_n1271), .ZN(new_n1284));
  XOR2_X1   g1084(.A(KEYINPUT124), .B(KEYINPUT62), .Z(new_n1285));
  AOI22_X1  g1085(.A1(KEYINPUT125), .A2(new_n1284), .B1(new_n1272), .B2(new_n1285), .ZN(new_n1286));
  AND2_X1   g1086(.A1(new_n1271), .A2(KEYINPUT62), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1287), .A2(new_n1288), .A3(new_n1221), .A4(new_n1259), .ZN(new_n1289));
  AOI21_X1  g1089(.A(new_n1283), .B1(new_n1286), .B2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1269), .ZN(new_n1291));
  OAI21_X1  g1091(.A(new_n1278), .B1(new_n1290), .B2(new_n1291), .ZN(G405));
  OR2_X1    g1092(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G375), .A2(new_n1219), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1294), .A2(KEYINPUT126), .A3(new_n1250), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT126), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(G375), .A2(new_n1296), .A3(new_n1219), .ZN(new_n1297));
  AOI21_X1  g1097(.A(new_n1247), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1295), .A2(new_n1271), .A3(new_n1297), .ZN(new_n1301));
  NAND4_X1  g1101(.A1(new_n1293), .A2(new_n1299), .A3(new_n1300), .A4(new_n1301), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1301), .ZN(new_n1303));
  OAI211_X1 g1103(.A(KEYINPUT127), .B(new_n1269), .C1(new_n1303), .C2(new_n1298), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1302), .A2(new_n1304), .ZN(G402));
endmodule


