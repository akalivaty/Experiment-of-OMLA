//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 0 0 1 1 1 1 0 0 1 0 1 1 0 1 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 1 1 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:02 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n673, new_n674, new_n675, new_n676, new_n678, new_n679, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n767, new_n768, new_n769, new_n770, new_n772,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n877, new_n878, new_n879, new_n881, new_n882,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n895, new_n896, new_n898, new_n899,
    new_n900, new_n901, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n937, new_n938;
  INV_X1    g000(.A(KEYINPUT67), .ZN(new_n202));
  INV_X1    g001(.A(G113gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n203), .A2(G120gat), .ZN(new_n204));
  INV_X1    g003(.A(G120gat), .ZN(new_n205));
  NOR2_X1   g004(.A1(new_n205), .A2(G113gat), .ZN(new_n206));
  OAI21_X1  g005(.A(KEYINPUT65), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(G134gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(G127gat), .A2(G134gat), .ZN(new_n211));
  AOI21_X1  g010(.A(KEYINPUT1), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n205), .A2(G113gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n203), .A2(G120gat), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT65), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  NAND3_X1  g015(.A1(new_n207), .A2(new_n212), .A3(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G127gat), .A2(G134gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(G127gat), .A2(G134gat), .ZN(new_n219));
  OAI21_X1  g018(.A(KEYINPUT64), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n210), .A2(new_n221), .A3(new_n211), .ZN(new_n222));
  XNOR2_X1  g021(.A(G113gat), .B(G120gat), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n220), .B(new_n222), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AND3_X1   g023(.A1(new_n217), .A2(new_n224), .A3(KEYINPUT66), .ZN(new_n225));
  AOI21_X1  g024(.A(KEYINPUT66), .B1(new_n217), .B2(new_n224), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  XNOR2_X1  g026(.A(KEYINPUT27), .B(G183gat), .ZN(new_n228));
  INV_X1    g027(.A(G190gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(KEYINPUT28), .ZN(new_n231));
  INV_X1    g030(.A(G169gat), .ZN(new_n232));
  INV_X1    g031(.A(G176gat), .ZN(new_n233));
  NAND3_X1  g032(.A1(new_n232), .A2(new_n233), .A3(KEYINPUT26), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT28), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n228), .A2(new_n235), .A3(new_n229), .ZN(new_n236));
  NAND2_X1  g035(.A1(G183gat), .A2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI21_X1  g037(.A(KEYINPUT26), .B1(new_n232), .B2(new_n233), .ZN(new_n239));
  NAND2_X1  g038(.A1(G169gat), .A2(G176gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n238), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n231), .A2(new_n234), .A3(new_n236), .A4(new_n241), .ZN(new_n242));
  OR3_X1    g041(.A1(KEYINPUT23), .A2(G169gat), .A3(G176gat), .ZN(new_n243));
  OAI21_X1  g042(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OR2_X1    g044(.A1(G183gat), .A2(G190gat), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n246), .A2(KEYINPUT24), .A3(new_n237), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT24), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n238), .A2(new_n248), .ZN(new_n249));
  NAND4_X1  g048(.A1(new_n245), .A2(new_n247), .A3(new_n240), .A4(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT25), .ZN(new_n251));
  AOI22_X1  g050(.A1(new_n243), .A2(new_n244), .B1(new_n238), .B2(new_n248), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT25), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n252), .A2(new_n253), .A3(new_n240), .A4(new_n247), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n242), .A2(new_n251), .A3(new_n254), .ZN(new_n255));
  OAI21_X1  g054(.A(new_n202), .B1(new_n227), .B2(new_n255), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n242), .A2(new_n251), .A3(new_n254), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n217), .A2(new_n224), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT66), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n217), .A2(new_n224), .A3(KEYINPUT66), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n257), .A2(new_n262), .A3(KEYINPUT67), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n227), .A2(new_n255), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n256), .A2(new_n263), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G227gat), .A2(G233gat), .ZN(new_n266));
  INV_X1    g065(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n265), .A2(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT33), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n268), .B1(KEYINPUT32), .B2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G15gat), .B(G43gat), .ZN(new_n271));
  XNOR2_X1  g070(.A(G71gat), .B(G99gat), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n271), .B(new_n272), .Z(new_n273));
  NAND2_X1  g072(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT32), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(new_n265), .B2(new_n267), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT69), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT68), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n269), .B1(new_n273), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(new_n278), .B2(new_n273), .ZN(new_n280));
  AND3_X1   g079(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g080(.A(new_n277), .B1(new_n276), .B2(new_n280), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n274), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND4_X1  g082(.A1(new_n256), .A2(new_n263), .A3(new_n266), .A4(new_n264), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n284), .B(KEYINPUT34), .ZN(new_n285));
  INV_X1    g084(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n283), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g086(.A(new_n274), .B(new_n285), .C1(new_n281), .C2(new_n282), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n287), .A2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT90), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n287), .A2(KEYINPUT90), .A3(new_n288), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(G197gat), .B(G204gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(G211gat), .A2(G218gat), .ZN(new_n295));
  INV_X1    g094(.A(KEYINPUT22), .ZN(new_n296));
  AND3_X1   g095(.A1(new_n295), .A2(KEYINPUT71), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT71), .B1(new_n295), .B2(new_n296), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n294), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT72), .ZN(new_n300));
  INV_X1    g099(.A(G211gat), .ZN(new_n301));
  INV_X1    g100(.A(G218gat), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n303), .A2(new_n295), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n299), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n295), .A2(new_n296), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT71), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n295), .A2(KEYINPUT71), .A3(new_n296), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n304), .A2(new_n300), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n303), .A2(KEYINPUT72), .A3(new_n295), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .A4(new_n294), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT29), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n305), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  INV_X1    g114(.A(KEYINPUT3), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(G148gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n318), .A2(G141gat), .ZN(new_n319));
  INV_X1    g118(.A(G141gat), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(G148gat), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(KEYINPUT2), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g123(.A1(G155gat), .A2(G162gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G155gat), .A2(G162gat), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(G155gat), .ZN(new_n329));
  INV_X1    g128(.A(G162gat), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n323), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G155gat), .A2(G162gat), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT77), .ZN(new_n334));
  AND3_X1   g133(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n334), .B1(new_n333), .B2(new_n322), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n317), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g137(.A(new_n316), .B(new_n328), .C1(new_n335), .C2(new_n336), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n314), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n305), .A2(new_n313), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(KEYINPUT83), .A3(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT83), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n325), .B1(new_n323), .B2(new_n326), .ZN(new_n345));
  XNOR2_X1  g144(.A(G141gat), .B(G148gat), .ZN(new_n346));
  OAI21_X1  g145(.A(KEYINPUT77), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n333), .A2(new_n334), .A3(new_n322), .ZN(new_n348));
  AOI22_X1  g147(.A1(new_n347), .A2(new_n348), .B1(new_n324), .B2(new_n327), .ZN(new_n349));
  AOI21_X1  g148(.A(new_n349), .B1(new_n315), .B2(new_n316), .ZN(new_n350));
  AOI22_X1  g149(.A1(new_n339), .A2(new_n314), .B1(new_n305), .B2(new_n313), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n344), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(G228gat), .A2(G233gat), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n353), .ZN(new_n355));
  OAI211_X1 g154(.A(new_n344), .B(new_n355), .C1(new_n350), .C2(new_n351), .ZN(new_n356));
  AOI21_X1  g155(.A(G22gat), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  XOR2_X1   g156(.A(G78gat), .B(G106gat), .Z(new_n358));
  XNOR2_X1  g157(.A(new_n358), .B(KEYINPUT31), .ZN(new_n359));
  XOR2_X1   g158(.A(KEYINPUT82), .B(G50gat), .Z(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n354), .A2(G22gat), .A3(new_n356), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n363), .B1(new_n357), .B2(KEYINPUT84), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT84), .ZN(new_n367));
  AOI211_X1 g166(.A(new_n367), .B(G22gat), .C1(new_n354), .C2(new_n356), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n361), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n369), .A2(KEYINPUT85), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT85), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n371), .B(new_n361), .C1(new_n366), .C2(new_n368), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n365), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n293), .A2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(G226gat), .ZN(new_n375));
  INV_X1    g174(.A(G233gat), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n257), .B2(KEYINPUT29), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n255), .A2(new_n377), .ZN(new_n380));
  AOI22_X1  g179(.A1(new_n379), .A2(KEYINPUT73), .B1(KEYINPUT74), .B2(new_n380), .ZN(new_n381));
  OR2_X1    g180(.A1(new_n380), .A2(KEYINPUT74), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n377), .B1(new_n255), .B2(new_n314), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT73), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n381), .A2(new_n341), .A3(new_n382), .A4(new_n385), .ZN(new_n386));
  INV_X1    g185(.A(new_n341), .ZN(new_n387));
  INV_X1    g186(.A(new_n380), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n387), .B1(new_n388), .B2(new_n383), .ZN(new_n389));
  XOR2_X1   g188(.A(G8gat), .B(G36gat), .Z(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G92gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(KEYINPUT75), .B(G64gat), .ZN(new_n392));
  XOR2_X1   g191(.A(new_n391), .B(new_n392), .Z(new_n393));
  INV_X1    g192(.A(new_n393), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n386), .A2(new_n389), .A3(new_n394), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT76), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n386), .A2(new_n389), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(new_n393), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT30), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT30), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n398), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g201(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n403));
  XNOR2_X1  g202(.A(G57gat), .B(G85gat), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT79), .B(KEYINPUT0), .ZN(new_n405));
  XNOR2_X1  g204(.A(new_n404), .B(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G1gat), .B(G29gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n406), .B(new_n407), .Z(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(G225gat), .A2(G233gat), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n347), .A2(new_n348), .ZN(new_n412));
  NAND4_X1  g211(.A1(new_n412), .A2(new_n217), .A3(new_n224), .A4(new_n328), .ZN(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  AND2_X1   g213(.A1(new_n337), .A2(new_n258), .ZN(new_n415));
  OAI21_X1  g214(.A(new_n411), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT4), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n413), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n337), .A2(KEYINPUT3), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n420), .A2(new_n258), .A3(new_n339), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n349), .B(KEYINPUT4), .C1(new_n225), .C2(new_n226), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT78), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT78), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n419), .A2(new_n421), .A3(new_n422), .A4(new_n425), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n417), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n418), .B1(new_n227), .B2(new_n337), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(new_n421), .C1(new_n418), .C2(new_n413), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n411), .A2(KEYINPUT5), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI211_X1 g230(.A(KEYINPUT6), .B(new_n409), .C1(new_n427), .C2(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(new_n432), .B(KEYINPUT81), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n424), .A2(new_n426), .ZN(new_n434));
  INV_X1    g233(.A(new_n417), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n429), .A2(new_n430), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n408), .A3(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT6), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n409), .B1(new_n427), .B2(new_n431), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT35), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n374), .A2(new_n403), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n365), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n354), .A2(new_n356), .ZN(new_n445));
  INV_X1    g244(.A(G22gat), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(new_n367), .ZN(new_n448));
  NAND2_X1  g247(.A1(new_n357), .A2(KEYINPUT84), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n448), .A2(new_n449), .A3(new_n363), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n371), .B1(new_n450), .B2(new_n361), .ZN(new_n451));
  INV_X1    g250(.A(new_n372), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n444), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT80), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n441), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g254(.A1(new_n438), .A2(new_n440), .A3(KEYINPUT80), .A4(new_n439), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n433), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n276), .A2(new_n280), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(KEYINPUT69), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n276), .A2(new_n277), .A3(new_n280), .ZN(new_n461));
  AOI22_X1  g260(.A1(new_n460), .A2(new_n461), .B1(new_n273), .B2(new_n270), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n285), .B1(new_n462), .B2(KEYINPUT70), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT70), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n283), .A2(new_n464), .A3(new_n286), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n453), .A2(new_n458), .A3(new_n403), .A4(new_n466), .ZN(new_n467));
  AND3_X1   g266(.A1(new_n467), .A2(KEYINPUT91), .A3(KEYINPUT35), .ZN(new_n468));
  AOI21_X1  g267(.A(KEYINPUT91), .B1(new_n467), .B2(KEYINPUT35), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n443), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT81), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n432), .B(new_n471), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n472), .B1(new_n455), .B2(new_n456), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n396), .A2(new_n400), .A3(new_n402), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n373), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n463), .A2(KEYINPUT36), .A3(new_n465), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT36), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n289), .A2(new_n477), .ZN(new_n478));
  AND2_X1   g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n475), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT86), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n381), .A2(new_n382), .A3(new_n385), .ZN(new_n482));
  OR3_X1    g281(.A1(new_n482), .A2(KEYINPUT88), .A3(new_n341), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n341), .B1(new_n388), .B2(new_n383), .ZN(new_n484));
  OAI21_X1  g283(.A(KEYINPUT88), .B1(new_n482), .B2(new_n341), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n483), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(KEYINPUT37), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT38), .ZN(new_n488));
  XNOR2_X1  g287(.A(KEYINPUT89), .B(KEYINPUT37), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n397), .A2(new_n489), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n487), .A2(new_n488), .A3(new_n394), .A4(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  OAI211_X1 g291(.A(new_n490), .B(new_n394), .C1(new_n492), .C2(new_n397), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n399), .B1(new_n493), .B2(KEYINPUT38), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n491), .A2(new_n494), .A3(new_n433), .A4(new_n441), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n429), .A2(KEYINPUT87), .A3(new_n411), .ZN(new_n496));
  OR2_X1    g295(.A1(new_n414), .A2(new_n415), .ZN(new_n497));
  OAI211_X1 g296(.A(new_n496), .B(KEYINPUT39), .C1(new_n411), .C2(new_n497), .ZN(new_n498));
  OAI211_X1 g297(.A(new_n498), .B(new_n408), .C1(KEYINPUT39), .C2(new_n496), .ZN(new_n499));
  XNOR2_X1  g298(.A(new_n499), .B(KEYINPUT40), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n500), .A2(new_n440), .A3(new_n474), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n453), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT86), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n475), .A2(new_n479), .A3(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n481), .A2(new_n502), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n470), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(G15gat), .B(G22gat), .ZN(new_n507));
  INV_X1    g306(.A(G1gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(KEYINPUT16), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n510), .B1(G1gat), .B2(new_n507), .ZN(new_n511));
  INV_X1    g310(.A(G8gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(new_n511), .B(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT21), .ZN(new_n514));
  NAND2_X1  g313(.A1(G71gat), .A2(G78gat), .ZN(new_n515));
  XNOR2_X1  g314(.A(new_n515), .B(KEYINPUT99), .ZN(new_n516));
  AOI21_X1  g315(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(G57gat), .B(G64gat), .ZN(new_n518));
  OAI221_X1 g317(.A(new_n516), .B1(G71gat), .B2(G78gat), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(G64gat), .ZN(new_n520));
  OR3_X1    g319(.A1(new_n520), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n520), .A2(G57gat), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT100), .B1(new_n520), .B2(G57gat), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(G71gat), .ZN(new_n525));
  INV_X1    g324(.A(G78gat), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n525), .A2(new_n526), .A3(KEYINPUT9), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n519), .A2(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n513), .B1(new_n514), .B2(new_n530), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n531), .B(G183gat), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n530), .A2(new_n514), .ZN(new_n533));
  XOR2_X1   g332(.A(new_n532), .B(new_n533), .Z(new_n534));
  INV_X1    g333(.A(G231gat), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n535), .A2(new_n376), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n532), .B(new_n533), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(new_n536), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(G127gat), .B(G155gat), .ZN(new_n542));
  XNOR2_X1  g341(.A(new_n542), .B(G211gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(new_n543), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n538), .A2(new_n545), .A3(new_n540), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n544), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n544), .A2(new_n548), .A3(new_n546), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(G232gat), .A2(G233gat), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT41), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT101), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(G85gat), .A3(G92gat), .ZN(new_n558));
  XNOR2_X1  g357(.A(new_n558), .B(KEYINPUT7), .ZN(new_n559));
  XOR2_X1   g358(.A(KEYINPUT102), .B(G85gat), .Z(new_n560));
  XOR2_X1   g359(.A(KEYINPUT103), .B(G92gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(G99gat), .A2(G106gat), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT8), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n559), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(G99gat), .B(G106gat), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G43gat), .B(G50gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g368(.A1(G29gat), .A2(G36gat), .ZN(new_n570));
  INV_X1    g369(.A(G29gat), .ZN(new_n571));
  INV_X1    g370(.A(G36gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n571), .A2(new_n572), .A3(KEYINPUT14), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT14), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n574), .B1(G29gat), .B2(G36gat), .ZN(new_n575));
  AND2_X1   g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n569), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT93), .ZN(new_n578));
  XNOR2_X1  g377(.A(new_n577), .B(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(KEYINPUT17), .ZN(new_n580));
  OR2_X1    g379(.A1(new_n568), .A2(KEYINPUT15), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n581), .A2(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n583));
  OR2_X1    g382(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n570), .B(KEYINPUT95), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n582), .A2(new_n583), .A3(new_n584), .A4(new_n585), .ZN(new_n586));
  AND3_X1   g385(.A1(new_n579), .A2(new_n580), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(new_n580), .B1(new_n579), .B2(new_n586), .ZN(new_n588));
  OR2_X1    g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT104), .ZN(new_n590));
  AOI21_X1  g389(.A(new_n567), .B1(new_n589), .B2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n579), .A2(new_n586), .ZN(new_n592));
  INV_X1    g391(.A(new_n567), .ZN(new_n593));
  AOI211_X1 g392(.A(new_n592), .B(new_n593), .C1(KEYINPUT104), .C2(new_n580), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n553), .B(new_n556), .C1(new_n591), .C2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(new_n594), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n587), .A2(new_n588), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n593), .B1(new_n597), .B2(KEYINPUT104), .ZN(new_n598));
  NAND4_X1  g397(.A1(new_n596), .A2(new_n598), .A3(new_n555), .A4(new_n554), .ZN(new_n599));
  XOR2_X1   g398(.A(G134gat), .B(G162gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT105), .ZN(new_n601));
  XNOR2_X1  g400(.A(G190gat), .B(G218gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  AND3_X1   g402(.A1(new_n595), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n603), .B1(new_n595), .B2(new_n599), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(G230gat), .A2(G233gat), .ZN(new_n608));
  INV_X1    g407(.A(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n567), .B(new_n530), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT10), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND4_X1  g411(.A1(new_n567), .A2(KEYINPUT10), .A3(new_n529), .A4(new_n519), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  OR2_X1    g414(.A1(new_n610), .A2(new_n608), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(G120gat), .B(G148gat), .ZN(new_n618));
  XNOR2_X1  g417(.A(G176gat), .B(G204gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n620), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n615), .A2(new_n616), .A3(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR3_X1   g423(.A1(new_n552), .A2(new_n607), .A3(new_n624), .ZN(new_n625));
  AND2_X1   g424(.A1(new_n506), .A2(new_n625), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n513), .B1(new_n587), .B2(new_n588), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n627), .A2(KEYINPUT96), .ZN(new_n628));
  INV_X1    g427(.A(new_n592), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n629), .A2(new_n513), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT96), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n631), .B(new_n513), .C1(new_n587), .C2(new_n588), .ZN(new_n632));
  AND3_X1   g431(.A1(new_n628), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G229gat), .A2(G233gat), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(KEYINPUT97), .A3(KEYINPUT18), .A4(new_n634), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n592), .B(new_n513), .ZN(new_n636));
  XNOR2_X1  g435(.A(new_n634), .B(KEYINPUT13), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT97), .ZN(new_n639));
  NAND4_X1  g438(.A1(new_n628), .A2(new_n634), .A3(new_n630), .A4(new_n632), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT18), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n639), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g441(.A1(new_n635), .A2(new_n638), .A3(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n640), .A2(new_n641), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  XNOR2_X1  g444(.A(G113gat), .B(G141gat), .ZN(new_n646));
  INV_X1    g445(.A(G197gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT11), .B(G169gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT12), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n643), .A2(new_n645), .A3(new_n652), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT98), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n643), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g454(.A1(new_n635), .A2(KEYINPUT98), .A3(new_n642), .A4(new_n638), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n655), .A2(new_n644), .A3(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n651), .B(KEYINPUT92), .Z(new_n658));
  AOI21_X1  g457(.A(new_n653), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n626), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n458), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT106), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  INV_X1    g463(.A(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n665), .A2(new_n474), .ZN(new_n666));
  XNOR2_X1  g465(.A(KEYINPUT16), .B(G8gat), .ZN(new_n667));
  OAI21_X1  g466(.A(KEYINPUT107), .B1(new_n666), .B2(new_n667), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT42), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n666), .A2(G8gat), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n668), .A2(KEYINPUT42), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n669), .A2(new_n670), .A3(new_n671), .ZN(G1325gat));
  INV_X1    g471(.A(new_n479), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n665), .A2(G15gat), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n293), .ZN(new_n675));
  AOI21_X1  g474(.A(G15gat), .B1(new_n665), .B2(new_n675), .ZN(new_n676));
  NOR2_X1   g475(.A1(new_n674), .A2(new_n676), .ZN(G1326gat));
  NOR2_X1   g476(.A1(new_n661), .A2(new_n453), .ZN(new_n678));
  XOR2_X1   g477(.A(KEYINPUT43), .B(G22gat), .Z(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(G1327gat));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n681));
  AOI211_X1 g480(.A(new_n681), .B(new_n606), .C1(new_n470), .C2(new_n505), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT108), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n470), .A2(new_n683), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n502), .A2(new_n475), .A3(new_n479), .ZN(new_n685));
  OAI211_X1 g484(.A(new_n443), .B(KEYINPUT108), .C1(new_n468), .C2(new_n469), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n684), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(new_n607), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n682), .B1(new_n688), .B2(new_n681), .ZN(new_n689));
  INV_X1    g488(.A(new_n624), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n660), .A2(new_n552), .A3(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  OAI21_X1  g492(.A(G29gat), .B1(new_n693), .B2(new_n458), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n606), .B(new_n691), .C1(new_n470), .C2(new_n505), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n695), .A2(new_n571), .A3(new_n473), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT45), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n694), .A2(new_n697), .ZN(G1328gat));
  INV_X1    g497(.A(KEYINPUT109), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n403), .A2(G36gat), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n699), .B1(new_n695), .B2(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n606), .B1(new_n470), .B2(new_n505), .ZN(new_n702));
  AND4_X1   g501(.A1(new_n699), .A2(new_n702), .A3(new_n692), .A4(new_n700), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT110), .ZN(new_n704));
  OAI22_X1  g503(.A1(new_n701), .A2(new_n703), .B1(new_n704), .B2(KEYINPUT46), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(KEYINPUT46), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g506(.A(new_n704), .B(KEYINPUT46), .C1(new_n701), .C2(new_n703), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n687), .B2(new_n607), .ZN(new_n710));
  NOR3_X1   g509(.A1(new_n710), .A2(new_n682), .A3(new_n691), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n572), .B1(new_n711), .B2(new_n474), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT111), .B1(new_n709), .B2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G36gat), .B1(new_n693), .B2(new_n403), .ZN(new_n714));
  INV_X1    g513(.A(KEYINPUT111), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n715), .A3(new_n707), .A4(new_n708), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(G1329gat));
  INV_X1    g516(.A(KEYINPUT112), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT47), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(G43gat), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n695), .A2(new_n721), .A3(new_n675), .ZN(new_n722));
  NOR4_X1   g521(.A1(new_n710), .A2(new_n479), .A3(new_n682), .A4(new_n691), .ZN(new_n723));
  OAI211_X1 g522(.A(new_n720), .B(new_n722), .C1(new_n723), .C2(new_n721), .ZN(new_n724));
  NOR2_X1   g523(.A1(new_n718), .A2(new_n719), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(new_n725), .ZN(new_n727));
  INV_X1    g526(.A(new_n722), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n688), .A2(new_n681), .ZN(new_n729));
  INV_X1    g528(.A(new_n682), .ZN(new_n730));
  NAND4_X1  g529(.A1(new_n729), .A2(new_n673), .A3(new_n730), .A4(new_n692), .ZN(new_n731));
  AOI21_X1  g530(.A(new_n728), .B1(new_n731), .B2(G43gat), .ZN(new_n732));
  AOI21_X1  g531(.A(new_n727), .B1(new_n732), .B2(new_n720), .ZN(new_n733));
  NOR2_X1   g532(.A1(new_n726), .A2(new_n733), .ZN(G1330gat));
  INV_X1    g533(.A(KEYINPUT113), .ZN(new_n735));
  NOR4_X1   g534(.A1(new_n710), .A2(new_n453), .A3(new_n682), .A4(new_n691), .ZN(new_n736));
  INV_X1    g535(.A(G50gat), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n735), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n695), .A2(new_n737), .A3(new_n373), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(new_n740));
  INV_X1    g539(.A(KEYINPUT48), .ZN(new_n741));
  NAND3_X1  g540(.A1(new_n738), .A2(new_n740), .A3(new_n741), .ZN(new_n742));
  OAI221_X1 g541(.A(new_n739), .B1(new_n735), .B2(KEYINPUT48), .C1(new_n736), .C2(new_n737), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(G1331gat));
  OAI21_X1  g543(.A(new_n624), .B1(new_n604), .B2(new_n605), .ZN(new_n745));
  INV_X1    g544(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n660), .A2(new_n552), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n687), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n749), .A2(new_n473), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g550(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n748), .A2(KEYINPUT114), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT114), .ZN(new_n754));
  NAND4_X1  g553(.A1(new_n687), .A2(new_n754), .A3(new_n746), .A4(new_n747), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n752), .B1(new_n756), .B2(new_n474), .ZN(new_n757));
  XOR2_X1   g556(.A(KEYINPUT49), .B(G64gat), .Z(new_n758));
  AOI211_X1 g557(.A(new_n403), .B(new_n758), .C1(new_n753), .C2(new_n755), .ZN(new_n759));
  OAI21_X1  g558(.A(KEYINPUT115), .B1(new_n757), .B2(new_n759), .ZN(new_n760));
  INV_X1    g559(.A(new_n758), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n756), .A2(new_n474), .A3(new_n761), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT115), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n403), .B1(new_n753), .B2(new_n755), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n762), .B(new_n763), .C1(new_n764), .C2(new_n752), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n760), .A2(new_n765), .ZN(G1333gat));
  NAND3_X1  g565(.A1(new_n749), .A2(new_n525), .A3(new_n675), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n479), .B1(new_n753), .B2(new_n755), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n767), .B1(new_n768), .B2(new_n525), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT50), .ZN(new_n770));
  XNOR2_X1  g569(.A(new_n769), .B(new_n770), .ZN(G1334gat));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n373), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n772), .B(G78gat), .ZN(G1335gat));
  INV_X1    g572(.A(new_n552), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n774), .A2(new_n660), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n689), .A2(new_n624), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(new_n776), .A2(new_n458), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT51), .ZN(new_n778));
  INV_X1    g577(.A(new_n775), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n778), .B1(new_n688), .B2(new_n779), .ZN(new_n780));
  NAND4_X1  g579(.A1(new_n687), .A2(KEYINPUT51), .A3(new_n607), .A4(new_n775), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n780), .A2(KEYINPUT116), .A3(new_n781), .ZN(new_n782));
  OR2_X1    g581(.A1(new_n781), .A2(KEYINPUT116), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n473), .A2(new_n560), .A3(new_n624), .ZN(new_n785));
  XNOR2_X1  g584(.A(new_n785), .B(KEYINPUT117), .ZN(new_n786));
  OAI22_X1  g585(.A1(new_n777), .A2(new_n560), .B1(new_n784), .B2(new_n786), .ZN(G1336gat));
  NOR3_X1   g586(.A1(new_n403), .A2(new_n690), .A3(G92gat), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n782), .A2(new_n783), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n689), .A2(new_n624), .A3(new_n474), .A4(new_n775), .ZN(new_n790));
  INV_X1    g589(.A(new_n561), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n780), .A2(new_n781), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n790), .A2(new_n791), .B1(new_n795), .B2(new_n788), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n794), .B1(new_n793), .B2(new_n796), .ZN(G1337gat));
  XNOR2_X1  g596(.A(KEYINPUT118), .B(G99gat), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n776), .B2(new_n479), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n293), .A2(new_n690), .A3(new_n798), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n799), .B1(new_n784), .B2(new_n800), .ZN(G1338gat));
  NOR3_X1   g600(.A1(new_n453), .A2(G106gat), .A3(new_n690), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n782), .A2(new_n783), .A3(new_n802), .ZN(new_n803));
  NAND4_X1  g602(.A1(new_n689), .A2(new_n624), .A3(new_n373), .A4(new_n775), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(G106gat), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT53), .ZN(new_n806));
  NAND3_X1  g605(.A1(new_n803), .A2(new_n805), .A3(new_n806), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n804), .A2(G106gat), .B1(new_n795), .B2(new_n802), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n807), .B1(new_n806), .B2(new_n808), .ZN(G1339gat));
  INV_X1    g608(.A(KEYINPUT55), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n612), .A2(new_n613), .A3(new_n609), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n811), .A2(KEYINPUT54), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n812), .A2(new_n614), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n612), .A2(new_n613), .ZN(new_n814));
  INV_X1    g613(.A(KEYINPUT54), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n814), .A2(new_n815), .A3(new_n608), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n620), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n810), .B1(new_n813), .B2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n622), .B1(new_n614), .B2(new_n815), .ZN(new_n819));
  OAI211_X1 g618(.A(new_n819), .B(KEYINPUT55), .C1(new_n614), .C2(new_n812), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n818), .A2(new_n623), .A3(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n659), .A2(new_n607), .A3(new_n821), .ZN(new_n822));
  OAI21_X1  g621(.A(new_n745), .B1(new_n606), .B2(new_n821), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n636), .A2(new_n637), .ZN(new_n824));
  OAI21_X1  g623(.A(new_n824), .B1(new_n633), .B2(new_n634), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n825), .A2(new_n650), .ZN(new_n826));
  INV_X1    g625(.A(new_n653), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n823), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n552), .B1(new_n822), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n625), .A2(new_n659), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n373), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  AND2_X1   g630(.A1(new_n831), .A2(new_n466), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n458), .A2(new_n474), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n203), .B1(new_n834), .B2(new_n659), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n829), .A2(new_n830), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n374), .A3(new_n833), .ZN(new_n837));
  XNOR2_X1  g636(.A(new_n837), .B(KEYINPUT119), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n660), .A2(G113gat), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  XNOR2_X1  g639(.A(new_n840), .B(KEYINPUT120), .ZN(G1340gat));
  OAI21_X1  g640(.A(G120gat), .B1(new_n838), .B2(new_n690), .ZN(new_n842));
  INV_X1    g641(.A(new_n834), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n843), .A2(new_n205), .A3(new_n624), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(new_n844), .ZN(G1341gat));
  NOR3_X1   g644(.A1(new_n838), .A2(new_n208), .A3(new_n552), .ZN(new_n846));
  OR3_X1    g645(.A1(new_n834), .A2(KEYINPUT121), .A3(new_n552), .ZN(new_n847));
  OAI21_X1  g646(.A(KEYINPUT121), .B1(new_n834), .B2(new_n552), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n208), .ZN(G1342gat));
  NAND3_X1  g649(.A1(new_n843), .A2(new_n209), .A3(new_n607), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n852));
  OAI21_X1  g651(.A(G134gat), .B1(new_n838), .B2(new_n606), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(KEYINPUT56), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n853), .A3(new_n854), .ZN(G1343gat));
  NAND2_X1  g654(.A1(new_n836), .A2(new_n373), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT57), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NAND3_X1  g657(.A1(new_n836), .A2(KEYINPUT57), .A3(new_n373), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n479), .A2(new_n833), .ZN(new_n861));
  INV_X1    g660(.A(new_n861), .ZN(new_n862));
  NAND4_X1  g661(.A1(new_n860), .A2(G141gat), .A3(new_n660), .A4(new_n862), .ZN(new_n863));
  NAND3_X1  g662(.A1(new_n836), .A2(new_n373), .A3(new_n862), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n320), .B1(new_n864), .B2(new_n659), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n863), .A2(new_n865), .ZN(new_n866));
  XOR2_X1   g665(.A(new_n866), .B(KEYINPUT58), .Z(G1344gat));
  NOR3_X1   g666(.A1(new_n864), .A2(G148gat), .A3(new_n690), .ZN(new_n868));
  XNOR2_X1  g667(.A(new_n861), .B(KEYINPUT122), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n860), .A2(new_n624), .A3(new_n869), .ZN(new_n870));
  AND2_X1   g669(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n860), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n873), .A2(new_n861), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n318), .B1(new_n874), .B2(new_n624), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n872), .B1(new_n875), .B2(KEYINPUT59), .ZN(G1345gat));
  NAND4_X1  g675(.A1(new_n860), .A2(G155gat), .A3(new_n774), .A4(new_n862), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n329), .B1(new_n864), .B2(new_n552), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  XNOR2_X1  g678(.A(new_n879), .B(KEYINPUT123), .ZN(G1346gat));
  NOR2_X1   g679(.A1(new_n606), .A2(new_n330), .ZN(new_n881));
  OR2_X1    g680(.A1(new_n864), .A2(new_n606), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n874), .A2(new_n881), .B1(new_n330), .B2(new_n882), .ZN(G1347gat));
  NOR2_X1   g682(.A1(new_n473), .A2(new_n403), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n832), .A2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n232), .A3(new_n660), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n831), .A2(new_n675), .A3(new_n884), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT124), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT124), .ZN(new_n890));
  NAND4_X1  g689(.A1(new_n831), .A2(new_n890), .A3(new_n675), .A4(new_n884), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  AND2_X1   g691(.A1(new_n892), .A2(new_n660), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n887), .B1(new_n893), .B2(new_n232), .ZN(G1348gat));
  AOI21_X1  g693(.A(G176gat), .B1(new_n886), .B2(new_n624), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n690), .A2(new_n233), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n892), .B2(new_n896), .ZN(G1349gat));
  NAND3_X1  g696(.A1(new_n889), .A2(new_n774), .A3(new_n891), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n898), .A2(G183gat), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n774), .A2(new_n228), .ZN(new_n900));
  OAI21_X1  g699(.A(new_n899), .B1(new_n885), .B2(new_n900), .ZN(new_n901));
  XNOR2_X1  g700(.A(new_n901), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g701(.A1(new_n886), .A2(new_n229), .A3(new_n607), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT61), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n892), .A2(new_n607), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G190gat), .ZN(new_n906));
  AOI211_X1 g705(.A(KEYINPUT61), .B(new_n229), .C1(new_n892), .C2(new_n607), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n903), .B1(new_n906), .B2(new_n907), .ZN(G1351gat));
  NAND2_X1  g707(.A1(new_n479), .A2(new_n884), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n856), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n647), .A3(new_n660), .ZN(new_n911));
  XOR2_X1   g710(.A(new_n911), .B(KEYINPUT125), .Z(new_n912));
  NOR3_X1   g711(.A1(new_n873), .A2(new_n659), .A3(new_n909), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n912), .B1(new_n647), .B2(new_n913), .ZN(G1352gat));
  INV_X1    g713(.A(G204gat), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n915), .A3(new_n624), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n917));
  INV_X1    g716(.A(KEYINPUT62), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n916), .A2(KEYINPUT126), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n918), .B1(new_n917), .B2(new_n919), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n873), .A2(new_n690), .A3(new_n909), .ZN(new_n922));
  OAI22_X1  g721(.A1(new_n920), .A2(new_n921), .B1(new_n915), .B2(new_n922), .ZN(G1353gat));
  NAND3_X1  g722(.A1(new_n910), .A2(new_n301), .A3(new_n774), .ZN(new_n924));
  INV_X1    g723(.A(new_n909), .ZN(new_n925));
  NAND4_X1  g724(.A1(new_n860), .A2(KEYINPUT127), .A3(new_n774), .A4(new_n925), .ZN(new_n926));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n836), .B2(new_n373), .ZN(new_n927));
  AOI211_X1 g726(.A(new_n857), .B(new_n453), .C1(new_n829), .C2(new_n830), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n774), .B(new_n925), .C1(new_n927), .C2(new_n928), .ZN(new_n929));
  INV_X1    g728(.A(KEYINPUT127), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n926), .A2(new_n931), .A3(G211gat), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT63), .ZN(new_n933));
  AND2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  OAI21_X1  g734(.A(new_n924), .B1(new_n934), .B2(new_n935), .ZN(G1354gat));
  NAND3_X1  g735(.A1(new_n910), .A2(new_n302), .A3(new_n607), .ZN(new_n937));
  NOR3_X1   g736(.A1(new_n873), .A2(new_n606), .A3(new_n909), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n937), .B1(new_n938), .B2(new_n302), .ZN(G1355gat));
endmodule


