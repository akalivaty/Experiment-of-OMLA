

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714;

  AND2_X2 U364 ( .A1(n495), .A2(n494), .ZN(n388) );
  NOR2_X2 U365 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X2 U366 ( .A(n353), .B(n563), .ZN(n579) );
  INV_X2 U367 ( .A(G953), .ZN(n701) );
  NOR2_X1 U368 ( .A1(n625), .A2(n626), .ZN(n634) );
  NOR2_X1 U369 ( .A1(n686), .A2(n685), .ZN(n372) );
  NOR2_X1 U370 ( .A1(n354), .A2(n711), .ZN(n365) );
  NAND2_X1 U371 ( .A1(n392), .A2(n391), .ZN(n354) );
  NAND2_X1 U372 ( .A1(n393), .A2(n394), .ZN(n391) );
  AND2_X1 U373 ( .A1(n396), .A2(n395), .ZN(n392) );
  NOR2_X1 U374 ( .A1(n508), .A2(n505), .ZN(n507) );
  XNOR2_X1 U375 ( .A(n371), .B(n499), .ZN(n503) );
  NAND2_X1 U376 ( .A1(n608), .A2(n397), .ZN(n395) );
  XNOR2_X1 U377 ( .A(n697), .B(n408), .ZN(n438) );
  XNOR2_X1 U378 ( .A(n407), .B(n406), .ZN(n697) );
  XNOR2_X1 U379 ( .A(n479), .B(G131), .ZN(n407) );
  XNOR2_X1 U380 ( .A(n398), .B(n412), .ZN(n448) );
  XNOR2_X1 U381 ( .A(n379), .B(G101), .ZN(n398) );
  XNOR2_X1 U382 ( .A(n355), .B(G902), .ZN(n454) );
  XNOR2_X1 U383 ( .A(n445), .B(G134), .ZN(n479) );
  XNOR2_X2 U384 ( .A(n439), .B(KEYINPUT33), .ZN(n649) );
  XNOR2_X2 U385 ( .A(n388), .B(n387), .ZN(n709) );
  NOR2_X2 U386 ( .A1(n546), .A2(n468), .ZN(n512) );
  INV_X1 U387 ( .A(G146), .ZN(n408) );
  XNOR2_X1 U388 ( .A(n560), .B(n404), .ZN(n641) );
  XNOR2_X1 U389 ( .A(n405), .B(KEYINPUT38), .ZN(n404) );
  INV_X1 U390 ( .A(KEYINPUT71), .ZN(n405) );
  XNOR2_X1 U391 ( .A(n456), .B(n455), .ZN(n457) );
  INV_X1 U392 ( .A(KEYINPUT85), .ZN(n455) );
  XNOR2_X1 U393 ( .A(G110), .B(G107), .ZN(n412) );
  XNOR2_X1 U394 ( .A(n416), .B(KEYINPUT20), .ZN(n429) );
  AND2_X1 U395 ( .A1(n349), .A2(n348), .ZN(n569) );
  XNOR2_X1 U396 ( .A(n614), .B(KEYINPUT80), .ZN(n348) );
  XNOR2_X1 U397 ( .A(n621), .B(n356), .ZN(n496) );
  INV_X1 U398 ( .A(KEYINPUT93), .ZN(n356) );
  XNOR2_X1 U399 ( .A(G119), .B(G137), .ZN(n419) );
  XOR2_X1 U400 ( .A(KEYINPUT4), .B(KEYINPUT64), .Z(n452) );
  XOR2_X1 U401 ( .A(G125), .B(G146), .Z(n443) );
  XNOR2_X1 U402 ( .A(n359), .B(KEYINPUT102), .ZN(n642) );
  NOR2_X1 U403 ( .A1(n641), .A2(n640), .ZN(n645) );
  AND2_X1 U404 ( .A1(n642), .A2(n496), .ZN(n358) );
  XNOR2_X1 U405 ( .A(n512), .B(KEYINPUT0), .ZN(n497) );
  NAND2_X1 U406 ( .A1(n562), .A2(n561), .ZN(n353) );
  NOR2_X1 U407 ( .A1(n535), .A2(n640), .ZN(n352) );
  NAND2_X1 U408 ( .A1(n503), .A2(n502), .ZN(n508) );
  XNOR2_X1 U409 ( .A(n378), .B(n377), .ZN(n546) );
  INV_X1 U410 ( .A(KEYINPUT19), .ZN(n377) );
  OR2_X1 U411 ( .A1(n667), .A2(G902), .ZN(n389) );
  INV_X1 U412 ( .A(G472), .ZN(n399) );
  XNOR2_X1 U413 ( .A(n451), .B(n364), .ZN(n687) );
  XNOR2_X1 U414 ( .A(n448), .B(n447), .ZN(n364) );
  INV_X1 U415 ( .A(G122), .ZN(n449) );
  NAND2_X1 U416 ( .A1(n454), .A2(G475), .ZN(n401) );
  XNOR2_X1 U417 ( .A(n687), .B(n360), .ZN(n663) );
  XNOR2_X1 U418 ( .A(n362), .B(n361), .ZN(n360) );
  XNOR2_X1 U419 ( .A(n444), .B(n446), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n363), .B(n442), .ZN(n362) );
  NAND2_X1 U421 ( .A1(n454), .A2(G210), .ZN(n402) );
  NOR2_X1 U422 ( .A1(G952), .A2(n701), .ZN(n685) );
  XNOR2_X1 U423 ( .A(n357), .B(n417), .ZN(n621) );
  NAND2_X1 U424 ( .A1(n429), .A2(G221), .ZN(n357) );
  XNOR2_X1 U425 ( .A(n450), .B(G101), .ZN(n435) );
  INV_X1 U426 ( .A(KEYINPUT104), .ZN(n384) );
  OR2_X1 U427 ( .A1(n589), .A2(G902), .ZN(n346) );
  INV_X1 U428 ( .A(KEYINPUT16), .ZN(n447) );
  XNOR2_X1 U429 ( .A(n434), .B(n350), .ZN(n450) );
  XNOR2_X1 U430 ( .A(G119), .B(KEYINPUT3), .ZN(n434) );
  XNOR2_X1 U431 ( .A(n351), .B(G116), .ZN(n350) );
  INV_X1 U432 ( .A(G113), .ZN(n351) );
  XNOR2_X1 U433 ( .A(n369), .B(n420), .ZN(n422) );
  XNOR2_X1 U434 ( .A(n419), .B(n370), .ZN(n369) );
  INV_X1 U435 ( .A(KEYINPUT24), .ZN(n370) );
  XNOR2_X1 U436 ( .A(G128), .B(G110), .ZN(n421) );
  XNOR2_X1 U437 ( .A(KEYINPUT100), .B(KEYINPUT9), .ZN(n474) );
  XOR2_X1 U438 ( .A(KEYINPUT98), .B(KEYINPUT7), .Z(n475) );
  XNOR2_X1 U439 ( .A(G107), .B(G122), .ZN(n472) );
  XOR2_X1 U440 ( .A(KEYINPUT99), .B(G116), .Z(n473) );
  XOR2_X1 U441 ( .A(KEYINPUT8), .B(KEYINPUT66), .Z(n425) );
  XNOR2_X1 U442 ( .A(G113), .B(KEYINPUT11), .ZN(n485) );
  XNOR2_X1 U443 ( .A(G104), .B(G122), .ZN(n483) );
  XNOR2_X1 U444 ( .A(n438), .B(n390), .ZN(n667) );
  XNOR2_X1 U445 ( .A(n414), .B(n411), .ZN(n390) );
  XNOR2_X1 U446 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U447 ( .A(n453), .B(n443), .ZN(n363) );
  XNOR2_X1 U448 ( .A(KEYINPUT84), .B(KEYINPUT18), .ZN(n440) );
  INV_X1 U449 ( .A(KEYINPUT15), .ZN(n355) );
  AND2_X1 U450 ( .A1(n585), .A2(n584), .ZN(n700) );
  XNOR2_X1 U451 ( .A(n565), .B(n564), .ZN(n619) );
  NAND2_X1 U452 ( .A1(n645), .A2(n642), .ZN(n564) );
  INV_X1 U453 ( .A(KEYINPUT40), .ZN(n397) );
  AND2_X1 U454 ( .A1(n552), .A2(n341), .ZN(n562) );
  INV_X1 U455 ( .A(n554), .ZN(n555) );
  NAND2_X1 U456 ( .A1(n497), .A2(n358), .ZN(n371) );
  INV_X1 U457 ( .A(KEYINPUT22), .ZN(n498) );
  XNOR2_X1 U458 ( .A(n493), .B(n375), .ZN(n520) );
  XNOR2_X1 U459 ( .A(n376), .B(G475), .ZN(n375) );
  INV_X1 U460 ( .A(KEYINPUT13), .ZN(n376) );
  NOR2_X1 U461 ( .A1(n513), .A2(n626), .ZN(n518) );
  NAND2_X1 U462 ( .A1(n454), .A2(G217), .ZN(n400) );
  NAND2_X1 U463 ( .A1(n540), .A2(n539), .ZN(n614) );
  INV_X1 U464 ( .A(KEYINPUT35), .ZN(n387) );
  NOR2_X1 U465 ( .A1(n566), .A2(n546), .ZN(n547) );
  XNOR2_X1 U466 ( .A(n368), .B(n367), .ZN(n712) );
  INV_X1 U467 ( .A(KEYINPUT103), .ZN(n367) );
  NOR2_X1 U468 ( .A1(n592), .A2(n685), .ZN(n366) );
  NOR2_X1 U469 ( .A1(n677), .A2(n685), .ZN(n373) );
  NOR2_X1 U470 ( .A1(n666), .A2(n685), .ZN(n374) );
  AND2_X1 U471 ( .A1(n553), .A2(n555), .ZN(n341) );
  AND2_X1 U472 ( .A1(KEYINPUT77), .A2(n606), .ZN(n342) );
  AND2_X1 U473 ( .A1(n489), .A2(G210), .ZN(n343) );
  XOR2_X1 U474 ( .A(KEYINPUT95), .B(G472), .Z(n344) );
  OR2_X1 U475 ( .A1(n587), .A2(n399), .ZN(n345) );
  XNOR2_X2 U476 ( .A(n346), .B(n344), .ZN(n549) );
  XNOR2_X1 U477 ( .A(n438), .B(n347), .ZN(n589) );
  XNOR2_X1 U478 ( .A(n437), .B(n343), .ZN(n347) );
  NOR2_X1 U479 ( .A1(n559), .A2(n342), .ZN(n349) );
  NAND2_X1 U480 ( .A1(n352), .A2(n560), .ZN(n537) );
  NAND2_X1 U481 ( .A1(n352), .A2(n625), .ZN(n580) );
  XNOR2_X1 U482 ( .A(n354), .B(n714), .ZN(G33) );
  NOR2_X1 U483 ( .A1(n521), .A2(n523), .ZN(n359) );
  XNOR2_X1 U484 ( .A(n591), .B(n590), .ZN(n592) );
  XNOR2_X1 U485 ( .A(n665), .B(n664), .ZN(n666) );
  XNOR2_X1 U486 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U487 ( .A(n683), .B(n684), .ZN(n686) );
  XNOR2_X1 U488 ( .A(n365), .B(KEYINPUT46), .ZN(n568) );
  XNOR2_X1 U489 ( .A(n380), .B(KEYINPUT45), .ZN(n689) );
  XNOR2_X1 U490 ( .A(n385), .B(n384), .ZN(n383) );
  XNOR2_X1 U491 ( .A(n366), .B(n593), .ZN(G57) );
  NAND2_X1 U492 ( .A1(n511), .A2(n510), .ZN(n368) );
  XNOR2_X2 U493 ( .A(n433), .B(n432), .ZN(n620) );
  XNOR2_X1 U494 ( .A(n372), .B(KEYINPUT122), .ZN(G66) );
  XNOR2_X1 U495 ( .A(n373), .B(KEYINPUT60), .ZN(G60) );
  XNOR2_X1 U496 ( .A(n374), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U497 ( .A1(n536), .A2(n548), .ZN(n378) );
  XNOR2_X1 U498 ( .A(n458), .B(n457), .ZN(n536) );
  XNOR2_X2 U499 ( .A(G104), .B(KEYINPUT72), .ZN(n379) );
  NAND2_X1 U500 ( .A1(n383), .A2(n381), .ZN(n380) );
  XNOR2_X1 U501 ( .A(n382), .B(KEYINPUT44), .ZN(n381) );
  NOR2_X2 U502 ( .A1(n386), .A2(n709), .ZN(n382) );
  NAND2_X1 U503 ( .A1(n526), .A2(n712), .ZN(n385) );
  NAND2_X1 U504 ( .A1(n599), .A2(n713), .ZN(n386) );
  XNOR2_X2 U505 ( .A(n389), .B(G469), .ZN(n553) );
  AND2_X1 U506 ( .A1(n562), .A2(n560), .ZN(n556) );
  INV_X1 U507 ( .A(n579), .ZN(n393) );
  NAND2_X1 U508 ( .A1(n579), .A2(n397), .ZN(n396) );
  NOR2_X1 U509 ( .A1(n608), .A2(n397), .ZN(n394) );
  OR2_X2 U510 ( .A1(n618), .A2(n345), .ZN(n591) );
  OR2_X2 U511 ( .A1(n618), .A2(n401), .ZN(n676) );
  OR2_X2 U512 ( .A1(n618), .A2(n402), .ZN(n665) );
  NOR2_X1 U513 ( .A1(n618), .A2(n587), .ZN(n403) );
  OR2_X2 U514 ( .A1(n618), .A2(n400), .ZN(n683) );
  NAND2_X1 U515 ( .A1(n403), .A2(G469), .ZN(n670) );
  NAND2_X1 U516 ( .A1(n403), .A2(G478), .ZN(n681) );
  INV_X1 U517 ( .A(n452), .ZN(n453) );
  XNOR2_X2 U518 ( .A(n553), .B(n415), .ZN(n625) );
  XOR2_X2 U519 ( .A(n633), .B(KEYINPUT6), .Z(n534) );
  INV_X1 U520 ( .A(KEYINPUT74), .ZN(n409) );
  OR2_X1 U521 ( .A1(G902), .A2(G237), .ZN(n459) );
  INV_X1 U522 ( .A(n445), .ZN(n446) );
  INV_X1 U523 ( .A(n617), .ZN(n583) );
  XNOR2_X1 U524 ( .A(n448), .B(n413), .ZN(n414) );
  XNOR2_X1 U525 ( .A(n498), .B(KEYINPUT70), .ZN(n499) );
  NOR2_X1 U526 ( .A1(n615), .A2(n583), .ZN(n584) );
  XNOR2_X1 U527 ( .A(n674), .B(n673), .ZN(n675) );
  XNOR2_X1 U528 ( .A(KEYINPUT32), .B(KEYINPUT75), .ZN(n506) );
  XNOR2_X1 U529 ( .A(n507), .B(n506), .ZN(n713) );
  XNOR2_X2 U530 ( .A(G128), .B(G143), .ZN(n445) );
  XOR2_X1 U531 ( .A(G137), .B(n452), .Z(n406) );
  NAND2_X1 U532 ( .A1(G227), .A2(n701), .ZN(n410) );
  XNOR2_X1 U533 ( .A(G140), .B(KEYINPUT91), .ZN(n413) );
  XNOR2_X1 U534 ( .A(KEYINPUT1), .B(KEYINPUT65), .ZN(n415) );
  XOR2_X1 U535 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n417) );
  INV_X1 U536 ( .A(n454), .ZN(n587) );
  NAND2_X1 U537 ( .A1(G234), .A2(n587), .ZN(n416) );
  XNOR2_X1 U538 ( .A(n443), .B(KEYINPUT10), .ZN(n418) );
  XNOR2_X1 U539 ( .A(n418), .B(G140), .ZN(n698) );
  XOR2_X1 U540 ( .A(KEYINPUT67), .B(KEYINPUT23), .Z(n420) );
  XNOR2_X1 U541 ( .A(n422), .B(n421), .ZN(n423) );
  XOR2_X1 U542 ( .A(n698), .B(n423), .Z(n428) );
  NAND2_X1 U543 ( .A1(G234), .A2(n701), .ZN(n424) );
  XNOR2_X1 U544 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U545 ( .A(KEYINPUT79), .B(n426), .Z(n471) );
  NAND2_X1 U546 ( .A1(n471), .A2(G221), .ZN(n427) );
  XOR2_X1 U547 ( .A(n428), .B(n427), .Z(n684) );
  NOR2_X1 U548 ( .A1(n684), .A2(G902), .ZN(n433) );
  XOR2_X1 U549 ( .A(KEYINPUT25), .B(KEYINPUT73), .Z(n431) );
  NAND2_X1 U550 ( .A1(n429), .A2(G217), .ZN(n430) );
  XNOR2_X1 U551 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U552 ( .A1(n496), .A2(n620), .ZN(n626) );
  XOR2_X1 U553 ( .A(KEYINPUT94), .B(KEYINPUT5), .Z(n436) );
  XNOR2_X1 U554 ( .A(n436), .B(n435), .ZN(n437) );
  NOR2_X1 U555 ( .A1(G953), .A2(G237), .ZN(n489) );
  BUF_X4 U556 ( .A(n549), .Z(n633) );
  NAND2_X1 U557 ( .A1(n634), .A2(n534), .ZN(n439) );
  XOR2_X1 U558 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n441) );
  XNOR2_X1 U559 ( .A(n441), .B(n440), .ZN(n442) );
  NAND2_X1 U560 ( .A1(G224), .A2(n701), .ZN(n444) );
  XNOR2_X1 U561 ( .A(n450), .B(n449), .ZN(n451) );
  NOR2_X1 U562 ( .A1(n454), .A2(n663), .ZN(n458) );
  NAND2_X1 U563 ( .A1(G210), .A2(n459), .ZN(n456) );
  NAND2_X1 U564 ( .A1(G214), .A2(n459), .ZN(n460) );
  XNOR2_X1 U565 ( .A(KEYINPUT86), .B(n460), .ZN(n548) );
  NAND2_X1 U566 ( .A1(G237), .A2(G234), .ZN(n461) );
  XNOR2_X1 U567 ( .A(n461), .B(KEYINPUT87), .ZN(n462) );
  XOR2_X1 U568 ( .A(KEYINPUT14), .B(n462), .Z(n464) );
  NAND2_X1 U569 ( .A1(G902), .A2(n464), .ZN(n527) );
  NOR2_X1 U570 ( .A1(G898), .A2(n701), .ZN(n463) );
  XNOR2_X1 U571 ( .A(KEYINPUT89), .B(n463), .ZN(n688) );
  NOR2_X1 U572 ( .A1(n527), .A2(n688), .ZN(n466) );
  NAND2_X1 U573 ( .A1(G952), .A2(n464), .ZN(n654) );
  NOR2_X1 U574 ( .A1(G953), .A2(n654), .ZN(n465) );
  XNOR2_X1 U575 ( .A(KEYINPUT88), .B(n465), .ZN(n530) );
  NOR2_X1 U576 ( .A1(n466), .A2(n530), .ZN(n467) );
  XNOR2_X1 U577 ( .A(n467), .B(KEYINPUT90), .ZN(n468) );
  NAND2_X1 U578 ( .A1(n649), .A2(n497), .ZN(n470) );
  XNOR2_X1 U579 ( .A(KEYINPUT69), .B(KEYINPUT34), .ZN(n469) );
  XNOR2_X1 U580 ( .A(n470), .B(n469), .ZN(n495) );
  NAND2_X1 U581 ( .A1(G217), .A2(n471), .ZN(n481) );
  XNOR2_X1 U582 ( .A(n473), .B(n472), .ZN(n477) );
  XNOR2_X1 U583 ( .A(n475), .B(n474), .ZN(n476) );
  XNOR2_X1 U584 ( .A(n477), .B(n476), .ZN(n478) );
  XOR2_X1 U585 ( .A(n479), .B(n478), .Z(n480) );
  XNOR2_X1 U586 ( .A(n481), .B(n480), .ZN(n679) );
  NOR2_X1 U587 ( .A1(G902), .A2(n679), .ZN(n482) );
  XOR2_X1 U588 ( .A(G478), .B(n482), .Z(n521) );
  XOR2_X1 U589 ( .A(G131), .B(G143), .Z(n484) );
  XNOR2_X1 U590 ( .A(n484), .B(n483), .ZN(n488) );
  XOR2_X1 U591 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n486) );
  XNOR2_X1 U592 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U593 ( .A(n488), .B(n487), .Z(n491) );
  NAND2_X1 U594 ( .A1(n489), .A2(G214), .ZN(n490) );
  XNOR2_X1 U595 ( .A(n491), .B(n490), .ZN(n492) );
  XNOR2_X1 U596 ( .A(n492), .B(n698), .ZN(n674) );
  NOR2_X1 U597 ( .A1(G902), .A2(n674), .ZN(n493) );
  INV_X1 U598 ( .A(n520), .ZN(n523) );
  NAND2_X1 U599 ( .A1(n521), .A2(n523), .ZN(n558) );
  INV_X1 U600 ( .A(n558), .ZN(n494) );
  INV_X1 U601 ( .A(n620), .ZN(n509) );
  NAND2_X1 U602 ( .A1(n509), .A2(n503), .ZN(n500) );
  NOR2_X1 U603 ( .A1(n633), .A2(n500), .ZN(n501) );
  NAND2_X1 U604 ( .A1(n625), .A2(n501), .ZN(n599) );
  INV_X1 U605 ( .A(n534), .ZN(n502) );
  NOR2_X1 U606 ( .A1(n625), .A2(n620), .ZN(n504) );
  XNOR2_X1 U607 ( .A(n504), .B(KEYINPUT105), .ZN(n505) );
  XNOR2_X1 U608 ( .A(n508), .B(KEYINPUT81), .ZN(n511) );
  INV_X1 U609 ( .A(n625), .ZN(n539) );
  NOR2_X1 U610 ( .A1(n509), .A2(n539), .ZN(n510) );
  XOR2_X1 U611 ( .A(KEYINPUT0), .B(n512), .Z(n513) );
  NAND2_X1 U612 ( .A1(n633), .A2(n518), .ZN(n514) );
  NOR2_X1 U613 ( .A1(n514), .A2(n625), .ZN(n515) );
  XNOR2_X1 U614 ( .A(n515), .B(KEYINPUT31), .ZN(n610) );
  INV_X1 U615 ( .A(n553), .ZN(n516) );
  NOR2_X1 U616 ( .A1(n516), .A2(n633), .ZN(n517) );
  NAND2_X1 U617 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U618 ( .A(KEYINPUT96), .B(n519), .ZN(n595) );
  NAND2_X1 U619 ( .A1(n610), .A2(n595), .ZN(n525) );
  NAND2_X1 U620 ( .A1(n521), .A2(n520), .ZN(n611) );
  INV_X1 U621 ( .A(n611), .ZN(n600) );
  INV_X1 U622 ( .A(n521), .ZN(n522) );
  NAND2_X1 U623 ( .A1(n523), .A2(n522), .ZN(n608) );
  INV_X1 U624 ( .A(n608), .ZN(n605) );
  NOR2_X1 U625 ( .A1(n600), .A2(n605), .ZN(n524) );
  XNOR2_X1 U626 ( .A(n524), .B(KEYINPUT101), .ZN(n644) );
  NAND2_X1 U627 ( .A1(n525), .A2(n644), .ZN(n526) );
  XOR2_X1 U628 ( .A(KEYINPUT110), .B(KEYINPUT36), .Z(n538) );
  INV_X1 U629 ( .A(n548), .ZN(n640) );
  OR2_X1 U630 ( .A1(n701), .A2(n527), .ZN(n528) );
  XNOR2_X1 U631 ( .A(KEYINPUT106), .B(n528), .ZN(n529) );
  NOR2_X1 U632 ( .A1(G900), .A2(n529), .ZN(n531) );
  NOR2_X1 U633 ( .A1(n531), .A2(n530), .ZN(n554) );
  NOR2_X1 U634 ( .A1(n554), .A2(n620), .ZN(n532) );
  NAND2_X1 U635 ( .A1(n621), .A2(n532), .ZN(n541) );
  NOR2_X1 U636 ( .A1(n608), .A2(n541), .ZN(n533) );
  NAND2_X1 U637 ( .A1(n534), .A2(n533), .ZN(n535) );
  BUF_X1 U638 ( .A(n536), .Z(n560) );
  XNOR2_X1 U639 ( .A(n538), .B(n537), .ZN(n540) );
  XOR2_X1 U640 ( .A(KEYINPUT28), .B(KEYINPUT108), .Z(n544) );
  INV_X1 U641 ( .A(n541), .ZN(n542) );
  NAND2_X1 U642 ( .A1(n542), .A2(n633), .ZN(n543) );
  XNOR2_X1 U643 ( .A(n544), .B(n543), .ZN(n545) );
  NAND2_X1 U644 ( .A1(n553), .A2(n545), .ZN(n566) );
  XNOR2_X1 U645 ( .A(KEYINPUT76), .B(n547), .ZN(n606) );
  INV_X1 U646 ( .A(n560), .ZN(n581) );
  NAND2_X1 U647 ( .A1(n549), .A2(n548), .ZN(n550) );
  XNOR2_X1 U648 ( .A(KEYINPUT30), .B(n550), .ZN(n551) );
  NOR2_X1 U649 ( .A1(n626), .A2(n551), .ZN(n552) );
  XNOR2_X1 U650 ( .A(n556), .B(KEYINPUT107), .ZN(n557) );
  NOR2_X1 U651 ( .A1(n558), .A2(n557), .ZN(n603) );
  XNOR2_X1 U652 ( .A(n603), .B(KEYINPUT78), .ZN(n559) );
  XOR2_X1 U653 ( .A(KEYINPUT68), .B(KEYINPUT39), .Z(n563) );
  INV_X1 U654 ( .A(n641), .ZN(n561) );
  XNOR2_X1 U655 ( .A(KEYINPUT109), .B(KEYINPUT41), .ZN(n565) );
  NOR2_X1 U656 ( .A1(n619), .A2(n566), .ZN(n567) );
  XNOR2_X1 U657 ( .A(n567), .B(KEYINPUT42), .ZN(n711) );
  NAND2_X1 U658 ( .A1(n569), .A2(n568), .ZN(n577) );
  NAND2_X1 U659 ( .A1(n606), .A2(n644), .ZN(n570) );
  XNOR2_X1 U660 ( .A(n570), .B(KEYINPUT47), .ZN(n572) );
  INV_X1 U661 ( .A(KEYINPUT77), .ZN(n571) );
  NAND2_X1 U662 ( .A1(n572), .A2(n571), .ZN(n575) );
  NAND2_X1 U663 ( .A1(KEYINPUT47), .A2(n644), .ZN(n573) );
  NAND2_X1 U664 ( .A1(n573), .A2(KEYINPUT77), .ZN(n574) );
  NAND2_X1 U665 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U666 ( .A(n578), .B(KEYINPUT48), .ZN(n585) );
  NOR2_X1 U667 ( .A1(n579), .A2(n611), .ZN(n615) );
  XNOR2_X1 U668 ( .A(n580), .B(KEYINPUT43), .ZN(n582) );
  NAND2_X1 U669 ( .A1(n582), .A2(n581), .ZN(n617) );
  AND2_X2 U670 ( .A1(n689), .A2(n700), .ZN(n586) );
  XNOR2_X2 U671 ( .A(n586), .B(KEYINPUT2), .ZN(n618) );
  XOR2_X1 U672 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n588) );
  XNOR2_X1 U673 ( .A(n589), .B(n588), .ZN(n590) );
  XNOR2_X1 U674 ( .A(KEYINPUT83), .B(KEYINPUT63), .ZN(n593) );
  NOR2_X1 U675 ( .A1(n595), .A2(n608), .ZN(n594) );
  XOR2_X1 U676 ( .A(G104), .B(n594), .Z(G6) );
  NOR2_X1 U677 ( .A1(n595), .A2(n611), .ZN(n597) );
  XNOR2_X1 U678 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n596) );
  XNOR2_X1 U679 ( .A(n597), .B(n596), .ZN(n598) );
  XNOR2_X1 U680 ( .A(G107), .B(n598), .ZN(G9) );
  XNOR2_X1 U681 ( .A(G110), .B(n599), .ZN(G12) );
  XOR2_X1 U682 ( .A(G128), .B(KEYINPUT29), .Z(n602) );
  NAND2_X1 U683 ( .A1(n600), .A2(n606), .ZN(n601) );
  XNOR2_X1 U684 ( .A(n602), .B(n601), .ZN(G30) );
  XOR2_X1 U685 ( .A(G143), .B(n603), .Z(n604) );
  XNOR2_X1 U686 ( .A(KEYINPUT112), .B(n604), .ZN(G45) );
  NAND2_X1 U687 ( .A1(n606), .A2(n605), .ZN(n607) );
  XNOR2_X1 U688 ( .A(n607), .B(G146), .ZN(G48) );
  NOR2_X1 U689 ( .A1(n608), .A2(n610), .ZN(n609) );
  XOR2_X1 U690 ( .A(G113), .B(n609), .Z(G15) );
  NOR2_X1 U691 ( .A1(n611), .A2(n610), .ZN(n612) );
  XOR2_X1 U692 ( .A(G116), .B(n612), .Z(G18) );
  XOR2_X1 U693 ( .A(G125), .B(KEYINPUT37), .Z(n613) );
  XNOR2_X1 U694 ( .A(n614), .B(n613), .ZN(G27) );
  XOR2_X1 U695 ( .A(G134), .B(n615), .Z(G36) );
  XOR2_X1 U696 ( .A(G140), .B(KEYINPUT113), .Z(n616) );
  XNOR2_X1 U697 ( .A(n617), .B(n616), .ZN(G42) );
  NAND2_X1 U698 ( .A1(n701), .A2(n618), .ZN(n660) );
  INV_X1 U699 ( .A(n619), .ZN(n639) );
  AND2_X1 U700 ( .A1(n639), .A2(n649), .ZN(n657) );
  NOR2_X1 U701 ( .A1(n621), .A2(n620), .ZN(n623) );
  XNOR2_X1 U702 ( .A(KEYINPUT115), .B(KEYINPUT49), .ZN(n622) );
  XNOR2_X1 U703 ( .A(n623), .B(n622), .ZN(n624) );
  XOR2_X1 U704 ( .A(KEYINPUT114), .B(n624), .Z(n630) );
  NAND2_X1 U705 ( .A1(n626), .A2(n625), .ZN(n627) );
  XNOR2_X1 U706 ( .A(n627), .B(KEYINPUT116), .ZN(n628) );
  XNOR2_X1 U707 ( .A(KEYINPUT50), .B(n628), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  NOR2_X1 U709 ( .A1(n633), .A2(n631), .ZN(n632) );
  XNOR2_X1 U710 ( .A(n632), .B(KEYINPUT117), .ZN(n636) );
  NAND2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(n637) );
  XOR2_X1 U713 ( .A(KEYINPUT51), .B(n637), .Z(n638) );
  NAND2_X1 U714 ( .A1(n639), .A2(n638), .ZN(n651) );
  NAND2_X1 U715 ( .A1(n641), .A2(n640), .ZN(n643) );
  NAND2_X1 U716 ( .A1(n643), .A2(n642), .ZN(n647) );
  NAND2_X1 U717 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U718 ( .A1(n647), .A2(n646), .ZN(n648) );
  NAND2_X1 U719 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U720 ( .A1(n651), .A2(n650), .ZN(n653) );
  XOR2_X1 U721 ( .A(KEYINPUT118), .B(KEYINPUT52), .Z(n652) );
  XNOR2_X1 U722 ( .A(n653), .B(n652), .ZN(n655) );
  NOR2_X1 U723 ( .A1(n655), .A2(n654), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  XNOR2_X1 U725 ( .A(n658), .B(KEYINPUT119), .ZN(n659) );
  NOR2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U727 ( .A(KEYINPUT53), .B(n661), .ZN(G75) );
  XOR2_X1 U728 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n662) );
  XNOR2_X1 U729 ( .A(n663), .B(n662), .ZN(n664) );
  XNOR2_X1 U730 ( .A(KEYINPUT58), .B(KEYINPUT120), .ZN(n669) );
  XNOR2_X1 U731 ( .A(n667), .B(KEYINPUT57), .ZN(n668) );
  XNOR2_X1 U732 ( .A(n669), .B(n668), .ZN(n671) );
  XOR2_X1 U733 ( .A(n671), .B(n670), .Z(n672) );
  NOR2_X1 U734 ( .A1(n685), .A2(n672), .ZN(G54) );
  INV_X1 U735 ( .A(KEYINPUT59), .ZN(n673) );
  INV_X1 U736 ( .A(KEYINPUT121), .ZN(n678) );
  XNOR2_X1 U737 ( .A(n679), .B(n678), .ZN(n680) );
  XNOR2_X1 U738 ( .A(n681), .B(n680), .ZN(n682) );
  NOR2_X1 U739 ( .A1(n685), .A2(n682), .ZN(G63) );
  NAND2_X1 U740 ( .A1(n688), .A2(n687), .ZN(n696) );
  NAND2_X1 U741 ( .A1(n689), .A2(n701), .ZN(n690) );
  XOR2_X1 U742 ( .A(KEYINPUT123), .B(n690), .Z(n694) );
  NAND2_X1 U743 ( .A1(G953), .A2(G224), .ZN(n691) );
  XNOR2_X1 U744 ( .A(KEYINPUT61), .B(n691), .ZN(n692) );
  NAND2_X1 U745 ( .A1(n692), .A2(G898), .ZN(n693) );
  NAND2_X1 U746 ( .A1(n694), .A2(n693), .ZN(n695) );
  XOR2_X1 U747 ( .A(n696), .B(n695), .Z(G69) );
  XOR2_X1 U748 ( .A(n698), .B(n697), .Z(n699) );
  XOR2_X1 U749 ( .A(KEYINPUT124), .B(n699), .Z(n703) );
  XOR2_X1 U750 ( .A(n703), .B(n700), .Z(n702) );
  NAND2_X1 U751 ( .A1(n702), .A2(n701), .ZN(n708) );
  XNOR2_X1 U752 ( .A(G227), .B(n703), .ZN(n704) );
  NAND2_X1 U753 ( .A1(n704), .A2(G900), .ZN(n705) );
  XOR2_X1 U754 ( .A(KEYINPUT125), .B(n705), .Z(n706) );
  NAND2_X1 U755 ( .A1(G953), .A2(n706), .ZN(n707) );
  NAND2_X1 U756 ( .A1(n708), .A2(n707), .ZN(G72) );
  XOR2_X1 U757 ( .A(n709), .B(G122), .Z(G24) );
  XOR2_X1 U758 ( .A(G137), .B(KEYINPUT126), .Z(n710) );
  XNOR2_X1 U759 ( .A(n711), .B(n710), .ZN(G39) );
  XNOR2_X1 U760 ( .A(n712), .B(G101), .ZN(G3) );
  XNOR2_X1 U761 ( .A(G119), .B(n713), .ZN(G21) );
  XNOR2_X1 U762 ( .A(G131), .B(KEYINPUT127), .ZN(n714) );
endmodule

