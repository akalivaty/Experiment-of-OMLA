//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n484, new_n485, new_n486,
    new_n487, new_n488, new_n489, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n540, new_n541, new_n542, new_n543, new_n544, new_n545, new_n546,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n568, new_n570, new_n571, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n579, new_n580, new_n582,
    new_n583, new_n584, new_n586, new_n587, new_n588, new_n589, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n621, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(new_n436));
  XNOR2_X1  g011(.A(new_n436), .B(KEYINPUT65), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  AND2_X1   g017(.A1(G2072), .A2(G2078), .ZN(new_n443));
  NAND3_X1  g018(.A1(new_n443), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR4_X1   g029(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n454), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n454), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  XNOR2_X1  g038(.A(new_n463), .B(KEYINPUT68), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n466));
  XNOR2_X1  g041(.A(KEYINPUT3), .B(G2104), .ZN(new_n467));
  AOI21_X1  g042(.A(new_n466), .B1(new_n467), .B2(G125), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  AND4_X1   g047(.A1(new_n466), .A2(new_n470), .A3(new_n472), .A4(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n465), .B1(new_n468), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NOR2_X1   g050(.A1(new_n469), .A2(G2105), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G101), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT69), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n479), .A2(new_n469), .A3(KEYINPUT3), .ZN(new_n480));
  AND2_X1   g055(.A1(new_n480), .A2(new_n472), .ZN(new_n481));
  INV_X1    g056(.A(KEYINPUT70), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT69), .B1(new_n471), .B2(G2104), .ZN(new_n483));
  INV_X1    g058(.A(G137), .ZN(new_n484));
  NOR2_X1   g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  NAND4_X1  g060(.A1(new_n481), .A2(new_n482), .A3(new_n483), .A4(new_n485), .ZN(new_n486));
  NAND4_X1  g061(.A1(new_n483), .A2(new_n480), .A3(new_n472), .A4(new_n485), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n488));
  AOI21_X1  g063(.A(new_n478), .B1(new_n486), .B2(new_n488), .ZN(new_n489));
  AND2_X1   g064(.A1(new_n475), .A2(new_n489), .ZN(G160));
  NAND4_X1  g065(.A1(new_n483), .A2(new_n480), .A3(G2105), .A4(new_n472), .ZN(new_n491));
  XNOR2_X1  g066(.A(new_n491), .B(KEYINPUT71), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n493), .A2(G124), .ZN(new_n494));
  OR2_X1    g069(.A1(G100), .A2(G2105), .ZN(new_n495));
  INV_X1    g070(.A(G2105), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n495), .B(G2104), .C1(G112), .C2(new_n496), .ZN(new_n497));
  XNOR2_X1  g072(.A(new_n497), .B(KEYINPUT72), .ZN(new_n498));
  AND3_X1   g073(.A1(new_n483), .A2(new_n480), .A3(new_n472), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n496), .ZN(new_n500));
  INV_X1    g075(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n498), .B1(G136), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n494), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(new_n503), .ZN(G162));
  NAND4_X1  g079(.A1(new_n499), .A2(KEYINPUT73), .A3(G126), .A4(G2105), .ZN(new_n505));
  INV_X1    g080(.A(G114), .ZN(new_n506));
  AND2_X1   g081(.A1(new_n506), .A2(KEYINPUT74), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(KEYINPUT74), .ZN(new_n508));
  OAI21_X1  g083(.A(G2105), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  OAI21_X1  g084(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(new_n511));
  INV_X1    g086(.A(G138), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n512), .A2(G2105), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(new_n470), .A3(new_n472), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT4), .ZN(new_n515));
  AOI22_X1  g090(.A1(new_n509), .A2(new_n511), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  INV_X1    g092(.A(G126), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n517), .B1(new_n491), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n483), .A4(new_n513), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n505), .A2(new_n516), .A3(new_n519), .A4(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(new_n521), .ZN(G164));
  XNOR2_X1  g097(.A(KEYINPUT5), .B(G543), .ZN(new_n523));
  XNOR2_X1  g098(.A(KEYINPUT75), .B(G651), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(KEYINPUT6), .A2(G651), .ZN(new_n527));
  OAI211_X1 g102(.A(G88), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(G50), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(KEYINPUT76), .ZN(new_n531));
  INV_X1    g106(.A(KEYINPUT76), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(G75), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n523), .ZN(new_n535));
  INV_X1    g110(.A(G62), .ZN(new_n536));
  OAI21_X1  g111(.A(new_n534), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(new_n524), .ZN(new_n538));
  AOI22_X1  g113(.A1(new_n531), .A2(new_n533), .B1(new_n537), .B2(new_n538), .ZN(G166));
  NAND3_X1  g114(.A1(new_n523), .A2(G63), .A3(G651), .ZN(new_n540));
  XOR2_X1   g115(.A(new_n540), .B(KEYINPUT77), .Z(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  XOR2_X1   g117(.A(new_n542), .B(KEYINPUT7), .Z(new_n543));
  NOR2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n526), .A2(new_n527), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n535), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G89), .ZN(new_n547));
  INV_X1    g122(.A(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n545), .A2(new_n548), .ZN(new_n549));
  XOR2_X1   g124(.A(KEYINPUT78), .B(G51), .Z(new_n550));
  NAND2_X1  g125(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n544), .A2(new_n547), .A3(new_n551), .ZN(G286));
  INV_X1    g127(.A(G286), .ZN(G168));
  AOI22_X1  g128(.A1(G52), .A2(new_n549), .B1(new_n546), .B2(G90), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n523), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n555));
  OR2_X1    g130(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n555), .A2(KEYINPUT79), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n556), .A2(new_n538), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n554), .A2(new_n558), .ZN(G301));
  INV_X1    g134(.A(G301), .ZN(G171));
  NAND2_X1  g135(.A1(new_n546), .A2(G81), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n549), .A2(G43), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n523), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n563));
  OR2_X1    g138(.A1(new_n563), .A2(new_n524), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n561), .A2(new_n562), .A3(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT80), .ZN(G176));
  NAND2_X1  g144(.A1(G1), .A2(G3), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT8), .ZN(new_n571));
  NAND4_X1  g146(.A1(G319), .A2(G483), .A3(G661), .A4(new_n571), .ZN(G188));
  OAI211_X1 g147(.A(G53), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n573));
  XNOR2_X1  g148(.A(new_n573), .B(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n535), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n546), .A2(G91), .B1(G651), .B2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  INV_X1    g154(.A(KEYINPUT81), .ZN(new_n580));
  XNOR2_X1  g155(.A(new_n579), .B(new_n580), .ZN(G299));
  NAND2_X1  g156(.A1(new_n537), .A2(new_n538), .ZN(new_n582));
  INV_X1    g157(.A(new_n533), .ZN(new_n583));
  AOI21_X1  g158(.A(new_n532), .B1(new_n528), .B2(new_n529), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n582), .B1(new_n583), .B2(new_n584), .ZN(G303));
  NAND2_X1  g160(.A1(new_n549), .A2(G49), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n546), .A2(G87), .ZN(new_n587));
  OAI21_X1  g162(.A(G651), .B1(new_n523), .B2(G74), .ZN(new_n588));
  AND3_X1   g163(.A1(new_n586), .A2(new_n587), .A3(new_n588), .ZN(new_n589));
  INV_X1    g164(.A(new_n589), .ZN(G288));
  AND2_X1   g165(.A1(new_n523), .A2(G61), .ZN(new_n591));
  NAND2_X1  g166(.A1(G73), .A2(G543), .ZN(new_n592));
  XNOR2_X1  g167(.A(new_n592), .B(KEYINPUT82), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n538), .B1(new_n591), .B2(new_n593), .ZN(new_n594));
  OAI211_X1 g169(.A(G48), .B(G543), .C1(new_n526), .C2(new_n527), .ZN(new_n595));
  OAI211_X1 g170(.A(G86), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G305));
  NAND2_X1  g172(.A1(new_n546), .A2(G85), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n549), .A2(G47), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n523), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  OR2_X1    g175(.A1(new_n600), .A2(new_n524), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n598), .A2(new_n599), .A3(new_n601), .ZN(G290));
  INV_X1    g177(.A(G868), .ZN(new_n603));
  NOR2_X1   g178(.A1(G301), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g179(.A1(G79), .A2(G543), .ZN(new_n605));
  INV_X1    g180(.A(G66), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n605), .B1(new_n535), .B2(new_n606), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT83), .ZN(new_n608));
  OR2_X1    g183(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(G651), .ZN(new_n610));
  AOI21_X1  g185(.A(new_n610), .B1(new_n607), .B2(new_n608), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n609), .A2(new_n611), .B1(new_n549), .B2(G54), .ZN(new_n612));
  OAI211_X1 g187(.A(G92), .B(new_n523), .C1(new_n526), .C2(new_n527), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n613), .B(new_n614), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT84), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n616), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g193(.A(new_n604), .B1(new_n618), .B2(new_n603), .ZN(G284));
  AOI21_X1  g194(.A(new_n604), .B1(new_n618), .B2(new_n603), .ZN(G321));
  NAND2_X1  g195(.A1(G286), .A2(G868), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n579), .B(KEYINPUT81), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n621), .B1(new_n622), .B2(G868), .ZN(G297));
  XNOR2_X1  g198(.A(G297), .B(KEYINPUT85), .ZN(G280));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n618), .B1(new_n625), .B2(G860), .ZN(G148));
  NAND2_X1  g201(.A1(new_n565), .A2(new_n603), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n618), .A2(new_n625), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n627), .B1(new_n629), .B2(new_n603), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n467), .A2(new_n476), .ZN(new_n632));
  XNOR2_X1  g207(.A(KEYINPUT86), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  INV_X1    g209(.A(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(KEYINPUT13), .ZN(new_n636));
  INV_X1    g211(.A(KEYINPUT87), .ZN(new_n637));
  INV_X1    g212(.A(G2100), .ZN(new_n638));
  OAI22_X1  g213(.A1(new_n635), .A2(new_n636), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  AOI21_X1  g214(.A(new_n639), .B1(new_n636), .B2(new_n635), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n637), .A2(new_n638), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n501), .A2(G135), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n496), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  INV_X1    g220(.A(G123), .ZN(new_n646));
  OAI221_X1 g221(.A(new_n643), .B1(new_n644), .B2(new_n645), .C1(new_n492), .C2(new_n646), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n647), .A2(G2096), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n647), .A2(G2096), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n642), .A2(new_n648), .A3(new_n649), .ZN(G156));
  XNOR2_X1  g225(.A(KEYINPUT15), .B(G2435), .ZN(new_n651));
  XNOR2_X1  g226(.A(KEYINPUT88), .B(G2438), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n651), .B(new_n652), .ZN(new_n653));
  XOR2_X1   g228(.A(G2427), .B(G2430), .Z(new_n654));
  OR2_X1    g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n653), .A2(new_n654), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n655), .A2(KEYINPUT14), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2451), .B(G2454), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT16), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n657), .B(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2443), .B(G2446), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XNOR2_X1  g237(.A(G1341), .B(G1348), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(new_n664), .B(KEYINPUT89), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n662), .A2(new_n663), .ZN(new_n666));
  AND3_X1   g241(.A1(new_n665), .A2(G14), .A3(new_n666), .ZN(G401));
  XOR2_X1   g242(.A(G2084), .B(G2090), .Z(new_n668));
  XNOR2_X1  g243(.A(G2067), .B(G2678), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT90), .Z(new_n670));
  NOR2_X1   g245(.A1(G2072), .A2(G2078), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n443), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g247(.A(new_n668), .B1(new_n670), .B2(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(KEYINPUT17), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n673), .B1(new_n670), .B2(new_n674), .ZN(new_n675));
  OAI211_X1 g250(.A(new_n668), .B(new_n669), .C1(new_n443), .C2(new_n671), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT18), .Z(new_n677));
  NAND3_X1  g252(.A1(new_n670), .A2(new_n674), .A3(new_n668), .ZN(new_n678));
  NAND3_X1  g253(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(G2096), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT91), .B(G2100), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(G227));
  XOR2_X1   g257(.A(G1971), .B(G1976), .Z(new_n683));
  XNOR2_X1  g258(.A(new_n683), .B(KEYINPUT19), .ZN(new_n684));
  XOR2_X1   g259(.A(G1956), .B(G2474), .Z(new_n685));
  XOR2_X1   g260(.A(G1961), .B(G1966), .Z(new_n686));
  AND2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT20), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n685), .A2(new_n686), .ZN(new_n690));
  NOR3_X1   g265(.A1(new_n684), .A2(new_n687), .A3(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n691), .B1(new_n684), .B2(new_n690), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g268(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G23), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(new_n589), .B2(new_n700), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT33), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n703), .B(G1976), .ZN(new_n704));
  MUX2_X1   g279(.A(G6), .B(G305), .S(G16), .Z(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT94), .ZN(new_n706));
  XOR2_X1   g281(.A(KEYINPUT32), .B(G1981), .Z(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NOR2_X1   g283(.A1(G16), .A2(G22), .ZN(new_n709));
  AOI21_X1  g284(.A(new_n709), .B1(G166), .B2(G16), .ZN(new_n710));
  XOR2_X1   g285(.A(new_n710), .B(G1971), .Z(new_n711));
  NAND3_X1  g286(.A1(new_n704), .A2(new_n708), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT34), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n501), .A2(G131), .ZN(new_n715));
  NOR2_X1   g290(.A1(new_n496), .A2(G107), .ZN(new_n716));
  OAI21_X1  g291(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n717));
  INV_X1    g292(.A(G119), .ZN(new_n718));
  OAI221_X1 g293(.A(new_n715), .B1(new_n716), .B2(new_n717), .C1(new_n492), .C2(new_n718), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n719), .B(KEYINPUT92), .ZN(new_n720));
  MUX2_X1   g295(.A(G25), .B(new_n720), .S(G29), .Z(new_n721));
  XNOR2_X1  g296(.A(KEYINPUT35), .B(G1991), .ZN(new_n722));
  XOR2_X1   g297(.A(new_n721), .B(new_n722), .Z(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G24), .ZN(new_n724));
  XOR2_X1   g299(.A(G290), .B(KEYINPUT93), .Z(new_n725));
  AOI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(G16), .ZN(new_n726));
  INV_X1    g301(.A(G1986), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NAND4_X1  g303(.A1(new_n713), .A2(new_n714), .A3(new_n723), .A4(new_n728), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n700), .A2(G19), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT96), .Z(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n566), .B2(new_n700), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1341), .ZN(new_n736));
  INV_X1    g311(.A(G29), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n737), .A2(G26), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT28), .Z(new_n739));
  AND3_X1   g314(.A1(new_n499), .A2(G140), .A3(new_n496), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT97), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n493), .A2(G128), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n496), .A2(G116), .ZN(new_n743));
  OAI21_X1  g318(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n744));
  OAI211_X1 g319(.A(new_n741), .B(new_n742), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n739), .B1(new_n745), .B2(G29), .ZN(new_n746));
  INV_X1    g321(.A(G2067), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n746), .B(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n737), .A2(G35), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT102), .Z(new_n750));
  AOI21_X1  g325(.A(new_n750), .B1(new_n503), .B2(G29), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT29), .ZN(new_n752));
  INV_X1    g327(.A(new_n752), .ZN(new_n753));
  AOI211_X1 g328(.A(new_n736), .B(new_n748), .C1(G2090), .C2(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n700), .A2(G20), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT23), .Z(new_n756));
  AOI21_X1  g331(.A(new_n756), .B1(G299), .B2(G16), .ZN(new_n757));
  INV_X1    g332(.A(G1956), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n753), .A2(G2090), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n759), .B1(KEYINPUT103), .B2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(G4), .A2(G16), .ZN(new_n762));
  AOI21_X1  g337(.A(new_n762), .B1(new_n618), .B2(G16), .ZN(new_n763));
  INV_X1    g338(.A(G1348), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n763), .B(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n760), .A2(KEYINPUT103), .ZN(new_n766));
  AND4_X1   g341(.A1(new_n754), .A2(new_n761), .A3(new_n765), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n700), .A2(G5), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G171), .B2(new_n700), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n769), .A2(G1961), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(KEYINPUT100), .Z(new_n771));
  AND2_X1   g346(.A1(new_n700), .A2(G21), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G286), .B2(G16), .ZN(new_n773));
  INV_X1    g348(.A(G1966), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT99), .Z(new_n776));
  XNOR2_X1  g351(.A(KEYINPUT30), .B(G28), .ZN(new_n777));
  OR2_X1    g352(.A1(KEYINPUT31), .A2(G11), .ZN(new_n778));
  NAND2_X1  g353(.A1(KEYINPUT31), .A2(G11), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n777), .A2(new_n737), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(new_n647), .B2(new_n737), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n781), .B(KEYINPUT98), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n771), .A2(new_n776), .A3(new_n782), .ZN(new_n783));
  NOR2_X1   g358(.A1(G160), .A2(new_n737), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n737), .B1(KEYINPUT24), .B2(G34), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(KEYINPUT24), .B2(G34), .ZN(new_n786));
  NOR2_X1   g361(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G2084), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n737), .A2(G32), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n501), .A2(G141), .ZN(new_n790));
  NAND3_X1  g365(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n791));
  INV_X1    g366(.A(KEYINPUT26), .ZN(new_n792));
  OR2_X1    g367(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  AOI22_X1  g369(.A1(new_n793), .A2(new_n794), .B1(G105), .B2(new_n476), .ZN(new_n795));
  INV_X1    g370(.A(G129), .ZN(new_n796));
  OAI211_X1 g371(.A(new_n790), .B(new_n795), .C1(new_n492), .C2(new_n796), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n789), .B1(new_n798), .B2(new_n737), .ZN(new_n799));
  XNOR2_X1  g374(.A(KEYINPUT27), .B(G1996), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n737), .A2(G27), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G164), .B2(new_n737), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G2078), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n737), .A2(G33), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n501), .A2(G139), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n496), .A2(G103), .A3(G2104), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(KEYINPUT25), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n467), .A2(G127), .ZN(new_n810));
  INV_X1    g385(.A(G115), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n810), .B1(new_n811), .B2(new_n469), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n809), .B1(new_n812), .B2(G2105), .ZN(new_n813));
  AND2_X1   g388(.A1(new_n807), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g389(.A(new_n806), .B1(new_n814), .B2(new_n737), .ZN(new_n815));
  XOR2_X1   g390(.A(new_n815), .B(G2072), .Z(new_n816));
  OAI221_X1 g391(.A(new_n816), .B1(G1961), .B2(new_n769), .C1(new_n774), .C2(new_n773), .ZN(new_n817));
  NOR4_X1   g392(.A1(new_n783), .A2(new_n802), .A3(new_n805), .A4(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n818), .B(KEYINPUT101), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n731), .A2(new_n732), .A3(new_n767), .A4(new_n819), .ZN(G150));
  INV_X1    g395(.A(G150), .ZN(G311));
  XNOR2_X1  g396(.A(KEYINPUT105), .B(G93), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n546), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n549), .A2(G55), .ZN(new_n824));
  AOI22_X1  g399(.A1(new_n523), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n825));
  OAI211_X1 g400(.A(new_n823), .B(new_n824), .C1(new_n524), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g401(.A1(new_n826), .A2(G860), .ZN(new_n827));
  XOR2_X1   g402(.A(KEYINPUT108), .B(KEYINPUT37), .Z(new_n828));
  XNOR2_X1  g403(.A(new_n827), .B(new_n828), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n618), .A2(G559), .ZN(new_n830));
  XNOR2_X1  g405(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n830), .B(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n826), .A2(KEYINPUT106), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n826), .A2(KEYINPUT106), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n833), .A2(new_n566), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n566), .B1(new_n833), .B2(new_n834), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n832), .B(new_n837), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n838), .A2(KEYINPUT39), .ZN(new_n839));
  XOR2_X1   g414(.A(new_n839), .B(KEYINPUT107), .Z(new_n840));
  INV_X1    g415(.A(G860), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n841), .B1(new_n838), .B2(KEYINPUT39), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n829), .B1(new_n840), .B2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n720), .B(new_n635), .ZN(new_n844));
  OR2_X1    g419(.A1(G106), .A2(G2105), .ZN(new_n845));
  OAI211_X1 g420(.A(new_n845), .B(G2104), .C1(G118), .C2(new_n496), .ZN(new_n846));
  INV_X1    g421(.A(G142), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n846), .B1(new_n500), .B2(new_n847), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(new_n493), .B2(G130), .ZN(new_n849));
  OR2_X1    g424(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n814), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n745), .B(new_n521), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(new_n798), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n798), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n851), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n852), .A2(new_n798), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n852), .A2(new_n798), .ZN(new_n857));
  NAND3_X1  g432(.A1(new_n856), .A2(new_n814), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g433(.A1(new_n844), .A2(new_n849), .ZN(new_n859));
  NAND4_X1  g434(.A1(new_n850), .A2(new_n855), .A3(new_n858), .A4(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT109), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n850), .A2(new_n859), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n858), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n861), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n503), .B(G160), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n869), .B(new_n647), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n860), .A2(new_n872), .ZN(new_n873));
  AOI21_X1  g448(.A(G37), .B1(new_n873), .B2(new_n865), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n871), .A2(KEYINPUT40), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(KEYINPUT40), .B1(new_n871), .B2(new_n874), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(G395));
  NAND2_X1  g452(.A1(new_n629), .A2(KEYINPUT110), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n835), .A2(new_n836), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT110), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n628), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(new_n881), .ZN(new_n883));
  NOR2_X1   g458(.A1(new_n628), .A2(new_n880), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n837), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT111), .ZN(new_n886));
  NAND2_X1  g461(.A1(G299), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n622), .A2(KEYINPUT111), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n887), .A2(new_n888), .A3(new_n616), .ZN(new_n889));
  NAND4_X1  g464(.A1(new_n622), .A2(KEYINPUT111), .A3(new_n615), .A4(new_n612), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT41), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n889), .A2(KEYINPUT41), .A3(new_n890), .ZN(new_n894));
  AOI22_X1  g469(.A1(new_n882), .A2(new_n885), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n897));
  NAND3_X1  g472(.A1(new_n885), .A2(new_n882), .A3(new_n891), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n896), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  INV_X1    g474(.A(new_n898), .ZN(new_n900));
  OAI21_X1  g475(.A(KEYINPUT42), .B1(new_n895), .B2(new_n900), .ZN(new_n901));
  XOR2_X1   g476(.A(new_n589), .B(G305), .Z(new_n902));
  XNOR2_X1  g477(.A(G303), .B(G290), .ZN(new_n903));
  XNOR2_X1  g478(.A(new_n902), .B(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(new_n904), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n899), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n899), .B2(new_n901), .ZN(new_n907));
  OAI21_X1  g482(.A(G868), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n826), .A2(new_n603), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n908), .A2(new_n909), .ZN(G295));
  NAND2_X1  g485(.A1(new_n908), .A2(new_n909), .ZN(G331));
  INV_X1    g486(.A(KEYINPUT44), .ZN(new_n912));
  NOR2_X1   g487(.A1(G286), .A2(KEYINPUT112), .ZN(new_n913));
  NAND2_X1  g488(.A1(G286), .A2(KEYINPUT112), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT113), .ZN(new_n915));
  AND3_X1   g490(.A1(new_n914), .A2(new_n915), .A3(G301), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n915), .B1(new_n914), .B2(G301), .ZN(new_n917));
  OAI21_X1  g492(.A(new_n913), .B1(new_n916), .B2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n914), .A2(G301), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT113), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n914), .A2(new_n915), .A3(G301), .ZN(new_n921));
  INV_X1    g496(.A(new_n913), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(new_n837), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n879), .A2(new_n918), .A3(new_n923), .ZN(new_n926));
  NAND4_X1  g501(.A1(new_n925), .A2(new_n890), .A3(new_n889), .A4(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n893), .A2(new_n894), .ZN(new_n928));
  AND3_X1   g503(.A1(new_n918), .A2(new_n879), .A3(new_n923), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n879), .B1(new_n918), .B2(new_n923), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n927), .B1(new_n928), .B2(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(G37), .B1(new_n932), .B2(new_n905), .ZN(new_n933));
  INV_X1    g508(.A(KEYINPUT43), .ZN(new_n934));
  OAI211_X1 g509(.A(new_n927), .B(new_n904), .C1(new_n928), .C2(new_n931), .ZN(new_n935));
  AND3_X1   g510(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n933), .B2(new_n935), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n912), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n932), .A2(new_n905), .ZN(new_n939));
  INV_X1    g514(.A(G37), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n939), .A2(new_n940), .A3(new_n935), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n941), .A2(KEYINPUT43), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n933), .A2(new_n934), .A3(new_n935), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n942), .A2(KEYINPUT44), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n938), .A2(new_n944), .ZN(G397));
  INV_X1    g520(.A(G1384), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n521), .A2(new_n946), .ZN(new_n947));
  OR2_X1    g522(.A1(new_n947), .A2(KEYINPUT114), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n470), .A2(new_n472), .A3(G125), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(KEYINPUT67), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n470), .A2(new_n472), .A3(new_n466), .A4(G125), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n464), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g527(.A(G40), .B1(new_n952), .B2(new_n496), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n487), .A2(KEYINPUT70), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n477), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g531(.A(KEYINPUT115), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT115), .ZN(new_n958));
  NAND4_X1  g533(.A1(new_n475), .A2(new_n489), .A3(new_n958), .A4(G40), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g535(.A(KEYINPUT45), .B1(new_n947), .B2(KEYINPUT114), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n948), .A2(new_n960), .A3(new_n961), .ZN(new_n962));
  XNOR2_X1  g537(.A(new_n745), .B(new_n747), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n962), .B1(new_n963), .B2(new_n798), .ZN(new_n964));
  OR3_X1    g539(.A1(new_n962), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n965));
  OAI21_X1  g540(.A(KEYINPUT46), .B1(new_n962), .B2(G1996), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n964), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  XOR2_X1   g542(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n968));
  XNOR2_X1  g543(.A(new_n967), .B(new_n968), .ZN(new_n969));
  INV_X1    g544(.A(new_n962), .ZN(new_n970));
  INV_X1    g545(.A(G1996), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n798), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n972), .B(KEYINPUT117), .Z(new_n973));
  OAI21_X1  g548(.A(new_n963), .B1(new_n971), .B2(new_n798), .ZN(new_n974));
  AOI21_X1  g549(.A(new_n973), .B1(new_n970), .B2(new_n974), .ZN(new_n975));
  AND2_X1   g550(.A1(new_n720), .A2(new_n722), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n720), .A2(new_n722), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(G290), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n727), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT116), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n982), .A2(new_n962), .ZN(new_n983));
  XNOR2_X1  g558(.A(new_n983), .B(KEYINPUT48), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n969), .B1(new_n979), .B2(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n975), .A2(new_n977), .ZN(new_n986));
  OR2_X1    g561(.A1(new_n745), .A2(G2067), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n962), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT126), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n982), .B1(new_n727), .B2(new_n980), .ZN(new_n991));
  AND2_X1   g566(.A1(new_n991), .A2(new_n970), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n979), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT45), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n947), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n521), .A2(KEYINPUT45), .A3(new_n946), .ZN(new_n996));
  AND4_X1   g571(.A1(new_n971), .A2(new_n960), .A3(new_n995), .A4(new_n996), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n947), .B1(new_n957), .B2(new_n959), .ZN(new_n998));
  XNOR2_X1  g573(.A(KEYINPUT58), .B(G1341), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OAI21_X1  g575(.A(new_n566), .B1(new_n997), .B2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT59), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT59), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n1003), .B(new_n566), .C1(new_n997), .C2(new_n1000), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1002), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n947), .A2(KEYINPUT50), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT50), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n521), .A2(new_n1007), .A3(new_n946), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n953), .A2(new_n956), .A3(KEYINPUT115), .ZN(new_n1009));
  INV_X1    g584(.A(G40), .ZN(new_n1010));
  AOI21_X1  g585(.A(new_n1010), .B1(new_n474), .B2(G2105), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n958), .B1(new_n1011), .B2(new_n489), .ZN(new_n1012));
  OAI211_X1 g587(.A(new_n1006), .B(new_n1008), .C1(new_n1009), .C2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n764), .ZN(new_n1014));
  NAND2_X1  g589(.A1(new_n998), .A2(new_n747), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1014), .A2(KEYINPUT60), .A3(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n616), .B(KEYINPUT84), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT60), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND4_X1  g596(.A1(new_n618), .A2(KEYINPUT60), .A3(new_n1014), .A4(new_n1015), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1018), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1013), .A2(new_n758), .ZN(new_n1024));
  XNOR2_X1  g599(.A(KEYINPUT56), .B(G2072), .ZN(new_n1025));
  NAND4_X1  g600(.A1(new_n960), .A2(new_n995), .A3(new_n996), .A4(new_n1025), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n1024), .A2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT57), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n579), .A2(new_n1028), .ZN(new_n1029));
  NAND3_X1  g604(.A1(new_n574), .A2(KEYINPUT57), .A3(new_n578), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1027), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1024), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n1033), .A2(KEYINPUT61), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT61), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n1024), .A2(new_n1031), .A3(new_n1026), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1031), .B1(new_n1024), .B2(new_n1026), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1036), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  NAND4_X1  g614(.A1(new_n1005), .A2(new_n1023), .A3(new_n1035), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1017), .B1(new_n1015), .B2(new_n1014), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n1034), .B1(new_n1041), .B2(new_n1038), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n1040), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(G1976), .ZN(new_n1044));
  NOR2_X1   g619(.A1(G288), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(new_n947), .ZN(new_n1046));
  OAI21_X1  g621(.A(new_n1046), .B1(new_n1009), .B2(new_n1012), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT119), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1047), .A2(new_n1048), .A3(G8), .ZN(new_n1049));
  INV_X1    g624(.A(G8), .ZN(new_n1050));
  OAI21_X1  g625(.A(KEYINPUT119), .B1(new_n998), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1045), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1052));
  XOR2_X1   g627(.A(KEYINPUT120), .B(G1976), .Z(new_n1053));
  AOI21_X1  g628(.A(KEYINPUT52), .B1(G288), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1055));
  NAND2_X1  g630(.A1(G305), .A2(G1981), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT49), .ZN(new_n1057));
  INV_X1    g632(.A(G1981), .ZN(new_n1058));
  NAND4_X1  g633(.A1(new_n595), .A2(new_n594), .A3(new_n596), .A4(new_n1058), .ZN(new_n1059));
  AND3_X1   g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1057), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1061));
  NOR2_X1   g636(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(new_n1062), .ZN(new_n1063));
  AOI22_X1  g638(.A1(new_n1052), .A2(new_n1054), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1048), .B1(new_n1047), .B2(G8), .ZN(new_n1065));
  NOR3_X1   g640(.A1(new_n998), .A2(KEYINPUT119), .A3(new_n1050), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT52), .B1(new_n1067), .B2(new_n1045), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT55), .ZN(new_n1069));
  OAI21_X1  g644(.A(new_n1069), .B1(G166), .B2(new_n1050), .ZN(new_n1070));
  NAND3_X1  g645(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1071));
  AND2_X1   g646(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n960), .A2(new_n1008), .A3(new_n1006), .ZN(new_n1073));
  INV_X1    g648(.A(G2090), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n960), .A2(new_n995), .A3(new_n996), .ZN(new_n1075));
  XOR2_X1   g650(.A(KEYINPUT118), .B(G1971), .Z(new_n1076));
  AOI22_X1  g651(.A1(new_n1073), .A2(new_n1074), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1077));
  OAI21_X1  g652(.A(new_n1072), .B1(new_n1077), .B2(new_n1050), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1079));
  AOI22_X1  g654(.A1(new_n957), .A2(new_n959), .B1(new_n947), .B2(KEYINPUT50), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(new_n1074), .A3(new_n1008), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1082), .A2(G8), .A3(new_n1083), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1064), .A2(new_n1068), .A3(new_n1078), .A4(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(G2084), .ZN(new_n1087));
  AOI22_X1  g662(.A1(new_n1073), .A2(new_n1087), .B1(new_n1075), .B2(new_n774), .ZN(new_n1088));
  NAND2_X1  g663(.A1(G286), .A2(G8), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT51), .ZN(new_n1091));
  AOI21_X1  g666(.A(new_n1091), .B1(new_n1089), .B2(KEYINPUT123), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1092), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1093), .B(new_n1089), .C1(new_n1088), .C2(new_n1050), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1075), .A2(new_n774), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1080), .A2(new_n1087), .A3(new_n1008), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g672(.A(G8), .B(new_n1092), .C1(new_n1097), .C2(G286), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n1090), .B1(new_n1094), .B2(new_n1098), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT53), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1100), .B1(new_n1075), .B2(G2078), .ZN(new_n1101));
  AOI22_X1  g676(.A1(KEYINPUT45), .A2(new_n1046), .B1(new_n957), .B2(new_n959), .ZN(new_n1102));
  NOR2_X1   g677(.A1(new_n1100), .A2(G2078), .ZN(new_n1103));
  NAND3_X1  g678(.A1(new_n1102), .A2(new_n995), .A3(new_n1103), .ZN(new_n1104));
  OAI211_X1 g679(.A(new_n1101), .B(new_n1104), .C1(G1961), .C2(new_n1073), .ZN(new_n1105));
  NAND2_X1  g680(.A1(G171), .A2(KEYINPUT54), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT54), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G301), .A2(new_n1107), .ZN(new_n1108));
  AND2_X1   g683(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1105), .A2(new_n1109), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n948), .A2(new_n961), .ZN(new_n1111));
  AOI21_X1  g686(.A(new_n496), .B1(new_n474), .B2(KEYINPUT124), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1112), .B1(KEYINPUT124), .B2(new_n474), .ZN(new_n1113));
  AND3_X1   g688(.A1(new_n489), .A2(G40), .A3(new_n1103), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n996), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1106), .A2(new_n1108), .B1(new_n1111), .B2(new_n1115), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n1116), .B(new_n1101), .C1(G1961), .C2(new_n1073), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1110), .A2(new_n1117), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1099), .A2(new_n1118), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1043), .A2(new_n1086), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n589), .A2(new_n1044), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1121), .B1(new_n1055), .B2(new_n1063), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1059), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT121), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT121), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n1062), .B1(new_n1049), .B2(new_n1051), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1125), .B(new_n1059), .C1(new_n1126), .C2(new_n1121), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1124), .A2(new_n1055), .A3(new_n1127), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1077), .A2(new_n1050), .A3(new_n1072), .ZN(new_n1129));
  NAND3_X1  g704(.A1(new_n1064), .A2(new_n1129), .A3(new_n1068), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1128), .A2(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT122), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT63), .ZN(new_n1134));
  AOI21_X1  g709(.A(G1966), .B1(new_n1102), .B2(new_n995), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n1013), .A2(G2084), .ZN(new_n1136));
  OAI21_X1  g711(.A(G8), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(new_n1137), .A2(G286), .ZN(new_n1138));
  INV_X1    g713(.A(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1134), .B1(new_n1085), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1045), .ZN(new_n1141));
  OAI211_X1 g716(.A(new_n1141), .B(new_n1054), .C1(new_n1065), .C2(new_n1066), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1055), .A2(new_n1063), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT52), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n1052), .A2(new_n1145), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1144), .A2(new_n1146), .ZN(new_n1147));
  AOI21_X1  g722(.A(new_n1083), .B1(new_n1082), .B2(G8), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1129), .A2(new_n1148), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1147), .A2(new_n1149), .A3(KEYINPUT63), .A4(new_n1138), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1140), .A2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1128), .A2(KEYINPUT122), .A3(new_n1130), .ZN(new_n1152));
  NAND4_X1  g727(.A1(new_n1120), .A2(new_n1133), .A3(new_n1151), .A4(new_n1152), .ZN(new_n1153));
  AOI211_X1 g728(.A(KEYINPUT62), .B(new_n1090), .C1(new_n1094), .C2(new_n1098), .ZN(new_n1154));
  AND2_X1   g729(.A1(new_n1105), .A2(G171), .ZN(new_n1155));
  NAND3_X1  g730(.A1(new_n1147), .A2(new_n1149), .A3(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n1090), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1093), .B1(new_n1137), .B2(new_n1089), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1050), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1089), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1092), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n1157), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1162), .A2(KEYINPUT125), .A3(KEYINPUT62), .ZN(new_n1163));
  INV_X1    g738(.A(KEYINPUT125), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1164), .B1(new_n1099), .B2(new_n1165), .ZN(new_n1166));
  AOI211_X1 g741(.A(new_n1154), .B(new_n1156), .C1(new_n1163), .C2(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n990), .B(new_n993), .C1(new_n1153), .C2(new_n1167), .ZN(new_n1168));
  INV_X1    g743(.A(new_n1168), .ZN(new_n1169));
  NOR3_X1   g744(.A1(new_n1085), .A2(new_n1099), .A3(new_n1118), .ZN(new_n1170));
  OAI21_X1  g745(.A(new_n1059), .B1(new_n1126), .B2(new_n1121), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1067), .B1(new_n1171), .B2(KEYINPUT121), .ZN(new_n1172));
  AOI22_X1  g747(.A1(new_n1172), .A2(new_n1127), .B1(new_n1147), .B2(new_n1129), .ZN(new_n1173));
  AOI22_X1  g748(.A1(new_n1043), .A2(new_n1170), .B1(new_n1173), .B2(KEYINPUT122), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1163), .A2(new_n1166), .ZN(new_n1175));
  NOR2_X1   g750(.A1(new_n1156), .A2(new_n1154), .ZN(new_n1176));
  NAND2_X1  g751(.A1(new_n1175), .A2(new_n1176), .ZN(new_n1177));
  AOI22_X1  g752(.A1(new_n1132), .A2(new_n1131), .B1(new_n1140), .B2(new_n1150), .ZN(new_n1178));
  NAND3_X1  g753(.A1(new_n1174), .A2(new_n1177), .A3(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n990), .B1(new_n1179), .B2(new_n993), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n989), .B1(new_n1169), .B2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  NOR4_X1   g756(.A1(G401), .A2(G229), .A3(new_n461), .A4(G227), .ZN(new_n1183));
  AOI21_X1  g757(.A(new_n872), .B1(new_n866), .B2(new_n867), .ZN(new_n1184));
  NAND2_X1  g758(.A1(new_n873), .A2(new_n865), .ZN(new_n1185));
  NAND2_X1  g759(.A1(new_n1185), .A2(new_n940), .ZN(new_n1186));
  OAI21_X1  g760(.A(new_n1183), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  AOI21_X1  g761(.A(new_n1187), .B1(new_n942), .B2(new_n943), .ZN(G308));
  OAI221_X1 g762(.A(new_n1183), .B1(new_n1184), .B2(new_n1186), .C1(new_n936), .C2(new_n937), .ZN(G225));
endmodule


