//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 1 1 1 0 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1 1 1 1 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:50 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n948, new_n949, new_n950, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035;
  OAI21_X1  g000(.A(G210), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  XOR2_X1   g002(.A(G110), .B(G122), .Z(new_n189));
  XNOR2_X1  g003(.A(G116), .B(G119), .ZN(new_n190));
  XNOR2_X1  g004(.A(KEYINPUT2), .B(G113), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT3), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n193), .B1(new_n194), .B2(G107), .ZN(new_n195));
  INV_X1    g009(.A(G107), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n196), .A2(KEYINPUT3), .A3(G104), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n195), .A2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(KEYINPUT79), .A2(G101), .ZN(new_n199));
  NOR2_X1   g013(.A1(KEYINPUT79), .A2(G101), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n199), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(KEYINPUT78), .B1(new_n196), .B2(G104), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT78), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n194), .A3(G107), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n201), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  AND2_X1   g021(.A1(new_n202), .A2(new_n204), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n207), .B1(new_n208), .B2(new_n198), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT4), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n198), .A2(new_n202), .A3(new_n204), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G101), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT4), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n192), .B1(new_n210), .B2(new_n214), .ZN(new_n215));
  XOR2_X1   g029(.A(G116), .B(G119), .Z(new_n216));
  OR2_X1    g030(.A1(new_n216), .A2(new_n191), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n194), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n196), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n205), .A2(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT5), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT82), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT82), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n224), .A2(KEYINPUT5), .ZN(new_n225));
  INV_X1    g039(.A(G119), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n223), .A2(new_n225), .A3(G116), .A4(new_n226), .ZN(new_n227));
  XNOR2_X1  g041(.A(KEYINPUT82), .B(KEYINPUT5), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n227), .B(G113), .C1(new_n216), .C2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(KEYINPUT83), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n228), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n232), .A2(new_n190), .ZN(new_n233));
  NAND4_X1  g047(.A1(new_n233), .A2(KEYINPUT83), .A3(G113), .A4(new_n227), .ZN(new_n234));
  AND4_X1   g048(.A1(new_n217), .A2(new_n221), .A3(new_n231), .A4(new_n234), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n189), .B1(new_n215), .B2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n192), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n213), .B1(new_n212), .B2(new_n205), .ZN(new_n238));
  NOR2_X1   g052(.A1(new_n209), .A2(KEYINPUT4), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n237), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND4_X1  g054(.A1(new_n221), .A2(new_n231), .A3(new_n234), .A4(new_n217), .ZN(new_n241));
  INV_X1    g055(.A(new_n189), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n240), .A2(new_n241), .A3(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n236), .A2(KEYINPUT6), .A3(new_n243), .ZN(new_n244));
  NOR2_X1   g058(.A1(KEYINPUT0), .A2(G128), .ZN(new_n245));
  NAND2_X1  g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(KEYINPUT65), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT65), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n248), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n245), .B1(new_n247), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(G143), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT66), .B1(new_n251), .B2(G146), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT66), .ZN(new_n253));
  INV_X1    g067(.A(G146), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n253), .A2(new_n254), .A3(G143), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT67), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n257), .B1(new_n254), .B2(G143), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n251), .A2(KEYINPUT67), .A3(G146), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n250), .B1(new_n256), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n254), .A2(G143), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n251), .A2(G146), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(new_n246), .ZN(new_n265));
  INV_X1    g079(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G125), .ZN(new_n268));
  INV_X1    g082(.A(G128), .ZN(new_n269));
  NOR2_X1   g083(.A1(new_n269), .A2(KEYINPUT1), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n270), .A2(new_n262), .A3(new_n263), .ZN(new_n271));
  INV_X1    g085(.A(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n253), .B1(G143), .B2(new_n254), .ZN(new_n273));
  NOR3_X1   g087(.A1(new_n251), .A2(KEYINPUT66), .A3(G146), .ZN(new_n274));
  OAI211_X1 g088(.A(new_n258), .B(new_n259), .C1(new_n273), .C2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n251), .A2(G146), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT1), .ZN(new_n277));
  OAI21_X1  g091(.A(G128), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(new_n272), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(G125), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n268), .A2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G224), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n283), .A2(G953), .ZN(new_n284));
  XNOR2_X1  g098(.A(new_n282), .B(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(KEYINPUT6), .ZN(new_n286));
  OAI211_X1 g100(.A(new_n286), .B(new_n189), .C1(new_n215), .C2(new_n235), .ZN(new_n287));
  AND3_X1   g101(.A1(new_n244), .A2(new_n285), .A3(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G902), .ZN(new_n289));
  INV_X1    g103(.A(new_n284), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(KEYINPUT7), .ZN(new_n291));
  AOI21_X1  g105(.A(new_n265), .B1(new_n275), .B2(new_n250), .ZN(new_n292));
  NOR2_X1   g106(.A1(new_n292), .A2(new_n280), .ZN(new_n293));
  AOI211_X1 g107(.A(G125), .B(new_n272), .C1(new_n275), .C2(new_n278), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n291), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(KEYINPUT86), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT86), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n282), .A2(new_n297), .A3(new_n291), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n268), .A2(KEYINPUT7), .A3(new_n290), .A4(new_n281), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n300));
  OAI211_X1 g114(.A(new_n227), .B(G113), .C1(new_n216), .C2(new_n222), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(new_n217), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT85), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n301), .A2(new_n217), .A3(KEYINPUT85), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n304), .A2(new_n221), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n205), .A2(new_n220), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n231), .A2(new_n234), .A3(new_n217), .A4(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT84), .B(KEYINPUT8), .ZN(new_n309));
  XNOR2_X1  g123(.A(new_n189), .B(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n306), .A2(new_n308), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n243), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n289), .B1(new_n300), .B2(new_n312), .ZN(new_n313));
  OAI21_X1  g127(.A(new_n188), .B1(new_n288), .B2(new_n313), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n296), .A2(new_n298), .A3(new_n299), .ZN(new_n315));
  AND2_X1   g129(.A1(new_n243), .A2(new_n311), .ZN(new_n316));
  AOI21_X1  g130(.A(G902), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n244), .A2(new_n285), .A3(new_n287), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n317), .A2(new_n318), .A3(new_n187), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n314), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(G234), .A2(G237), .ZN(new_n321));
  INV_X1    g135(.A(G953), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n321), .A2(G952), .A3(new_n322), .ZN(new_n323));
  XOR2_X1   g137(.A(new_n323), .B(KEYINPUT93), .Z(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(KEYINPUT21), .B(G898), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n321), .A2(G902), .A3(G953), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n325), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(G214), .B1(G237), .B2(G902), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n320), .A2(new_n330), .A3(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n279), .A2(new_n333), .A3(new_n307), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n333), .B1(new_n279), .B2(new_n307), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n272), .B1(new_n278), .B2(new_n264), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n336), .A2(new_n307), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT11), .ZN(new_n339));
  INV_X1    g153(.A(G134), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n339), .B1(new_n340), .B2(G137), .ZN(new_n341));
  INV_X1    g155(.A(G137), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n342), .A2(KEYINPUT11), .A3(G134), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n340), .A2(G137), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n341), .A2(new_n343), .A3(new_n344), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n345), .A2(G131), .ZN(new_n346));
  INV_X1    g160(.A(G131), .ZN(new_n347));
  NAND4_X1  g161(.A1(new_n341), .A2(new_n343), .A3(new_n347), .A4(new_n344), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT12), .B1(new_n338), .B2(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n335), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n278), .A2(new_n264), .ZN(new_n353));
  OAI211_X1 g167(.A(new_n205), .B(new_n220), .C1(new_n353), .C2(new_n272), .ZN(new_n354));
  NAND3_X1  g168(.A1(new_n279), .A2(new_n307), .A3(new_n333), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n352), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT12), .ZN(new_n357));
  NAND3_X1  g171(.A1(new_n356), .A2(new_n357), .A3(new_n349), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n359));
  NOR2_X1   g173(.A1(new_n279), .A2(new_n359), .ZN(new_n360));
  XNOR2_X1  g174(.A(KEYINPUT80), .B(KEYINPUT10), .ZN(new_n361));
  AOI22_X1  g175(.A1(new_n360), .A2(new_n221), .B1(new_n354), .B2(new_n361), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n292), .B1(new_n238), .B2(new_n239), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n350), .A3(new_n363), .ZN(new_n364));
  XNOR2_X1  g178(.A(G110), .B(G140), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n322), .A2(G227), .ZN(new_n366));
  XOR2_X1   g180(.A(new_n365), .B(new_n366), .Z(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND4_X1  g182(.A1(new_n351), .A2(new_n358), .A3(new_n364), .A4(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n364), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n350), .B1(new_n362), .B2(new_n363), .ZN(new_n371));
  OAI21_X1  g185(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(G469), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n373), .A2(new_n374), .A3(new_n289), .ZN(new_n375));
  NAND2_X1  g189(.A1(G469), .A2(G902), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n351), .A2(new_n364), .A3(new_n358), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(new_n367), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n362), .A2(new_n363), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(new_n349), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n380), .A2(new_n364), .A3(new_n368), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n378), .A2(G469), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n375), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  INV_X1    g197(.A(G221), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT9), .B(G234), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n386), .B2(new_n289), .ZN(new_n387));
  INV_X1    g201(.A(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT92), .ZN(new_n390));
  INV_X1    g204(.A(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n391), .A2(G116), .ZN(new_n392));
  INV_X1    g206(.A(G116), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(G122), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(KEYINPUT14), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT14), .ZN(new_n397));
  OAI21_X1  g211(.A(G107), .B1(new_n394), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n390), .B1(new_n396), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n398), .ZN(new_n400));
  XNOR2_X1  g214(.A(G116), .B(G122), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(new_n397), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n400), .A2(new_n402), .A3(KEYINPUT92), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n399), .A2(new_n403), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n395), .A2(G107), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n251), .A2(G128), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n269), .A2(G143), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n406), .A2(new_n407), .A3(new_n340), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n406), .A2(new_n407), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n409), .A2(G134), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n405), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n401), .A2(new_n196), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n408), .B1(new_n405), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(KEYINPUT13), .B1(new_n251), .B2(G128), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n415), .B1(new_n269), .B2(G143), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n251), .A2(KEYINPUT13), .A3(G128), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n340), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  OR2_X1    g232(.A1(new_n414), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n412), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT73), .B(G217), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n421), .A2(new_n385), .A3(G953), .ZN(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  XNOR2_X1  g237(.A(new_n420), .B(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(new_n289), .ZN(new_n425));
  INV_X1    g239(.A(G478), .ZN(new_n426));
  NOR2_X1   g240(.A1(new_n426), .A2(KEYINPUT15), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n425), .B(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G475), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT90), .ZN(new_n431));
  INV_X1    g245(.A(G140), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(G125), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n280), .A2(G140), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n433), .A2(new_n434), .A3(KEYINPUT16), .ZN(new_n435));
  OR3_X1    g249(.A1(new_n280), .A2(KEYINPUT16), .A3(G140), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(G146), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(G146), .B1(new_n435), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NOR2_X1   g253(.A1(G237), .A2(G953), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n440), .A2(G143), .A3(G214), .ZN(new_n441));
  AOI21_X1  g255(.A(G143), .B1(new_n440), .B2(G214), .ZN(new_n442));
  OAI21_X1  g256(.A(G131), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n440), .A2(G214), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(new_n251), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n440), .A2(G143), .A3(G214), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n445), .A2(new_n347), .A3(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT17), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n443), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  OAI211_X1 g263(.A(KEYINPUT17), .B(G131), .C1(new_n441), .C2(new_n442), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n439), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  XNOR2_X1  g265(.A(G125), .B(G140), .ZN(new_n452));
  XNOR2_X1  g266(.A(new_n452), .B(new_n254), .ZN(new_n453));
  OAI211_X1 g267(.A(KEYINPUT18), .B(G131), .C1(new_n441), .C2(new_n442), .ZN(new_n454));
  NAND2_X1  g268(.A1(KEYINPUT18), .A2(G131), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n445), .A2(new_n446), .A3(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n451), .A2(new_n457), .ZN(new_n458));
  XNOR2_X1  g272(.A(G113), .B(G122), .ZN(new_n459));
  XNOR2_X1  g273(.A(new_n459), .B(new_n194), .ZN(new_n460));
  INV_X1    g274(.A(new_n460), .ZN(new_n461));
  OAI21_X1  g275(.A(new_n431), .B1(new_n458), .B2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n451), .A2(KEYINPUT90), .A3(new_n460), .A4(new_n457), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT91), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n458), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n451), .A2(KEYINPUT91), .A3(new_n457), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n466), .A2(new_n461), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n464), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n430), .B1(new_n469), .B2(new_n289), .ZN(new_n470));
  AND3_X1   g284(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT87), .B(KEYINPUT19), .ZN(new_n472));
  OR2_X1    g286(.A1(new_n452), .A2(new_n472), .ZN(new_n473));
  INV_X1    g287(.A(KEYINPUT19), .ZN(new_n474));
  OAI211_X1 g288(.A(new_n433), .B(new_n434), .C1(KEYINPUT87), .C2(new_n474), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n473), .A2(KEYINPUT88), .A3(new_n254), .A4(new_n475), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n475), .B(new_n254), .C1(new_n452), .C2(new_n472), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT88), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n476), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n437), .B1(new_n443), .B2(new_n447), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n471), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n460), .B1(new_n482), .B2(KEYINPUT89), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT89), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n480), .A2(new_n481), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n484), .B1(new_n485), .B2(new_n471), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(new_n464), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT20), .ZN(new_n489));
  NOR2_X1   g303(.A1(G475), .A2(G902), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n488), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  AOI22_X1  g305(.A1(new_n483), .A2(new_n486), .B1(new_n462), .B2(new_n463), .ZN(new_n492));
  INV_X1    g306(.A(new_n490), .ZN(new_n493));
  OAI21_X1  g307(.A(KEYINPUT20), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n470), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n429), .A2(new_n495), .ZN(new_n496));
  NOR3_X1   g310(.A1(new_n332), .A2(new_n389), .A3(new_n496), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n421), .B1(G234), .B2(new_n289), .ZN(new_n498));
  INV_X1    g312(.A(KEYINPUT23), .ZN(new_n499));
  OAI21_X1  g313(.A(new_n499), .B1(new_n226), .B2(G128), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n226), .A2(G128), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n269), .A2(KEYINPUT23), .A3(G119), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G119), .B(G128), .ZN(new_n504));
  INV_X1    g318(.A(G110), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n505), .A2(KEYINPUT24), .ZN(new_n506));
  INV_X1    g320(.A(KEYINPUT24), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n507), .A2(G110), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  AOI22_X1  g323(.A1(new_n503), .A2(G110), .B1(new_n504), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n437), .B2(new_n438), .ZN(new_n511));
  XOR2_X1   g325(.A(KEYINPUT74), .B(G110), .Z(new_n512));
  OAI22_X1  g326(.A1(new_n503), .A2(new_n512), .B1(new_n504), .B2(new_n509), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n435), .A2(new_n436), .A3(G146), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n452), .A2(new_n254), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n342), .A2(KEYINPUT22), .ZN(new_n518));
  INV_X1    g332(.A(KEYINPUT22), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n519), .A2(G137), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n518), .A2(new_n520), .A3(KEYINPUT75), .ZN(new_n521));
  INV_X1    g335(.A(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(KEYINPUT75), .B1(new_n518), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g337(.A(KEYINPUT76), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n525));
  NOR2_X1   g339(.A1(new_n519), .A2(G137), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n342), .A2(KEYINPUT22), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n525), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT76), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n521), .ZN(new_n530));
  INV_X1    g344(.A(G234), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n384), .A2(new_n531), .A3(G953), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n524), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  INV_X1    g347(.A(new_n533), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n532), .B1(new_n524), .B2(new_n530), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n517), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n532), .ZN(new_n537));
  INV_X1    g351(.A(new_n530), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n529), .B1(new_n528), .B2(new_n521), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n540), .A2(new_n511), .A3(new_n516), .A4(new_n533), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(KEYINPUT25), .B1(new_n542), .B2(new_n289), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT25), .ZN(new_n544));
  AOI211_X1 g358(.A(new_n544), .B(G902), .C1(new_n536), .C2(new_n541), .ZN(new_n545));
  OAI21_X1  g359(.A(new_n498), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(KEYINPUT77), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT77), .ZN(new_n548));
  OAI211_X1 g362(.A(new_n548), .B(new_n498), .C1(new_n543), .C2(new_n545), .ZN(new_n549));
  NOR2_X1   g363(.A1(new_n498), .A2(G902), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n542), .A2(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n547), .A2(new_n549), .A3(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n344), .ZN(new_n554));
  NOR2_X1   g368(.A1(new_n340), .A2(G137), .ZN(new_n555));
  OAI21_X1  g369(.A(G131), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(new_n348), .ZN(new_n557));
  OR2_X1    g371(.A1(new_n279), .A2(new_n557), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n349), .A2(new_n261), .A3(new_n266), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n558), .A2(new_n192), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n440), .A2(G210), .ZN(new_n561));
  XOR2_X1   g375(.A(new_n561), .B(KEYINPUT27), .Z(new_n562));
  XNOR2_X1  g376(.A(KEYINPUT26), .B(G101), .ZN(new_n563));
  XOR2_X1   g377(.A(new_n562), .B(new_n563), .Z(new_n564));
  AND2_X1   g378(.A1(new_n560), .A2(new_n564), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n566));
  NOR2_X1   g380(.A1(new_n279), .A2(new_n557), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n559), .A2(KEYINPUT68), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT68), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n292), .A2(new_n569), .A3(new_n349), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n567), .B1(new_n568), .B2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT64), .B(KEYINPUT30), .ZN(new_n572));
  OAI21_X1  g386(.A(KEYINPUT69), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n292), .A2(new_n569), .A3(new_n349), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n569), .B1(new_n292), .B2(new_n349), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n558), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT69), .ZN(new_n577));
  INV_X1    g391(.A(new_n572), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n573), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n558), .A2(KEYINPUT30), .A3(new_n559), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n237), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n566), .B1(new_n580), .B2(new_n583), .ZN(new_n584));
  AOI211_X1 g398(.A(KEYINPUT70), .B(new_n582), .C1(new_n573), .C2(new_n579), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n565), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT31), .ZN(new_n587));
  XNOR2_X1  g401(.A(new_n560), .B(KEYINPUT28), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n576), .A2(new_n237), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n564), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT71), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT31), .ZN(new_n593));
  OAI211_X1 g407(.A(new_n593), .B(new_n565), .C1(new_n584), .C2(new_n585), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n592), .A3(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT32), .ZN(new_n596));
  NOR3_X1   g410(.A1(new_n596), .A2(G472), .A3(G902), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n595), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n588), .A2(new_n589), .A3(new_n564), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT29), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n560), .B1(new_n584), .B2(new_n585), .ZN(new_n602));
  INV_X1    g416(.A(new_n564), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n567), .B1(new_n349), .B2(new_n292), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n605), .A2(new_n192), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n588), .A2(new_n607), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n608), .A2(KEYINPUT29), .A3(new_n564), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n609), .A2(new_n289), .ZN(new_n610));
  OAI21_X1  g424(.A(G472), .B1(new_n604), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n598), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT72), .B(KEYINPUT32), .Z(new_n613));
  NOR2_X1   g427(.A1(G472), .A2(G902), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n613), .B1(new_n595), .B2(new_n614), .ZN(new_n615));
  OAI211_X1 g429(.A(new_n497), .B(new_n553), .C1(new_n612), .C2(new_n615), .ZN(new_n616));
  XOR2_X1   g430(.A(new_n616), .B(new_n201), .Z(G3));
  INV_X1    g431(.A(G472), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n618), .B1(new_n595), .B2(new_n289), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n619), .B1(new_n595), .B2(new_n614), .ZN(new_n620));
  INV_X1    g434(.A(new_n470), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n489), .B1(new_n488), .B2(new_n490), .ZN(new_n622));
  NOR3_X1   g436(.A1(new_n492), .A2(KEYINPUT20), .A3(new_n493), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n621), .B1(new_n622), .B2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n420), .A2(new_n423), .ZN(new_n625));
  INV_X1    g439(.A(KEYINPUT33), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  AOI21_X1  g441(.A(new_n422), .B1(new_n420), .B2(KEYINPUT95), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT95), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n412), .A2(new_n419), .A3(new_n629), .ZN(new_n630));
  AOI21_X1  g444(.A(KEYINPUT96), .B1(new_n628), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n410), .A2(new_n408), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n401), .A2(new_n196), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n634), .B1(new_n403), .B2(new_n399), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n414), .A2(new_n418), .ZN(new_n636));
  OAI21_X1  g450(.A(KEYINPUT95), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  AND4_X1   g451(.A1(KEYINPUT96), .A2(new_n637), .A3(new_n630), .A4(new_n423), .ZN(new_n638));
  OAI21_X1  g452(.A(new_n627), .B1(new_n631), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n424), .A2(new_n626), .ZN(new_n640));
  NOR2_X1   g454(.A1(new_n426), .A2(G902), .ZN(new_n641));
  NAND3_X1  g455(.A1(new_n639), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n425), .A2(new_n426), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n624), .A2(new_n644), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n317), .A2(new_n318), .A3(new_n187), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n187), .B1(new_n317), .B2(new_n318), .ZN(new_n647));
  OAI21_X1  g461(.A(new_n331), .B1(new_n646), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n648), .A2(KEYINPUT94), .ZN(new_n649));
  INV_X1    g463(.A(KEYINPUT94), .ZN(new_n650));
  OAI211_X1 g464(.A(new_n650), .B(new_n331), .C1(new_n646), .C2(new_n647), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n329), .B(new_n645), .C1(new_n649), .C2(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n389), .A2(new_n552), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n620), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(KEYINPUT34), .B(G104), .Z(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G6));
  AOI21_X1  g470(.A(new_n470), .B1(new_n622), .B2(KEYINPUT97), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT97), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n491), .A2(new_n494), .A3(new_n658), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n657), .A2(new_n428), .A3(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n329), .B(new_n660), .C1(new_n649), .C2(new_n651), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n620), .A2(new_n653), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT35), .B(G107), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G9));
  INV_X1    g478(.A(KEYINPUT98), .ZN(new_n665));
  INV_X1    g479(.A(KEYINPUT36), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n666), .B1(new_n534), .B2(new_n535), .ZN(new_n667));
  XOR2_X1   g481(.A(new_n667), .B(new_n517), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n550), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n547), .A2(new_n669), .A3(new_n549), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n620), .A2(new_n665), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n595), .A2(new_n289), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n672), .A2(G472), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n595), .A2(new_n614), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n673), .A2(new_n674), .A3(new_n670), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n675), .A2(KEYINPUT98), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n671), .A2(new_n497), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g491(.A(KEYINPUT37), .B(G110), .Z(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(KEYINPUT99), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n677), .B(new_n679), .ZN(G12));
  INV_X1    g494(.A(new_n613), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n674), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n682), .A2(new_n598), .A3(new_n611), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n383), .A2(new_n388), .A3(new_n670), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n684), .B1(new_n649), .B2(new_n651), .ZN(new_n685));
  INV_X1    g499(.A(G900), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n325), .B1(new_n686), .B2(new_n328), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n660), .A2(new_n687), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G128), .ZN(G30));
  XOR2_X1   g504(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n691));
  XNOR2_X1  g505(.A(new_n320), .B(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n624), .A2(new_n428), .ZN(new_n693));
  INV_X1    g507(.A(new_n331), .ZN(new_n694));
  NOR3_X1   g508(.A1(new_n693), .A2(new_n694), .A3(new_n670), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT40), .ZN(new_n697));
  AND2_X1   g511(.A1(new_n383), .A2(new_n388), .ZN(new_n698));
  XOR2_X1   g512(.A(new_n687), .B(KEYINPUT39), .Z(new_n699));
  NAND2_X1  g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(new_n700), .ZN(new_n701));
  AOI21_X1  g515(.A(new_n696), .B1(new_n697), .B2(new_n701), .ZN(new_n702));
  AND2_X1   g516(.A1(new_n602), .A2(new_n564), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n603), .A2(new_n560), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n289), .B1(new_n704), .B2(new_n606), .ZN(new_n705));
  OAI21_X1  g519(.A(G472), .B1(new_n703), .B2(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n682), .A2(new_n598), .A3(new_n706), .ZN(new_n707));
  OAI211_X1 g521(.A(new_n702), .B(new_n707), .C1(new_n697), .C2(new_n701), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G143), .ZN(G45));
  INV_X1    g523(.A(new_n687), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n624), .A2(new_n644), .A3(new_n710), .ZN(new_n711));
  INV_X1    g525(.A(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n683), .A2(new_n685), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G146), .ZN(G48));
  INV_X1    g528(.A(new_n375), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n374), .B1(new_n373), .B2(new_n289), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n715), .A2(new_n387), .A3(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(new_n717), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n718), .A2(new_n552), .ZN(new_n719));
  OAI211_X1 g533(.A(new_n652), .B(new_n719), .C1(new_n612), .C2(new_n615), .ZN(new_n720));
  XNOR2_X1  g534(.A(KEYINPUT41), .B(G113), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(KEYINPUT101), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n720), .B(new_n722), .ZN(G15));
  OAI211_X1 g537(.A(new_n661), .B(new_n719), .C1(new_n612), .C2(new_n615), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  AOI21_X1  g539(.A(new_n329), .B1(new_n649), .B2(new_n651), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n373), .A2(new_n289), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n727), .A2(G469), .ZN(new_n728));
  NAND4_X1  g542(.A1(new_n728), .A2(new_n670), .A3(new_n388), .A4(new_n375), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n729), .A2(new_n496), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n726), .B(new_n730), .C1(new_n612), .C2(new_n615), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(G119), .ZN(G21));
  OR2_X1    g546(.A1(new_n608), .A2(new_n564), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n587), .A2(new_n594), .A3(new_n733), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(KEYINPUT102), .A3(new_n614), .ZN(new_n735));
  INV_X1    g549(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT102), .B1(new_n734), .B2(new_n614), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n736), .A2(new_n619), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n693), .B1(new_n649), .B2(new_n651), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n718), .A2(new_n329), .ZN(new_n740));
  NAND4_X1  g554(.A1(new_n738), .A2(new_n553), .A3(new_n739), .A4(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(G122), .ZN(G24));
  NOR2_X1   g556(.A1(new_n619), .A2(new_n737), .ZN(new_n743));
  AOI211_X1 g557(.A(new_n711), .B(new_n729), .C1(new_n649), .C2(new_n651), .ZN(new_n744));
  NAND3_X1  g558(.A1(new_n743), .A2(new_n744), .A3(new_n735), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G125), .ZN(G27));
  INV_X1    g560(.A(KEYINPUT105), .ZN(new_n747));
  INV_X1    g561(.A(KEYINPUT103), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n381), .A2(new_n748), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n380), .A2(KEYINPUT103), .A3(new_n364), .A4(new_n368), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n378), .A2(new_n749), .A3(G469), .A4(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(new_n375), .A3(new_n376), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n752), .A2(new_n388), .ZN(new_n753));
  NAND3_X1  g567(.A1(new_n314), .A2(new_n331), .A3(new_n319), .ZN(new_n754));
  NOR3_X1   g568(.A1(new_n753), .A2(new_n711), .A3(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT42), .ZN(new_n756));
  AOI21_X1  g570(.A(KEYINPUT32), .B1(new_n595), .B2(new_n614), .ZN(new_n757));
  OAI211_X1 g571(.A(new_n598), .B(new_n611), .C1(new_n757), .C2(KEYINPUT104), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n757), .A2(KEYINPUT104), .ZN(new_n759));
  OAI211_X1 g573(.A(new_n553), .B(new_n756), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  OAI211_X1 g574(.A(new_n553), .B(new_n755), .C1(new_n612), .C2(new_n615), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT42), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g577(.A(new_n747), .B1(new_n760), .B2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n760), .A2(new_n747), .A3(new_n763), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(new_n767), .B(new_n347), .ZN(G33));
  NOR3_X1   g582(.A1(new_n753), .A2(new_n754), .A3(new_n552), .ZN(new_n769));
  OAI211_X1 g583(.A(new_n688), .B(new_n769), .C1(new_n612), .C2(new_n615), .ZN(new_n770));
  XNOR2_X1  g584(.A(new_n770), .B(G134), .ZN(G36));
  AND2_X1   g585(.A1(new_n642), .A2(new_n643), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n624), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT43), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n774), .A2(new_n670), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n775), .A2(new_n620), .ZN(new_n776));
  AOI21_X1  g590(.A(new_n754), .B1(new_n776), .B2(KEYINPUT44), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n378), .A2(new_n749), .A3(new_n750), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n374), .B1(new_n778), .B2(KEYINPUT45), .ZN(new_n779));
  AND2_X1   g593(.A1(new_n378), .A2(new_n381), .ZN(new_n780));
  OAI21_X1  g594(.A(new_n779), .B1(KEYINPUT45), .B2(new_n780), .ZN(new_n781));
  AOI21_X1  g595(.A(KEYINPUT46), .B1(new_n781), .B2(new_n376), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n782), .A2(new_n715), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n781), .A2(KEYINPUT46), .A3(new_n376), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n387), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AND2_X1   g599(.A1(new_n785), .A2(new_n699), .ZN(new_n786));
  OAI211_X1 g600(.A(new_n777), .B(new_n786), .C1(KEYINPUT44), .C2(new_n776), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G137), .ZN(G39));
  XNOR2_X1  g602(.A(KEYINPUT106), .B(KEYINPUT47), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n785), .A2(new_n789), .ZN(new_n790));
  NOR4_X1   g604(.A1(new_n683), .A2(new_n553), .A3(new_n711), .A4(new_n754), .ZN(new_n791));
  NOR2_X1   g605(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n792));
  OAI211_X1 g606(.A(new_n790), .B(new_n791), .C1(new_n785), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g607(.A(new_n793), .B(G140), .ZN(G42));
  NOR2_X1   g608(.A1(new_n715), .A2(new_n716), .ZN(new_n795));
  XOR2_X1   g609(.A(new_n795), .B(KEYINPUT49), .Z(new_n796));
  NAND4_X1  g610(.A1(new_n773), .A2(new_n553), .A3(new_n388), .A4(new_n331), .ZN(new_n797));
  OR4_X1    g611(.A1(new_n707), .A2(new_n796), .A3(new_n692), .A4(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n598), .A2(new_n706), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n799), .A2(new_n615), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n491), .A2(new_n494), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n801), .A2(new_n621), .B1(new_n642), .B2(new_n643), .ZN(new_n802));
  INV_X1    g616(.A(new_n754), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n717), .A2(new_n803), .ZN(new_n804));
  NOR3_X1   g618(.A1(new_n804), .A2(new_n552), .A3(new_n324), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n800), .A2(new_n802), .A3(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n806), .A2(G952), .A3(new_n322), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n758), .A2(new_n759), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n808), .A2(new_n552), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n774), .A2(new_n325), .ZN(new_n810));
  NOR2_X1   g624(.A1(new_n810), .A2(new_n804), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  XOR2_X1   g626(.A(KEYINPUT114), .B(KEYINPUT48), .Z(new_n813));
  AOI21_X1  g627(.A(new_n807), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n734), .A2(new_n614), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT102), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n673), .A2(new_n817), .A3(new_n553), .A4(new_n735), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n810), .A3(new_n718), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  AOI21_X1  g634(.A(new_n650), .B1(new_n320), .B2(new_n331), .ZN(new_n821));
  AOI211_X1 g635(.A(KEYINPUT94), .B(new_n694), .C1(new_n314), .C2(new_n319), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g637(.A(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n819), .A2(new_n820), .A3(new_n824), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n820), .B1(new_n819), .B2(new_n824), .ZN(new_n826));
  OAI221_X1 g640(.A(new_n814), .B1(new_n825), .B2(new_n826), .C1(new_n812), .C2(new_n813), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n811), .A2(new_n670), .A3(new_n738), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n800), .A2(new_n495), .A3(new_n772), .A4(new_n805), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT112), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n829), .A2(new_n830), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n828), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n790), .B1(new_n785), .B2(new_n792), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n795), .A2(new_n387), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n818), .A2(new_n810), .A3(new_n754), .ZN(new_n837));
  AOI21_X1  g651(.A(new_n833), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n692), .A2(new_n331), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n819), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT50), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n840), .A2(KEYINPUT110), .A3(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(KEYINPUT110), .B1(new_n840), .B2(new_n841), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NAND3_X1  g658(.A1(new_n819), .A2(KEYINPUT50), .A3(new_n839), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT111), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n845), .B(new_n846), .ZN(new_n847));
  OAI21_X1  g661(.A(new_n838), .B1(new_n844), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n848), .A2(KEYINPUT51), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT51), .ZN(new_n850));
  OAI211_X1 g664(.A(new_n838), .B(new_n850), .C1(new_n844), .C2(new_n847), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n827), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT107), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n802), .A2(new_n853), .B1(new_n495), .B2(new_n428), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n645), .A2(KEYINPUT107), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n332), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n856), .A2(new_n674), .A3(new_n673), .A4(new_n653), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n720), .A2(new_n724), .A3(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n740), .A2(new_n739), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n616), .B(new_n731), .C1(new_n818), .C2(new_n859), .ZN(new_n860));
  NOR2_X1   g674(.A1(new_n858), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g675(.A1(new_n743), .A2(new_n670), .A3(new_n735), .A4(new_n755), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n657), .A2(new_n429), .A3(new_n659), .A4(new_n710), .ZN(new_n863));
  NOR3_X1   g677(.A1(new_n684), .A2(new_n863), .A3(new_n754), .ZN(new_n864));
  OAI21_X1  g678(.A(new_n864), .B1(new_n612), .B2(new_n615), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n862), .A2(new_n770), .A3(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(new_n866), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n861), .A2(new_n677), .A3(new_n867), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n767), .A2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  OAI221_X1 g684(.A(new_n685), .B1(new_n688), .B2(new_n712), .C1(new_n612), .C2(new_n615), .ZN(new_n871));
  INV_X1    g685(.A(new_n670), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n752), .A2(new_n872), .A3(new_n388), .A4(new_n710), .ZN(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  OAI211_X1 g688(.A(new_n739), .B(new_n874), .C1(new_n799), .C2(new_n615), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n871), .A2(new_n745), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT52), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n871), .A2(new_n745), .A3(KEYINPUT52), .A4(new_n875), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n869), .A2(new_n870), .A3(new_n880), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n616), .A2(new_n731), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n683), .B(new_n719), .C1(new_n652), .C2(new_n661), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n882), .A2(new_n741), .A3(new_n857), .A4(new_n883), .ZN(new_n884));
  INV_X1    g698(.A(new_n677), .ZN(new_n885));
  NOR3_X1   g699(.A1(new_n884), .A2(new_n885), .A3(new_n866), .ZN(new_n886));
  INV_X1    g700(.A(new_n766), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n764), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n879), .ZN(new_n889));
  AOI21_X1  g703(.A(KEYINPUT108), .B1(new_n878), .B2(new_n879), .ZN(new_n890));
  OAI211_X1 g704(.A(new_n886), .B(new_n888), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  OAI211_X1 g706(.A(KEYINPUT54), .B(new_n881), .C1(new_n892), .C2(new_n870), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT109), .ZN(new_n894));
  NAND4_X1  g708(.A1(new_n862), .A2(KEYINPUT53), .A3(new_n770), .A4(new_n865), .ZN(new_n895));
  INV_X1    g709(.A(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n760), .A2(new_n763), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n861), .A2(new_n896), .A3(new_n677), .A4(new_n897), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n823), .A2(new_n693), .A3(new_n873), .ZN(new_n899));
  AOI22_X1  g713(.A1(new_n738), .A2(new_n744), .B1(new_n707), .B2(new_n899), .ZN(new_n900));
  AOI21_X1  g714(.A(KEYINPUT52), .B1(new_n900), .B2(new_n871), .ZN(new_n901));
  INV_X1    g715(.A(new_n879), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n894), .B1(new_n898), .B2(new_n903), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n884), .A2(new_n885), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n895), .B1(new_n763), .B2(new_n760), .ZN(new_n906));
  NAND4_X1  g720(.A1(new_n905), .A2(KEYINPUT109), .A3(new_n880), .A4(new_n906), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n891), .A2(new_n870), .B1(new_n904), .B2(new_n907), .ZN(new_n908));
  INV_X1    g722(.A(KEYINPUT54), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n852), .A2(new_n893), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n911), .A2(KEYINPUT115), .ZN(new_n912));
  OR2_X1    g726(.A1(G952), .A2(G953), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g728(.A1(new_n911), .A2(KEYINPUT115), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n798), .B1(new_n914), .B2(new_n915), .ZN(G75));
  NOR2_X1   g730(.A1(new_n322), .A2(G952), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n908), .A2(new_n289), .ZN(new_n919));
  AOI21_X1  g733(.A(KEYINPUT56), .B1(new_n919), .B2(G210), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n244), .A2(new_n287), .ZN(new_n921));
  XNOR2_X1  g735(.A(new_n921), .B(new_n285), .ZN(new_n922));
  XNOR2_X1  g736(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n922), .B(new_n923), .Z(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  OAI21_X1  g739(.A(new_n918), .B1(new_n920), .B2(new_n925), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n926), .B1(new_n920), .B2(new_n925), .ZN(G51));
  INV_X1    g741(.A(new_n373), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n904), .A2(new_n907), .ZN(new_n929));
  INV_X1    g743(.A(KEYINPUT108), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n880), .A2(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n878), .A2(KEYINPUT108), .A3(new_n879), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g747(.A(KEYINPUT53), .B1(new_n933), .B2(new_n869), .ZN(new_n934));
  OAI21_X1  g748(.A(KEYINPUT54), .B1(new_n929), .B2(new_n934), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n935), .A2(new_n910), .ZN(new_n936));
  XOR2_X1   g750(.A(new_n376), .B(KEYINPUT117), .Z(new_n937));
  XOR2_X1   g751(.A(new_n937), .B(KEYINPUT57), .Z(new_n938));
  AOI21_X1  g752(.A(new_n928), .B1(new_n936), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT118), .ZN(new_n940));
  INV_X1    g754(.A(new_n781), .ZN(new_n941));
  AOI22_X1  g755(.A1(new_n939), .A2(new_n940), .B1(new_n941), .B2(new_n919), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n935), .A2(new_n910), .ZN(new_n943));
  INV_X1    g757(.A(new_n938), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n373), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT118), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n917), .B1(new_n942), .B2(new_n946), .ZN(G54));
  NAND3_X1  g761(.A1(new_n919), .A2(KEYINPUT58), .A3(G475), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n948), .A2(new_n492), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n948), .A2(new_n492), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(new_n917), .ZN(G60));
  AND2_X1   g765(.A1(new_n639), .A2(new_n640), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n910), .A2(new_n893), .ZN(new_n953));
  NAND2_X1  g767(.A1(G478), .A2(G902), .ZN(new_n954));
  XNOR2_X1  g768(.A(new_n954), .B(KEYINPUT59), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n953), .B2(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n952), .A2(new_n955), .ZN(new_n957));
  AOI211_X1 g771(.A(new_n917), .B(new_n956), .C1(new_n936), .C2(new_n957), .ZN(G63));
  INV_X1    g772(.A(new_n542), .ZN(new_n959));
  NAND2_X1  g773(.A1(G217), .A2(G902), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT60), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n959), .B1(new_n908), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n961), .ZN(new_n963));
  OAI211_X1 g777(.A(new_n668), .B(new_n963), .C1(new_n929), .C2(new_n934), .ZN(new_n964));
  NAND3_X1  g778(.A1(new_n962), .A2(new_n964), .A3(new_n918), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n965), .A2(KEYINPUT120), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT119), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT61), .B1(new_n964), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(KEYINPUT120), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n962), .A2(new_n964), .A3(new_n969), .A4(new_n918), .ZN(new_n970));
  AND3_X1   g784(.A1(new_n966), .A2(new_n968), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n968), .B1(new_n966), .B2(new_n970), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n971), .A2(new_n972), .ZN(G66));
  OAI21_X1  g787(.A(G953), .B1(new_n326), .B2(new_n283), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n974), .B1(new_n905), .B2(G953), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n921), .B1(G898), .B2(new_n322), .ZN(new_n976));
  XNOR2_X1  g790(.A(new_n975), .B(new_n976), .ZN(G69));
  AND2_X1   g791(.A1(new_n871), .A2(new_n745), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n978), .A2(new_n708), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT121), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  OR2_X1    g796(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n854), .A2(new_n855), .ZN(new_n984));
  NOR2_X1   g798(.A1(new_n700), .A2(new_n754), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n683), .A2(new_n553), .A3(new_n984), .A4(new_n985), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n983), .A2(new_n787), .A3(new_n793), .A4(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(KEYINPUT122), .B1(new_n982), .B2(new_n987), .ZN(new_n988));
  INV_X1    g802(.A(new_n987), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT122), .ZN(new_n990));
  NAND3_X1  g804(.A1(new_n989), .A2(new_n990), .A3(new_n981), .ZN(new_n991));
  AOI21_X1  g805(.A(G953), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n580), .A2(new_n581), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n473), .A2(new_n475), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n994), .B(new_n995), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  NAND3_X1  g811(.A1(new_n993), .A2(KEYINPUT123), .A3(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n787), .A2(new_n770), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n786), .A2(new_n739), .A3(new_n809), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n1000), .A2(new_n793), .A3(new_n978), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  AOI21_X1  g816(.A(G953), .B1(new_n1002), .B2(new_n888), .ZN(new_n1003));
  INV_X1    g817(.A(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(KEYINPUT125), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n322), .A2(G900), .ZN(new_n1006));
  INV_X1    g820(.A(new_n1006), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n1004), .A2(new_n1005), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(KEYINPUT125), .B1(new_n1003), .B2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n996), .ZN(new_n1011));
  INV_X1    g825(.A(KEYINPUT123), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1012), .B1(new_n992), .B2(new_n996), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n322), .B1(G227), .B2(G900), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1014), .B(KEYINPUT124), .ZN(new_n1015));
  NAND4_X1  g829(.A1(new_n998), .A2(new_n1011), .A3(new_n1013), .A4(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n997), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1017));
  NOR2_X1   g831(.A1(new_n992), .A2(new_n996), .ZN(new_n1018));
  OAI21_X1  g832(.A(new_n1014), .B1(new_n1017), .B2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1016), .A2(new_n1019), .ZN(G72));
  OAI21_X1  g834(.A(new_n881), .B1(new_n892), .B2(new_n870), .ZN(new_n1021));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  INV_X1    g838(.A(new_n584), .ZN(new_n1025));
  INV_X1    g839(.A(new_n585), .ZN(new_n1026));
  AOI21_X1  g840(.A(new_n704), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NOR3_X1   g841(.A1(new_n703), .A2(new_n1024), .A3(new_n1027), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT127), .Z(new_n1029));
  NAND3_X1  g843(.A1(new_n1002), .A2(new_n888), .A3(new_n905), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(new_n1023), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1027), .B(KEYINPUT126), .Z(new_n1032));
  OAI221_X1 g846(.A(new_n918), .B1(new_n1021), .B2(new_n1029), .C1(new_n1031), .C2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n988), .A2(new_n905), .A3(new_n991), .ZN(new_n1034));
  NAND2_X1  g848(.A1(new_n1034), .A2(new_n1023), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1033), .B1(new_n703), .B2(new_n1035), .ZN(G57));
endmodule


