//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 0 1 0 0 1 0 0 0 0 0 1 0 0 1 0 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 0 1 0 1 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:53 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n706, new_n708, new_n709, new_n711, new_n712, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n956, new_n957, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  XNOR2_X1  g000(.A(G113), .B(G122), .ZN(new_n187));
  INV_X1    g001(.A(G104), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n187), .B(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(G237), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n190), .A2(new_n191), .A3(G214), .ZN(new_n192));
  INV_X1    g006(.A(G143), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n190), .A2(new_n191), .A3(G143), .A4(G214), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G131), .ZN(new_n197));
  INV_X1    g011(.A(G131), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n194), .A2(new_n198), .A3(new_n195), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT17), .ZN(new_n201));
  MUX2_X1   g015(.A(new_n197), .B(new_n200), .S(new_n201), .Z(new_n202));
  INV_X1    g016(.A(G125), .ZN(new_n203));
  OAI21_X1  g017(.A(G140), .B1(new_n203), .B2(KEYINPUT74), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  INV_X1    g019(.A(G140), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G125), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n204), .A2(new_n207), .A3(KEYINPUT16), .ZN(new_n208));
  OR3_X1    g022(.A1(new_n203), .A2(KEYINPUT16), .A3(G140), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(G146), .A3(new_n209), .ZN(new_n210));
  AOI21_X1  g024(.A(G146), .B1(new_n208), .B2(new_n209), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT75), .ZN(new_n212));
  OAI21_X1  g026(.A(new_n210), .B1(new_n211), .B2(new_n212), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n213), .B1(new_n212), .B2(new_n211), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n202), .A2(new_n214), .ZN(new_n215));
  AND2_X1   g029(.A1(new_n204), .A2(new_n207), .ZN(new_n216));
  INV_X1    g030(.A(G146), .ZN(new_n217));
  OR2_X1    g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(KEYINPUT65), .B(G146), .ZN(new_n219));
  XNOR2_X1  g033(.A(G125), .B(G140), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT76), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n219), .A2(new_n220), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n221), .B1(new_n219), .B2(new_n220), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n218), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(KEYINPUT18), .A2(G131), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI21_X1  g041(.A(KEYINPUT91), .B1(new_n196), .B2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT91), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n194), .A2(new_n229), .A3(new_n195), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n196), .A2(new_n227), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n225), .A2(new_n231), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT92), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  INV_X1    g049(.A(new_n224), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n236), .A2(new_n222), .ZN(new_n237));
  AOI22_X1  g051(.A1(new_n237), .A2(new_n218), .B1(new_n196), .B2(new_n227), .ZN(new_n238));
  AOI21_X1  g052(.A(KEYINPUT92), .B1(new_n238), .B2(new_n231), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n189), .B(new_n215), .C1(new_n235), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT93), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n233), .A2(new_n234), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n238), .A2(KEYINPUT92), .A3(new_n231), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n243), .A2(new_n244), .B1(new_n214), .B2(new_n202), .ZN(new_n245));
  AOI21_X1  g059(.A(KEYINPUT93), .B1(new_n245), .B2(new_n189), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n244), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n217), .A2(KEYINPUT65), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT65), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G146), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n248), .A2(new_n250), .ZN(new_n251));
  NOR2_X1   g065(.A1(new_n220), .A2(KEYINPUT19), .ZN(new_n252));
  AOI21_X1  g066(.A(new_n252), .B1(new_n216), .B2(KEYINPUT19), .ZN(new_n253));
  OAI211_X1 g067(.A(new_n200), .B(new_n210), .C1(new_n251), .C2(new_n253), .ZN(new_n254));
  AND2_X1   g068(.A1(new_n247), .A2(new_n254), .ZN(new_n255));
  OAI22_X1  g069(.A1(new_n242), .A2(new_n246), .B1(new_n189), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT20), .ZN(new_n257));
  NOR2_X1   g071(.A1(G475), .A2(G902), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n189), .B1(new_n247), .B2(new_n254), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n240), .A2(new_n241), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n245), .A2(KEYINPUT93), .A3(new_n189), .ZN(new_n262));
  AOI21_X1  g076(.A(new_n260), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(new_n258), .ZN(new_n264));
  OAI21_X1  g078(.A(KEYINPUT20), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n259), .A2(new_n265), .ZN(new_n266));
  NOR2_X1   g080(.A1(new_n245), .A2(new_n189), .ZN(new_n267));
  AOI21_X1  g081(.A(new_n267), .B1(new_n261), .B2(new_n262), .ZN(new_n268));
  OAI21_X1  g082(.A(G475), .B1(new_n268), .B2(G902), .ZN(new_n269));
  INV_X1    g083(.A(G902), .ZN(new_n270));
  INV_X1    g084(.A(G122), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n271), .A2(G116), .ZN(new_n272));
  INV_X1    g086(.A(G116), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G122), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n272), .A2(new_n274), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n275), .A2(G107), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n273), .A2(KEYINPUT14), .A3(G122), .ZN(new_n277));
  OAI211_X1 g091(.A(G107), .B(new_n277), .C1(new_n275), .C2(KEYINPUT14), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT94), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n276), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(KEYINPUT66), .B(G128), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G143), .ZN(new_n282));
  INV_X1    g096(.A(G134), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n193), .A2(G128), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n283), .B1(new_n282), .B2(new_n284), .ZN(new_n287));
  OAI221_X1 g101(.A(new_n280), .B1(new_n279), .B2(new_n278), .C1(new_n286), .C2(new_n287), .ZN(new_n288));
  XOR2_X1   g102(.A(new_n284), .B(KEYINPUT13), .Z(new_n289));
  INV_X1    g103(.A(new_n282), .ZN(new_n290));
  OAI21_X1  g104(.A(G134), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(G107), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n292), .B1(new_n272), .B2(new_n274), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n291), .B(new_n285), .C1(new_n293), .C2(new_n276), .ZN(new_n294));
  XNOR2_X1  g108(.A(KEYINPUT9), .B(G234), .ZN(new_n295));
  INV_X1    g109(.A(G217), .ZN(new_n296));
  NOR3_X1   g110(.A1(new_n295), .A2(new_n296), .A3(G953), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n288), .A2(new_n294), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n297), .B1(new_n288), .B2(new_n294), .ZN(new_n300));
  OAI21_X1  g114(.A(new_n270), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G478), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n302), .A2(KEYINPUT15), .ZN(new_n303));
  AND2_X1   g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g118(.A1(new_n301), .A2(new_n303), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  XNOR2_X1  g120(.A(KEYINPUT95), .B(G952), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n307), .A2(G953), .ZN(new_n308));
  NAND2_X1  g122(.A1(G234), .A2(G237), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT21), .B(G898), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n309), .A2(G902), .A3(G953), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(new_n311), .B1(new_n312), .B2(new_n314), .ZN(new_n315));
  INV_X1    g129(.A(new_n315), .ZN(new_n316));
  NAND4_X1  g130(.A1(new_n266), .A2(new_n269), .A3(new_n306), .A4(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT80), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n319), .A2(new_n292), .A3(G104), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(KEYINPUT3), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT3), .ZN(new_n322));
  NAND4_X1  g136(.A1(new_n319), .A2(new_n322), .A3(new_n292), .A4(G104), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n292), .A2(G104), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n321), .A2(new_n323), .A3(new_n325), .ZN(new_n326));
  AND2_X1   g140(.A1(new_n326), .A2(G101), .ZN(new_n327));
  AOI21_X1  g141(.A(G101), .B1(new_n188), .B2(G107), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n321), .A2(new_n323), .A3(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT81), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n329), .A2(KEYINPUT4), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT81), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n326), .A2(G101), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n332), .A2(new_n333), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n248), .A2(new_n250), .A3(G143), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n193), .A2(G146), .ZN(new_n338));
  AND2_X1   g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AND2_X1   g153(.A1(KEYINPUT0), .A2(G128), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n193), .A2(G146), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n342), .B1(new_n219), .B2(G143), .ZN(new_n343));
  NOR2_X1   g157(.A1(KEYINPUT0), .A2(G128), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n340), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g159(.A1(new_n339), .A2(new_n340), .B1(new_n343), .B2(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(G101), .ZN(new_n347));
  NOR2_X1   g161(.A1(new_n347), .A2(KEYINPUT4), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n326), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT82), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n326), .A2(KEYINPUT82), .A3(new_n348), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n336), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT11), .ZN(new_n355));
  OAI21_X1  g169(.A(new_n355), .B1(new_n283), .B2(G137), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n283), .A2(G137), .ZN(new_n357));
  INV_X1    g171(.A(G137), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n358), .A2(KEYINPUT11), .A3(G134), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n356), .A2(new_n357), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(G131), .ZN(new_n361));
  NAND4_X1  g175(.A1(new_n356), .A2(new_n359), .A3(new_n198), .A4(new_n357), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n188), .A2(G107), .ZN(new_n364));
  OAI21_X1  g178(.A(G101), .B1(new_n364), .B2(new_n324), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n329), .A2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(KEYINPUT10), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT1), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n337), .A2(new_n369), .A3(G128), .A4(new_n338), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n281), .B1(new_n337), .B2(KEYINPUT1), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n341), .B1(new_n251), .B2(new_n193), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n368), .A2(new_n373), .ZN(new_n374));
  OR2_X1    g188(.A1(new_n370), .A2(KEYINPUT83), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n337), .A2(new_n338), .ZN(new_n376));
  OAI21_X1  g190(.A(G128), .B1(new_n341), .B2(new_n369), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n370), .A2(KEYINPUT83), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n366), .B1(new_n375), .B2(new_n378), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n374), .B1(new_n379), .B2(KEYINPUT10), .ZN(new_n380));
  NOR3_X1   g194(.A1(new_n354), .A2(new_n363), .A3(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n363), .ZN(new_n382));
  INV_X1    g196(.A(new_n380), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n336), .A2(new_n346), .A3(new_n353), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g199(.A(G110), .B(G140), .ZN(new_n386));
  INV_X1    g200(.A(G227), .ZN(new_n387));
  NOR2_X1   g201(.A1(new_n387), .A2(G953), .ZN(new_n388));
  XNOR2_X1  g202(.A(new_n386), .B(new_n388), .ZN(new_n389));
  NOR3_X1   g203(.A1(new_n381), .A2(new_n385), .A3(new_n389), .ZN(new_n390));
  XNOR2_X1  g204(.A(new_n389), .B(KEYINPUT79), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n383), .A2(new_n382), .A3(new_n384), .ZN(new_n393));
  INV_X1    g207(.A(new_n366), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n394), .A2(new_n373), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n363), .B1(new_n379), .B2(new_n395), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT84), .ZN(new_n397));
  AOI21_X1  g211(.A(KEYINPUT12), .B1(new_n363), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  OAI221_X1 g213(.A(new_n363), .B1(new_n397), .B2(KEYINPUT12), .C1(new_n379), .C2(new_n395), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n392), .B1(new_n393), .B2(new_n401), .ZN(new_n402));
  OAI21_X1  g216(.A(new_n270), .B1(new_n390), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(G469), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT85), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT85), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n403), .A2(new_n406), .A3(G469), .ZN(new_n407));
  OAI21_X1  g221(.A(new_n389), .B1(new_n381), .B2(new_n385), .ZN(new_n408));
  INV_X1    g222(.A(new_n389), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n393), .A2(new_n401), .A3(new_n409), .ZN(new_n410));
  AOI21_X1  g224(.A(G902), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  XOR2_X1   g225(.A(KEYINPUT86), .B(G469), .Z(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n405), .A2(new_n407), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g228(.A(G221), .B1(new_n295), .B2(G902), .ZN(new_n415));
  AND3_X1   g229(.A1(new_n318), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT32), .ZN(new_n417));
  AND2_X1   g231(.A1(G116), .A2(G119), .ZN(new_n418));
  NOR2_X1   g232(.A1(G116), .A2(G119), .ZN(new_n419));
  NOR2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT2), .B(G113), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT67), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  XNOR2_X1  g236(.A(G116), .B(G119), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT67), .ZN(new_n424));
  OR2_X1    g238(.A1(KEYINPUT2), .A2(G113), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT2), .A2(G113), .ZN(new_n426));
  NAND4_X1  g240(.A1(new_n423), .A2(new_n424), .A3(new_n425), .A4(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n422), .A2(new_n427), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n420), .A2(new_n421), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT69), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n346), .A2(new_n363), .ZN(new_n433));
  INV_X1    g247(.A(new_n357), .ZN(new_n434));
  NOR2_X1   g248(.A1(new_n283), .A2(G137), .ZN(new_n435));
  OAI21_X1  g249(.A(G131), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  AND2_X1   g250(.A1(new_n436), .A2(new_n362), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n373), .A2(new_n437), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n422), .A2(new_n427), .B1(new_n421), .B2(new_n420), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n439), .A2(KEYINPUT69), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n432), .A2(new_n433), .A3(new_n438), .A4(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT28), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n442), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n363), .A2(new_n346), .B1(new_n373), .B2(new_n437), .ZN(new_n445));
  OAI211_X1 g259(.A(new_n443), .B(new_n444), .C1(new_n439), .C2(new_n445), .ZN(new_n446));
  XNOR2_X1  g260(.A(KEYINPUT70), .B(KEYINPUT27), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n190), .A2(new_n191), .A3(G210), .ZN(new_n448));
  XNOR2_X1  g262(.A(new_n447), .B(new_n448), .ZN(new_n449));
  XNOR2_X1  g263(.A(KEYINPUT26), .B(G101), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n446), .A2(new_n452), .ZN(new_n453));
  AND3_X1   g267(.A1(new_n441), .A2(KEYINPUT71), .A3(new_n451), .ZN(new_n454));
  AOI21_X1  g268(.A(KEYINPUT71), .B1(new_n441), .B2(new_n451), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT68), .ZN(new_n457));
  OAI211_X1 g271(.A(new_n457), .B(KEYINPUT30), .C1(new_n445), .C2(KEYINPUT64), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n433), .A2(new_n438), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT64), .ZN(new_n460));
  AOI21_X1  g274(.A(KEYINPUT68), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT30), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n462), .B1(new_n459), .B2(KEYINPUT68), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n430), .B(new_n458), .C1(new_n461), .C2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT31), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n456), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n453), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n456), .A2(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT31), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT72), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n468), .A2(KEYINPUT72), .A3(KEYINPUT31), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n467), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g287(.A1(G472), .A2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  OAI21_X1  g289(.A(new_n417), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n464), .A2(new_n441), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(new_n451), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n446), .A2(new_n452), .ZN(new_n480));
  NOR3_X1   g294(.A1(new_n479), .A2(KEYINPUT29), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n432), .A2(new_n440), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n459), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n443), .A2(new_n444), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n451), .A2(KEYINPUT29), .ZN(new_n485));
  OAI21_X1  g299(.A(new_n270), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G472), .B1(new_n481), .B2(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(KEYINPUT72), .B1(new_n468), .B2(KEYINPUT31), .ZN(new_n488));
  AOI211_X1 g302(.A(new_n470), .B(new_n465), .C1(new_n456), .C2(new_n464), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n466), .B(new_n453), .C1(new_n488), .C2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n490), .A2(KEYINPUT32), .A3(new_n474), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n476), .A2(new_n487), .A3(new_n491), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n296), .B1(G234), .B2(new_n270), .ZN(new_n493));
  INV_X1    g307(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n281), .A2(G119), .ZN(new_n495));
  INV_X1    g309(.A(G128), .ZN(new_n496));
  OAI21_X1  g310(.A(new_n495), .B1(G119), .B2(new_n496), .ZN(new_n497));
  XNOR2_X1  g311(.A(KEYINPUT24), .B(G110), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(KEYINPUT23), .ZN(new_n500));
  INV_X1    g314(.A(G119), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n500), .B1(new_n501), .B2(G128), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT73), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  OAI22_X1  g319(.A1(new_n502), .A2(new_n503), .B1(new_n501), .B2(G128), .ZN(new_n506));
  OAI22_X1  g320(.A1(new_n505), .A2(new_n506), .B1(new_n500), .B2(new_n495), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n499), .B1(new_n507), .B2(G110), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n508), .A2(new_n210), .A3(new_n237), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(G110), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n497), .B2(new_n498), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n509), .B1(new_n214), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n512), .A2(KEYINPUT77), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(KEYINPUT22), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(G137), .ZN(new_n516));
  INV_X1    g330(.A(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT77), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n509), .B(new_n518), .C1(new_n214), .C2(new_n511), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n513), .A2(new_n517), .A3(new_n519), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n520), .A2(KEYINPUT78), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT78), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n513), .A2(new_n522), .A3(new_n517), .A4(new_n519), .ZN(new_n523));
  INV_X1    g337(.A(new_n512), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(new_n516), .ZN(new_n525));
  NAND4_X1  g339(.A1(new_n521), .A2(new_n270), .A3(new_n523), .A4(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n494), .B1(new_n526), .B2(KEYINPUT25), .ZN(new_n527));
  AND2_X1   g341(.A1(new_n521), .A2(new_n525), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT25), .ZN(new_n529));
  NAND4_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n270), .A4(new_n523), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n528), .A2(new_n523), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n493), .A2(G902), .ZN(new_n532));
  AOI22_X1  g346(.A1(new_n527), .A2(new_n530), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  OAI21_X1  g347(.A(G214), .B1(G237), .B2(G902), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT6), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n439), .B1(new_n351), .B2(new_n352), .ZN(new_n537));
  NOR3_X1   g351(.A1(new_n327), .A2(KEYINPUT81), .A3(new_n330), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n333), .B1(new_n332), .B2(new_n334), .ZN(new_n539));
  OAI21_X1  g353(.A(new_n537), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT5), .B1(new_n418), .B2(new_n419), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT5), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n542), .A2(new_n501), .A3(G116), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(G113), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  AOI22_X1  g359(.A1(new_n422), .A2(new_n427), .B1(new_n541), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n394), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G110), .B(G122), .ZN(new_n549));
  INV_X1    g363(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g364(.A(new_n536), .B1(new_n548), .B2(new_n550), .ZN(new_n551));
  INV_X1    g365(.A(KEYINPUT87), .ZN(new_n552));
  AND4_X1   g366(.A1(new_n552), .A2(new_n540), .A3(new_n547), .A4(new_n549), .ZN(new_n553));
  INV_X1    g367(.A(new_n547), .ZN(new_n554));
  AOI21_X1  g368(.A(new_n554), .B1(new_n336), .B2(new_n537), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n552), .B1(new_n555), .B2(new_n549), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n551), .B1(new_n553), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n191), .A2(G224), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n339), .A2(new_n340), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n343), .A2(new_n345), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n203), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n203), .B(new_n370), .C1(new_n371), .C2(new_n372), .ZN(new_n563));
  INV_X1    g377(.A(new_n563), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n559), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  OAI211_X1 g379(.A(new_n563), .B(new_n558), .C1(new_n346), .C2(new_n203), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n548), .A2(new_n536), .A3(new_n550), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n557), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT88), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n557), .A2(KEYINPUT88), .A3(new_n567), .A4(new_n568), .ZN(new_n572));
  XOR2_X1   g386(.A(new_n549), .B(KEYINPUT8), .Z(new_n573));
  AOI21_X1  g387(.A(new_n573), .B1(new_n546), .B2(new_n366), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n544), .B1(KEYINPUT89), .B2(new_n541), .ZN(new_n575));
  INV_X1    g389(.A(KEYINPUT89), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n423), .A2(new_n576), .A3(KEYINPUT5), .ZN(new_n577));
  AOI22_X1  g391(.A1(new_n575), .A2(new_n577), .B1(new_n422), .B2(new_n427), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT90), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n394), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n575), .A2(new_n577), .ZN(new_n581));
  AND3_X1   g395(.A1(new_n581), .A2(new_n579), .A3(new_n428), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n574), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n559), .A2(KEYINPUT7), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n584), .B1(new_n562), .B2(new_n564), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n584), .B1(new_n565), .B2(new_n566), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n588), .B1(new_n553), .B2(new_n556), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n589), .A2(new_n270), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n571), .A2(new_n572), .A3(new_n591), .ZN(new_n592));
  OAI21_X1  g406(.A(G210), .B1(G237), .B2(G902), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n590), .B1(new_n569), .B2(new_n570), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n596), .A2(new_n593), .A3(new_n572), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n535), .B1(new_n595), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n416), .A2(new_n492), .A3(new_n533), .A4(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  AND3_X1   g414(.A1(new_n596), .A2(new_n593), .A3(new_n572), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n593), .B1(new_n596), .B2(new_n572), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n534), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(KEYINPUT96), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT96), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT33), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n608), .B1(new_n299), .B2(new_n300), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n288), .A2(new_n294), .ZN(new_n610));
  INV_X1    g424(.A(new_n297), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n612), .A2(KEYINPUT33), .A3(new_n298), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n302), .A2(G902), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n609), .A2(new_n613), .A3(new_n614), .ZN(new_n615));
  INV_X1    g429(.A(KEYINPUT97), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n301), .A2(new_n302), .ZN(new_n617));
  AND3_X1   g431(.A1(new_n615), .A2(new_n616), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(new_n615), .B2(new_n617), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n266), .B2(new_n269), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NOR2_X1   g436(.A1(new_n622), .A2(new_n315), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n607), .A2(new_n623), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n490), .B2(new_n270), .ZN(new_n626));
  NOR2_X1   g440(.A1(new_n473), .A2(new_n475), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(new_n415), .ZN(new_n629));
  INV_X1    g443(.A(new_n412), .ZN(new_n630));
  AOI211_X1 g444(.A(G902), .B(new_n630), .C1(new_n408), .C2(new_n410), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n631), .B1(new_n404), .B2(KEYINPUT85), .ZN(new_n632));
  AOI21_X1  g446(.A(new_n629), .B1(new_n632), .B2(new_n407), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n628), .A2(new_n633), .A3(new_n533), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n624), .A2(new_n634), .ZN(new_n635));
  XNOR2_X1  g449(.A(KEYINPUT34), .B(G104), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(G6));
  XNOR2_X1  g451(.A(new_n269), .B(KEYINPUT98), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n266), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n639), .A2(new_n306), .A3(new_n315), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n607), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n641), .A2(new_n634), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT35), .B(G107), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  NAND2_X1  g458(.A1(new_n513), .A2(new_n519), .ZN(new_n645));
  NOR3_X1   g459(.A1(new_n645), .A2(KEYINPUT36), .A3(new_n517), .ZN(new_n646));
  NOR2_X1   g460(.A1(new_n517), .A2(KEYINPUT36), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n647), .B1(new_n513), .B2(new_n519), .ZN(new_n648));
  OR2_X1    g462(.A1(new_n646), .A2(new_n648), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n530), .A2(new_n527), .B1(new_n532), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n650), .A2(new_n626), .A3(new_n627), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n416), .A2(new_n598), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n652), .B(G110), .ZN(new_n653));
  XOR2_X1   g467(.A(KEYINPUT99), .B(KEYINPUT37), .Z(new_n654));
  XNOR2_X1  g468(.A(new_n653), .B(new_n654), .ZN(G12));
  INV_X1    g469(.A(new_n650), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n492), .A2(new_n633), .A3(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n306), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n314), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n310), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n638), .A2(new_n266), .A3(new_n658), .A4(new_n661), .ZN(new_n662));
  INV_X1    g476(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n595), .A2(new_n597), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n605), .B1(new_n664), .B2(new_n534), .ZN(new_n665));
  AOI211_X1 g479(.A(KEYINPUT96), .B(new_n535), .C1(new_n595), .C2(new_n597), .ZN(new_n666));
  OAI21_X1  g480(.A(new_n663), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  INV_X1    g481(.A(KEYINPUT100), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n657), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  NAND3_X1  g483(.A1(new_n607), .A2(KEYINPUT100), .A3(new_n663), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  XNOR2_X1  g485(.A(new_n671), .B(G128), .ZN(G30));
  AND2_X1   g486(.A1(new_n476), .A2(new_n491), .ZN(new_n673));
  INV_X1    g487(.A(new_n468), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n451), .B1(new_n483), .B2(new_n441), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n270), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n676), .A2(G472), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n242), .A2(new_n246), .ZN(new_n680));
  OAI21_X1  g494(.A(new_n270), .B1(new_n680), .B2(new_n267), .ZN(new_n681));
  AOI22_X1  g495(.A1(new_n259), .A2(new_n265), .B1(new_n681), .B2(G475), .ZN(new_n682));
  NOR2_X1   g496(.A1(new_n682), .A2(new_n306), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  NOR4_X1   g498(.A1(new_n679), .A2(new_n535), .A3(new_n656), .A4(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n661), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n633), .A2(new_n686), .ZN(new_n687));
  XOR2_X1   g501(.A(new_n687), .B(KEYINPUT40), .Z(new_n688));
  XNOR2_X1  g502(.A(new_n664), .B(KEYINPUT38), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n685), .A2(new_n688), .A3(new_n689), .ZN(new_n690));
  XNOR2_X1  g504(.A(new_n690), .B(G143), .ZN(G45));
  NOR2_X1   g505(.A1(new_n665), .A2(new_n666), .ZN(new_n692));
  INV_X1    g506(.A(new_n661), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n622), .A2(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g509(.A1(new_n692), .A2(new_n657), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(new_n217), .ZN(G48));
  INV_X1    g511(.A(new_n411), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n631), .B1(G469), .B2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n699), .A2(new_n415), .ZN(new_n700));
  AND3_X1   g514(.A1(new_n492), .A2(new_n533), .A3(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n624), .A2(new_n702), .ZN(new_n703));
  XOR2_X1   g517(.A(KEYINPUT41), .B(G113), .Z(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(G15));
  NOR2_X1   g519(.A1(new_n641), .A2(new_n702), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(new_n273), .ZN(G18));
  AND3_X1   g521(.A1(new_n492), .A2(new_n318), .A3(new_n656), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n607), .A2(new_n708), .A3(new_n700), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(G119), .ZN(G21));
  NAND2_X1  g524(.A1(new_n700), .A2(new_n316), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n484), .A2(new_n452), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n469), .A3(new_n466), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n626), .B1(new_n474), .B2(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n533), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(KEYINPUT101), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT101), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n714), .A2(new_n717), .A3(new_n533), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n711), .B1(new_n716), .B2(new_n718), .ZN(new_n719));
  AOI21_X1  g533(.A(KEYINPUT102), .B1(new_n607), .B2(new_n683), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n721));
  AOI211_X1 g535(.A(new_n721), .B(new_n684), .C1(new_n604), .C2(new_n606), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n719), .B1(new_n720), .B2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(KEYINPUT103), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G122), .ZN(G24));
  INV_X1    g539(.A(new_n700), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n692), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(new_n626), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n713), .A2(new_n474), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n656), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(KEYINPUT104), .B1(new_n621), .B2(new_n661), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT104), .ZN(new_n732));
  NOR4_X1   g546(.A1(new_n682), .A2(new_n732), .A3(new_n620), .A4(new_n693), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n730), .A2(new_n731), .A3(new_n733), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n727), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G125), .ZN(G27));
  AND2_X1   g550(.A1(new_n492), .A2(new_n533), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n733), .A2(new_n731), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n629), .B1(new_n404), .B2(new_n413), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n595), .A2(new_n739), .A3(new_n534), .A4(new_n597), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n742));
  OAI211_X1 g556(.A(new_n737), .B(new_n738), .C1(new_n741), .C2(new_n742), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT42), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n492), .A2(new_n533), .ZN(new_n746));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n492), .A2(KEYINPUT106), .A3(new_n533), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g564(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n740), .A2(KEYINPUT105), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NOR3_X1   g567(.A1(new_n733), .A2(new_n731), .A3(new_n744), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n745), .A2(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G131), .ZN(G33));
  AOI21_X1  g571(.A(new_n746), .B1(new_n751), .B2(new_n752), .ZN(new_n758));
  XOR2_X1   g572(.A(new_n662), .B(KEYINPUT107), .Z(new_n759));
  NAND2_X1  g573(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NOR2_X1   g575(.A1(new_n628), .A2(new_n650), .ZN(new_n762));
  OR2_X1    g576(.A1(new_n618), .A2(new_n619), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT108), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n682), .B(new_n763), .C1(new_n764), .C2(KEYINPUT43), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n763), .A2(new_n266), .A3(new_n269), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  XNOR2_X1  g581(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n765), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n762), .A2(new_n769), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT44), .ZN(new_n771));
  OAI21_X1  g585(.A(KEYINPUT109), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n595), .A2(new_n534), .A3(new_n597), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT109), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n762), .A2(new_n769), .A3(new_n775), .A4(KEYINPUT44), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n774), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n777), .A2(KEYINPUT110), .ZN(new_n778));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n772), .A2(new_n779), .A3(new_n774), .A4(new_n776), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n770), .A2(new_n771), .ZN(new_n781));
  INV_X1    g595(.A(new_n402), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n393), .A2(new_n409), .ZN(new_n783));
  OAI211_X1 g597(.A(new_n782), .B(KEYINPUT45), .C1(new_n385), .C2(new_n783), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT45), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n785), .B1(new_n390), .B2(new_n402), .ZN(new_n786));
  NAND3_X1  g600(.A1(new_n784), .A2(G469), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(G469), .A2(G902), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT46), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n791), .A2(new_n413), .ZN(new_n792));
  NOR2_X1   g606(.A1(new_n789), .A2(new_n790), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n415), .B1(new_n792), .B2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n686), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n794), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g610(.A1(new_n778), .A2(new_n780), .A3(new_n781), .A4(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(new_n797), .B(KEYINPUT111), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n798), .B(G137), .ZN(G39));
  AND2_X1   g613(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n794), .A2(KEYINPUT47), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR3_X1   g616(.A1(new_n695), .A2(new_n492), .A3(new_n533), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n802), .A2(new_n774), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  OAI211_X1 g619(.A(new_n607), .B(new_n701), .C1(new_n623), .C2(new_n640), .ZN(new_n806));
  AND2_X1   g620(.A1(new_n806), .A2(new_n709), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n756), .A2(new_n723), .A3(new_n807), .ZN(new_n808));
  AOI22_X1  g622(.A1(new_n758), .A2(new_n759), .B1(new_n753), .B2(new_n734), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n599), .A2(new_n652), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n598), .A2(new_n316), .ZN(new_n811));
  NOR3_X1   g625(.A1(new_n634), .A2(new_n811), .A3(new_n622), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n810), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT112), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n682), .A2(new_n658), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n811), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  INV_X1    g630(.A(new_n634), .ZN(new_n817));
  OAI21_X1  g631(.A(new_n814), .B1(new_n811), .B2(new_n815), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT113), .ZN(new_n820));
  NAND4_X1  g634(.A1(new_n638), .A2(new_n266), .A3(new_n306), .A4(new_n661), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n821), .A2(new_n773), .ZN(new_n822));
  INV_X1    g636(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g637(.A(new_n820), .B1(new_n823), .B2(new_n657), .ZN(new_n824));
  INV_X1    g638(.A(new_n657), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(KEYINPUT113), .A3(new_n822), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n824), .A2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n809), .A2(new_n813), .A3(new_n819), .A4(new_n827), .ZN(new_n828));
  NOR2_X1   g642(.A1(new_n808), .A2(new_n828), .ZN(new_n829));
  OAI21_X1  g643(.A(new_n683), .B1(new_n665), .B2(new_n666), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(new_n721), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n607), .A2(KEYINPUT102), .A3(new_n683), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  AND4_X1   g647(.A1(new_n650), .A2(new_n678), .A3(new_n661), .A4(new_n739), .ZN(new_n834));
  AOI21_X1  g648(.A(new_n696), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  AOI22_X1  g649(.A1(new_n669), .A2(new_n670), .B1(new_n727), .B2(new_n734), .ZN(new_n836));
  AOI21_X1  g650(.A(KEYINPUT52), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT114), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n837), .B1(new_n838), .B2(new_n839), .ZN(new_n840));
  AOI211_X1 g654(.A(KEYINPUT114), .B(KEYINPUT52), .C1(new_n835), .C2(new_n836), .ZN(new_n841));
  OAI211_X1 g655(.A(KEYINPUT53), .B(new_n829), .C1(new_n840), .C2(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT54), .ZN(new_n843));
  AND3_X1   g657(.A1(new_n835), .A2(KEYINPUT52), .A3(new_n836), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n829), .B1(new_n844), .B2(new_n837), .ZN(new_n845));
  INV_X1    g659(.A(KEYINPUT53), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n842), .A2(new_n843), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n769), .A2(new_n311), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n726), .A2(new_n773), .ZN(new_n851));
  AND2_X1   g665(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g666(.A1(new_n852), .A2(new_n656), .A3(new_n714), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n679), .A2(new_n851), .A3(new_n533), .A4(new_n311), .ZN(new_n854));
  OR2_X1    g668(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(KEYINPUT116), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n855), .A2(new_n682), .A3(new_n620), .A4(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n716), .A2(new_n718), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n858), .A2(new_n850), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n689), .A2(new_n726), .A3(new_n534), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(KEYINPUT50), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g677(.A(KEYINPUT50), .B1(new_n859), .B2(new_n860), .ZN(new_n864));
  OAI211_X1 g678(.A(new_n853), .B(new_n857), .C1(new_n863), .C2(new_n864), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n859), .A2(KEYINPUT115), .A3(new_n774), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n699), .A2(new_n629), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n867), .B1(new_n800), .B2(new_n801), .ZN(new_n868));
  INV_X1    g682(.A(KEYINPUT115), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n858), .A2(new_n850), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n869), .B1(new_n870), .B2(new_n773), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n866), .A2(new_n868), .A3(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n849), .B1(new_n865), .B2(new_n873), .ZN(new_n874));
  XNOR2_X1  g688(.A(new_n861), .B(new_n862), .ZN(new_n875));
  AND2_X1   g689(.A1(new_n857), .A2(new_n853), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n875), .A2(new_n876), .A3(KEYINPUT51), .A4(new_n872), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n852), .A2(new_n750), .ZN(new_n878));
  XNOR2_X1  g692(.A(new_n878), .B(KEYINPUT48), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n855), .A2(new_n621), .A3(new_n856), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n859), .A2(new_n727), .ZN(new_n881));
  AND4_X1   g695(.A1(new_n308), .A2(new_n879), .A3(new_n880), .A4(new_n881), .ZN(new_n882));
  AND3_X1   g696(.A1(new_n874), .A2(new_n877), .A3(new_n882), .ZN(new_n883));
  OAI211_X1 g697(.A(new_n829), .B(KEYINPUT53), .C1(new_n844), .C2(new_n837), .ZN(new_n884));
  INV_X1    g698(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n885), .B1(new_n886), .B2(new_n846), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n848), .B(new_n883), .C1(new_n887), .C2(new_n843), .ZN(new_n888));
  OR2_X1    g702(.A1(G952), .A2(G953), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  XOR2_X1   g704(.A(new_n699), .B(KEYINPUT49), .Z(new_n891));
  NOR4_X1   g705(.A1(new_n891), .A2(new_n535), .A3(new_n629), .A4(new_n766), .ZN(new_n892));
  INV_X1    g706(.A(new_n689), .ZN(new_n893));
  NAND4_X1  g707(.A1(new_n892), .A2(new_n533), .A3(new_n893), .A4(new_n679), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n890), .A2(new_n894), .ZN(new_n895));
  INV_X1    g709(.A(KEYINPUT117), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n890), .A2(KEYINPUT117), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(G75));
  INV_X1    g713(.A(KEYINPUT56), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n557), .A2(new_n568), .ZN(new_n901));
  XNOR2_X1  g715(.A(new_n901), .B(new_n567), .ZN(new_n902));
  XNOR2_X1  g716(.A(new_n902), .B(KEYINPUT55), .ZN(new_n903));
  XOR2_X1   g717(.A(new_n903), .B(KEYINPUT118), .Z(new_n904));
  AND2_X1   g718(.A1(new_n842), .A2(new_n847), .ZN(new_n905));
  NAND2_X1  g719(.A1(G210), .A2(G902), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n900), .B(new_n904), .C1(new_n905), .C2(new_n906), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n191), .A2(G952), .ZN(new_n908));
  INV_X1    g722(.A(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(new_n903), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n842), .A2(new_n847), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n912), .A2(G210), .A3(G902), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n911), .B1(new_n913), .B2(new_n900), .ZN(new_n914));
  OAI21_X1  g728(.A(KEYINPUT119), .B1(new_n910), .B2(new_n914), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n913), .A2(new_n900), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n916), .A2(new_n903), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT119), .ZN(new_n918));
  NAND4_X1  g732(.A1(new_n917), .A2(new_n918), .A3(new_n907), .A4(new_n909), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G51));
  XOR2_X1   g734(.A(new_n788), .B(KEYINPUT57), .Z(new_n921));
  INV_X1    g735(.A(new_n848), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n843), .B1(new_n842), .B2(new_n847), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n921), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n408), .A2(new_n410), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OR3_X1    g740(.A1(new_n905), .A2(new_n270), .A3(new_n787), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n908), .B1(new_n926), .B2(new_n927), .ZN(G54));
  AND2_X1   g742(.A1(KEYINPUT58), .A2(G475), .ZN(new_n929));
  NAND4_X1  g743(.A1(new_n912), .A2(G902), .A3(new_n256), .A4(new_n929), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT120), .ZN(new_n931));
  OR2_X1    g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n930), .A2(new_n931), .ZN(new_n933));
  NAND3_X1  g747(.A1(new_n912), .A2(G902), .A3(new_n929), .ZN(new_n934));
  AOI21_X1  g748(.A(new_n908), .B1(new_n934), .B2(new_n263), .ZN(new_n935));
  AND3_X1   g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(G60));
  NAND2_X1  g750(.A1(new_n609), .A2(new_n613), .ZN(new_n937));
  NAND2_X1  g751(.A1(G478), .A2(G902), .ZN(new_n938));
  XOR2_X1   g752(.A(new_n938), .B(KEYINPUT59), .Z(new_n939));
  NOR2_X1   g753(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n922), .B2(new_n923), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT121), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT121), .B(new_n940), .C1(new_n922), .C2(new_n923), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  INV_X1    g759(.A(new_n829), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n835), .A2(new_n836), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT52), .ZN(new_n948));
  NAND2_X1  g762(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n949), .B1(new_n844), .B2(KEYINPUT114), .ZN(new_n950));
  INV_X1    g764(.A(new_n841), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n946), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n884), .B1(new_n952), .B2(KEYINPUT53), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(KEYINPUT54), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n939), .B1(new_n954), .B2(new_n848), .ZN(new_n955));
  INV_X1    g769(.A(new_n937), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n909), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n945), .A2(new_n957), .ZN(G63));
  INV_X1    g772(.A(KEYINPUT61), .ZN(new_n959));
  INV_X1    g773(.A(new_n531), .ZN(new_n960));
  NAND2_X1  g774(.A1(G217), .A2(G902), .ZN(new_n961));
  XOR2_X1   g775(.A(new_n961), .B(KEYINPUT122), .Z(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n960), .B1(new_n905), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n909), .ZN(new_n965));
  INV_X1    g779(.A(new_n649), .ZN(new_n966));
  NOR3_X1   g780(.A1(new_n905), .A2(new_n966), .A3(new_n963), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n959), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g782(.A(new_n967), .ZN(new_n969));
  NAND4_X1  g783(.A1(new_n969), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n964), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n968), .A2(new_n970), .ZN(G66));
  NAND4_X1  g785(.A1(new_n807), .A2(new_n723), .A3(new_n819), .A4(new_n813), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT123), .Z(new_n973));
  NAND2_X1  g787(.A1(G224), .A2(G953), .ZN(new_n974));
  OAI22_X1  g788(.A1(new_n973), .A2(G953), .B1(new_n312), .B2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(G898), .ZN(new_n976));
  AOI21_X1  g790(.A(new_n901), .B1(new_n976), .B2(G953), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n975), .B(new_n977), .ZN(G69));
  INV_X1    g792(.A(new_n696), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n836), .A2(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n797), .A2(new_n981), .ZN(new_n982));
  AND2_X1   g796(.A1(new_n796), .A2(new_n750), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(new_n833), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g799(.A(new_n804), .B1(new_n985), .B2(KEYINPUT124), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n983), .A2(new_n833), .A3(KEYINPUT124), .ZN(new_n987));
  INV_X1    g801(.A(new_n987), .ZN(new_n988));
  NOR3_X1   g802(.A1(new_n982), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n756), .A2(new_n760), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT125), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  NAND2_X1  g806(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n191), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n191), .A2(G900), .ZN(new_n995));
  INV_X1    g809(.A(new_n995), .ZN(new_n996));
  NAND3_X1  g810(.A1(new_n994), .A2(KEYINPUT126), .A3(new_n996), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT126), .ZN(new_n998));
  AOI21_X1  g812(.A(G953), .B1(new_n989), .B2(new_n992), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n998), .B1(new_n999), .B2(new_n995), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n997), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n461), .A2(new_n463), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(KEYINPUT30), .B2(new_n461), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(new_n253), .Z(new_n1004));
  NAND2_X1  g818(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n687), .B1(new_n622), .B2(new_n815), .ZN(new_n1006));
  NAND3_X1  g820(.A1(new_n1006), .A2(new_n737), .A3(new_n774), .ZN(new_n1007));
  NAND3_X1  g821(.A1(new_n797), .A2(new_n804), .A3(new_n1007), .ZN(new_n1008));
  NAND2_X1  g822(.A1(new_n981), .A2(new_n690), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n1008), .B1(KEYINPUT62), .B2(new_n1009), .ZN(new_n1010));
  OR2_X1    g824(.A1(new_n1009), .A2(KEYINPUT62), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1004), .ZN(new_n1013));
  NAND3_X1  g827(.A1(new_n1012), .A2(new_n191), .A3(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(G953), .B1(new_n387), .B2(new_n659), .ZN(new_n1015));
  INV_X1    g829(.A(new_n1015), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n1005), .A2(new_n1014), .A3(new_n1016), .ZN(new_n1017));
  AOI21_X1  g831(.A(new_n1013), .B1(new_n997), .B2(new_n1000), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1014), .ZN(new_n1019));
  OAI21_X1  g833(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1017), .A2(new_n1020), .ZN(G72));
  NAND2_X1  g835(.A1(G472), .A2(G902), .ZN(new_n1022));
  XOR2_X1   g836(.A(new_n1022), .B(KEYINPUT63), .Z(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(new_n1012), .B2(new_n973), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n451), .A3(new_n477), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1023), .B1(new_n993), .B2(new_n973), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n452), .A3(new_n478), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1025), .A2(new_n909), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1023), .ZN(new_n1029));
  INV_X1    g843(.A(new_n479), .ZN(new_n1030));
  AOI21_X1  g844(.A(new_n1029), .B1(new_n1030), .B2(new_n468), .ZN(new_n1031));
  AOI21_X1  g845(.A(new_n1028), .B1(new_n953), .B2(new_n1031), .ZN(G57));
endmodule


