//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 0 0 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 1 0 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:02 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n697, new_n698, new_n699, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n716, new_n717, new_n719, new_n720, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n761, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n782, new_n783, new_n784, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n956, new_n957, new_n958, new_n959, new_n960, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025;
  INV_X1    g000(.A(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G217), .B1(new_n187), .B2(G902), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT72), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT22), .B(G137), .ZN(new_n190));
  INV_X1    g004(.A(G953), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(G221), .A3(G234), .ZN(new_n192));
  XNOR2_X1  g006(.A(new_n190), .B(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G119), .ZN(new_n194));
  OAI21_X1  g008(.A(KEYINPUT73), .B1(new_n194), .B2(G128), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n196));
  INV_X1    g010(.A(G128), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(new_n197), .A3(G119), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n194), .A2(G128), .ZN(new_n199));
  AND3_X1   g013(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G110), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT24), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT24), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G110), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT74), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n202), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n203), .A2(G110), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n201), .A2(KEYINPUT24), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT74), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n200), .A2(new_n206), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n211), .B1(new_n194), .B2(G128), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n197), .A2(KEYINPUT23), .A3(G119), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(new_n199), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n214), .A2(G110), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G140), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(G125), .ZN(new_n218));
  INV_X1    g032(.A(G125), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(G140), .ZN(new_n220));
  NAND3_X1  g034(.A1(new_n218), .A2(new_n220), .A3(KEYINPUT16), .ZN(new_n221));
  OR3_X1    g035(.A1(new_n219), .A2(KEYINPUT16), .A3(G140), .ZN(new_n222));
  AND3_X1   g036(.A1(new_n221), .A2(G146), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(G146), .B1(new_n221), .B2(new_n222), .ZN(new_n224));
  NOR2_X1   g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  OAI21_X1  g039(.A(KEYINPUT75), .B1(new_n216), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n221), .A2(new_n222), .ZN(new_n227));
  INV_X1    g041(.A(G146), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n221), .A2(new_n222), .A3(G146), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT75), .ZN(new_n232));
  NAND4_X1  g046(.A1(new_n231), .A2(new_n232), .A3(new_n210), .A4(new_n215), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n226), .A2(new_n233), .ZN(new_n234));
  AND4_X1   g048(.A1(new_n201), .A2(new_n212), .A3(new_n213), .A4(new_n199), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n209), .A2(new_n206), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n195), .A2(new_n198), .A3(new_n199), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n235), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(G125), .B(G140), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n239), .A2(new_n228), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n230), .A2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(KEYINPUT76), .B1(new_n238), .B2(new_n241), .ZN(new_n242));
  AND2_X1   g056(.A1(new_n230), .A2(new_n240), .ZN(new_n243));
  INV_X1    g057(.A(KEYINPUT76), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n200), .B1(new_n206), .B2(new_n209), .ZN(new_n245));
  OAI211_X1 g059(.A(new_n243), .B(new_n244), .C1(new_n245), .C2(new_n235), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n242), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT77), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n234), .A2(new_n247), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n248), .B1(new_n234), .B2(new_n247), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n193), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G902), .ZN(new_n252));
  INV_X1    g066(.A(new_n193), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n234), .A2(new_n247), .ZN(new_n254));
  OAI21_X1  g068(.A(new_n253), .B1(new_n254), .B2(KEYINPUT77), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n251), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT78), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT25), .ZN(new_n258));
  AND3_X1   g072(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n256), .B2(new_n257), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n189), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g075(.A1(new_n251), .A2(new_n255), .ZN(new_n262));
  AOI21_X1  g076(.A(G902), .B1(new_n187), .B2(G217), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT84), .ZN(new_n266));
  XNOR2_X1  g080(.A(KEYINPUT9), .B(G234), .ZN(new_n267));
  OAI21_X1  g081(.A(G221), .B1(new_n267), .B2(G902), .ZN(new_n268));
  XOR2_X1   g082(.A(new_n268), .B(KEYINPUT79), .Z(new_n269));
  XOR2_X1   g083(.A(new_n269), .B(KEYINPUT80), .Z(new_n270));
  INV_X1    g084(.A(G104), .ZN(new_n271));
  OAI21_X1  g085(.A(KEYINPUT3), .B1(new_n271), .B2(G107), .ZN(new_n272));
  AOI21_X1  g086(.A(G101), .B1(new_n271), .B2(G107), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT3), .ZN(new_n274));
  INV_X1    g088(.A(G107), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n274), .A2(new_n275), .A3(G104), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n272), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT81), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  NAND4_X1  g093(.A1(new_n272), .A2(new_n273), .A3(new_n276), .A4(KEYINPUT81), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT4), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(G107), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n272), .A2(new_n276), .A3(new_n283), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n284), .B2(G101), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n228), .A2(G143), .ZN(new_n287));
  INV_X1    g101(.A(G143), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(G146), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(KEYINPUT0), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n291), .A2(new_n197), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(KEYINPUT64), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n294), .A2(new_n291), .A3(new_n197), .ZN(new_n295));
  OAI21_X1  g109(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n296));
  AOI22_X1  g110(.A1(new_n295), .A2(new_n296), .B1(new_n287), .B2(new_n289), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n297), .B2(new_n292), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n284), .A2(new_n282), .A3(G101), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G101), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n275), .A2(G104), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n301), .B1(new_n302), .B2(new_n283), .ZN(new_n303));
  INV_X1    g117(.A(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n305));
  AOI21_X1  g119(.A(new_n305), .B1(G143), .B2(new_n228), .ZN(new_n306));
  OAI21_X1  g120(.A(new_n290), .B1(new_n306), .B2(new_n197), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n287), .A2(new_n289), .A3(new_n305), .A4(G128), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n281), .A2(new_n304), .A3(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT10), .ZN(new_n311));
  AOI22_X1  g125(.A1(new_n286), .A2(new_n300), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n281), .A2(new_n304), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT82), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n313), .A2(new_n314), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n303), .B1(new_n279), .B2(new_n280), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(KEYINPUT82), .ZN(new_n317));
  INV_X1    g131(.A(KEYINPUT66), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n287), .A2(new_n318), .A3(KEYINPUT1), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G128), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n306), .A2(new_n318), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n290), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n311), .B1(new_n322), .B2(new_n308), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n315), .A2(new_n317), .A3(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(G134), .ZN(new_n325));
  OAI21_X1  g139(.A(KEYINPUT11), .B1(new_n325), .B2(G137), .ZN(new_n326));
  INV_X1    g140(.A(KEYINPUT11), .ZN(new_n327));
  INV_X1    g141(.A(G137), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(new_n328), .A3(G134), .ZN(new_n329));
  AND2_X1   g143(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  OAI21_X1  g144(.A(KEYINPUT65), .B1(new_n328), .B2(G134), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT65), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n332), .A2(new_n325), .A3(G137), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n331), .A2(new_n333), .ZN(new_n334));
  OAI21_X1  g148(.A(G131), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n326), .A2(new_n329), .ZN(new_n336));
  INV_X1    g150(.A(G131), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n336), .A2(new_n337), .A3(new_n331), .A4(new_n333), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n335), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n312), .A2(new_n324), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n322), .A2(new_n308), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n310), .B1(new_n342), .B2(new_n316), .ZN(new_n343));
  INV_X1    g157(.A(new_n338), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n331), .A2(new_n333), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n337), .B1(new_n345), .B2(new_n336), .ZN(new_n346));
  OAI21_X1  g160(.A(KEYINPUT83), .B1(new_n344), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(KEYINPUT12), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  AND3_X1   g163(.A1(new_n343), .A2(new_n339), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(new_n343), .B2(new_n339), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n341), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  XNOR2_X1  g166(.A(G110), .B(G140), .ZN(new_n353));
  INV_X1    g167(.A(G227), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n354), .A2(G953), .ZN(new_n355));
  XNOR2_X1  g169(.A(new_n353), .B(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n312), .A2(new_n324), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n358), .A2(new_n339), .ZN(new_n359));
  INV_X1    g173(.A(new_n356), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n359), .A2(new_n341), .A3(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(G469), .A3(new_n361), .ZN(new_n362));
  NAND2_X1  g176(.A1(G469), .A2(G902), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  AND3_X1   g178(.A1(new_n312), .A2(new_n324), .A3(new_n340), .ZN(new_n365));
  AOI21_X1  g179(.A(new_n340), .B1(new_n312), .B2(new_n324), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n356), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n341), .B(new_n360), .C1(new_n350), .C2(new_n351), .ZN(new_n368));
  AOI211_X1 g182(.A(G469), .B(G902), .C1(new_n367), .C2(new_n368), .ZN(new_n369));
  OAI211_X1 g183(.A(new_n266), .B(new_n270), .C1(new_n364), .C2(new_n369), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n270), .B1(new_n364), .B2(new_n369), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n371), .A2(KEYINPUT84), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n265), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n194), .A2(G116), .ZN(new_n374));
  INV_X1    g188(.A(G116), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(G119), .ZN(new_n376));
  AND2_X1   g190(.A1(new_n374), .A2(new_n376), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT2), .B(G113), .ZN(new_n378));
  XNOR2_X1  g192(.A(new_n377), .B(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n380), .B1(new_n339), .B2(new_n298), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n325), .A2(G137), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n328), .A2(G134), .ZN(new_n383));
  OAI21_X1  g197(.A(G131), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  AND3_X1   g198(.A1(new_n338), .A2(KEYINPUT69), .A3(new_n384), .ZN(new_n385));
  AOI21_X1  g199(.A(KEYINPUT69), .B1(new_n338), .B2(new_n384), .ZN(new_n386));
  OAI21_X1  g200(.A(new_n342), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(KEYINPUT28), .B1(new_n381), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  NOR2_X1   g203(.A1(G237), .A2(G953), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(G210), .ZN(new_n391));
  XOR2_X1   g205(.A(new_n391), .B(KEYINPUT27), .Z(new_n392));
  XNOR2_X1  g206(.A(KEYINPUT26), .B(G101), .ZN(new_n393));
  XNOR2_X1  g207(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT29), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  OAI211_X1 g210(.A(KEYINPUT68), .B(new_n298), .C1(new_n344), .C2(new_n346), .ZN(new_n397));
  INV_X1    g211(.A(new_n397), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT68), .B1(new_n339), .B2(new_n298), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(KEYINPUT70), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT70), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n402), .B(new_n342), .C1(new_n385), .C2(new_n386), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n400), .A2(new_n401), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n338), .A2(new_n384), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT69), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n338), .A2(KEYINPUT69), .A3(new_n384), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AOI21_X1  g223(.A(new_n402), .B1(new_n409), .B2(new_n342), .ZN(new_n410));
  INV_X1    g224(.A(new_n403), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NOR3_X1   g226(.A1(new_n398), .A2(new_n399), .A3(new_n380), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n380), .A2(new_n404), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT28), .ZN(new_n415));
  OAI211_X1 g229(.A(new_n389), .B(new_n396), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n416), .A2(new_n252), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n400), .A2(new_n401), .A3(new_n403), .A4(new_n379), .ZN(new_n418));
  AND2_X1   g232(.A1(new_n338), .A2(new_n384), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n342), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n339), .A2(new_n298), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n422), .A2(new_n380), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n418), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT28), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT71), .ZN(new_n426));
  INV_X1    g240(.A(new_n394), .ZN(new_n427));
  NAND4_X1  g241(.A1(new_n425), .A2(new_n426), .A3(new_n427), .A4(new_n389), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT67), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n342), .A2(new_n419), .B1(new_n339), .B2(new_n298), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n429), .B1(new_n430), .B2(KEYINPUT30), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT30), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n422), .A2(KEYINPUT67), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n431), .A2(new_n433), .ZN(new_n434));
  NAND4_X1  g248(.A1(new_n400), .A2(new_n401), .A3(KEYINPUT30), .A4(new_n403), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n434), .A2(new_n435), .A3(new_n380), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n418), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n394), .ZN(new_n438));
  AND3_X1   g252(.A1(new_n428), .A2(new_n438), .A3(new_n395), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n425), .A2(new_n389), .ZN(new_n440));
  OAI21_X1  g254(.A(KEYINPUT71), .B1(new_n440), .B2(new_n394), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n417), .B1(new_n439), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G472), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n415), .B1(new_n418), .B2(new_n423), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n394), .B1(new_n444), .B2(new_n388), .ZN(new_n445));
  AOI21_X1  g259(.A(new_n394), .B1(new_n412), .B2(new_n413), .ZN(new_n446));
  AND3_X1   g260(.A1(new_n436), .A2(KEYINPUT31), .A3(new_n446), .ZN(new_n447));
  AOI21_X1  g261(.A(KEYINPUT31), .B1(new_n436), .B2(new_n446), .ZN(new_n448));
  OAI21_X1  g262(.A(new_n445), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT32), .ZN(new_n450));
  NOR2_X1   g264(.A1(G472), .A2(G902), .ZN(new_n451));
  AND3_X1   g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g266(.A(new_n450), .B1(new_n449), .B2(new_n451), .ZN(new_n453));
  OAI22_X1  g267(.A1(new_n442), .A2(new_n443), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(G214), .B1(G237), .B2(G902), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  OAI21_X1  g270(.A(G210), .B1(G237), .B2(G902), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n459));
  OAI21_X1  g273(.A(new_n459), .B1(new_n342), .B2(G125), .ZN(new_n460));
  NAND4_X1  g274(.A1(new_n322), .A2(KEYINPUT89), .A3(new_n219), .A4(new_n308), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n191), .A2(G224), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n293), .B(G125), .C1(new_n297), .C2(new_n292), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n464), .B(KEYINPUT88), .ZN(new_n465));
  AND3_X1   g279(.A1(new_n462), .A2(new_n463), .A3(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n463), .B1(new_n462), .B2(new_n465), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n316), .A2(KEYINPUT82), .ZN(new_n469));
  AOI211_X1 g283(.A(new_n314), .B(new_n303), .C1(new_n279), .C2(new_n280), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n377), .A2(KEYINPUT5), .ZN(new_n471));
  NOR2_X1   g285(.A1(new_n374), .A2(KEYINPUT5), .ZN(new_n472));
  INV_X1    g286(.A(G113), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n377), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n378), .ZN(new_n477));
  NOR3_X1   g291(.A1(new_n469), .A2(new_n470), .A3(new_n477), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n380), .A2(new_n286), .A3(new_n299), .ZN(new_n479));
  INV_X1    g293(.A(new_n479), .ZN(new_n480));
  OAI21_X1  g294(.A(KEYINPUT85), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n477), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n315), .A2(new_n482), .A3(new_n317), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT85), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n483), .A2(new_n484), .A3(new_n479), .ZN(new_n485));
  XNOR2_X1  g299(.A(G110), .B(G122), .ZN(new_n486));
  XOR2_X1   g300(.A(new_n486), .B(KEYINPUT86), .Z(new_n487));
  NAND3_X1  g301(.A1(new_n481), .A2(new_n485), .A3(new_n487), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n478), .A2(new_n480), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n489), .B1(new_n490), .B2(new_n486), .ZN(new_n491));
  AND2_X1   g305(.A1(new_n487), .A2(new_n489), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n485), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT87), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n481), .A2(new_n485), .A3(KEYINPUT87), .A4(new_n492), .ZN(new_n496));
  AOI221_X4 g310(.A(new_n468), .B1(new_n488), .B2(new_n491), .C1(new_n495), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n462), .A2(new_n465), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n463), .A2(KEYINPUT7), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n490), .A2(new_n486), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n482), .A2(new_n313), .ZN(new_n502));
  XNOR2_X1  g316(.A(new_n486), .B(KEYINPUT8), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n477), .A2(new_n316), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  OAI21_X1  g320(.A(new_n252), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n458), .B1(new_n497), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n495), .A2(new_n496), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n488), .A2(new_n491), .ZN(new_n510));
  INV_X1    g324(.A(new_n468), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n507), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n512), .A2(new_n513), .A3(new_n457), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n456), .B1(new_n508), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g329(.A1(G475), .A2(G902), .ZN(new_n516));
  XNOR2_X1  g330(.A(G113), .B(G122), .ZN(new_n517));
  XNOR2_X1  g331(.A(new_n517), .B(new_n271), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n519));
  AOI21_X1  g333(.A(G143), .B1(new_n390), .B2(G214), .ZN(new_n520));
  OAI211_X1 g334(.A(KEYINPUT18), .B(G131), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n390), .A2(G214), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n288), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n390), .A2(G143), .A3(G214), .ZN(new_n524));
  NAND2_X1  g338(.A1(KEYINPUT18), .A2(G131), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n523), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(new_n240), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n239), .A2(new_n228), .ZN(new_n528));
  OAI211_X1 g342(.A(new_n521), .B(new_n526), .C1(new_n527), .C2(new_n528), .ZN(new_n529));
  OAI21_X1  g343(.A(G131), .B1(new_n519), .B2(new_n520), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n523), .A2(new_n337), .A3(new_n524), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  NOR2_X1   g346(.A1(new_n532), .A2(KEYINPUT17), .ZN(new_n533));
  INV_X1    g347(.A(KEYINPUT17), .ZN(new_n534));
  OAI211_X1 g348(.A(new_n229), .B(new_n230), .C1(new_n530), .C2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n518), .B(new_n529), .C1(new_n533), .C2(new_n535), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n239), .A2(KEYINPUT91), .A3(KEYINPUT19), .ZN(new_n538));
  INV_X1    g352(.A(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT19), .B1(new_n239), .B2(KEYINPUT91), .ZN(new_n540));
  OAI21_X1  g354(.A(new_n228), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n541), .A2(new_n230), .A3(new_n532), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n518), .B1(new_n542), .B2(new_n529), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n516), .B1(new_n537), .B2(new_n543), .ZN(new_n544));
  XNOR2_X1  g358(.A(KEYINPUT90), .B(KEYINPUT20), .ZN(new_n545));
  INV_X1    g359(.A(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n544), .A2(KEYINPUT92), .A3(new_n546), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n548));
  INV_X1    g362(.A(new_n516), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n532), .A2(new_n230), .ZN(new_n550));
  INV_X1    g364(.A(new_n540), .ZN(new_n551));
  AOI21_X1  g365(.A(G146), .B1(new_n551), .B2(new_n538), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n529), .B1(new_n550), .B2(new_n552), .ZN(new_n553));
  INV_X1    g367(.A(new_n518), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n549), .B1(new_n555), .B2(new_n536), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n548), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT20), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n547), .A2(new_n557), .A3(new_n559), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT94), .ZN(new_n561));
  OAI21_X1  g375(.A(new_n529), .B1(new_n533), .B2(new_n535), .ZN(new_n562));
  AND2_X1   g376(.A1(new_n562), .A2(new_n554), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n252), .B1(new_n563), .B2(new_n537), .ZN(new_n564));
  XOR2_X1   g378(.A(KEYINPUT93), .B(G475), .Z(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  AND3_X1   g380(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n561), .B1(new_n560), .B2(new_n566), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n288), .A2(G128), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n197), .A2(G143), .ZN(new_n571));
  AND2_X1   g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g386(.A(new_n572), .B(new_n325), .ZN(new_n573));
  XNOR2_X1  g387(.A(G116), .B(G122), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n574), .A2(new_n275), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n375), .A2(KEYINPUT14), .A3(G122), .ZN(new_n576));
  XOR2_X1   g390(.A(G116), .B(G122), .Z(new_n577));
  OAI211_X1 g391(.A(G107), .B(new_n576), .C1(new_n577), .C2(KEYINPUT14), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n573), .A2(new_n575), .A3(new_n578), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n577), .A2(G107), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n580), .A2(new_n575), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n572), .A2(new_n325), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n288), .A2(KEYINPUT13), .A3(G128), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n583), .A2(KEYINPUT95), .A3(new_n571), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT13), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n584), .B1(new_n585), .B2(new_n570), .ZN(new_n586));
  OAI21_X1  g400(.A(G134), .B1(new_n583), .B2(KEYINPUT95), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n581), .B(new_n582), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n579), .A2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(G217), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n267), .A2(new_n590), .A3(G953), .ZN(new_n591));
  XOR2_X1   g405(.A(new_n589), .B(new_n591), .Z(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n252), .ZN(new_n593));
  INV_X1    g407(.A(G478), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n594), .A2(KEYINPUT15), .ZN(new_n595));
  XOR2_X1   g409(.A(new_n593), .B(new_n595), .Z(new_n596));
  INV_X1    g410(.A(G952), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(G953), .ZN(new_n598));
  INV_X1    g412(.A(G237), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n598), .B1(new_n187), .B2(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(new_n600), .ZN(new_n601));
  OAI211_X1 g415(.A(G902), .B(G953), .C1(new_n187), .C2(new_n599), .ZN(new_n602));
  XNOR2_X1  g416(.A(new_n602), .B(KEYINPUT96), .ZN(new_n603));
  XNOR2_X1  g417(.A(KEYINPUT21), .B(G898), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n569), .A2(new_n596), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND4_X1  g422(.A1(new_n373), .A2(new_n454), .A3(new_n515), .A4(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(G101), .ZN(G3));
  AND3_X1   g424(.A1(new_n512), .A2(new_n513), .A3(new_n457), .ZN(new_n611));
  AOI21_X1  g425(.A(new_n457), .B1(new_n512), .B2(new_n513), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n455), .B(new_n606), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n594), .A2(new_n252), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n593), .B2(G478), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT33), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n592), .B(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n616), .B1(G478), .B2(new_n618), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n619), .B1(new_n567), .B2(new_n568), .ZN(new_n620));
  NOR2_X1   g434(.A1(new_n613), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n449), .A2(new_n252), .ZN(new_n622));
  AOI22_X1  g436(.A1(new_n622), .A2(G472), .B1(new_n451), .B2(new_n449), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n621), .A2(new_n373), .A3(new_n623), .ZN(new_n624));
  XOR2_X1   g438(.A(new_n624), .B(KEYINPUT97), .Z(new_n625));
  XNOR2_X1  g439(.A(KEYINPUT34), .B(G104), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n625), .B(new_n626), .ZN(G6));
  XNOR2_X1  g441(.A(new_n593), .B(new_n595), .ZN(new_n628));
  OAI211_X1 g442(.A(new_n547), .B(new_n557), .C1(new_n546), .C2(new_n544), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n628), .A2(new_n566), .A3(new_n629), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n613), .A2(new_n630), .ZN(new_n631));
  NAND3_X1  g445(.A1(new_n631), .A2(new_n373), .A3(new_n623), .ZN(new_n632));
  XOR2_X1   g446(.A(KEYINPUT35), .B(G107), .Z(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NAND2_X1  g448(.A1(new_n372), .A2(new_n370), .ZN(new_n635));
  AND3_X1   g449(.A1(new_n635), .A2(new_n515), .A3(new_n623), .ZN(new_n636));
  INV_X1    g450(.A(new_n189), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n256), .A2(new_n257), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(KEYINPUT25), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n256), .A2(new_n257), .A3(new_n258), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n637), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n253), .A2(KEYINPUT36), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n254), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n643), .A2(new_n263), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g459(.A(KEYINPUT98), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT98), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n261), .A2(new_n647), .A3(new_n644), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n607), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n636), .A2(new_n649), .ZN(new_n650));
  XNOR2_X1  g464(.A(KEYINPUT37), .B(G110), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT99), .ZN(new_n652));
  XNOR2_X1  g466(.A(new_n650), .B(new_n652), .ZN(G12));
  OAI21_X1  g467(.A(new_n455), .B1(new_n611), .B2(new_n612), .ZN(new_n654));
  NAND2_X1  g468(.A1(new_n449), .A2(new_n451), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n655), .A2(KEYINPUT32), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n416), .A2(new_n252), .ZN(new_n659));
  NAND3_X1  g473(.A1(new_n428), .A2(new_n438), .A3(new_n395), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n444), .A2(new_n388), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n426), .B1(new_n661), .B2(new_n427), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n659), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(G472), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n654), .B1(new_n658), .B2(new_n664), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n646), .A2(new_n648), .B1(new_n370), .B2(new_n372), .ZN(new_n666));
  AND2_X1   g480(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XOR2_X1   g481(.A(KEYINPUT100), .B(G900), .Z(new_n668));
  NAND2_X1  g482(.A1(new_n603), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(new_n600), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n630), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n667), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G128), .ZN(G30));
  NOR2_X1   g488(.A1(new_n611), .A2(new_n612), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(KEYINPUT38), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n437), .A2(new_n427), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n414), .A2(new_n394), .ZN(new_n678));
  NAND3_X1  g492(.A1(new_n677), .A2(new_n252), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g493(.A1(new_n679), .A2(G472), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n658), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n670), .B(KEYINPUT39), .ZN(new_n682));
  AND2_X1   g496(.A1(new_n635), .A2(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(KEYINPUT40), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n681), .B1(new_n683), .B2(new_n684), .ZN(new_n685));
  AOI211_X1 g499(.A(new_n676), .B(new_n685), .C1(new_n684), .C2(new_n683), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n646), .A2(new_n648), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n560), .A2(new_n566), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(KEYINPUT94), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n560), .A2(new_n561), .A3(new_n566), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n596), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  INV_X1    g505(.A(new_n691), .ZN(new_n692));
  NOR3_X1   g506(.A1(new_n687), .A2(new_n456), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(KEYINPUT101), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n686), .A2(new_n694), .ZN(new_n695));
  XNOR2_X1  g509(.A(new_n695), .B(G143), .ZN(G45));
  OAI211_X1 g510(.A(new_n619), .B(new_n670), .C1(new_n567), .C2(new_n568), .ZN(new_n697));
  INV_X1    g511(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n667), .A2(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G146), .ZN(G48));
  AOI21_X1  g514(.A(new_n265), .B1(new_n658), .B2(new_n664), .ZN(new_n701));
  INV_X1    g515(.A(new_n269), .ZN(new_n702));
  AOI21_X1  g516(.A(G902), .B1(new_n367), .B2(new_n368), .ZN(new_n703));
  INV_X1    g517(.A(G469), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT102), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n705), .A2(new_n369), .A3(new_n706), .ZN(new_n707));
  NOR3_X1   g521(.A1(new_n703), .A2(KEYINPUT102), .A3(new_n704), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n702), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n701), .A2(new_n621), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(KEYINPUT41), .B(G113), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n711), .B(new_n712), .ZN(G15));
  NAND3_X1  g527(.A1(new_n701), .A2(new_n631), .A3(new_n710), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(G116), .ZN(G18));
  NOR2_X1   g529(.A1(new_n654), .A2(new_n709), .ZN(new_n716));
  NAND4_X1  g530(.A1(new_n716), .A2(new_n687), .A3(new_n454), .A4(new_n608), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G119), .ZN(G21));
  INV_X1    g532(.A(new_n451), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n404), .A2(new_n380), .ZN(new_n720));
  AOI21_X1  g534(.A(new_n415), .B1(new_n720), .B2(new_n418), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT103), .B1(new_n721), .B2(new_n388), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT103), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n723), .B(new_n389), .C1(new_n414), .C2(new_n415), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n722), .A2(new_n394), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n436), .A2(new_n446), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT31), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n436), .A2(new_n446), .A3(KEYINPUT31), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  AOI21_X1  g544(.A(new_n719), .B1(new_n725), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g545(.A(G902), .B1(new_n730), .B2(new_n445), .ZN(new_n732));
  OAI21_X1  g546(.A(KEYINPUT104), .B1(new_n732), .B2(new_n443), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT104), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n622), .A2(new_n734), .A3(G472), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n731), .B1(new_n733), .B2(new_n735), .ZN(new_n736));
  INV_X1    g550(.A(new_n264), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n641), .A2(new_n737), .ZN(new_n738));
  AOI211_X1 g552(.A(new_n456), .B(new_n605), .C1(new_n508), .C2(new_n514), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n367), .A2(new_n368), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n740), .A2(new_n252), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(G469), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n706), .B1(new_n703), .B2(new_n704), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n708), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  AND3_X1   g560(.A1(new_n746), .A2(new_n691), .A3(new_n702), .ZN(new_n747));
  NAND4_X1  g561(.A1(new_n736), .A2(new_n738), .A3(new_n739), .A4(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(G122), .ZN(G24));
  NAND2_X1  g563(.A1(new_n716), .A2(new_n698), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT105), .ZN(new_n751));
  AND3_X1   g565(.A1(new_n261), .A2(new_n647), .A3(new_n644), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n647), .B1(new_n261), .B2(new_n644), .ZN(new_n753));
  NOR2_X1   g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g568(.A(new_n731), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n734), .B1(new_n622), .B2(G472), .ZN(new_n756));
  AOI211_X1 g570(.A(KEYINPUT104), .B(new_n443), .C1(new_n449), .C2(new_n252), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n755), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n751), .B1(new_n754), .B2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n736), .A2(new_n687), .A3(KEYINPUT105), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n750), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n761), .B(new_n219), .ZN(G27));
  INV_X1    g576(.A(KEYINPUT42), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n452), .A2(new_n453), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n441), .A2(new_n395), .A3(new_n428), .A4(new_n438), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n443), .B1(new_n765), .B2(new_n659), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n738), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NOR3_X1   g581(.A1(new_n611), .A2(new_n612), .A3(new_n456), .ZN(new_n768));
  AND2_X1   g582(.A1(new_n341), .A2(new_n360), .ZN(new_n769));
  AOI22_X1  g583(.A1(new_n359), .A2(new_n769), .B1(new_n352), .B2(new_n356), .ZN(new_n770));
  OAI21_X1  g584(.A(G469), .B1(new_n770), .B2(G902), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n740), .A2(new_n704), .A3(new_n252), .ZN(new_n772));
  AOI21_X1  g586(.A(new_n269), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g587(.A1(new_n768), .A2(new_n698), .A3(new_n773), .ZN(new_n774));
  OAI21_X1  g588(.A(new_n763), .B1(new_n767), .B2(new_n774), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n508), .A2(new_n455), .A3(new_n514), .ZN(new_n776));
  INV_X1    g590(.A(new_n773), .ZN(new_n777));
  NOR3_X1   g591(.A1(new_n776), .A2(new_n697), .A3(new_n777), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n701), .A2(new_n778), .A3(KEYINPUT42), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n775), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G131), .ZN(G33));
  AND4_X1   g595(.A1(new_n455), .A2(new_n508), .A3(new_n514), .A4(new_n773), .ZN(new_n782));
  NAND4_X1  g596(.A1(new_n454), .A2(new_n782), .A3(new_n738), .A4(new_n672), .ZN(new_n783));
  NAND2_X1  g597(.A1(new_n783), .A2(KEYINPUT106), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT106), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n701), .A2(new_n785), .A3(new_n672), .A4(new_n782), .ZN(new_n786));
  NAND2_X1  g600(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND2_X1  g602(.A1(new_n357), .A2(new_n361), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT45), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n704), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT107), .ZN(new_n792));
  OR2_X1    g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n792), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n795));
  NAND3_X1  g609(.A1(new_n793), .A2(new_n794), .A3(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n796), .A2(new_n363), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT46), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n369), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(KEYINPUT46), .A3(new_n363), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n269), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n776), .B(KEYINPUT111), .ZN(new_n802));
  NAND3_X1  g616(.A1(new_n801), .A2(new_n682), .A3(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(KEYINPUT44), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n689), .A2(new_n690), .ZN(new_n805));
  INV_X1    g619(.A(new_n619), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT43), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(KEYINPUT43), .ZN(new_n808));
  NAND3_X1  g622(.A1(new_n569), .A2(new_n808), .A3(new_n619), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g624(.A(new_n810), .B(KEYINPUT108), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT109), .ZN(new_n812));
  OAI21_X1  g626(.A(new_n812), .B1(new_n754), .B2(new_n623), .ZN(new_n813));
  INV_X1    g627(.A(new_n623), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n687), .A2(KEYINPUT109), .A3(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n811), .A2(new_n813), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n803), .B1(new_n804), .B2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n811), .A2(new_n813), .A3(KEYINPUT44), .A4(new_n815), .ZN(new_n818));
  INV_X1    g632(.A(KEYINPUT110), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n818), .A2(new_n819), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n817), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G137), .ZN(G39));
  NOR4_X1   g638(.A1(new_n454), .A2(new_n738), .A3(new_n697), .A4(new_n776), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n799), .A2(new_n800), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(KEYINPUT47), .A3(new_n702), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT47), .B1(new_n826), .B2(new_n702), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n825), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g643(.A(KEYINPUT112), .B(G140), .ZN(new_n830));
  XNOR2_X1  g644(.A(new_n829), .B(new_n830), .ZN(G42));
  NAND3_X1  g645(.A1(new_n738), .A2(new_n455), .A3(new_n270), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n832), .A2(new_n805), .A3(new_n806), .ZN(new_n833));
  INV_X1    g647(.A(new_n681), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n746), .B(KEYINPUT49), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n833), .A2(new_n834), .A3(new_n676), .A4(new_n835), .ZN(new_n836));
  NAND4_X1  g650(.A1(new_n596), .A2(new_n566), .A3(new_n629), .A4(new_n670), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n837), .B(new_n776), .C1(new_n658), .C2(new_n664), .ZN(new_n838));
  AOI22_X1  g652(.A1(new_n775), .A2(new_n779), .B1(new_n838), .B2(new_n666), .ZN(new_n839));
  AND3_X1   g653(.A1(new_n736), .A2(KEYINPUT105), .A3(new_n687), .ZN(new_n840));
  AOI21_X1  g654(.A(KEYINPUT105), .B1(new_n736), .B2(new_n687), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n778), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n839), .A2(new_n842), .A3(new_n787), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n714), .A2(new_n717), .ZN(new_n844));
  OAI211_X1 g658(.A(new_n738), .B(new_n755), .C1(new_n756), .C2(new_n757), .ZN(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n613), .A2(new_n709), .A3(new_n692), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n689), .A2(new_n690), .A3(new_n628), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n620), .A2(new_n848), .ZN(new_n849));
  AND4_X1   g663(.A1(new_n635), .A2(new_n738), .A3(new_n623), .A4(new_n849), .ZN(new_n850));
  AOI22_X1  g664(.A1(new_n846), .A2(new_n847), .B1(new_n850), .B2(new_n739), .ZN(new_n851));
  AND3_X1   g665(.A1(new_n608), .A2(new_n635), .A3(new_n738), .ZN(new_n852));
  AOI22_X1  g666(.A1(new_n852), .A2(new_n665), .B1(new_n636), .B2(new_n649), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n844), .A2(new_n711), .A3(new_n851), .A4(new_n853), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  INV_X1    g669(.A(new_n750), .ZN(new_n856));
  OAI21_X1  g670(.A(new_n856), .B1(new_n840), .B2(new_n841), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT52), .ZN(new_n858));
  OAI211_X1 g672(.A(new_n665), .B(new_n666), .C1(new_n672), .C2(new_n698), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n515), .A2(new_n691), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NOR4_X1   g675(.A1(new_n777), .A2(new_n641), .A3(new_n645), .A4(new_n671), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n861), .A2(new_n681), .A3(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n857), .A2(new_n858), .A3(new_n859), .A4(new_n863), .ZN(new_n864));
  XOR2_X1   g678(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n859), .A2(new_n863), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n866), .B1(new_n761), .B2(new_n867), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n864), .A4(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT53), .ZN(new_n870));
  OAI21_X1  g684(.A(KEYINPUT52), .B1(new_n761), .B2(new_n867), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n871), .A2(new_n864), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n373), .A2(new_n623), .A3(new_n739), .A4(new_n849), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n714), .A2(new_n717), .A3(new_n748), .A4(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n650), .A2(new_n711), .A3(new_n609), .ZN(new_n875));
  NOR2_X1   g689(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n759), .A2(new_n760), .ZN(new_n877));
  AOI22_X1  g691(.A1(new_n877), .A2(new_n778), .B1(new_n786), .B2(new_n784), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n876), .A2(new_n878), .A3(new_n839), .ZN(new_n879));
  OAI21_X1  g693(.A(new_n870), .B1(new_n872), .B2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT54), .ZN(new_n881));
  AND3_X1   g695(.A1(new_n869), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  NAND4_X1  g697(.A1(new_n855), .A2(KEYINPUT53), .A3(new_n864), .A4(new_n871), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n868), .A2(new_n864), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n885), .A2(new_n879), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n884), .B1(new_n886), .B2(KEYINPUT53), .ZN(new_n887));
  INV_X1    g701(.A(KEYINPUT114), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n887), .A2(new_n888), .A3(KEYINPUT54), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n883), .A2(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n887), .B2(KEYINPUT54), .ZN(new_n891));
  NOR3_X1   g705(.A1(new_n845), .A2(new_n810), .A3(new_n600), .ZN(new_n892));
  OR2_X1    g706(.A1(new_n827), .A2(new_n828), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n746), .A2(KEYINPUT115), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n270), .ZN(new_n896));
  OAI211_X1 g710(.A(new_n802), .B(new_n892), .C1(new_n893), .C2(new_n896), .ZN(new_n897));
  NAND3_X1  g711(.A1(new_n710), .A2(KEYINPUT116), .A3(new_n456), .ZN(new_n898));
  INV_X1    g712(.A(KEYINPUT116), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n899), .B1(new_n709), .B2(new_n455), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n892), .A2(new_n676), .A3(new_n898), .A4(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT50), .ZN(new_n902));
  OR3_X1    g716(.A1(new_n901), .A2(KEYINPUT118), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n901), .A2(new_n902), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT117), .ZN(new_n905));
  OAI21_X1  g719(.A(KEYINPUT118), .B1(new_n901), .B2(new_n902), .ZN(new_n906));
  INV_X1    g720(.A(KEYINPUT117), .ZN(new_n907));
  NAND3_X1  g721(.A1(new_n901), .A2(new_n907), .A3(new_n902), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n903), .A2(new_n905), .A3(new_n906), .A4(new_n908), .ZN(new_n909));
  NOR3_X1   g723(.A1(new_n681), .A2(new_n600), .A3(new_n265), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n910), .A2(new_n710), .A3(new_n768), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n911), .A2(new_n805), .A3(new_n619), .ZN(new_n912));
  NOR4_X1   g726(.A1(new_n810), .A2(new_n600), .A3(new_n709), .A4(new_n776), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n877), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n897), .A2(new_n909), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT51), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g731(.A1(new_n897), .A2(new_n909), .A3(KEYINPUT51), .A4(new_n914), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n598), .B1(new_n911), .B2(new_n620), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n913), .A2(new_n701), .ZN(new_n920));
  XOR2_X1   g734(.A(new_n920), .B(KEYINPUT48), .Z(new_n921));
  AOI211_X1 g735(.A(new_n919), .B(new_n921), .C1(new_n716), .C2(new_n892), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n917), .A2(new_n918), .A3(new_n922), .ZN(new_n923));
  NOR3_X1   g737(.A1(new_n890), .A2(new_n891), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n597), .A2(new_n191), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n925), .B(KEYINPUT119), .ZN(new_n926));
  OAI21_X1  g740(.A(new_n836), .B1(new_n924), .B2(new_n926), .ZN(G75));
  NOR2_X1   g741(.A1(new_n191), .A2(G952), .ZN(new_n928));
  INV_X1    g742(.A(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n252), .B1(new_n869), .B2(new_n880), .ZN(new_n930));
  AOI21_X1  g744(.A(KEYINPUT56), .B1(new_n930), .B2(G210), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n509), .A2(new_n510), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n932), .A2(new_n468), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n933), .A2(new_n512), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(KEYINPUT55), .ZN(new_n935));
  INV_X1    g749(.A(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n929), .B1(new_n931), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n937), .B1(new_n931), .B2(new_n936), .ZN(G51));
  XOR2_X1   g752(.A(new_n363), .B(KEYINPUT57), .Z(new_n939));
  AOI21_X1  g753(.A(new_n881), .B1(new_n869), .B2(new_n880), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n939), .B1(new_n882), .B2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(KEYINPUT120), .ZN(new_n942));
  NAND2_X1  g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT120), .B(new_n939), .C1(new_n882), .C2(new_n940), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n943), .A2(new_n740), .A3(new_n944), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n796), .B(KEYINPUT121), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n930), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n928), .B1(new_n945), .B2(new_n947), .ZN(G54));
  NOR2_X1   g762(.A1(new_n537), .A2(new_n543), .ZN(new_n949));
  INV_X1    g763(.A(new_n930), .ZN(new_n950));
  NAND2_X1  g764(.A1(KEYINPUT58), .A2(G475), .ZN(new_n951));
  OAI21_X1  g765(.A(new_n949), .B1(new_n950), .B2(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n929), .ZN(new_n953));
  NOR3_X1   g767(.A1(new_n950), .A2(new_n949), .A3(new_n951), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n953), .A2(new_n954), .ZN(G60));
  XNOR2_X1  g769(.A(new_n592), .B(KEYINPUT33), .ZN(new_n956));
  XOR2_X1   g770(.A(new_n614), .B(KEYINPUT59), .Z(new_n957));
  OAI211_X1 g771(.A(new_n956), .B(new_n957), .C1(new_n882), .C2(new_n940), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(new_n929), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n957), .B1(new_n890), .B2(new_n891), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n959), .B1(new_n960), .B2(new_n618), .ZN(G63));
  NAND2_X1  g775(.A1(G217), .A2(G902), .ZN(new_n962));
  XNOR2_X1  g776(.A(new_n962), .B(KEYINPUT60), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n963), .B1(new_n869), .B2(new_n880), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n964), .A2(new_n643), .ZN(new_n965));
  OAI211_X1 g779(.A(new_n965), .B(new_n929), .C1(new_n262), .C2(new_n964), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT122), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n965), .A2(new_n967), .A3(new_n929), .ZN(new_n968));
  NAND3_X1  g782(.A1(new_n966), .A2(KEYINPUT61), .A3(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n928), .B1(new_n964), .B2(new_n643), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT61), .ZN(new_n971));
  OAI221_X1 g785(.A(new_n970), .B1(new_n967), .B2(new_n971), .C1(new_n262), .C2(new_n964), .ZN(new_n972));
  AND2_X1   g786(.A1(new_n969), .A2(new_n972), .ZN(G66));
  INV_X1    g787(.A(G224), .ZN(new_n974));
  OAI21_X1  g788(.A(G953), .B1(new_n604), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n876), .B2(G953), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n932), .B1(G898), .B2(new_n191), .ZN(new_n977));
  XNOR2_X1  g791(.A(new_n976), .B(new_n977), .ZN(G69));
  NAND2_X1  g792(.A1(new_n434), .A2(new_n435), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n551), .A2(new_n538), .ZN(new_n980));
  XNOR2_X1  g794(.A(new_n980), .B(KEYINPUT123), .ZN(new_n981));
  XNOR2_X1  g795(.A(new_n981), .B(KEYINPUT124), .ZN(new_n982));
  XNOR2_X1  g796(.A(new_n979), .B(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n823), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n857), .A2(new_n859), .ZN(new_n986));
  NAND4_X1  g800(.A1(new_n801), .A2(new_n682), .A3(new_n701), .A4(new_n861), .ZN(new_n987));
  AND2_X1   g801(.A1(new_n787), .A2(new_n780), .ZN(new_n988));
  NAND4_X1  g802(.A1(new_n829), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n191), .B1(new_n985), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n191), .A2(G900), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(KEYINPUT125), .B1(new_n990), .B2(new_n992), .ZN(new_n993));
  AND4_X1   g807(.A1(new_n829), .A2(new_n986), .A3(new_n987), .A4(new_n988), .ZN(new_n994));
  AOI21_X1  g808(.A(G953), .B1(new_n994), .B2(new_n823), .ZN(new_n995));
  INV_X1    g809(.A(KEYINPUT125), .ZN(new_n996));
  NOR3_X1   g810(.A1(new_n995), .A2(new_n996), .A3(new_n991), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n984), .B1(new_n993), .B2(new_n997), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n695), .A2(new_n986), .ZN(new_n999));
  INV_X1    g813(.A(KEYINPUT62), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(new_n1001));
  NAND4_X1  g815(.A1(new_n701), .A2(new_n683), .A3(new_n768), .A4(new_n849), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n823), .A2(new_n829), .A3(new_n1002), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1001), .A2(new_n1003), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n984), .A2(G953), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n991), .B1(new_n354), .B2(G953), .ZN(new_n1007));
  XNOR2_X1  g821(.A(new_n1007), .B(KEYINPUT126), .ZN(new_n1008));
  NAND3_X1  g822(.A1(new_n998), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g823(.A(new_n1008), .ZN(new_n1010));
  NAND3_X1  g824(.A1(new_n990), .A2(KEYINPUT125), .A3(new_n992), .ZN(new_n1011));
  OAI21_X1  g825(.A(new_n996), .B1(new_n995), .B2(new_n991), .ZN(new_n1012));
  AOI21_X1  g826(.A(new_n983), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  AOI211_X1 g827(.A(G953), .B(new_n984), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1010), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n1009), .A2(new_n1015), .ZN(G72));
  NAND3_X1  g830(.A1(new_n1001), .A2(new_n876), .A3(new_n1003), .ZN(new_n1017));
  NAND2_X1  g831(.A1(G472), .A2(G902), .ZN(new_n1018));
  XOR2_X1   g832(.A(new_n1018), .B(KEYINPUT63), .Z(new_n1019));
  AOI21_X1  g833(.A(new_n677), .B1(new_n1017), .B2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g834(.A1(new_n994), .A2(new_n823), .A3(new_n876), .ZN(new_n1021));
  AOI211_X1 g835(.A(new_n427), .B(new_n437), .C1(new_n1021), .C2(new_n1019), .ZN(new_n1022));
  AOI22_X1  g836(.A1(new_n438), .A2(KEYINPUT127), .B1(new_n436), .B2(new_n446), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1023), .B1(KEYINPUT127), .B2(new_n438), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n887), .A2(new_n1019), .A3(new_n1024), .ZN(new_n1025));
  NOR4_X1   g839(.A1(new_n1020), .A2(new_n1022), .A3(new_n1025), .A4(new_n928), .ZN(G57));
endmodule


