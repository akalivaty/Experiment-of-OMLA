

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724;

  NOR2_X1 U366 ( .A1(G902), .A2(n679), .ZN(n484) );
  XNOR2_X1 U367 ( .A(n524), .B(KEYINPUT106), .ZN(n720) );
  AND2_X4 U368 ( .A1(n379), .A2(n411), .ZN(n687) );
  NOR2_X1 U369 ( .A1(n541), .A2(n525), .ZN(n526) );
  XNOR2_X2 U370 ( .A(n707), .B(G146), .ZN(n457) );
  NOR2_X1 U371 ( .A1(n722), .A2(n719), .ZN(n365) );
  INV_X1 U372 ( .A(n639), .ZN(n568) );
  AND2_X4 U373 ( .A1(n529), .A2(n528), .ZN(n530) );
  INV_X4 U374 ( .A(G143), .ZN(n419) );
  INV_X2 U375 ( .A(G125), .ZN(n378) );
  AND2_X1 U376 ( .A1(n533), .A2(n532), .ZN(n534) );
  AND2_X1 U377 ( .A1(n586), .A2(n587), .ZN(n361) );
  XNOR2_X1 U378 ( .A(n365), .B(n364), .ZN(n519) );
  NOR2_X1 U379 ( .A1(n514), .A2(n581), .ZN(n515) );
  NOR2_X1 U380 ( .A1(n640), .A2(n581), .ZN(n582) );
  NOR2_X1 U381 ( .A1(n654), .A2(n525), .ZN(n499) );
  AND2_X1 U382 ( .A1(n504), .A2(n503), .ZN(n520) );
  XNOR2_X1 U383 ( .A(n403), .B(KEYINPUT15), .ZN(n597) );
  XNOR2_X1 U384 ( .A(G137), .B(G140), .ZN(n438) );
  XOR2_X2 U385 ( .A(G116), .B(G107), .Z(n486) );
  XNOR2_X2 U386 ( .A(n466), .B(n410), .ZN(n707) );
  AND2_X1 U387 ( .A1(n613), .A2(n389), .ZN(n386) );
  XNOR2_X1 U388 ( .A(n402), .B(KEYINPUT20), .ZN(n448) );
  NAND2_X1 U389 ( .A1(n597), .A2(G234), .ZN(n402) );
  XNOR2_X1 U390 ( .A(n421), .B(G134), .ZN(n410) );
  XOR2_X1 U391 ( .A(G116), .B(G137), .Z(n455) );
  XNOR2_X1 U392 ( .A(KEYINPUT92), .B(KEYINPUT5), .ZN(n454) );
  NAND2_X1 U393 ( .A1(n353), .A2(n389), .ZN(n384) );
  AND2_X1 U394 ( .A1(n633), .A2(n380), .ZN(n451) );
  NOR2_X1 U395 ( .A1(n501), .A2(n381), .ZN(n380) );
  NOR2_X1 U396 ( .A1(G953), .A2(G237), .ZN(n474) );
  XNOR2_X1 U397 ( .A(KEYINPUT67), .B(G131), .ZN(n421) );
  XNOR2_X1 U398 ( .A(n357), .B(G104), .ZN(n479) );
  INV_X1 U399 ( .A(G122), .ZN(n357) );
  XNOR2_X1 U400 ( .A(n367), .B(n350), .ZN(n504) );
  XNOR2_X1 U401 ( .A(n498), .B(KEYINPUT87), .ZN(n525) );
  NOR2_X1 U402 ( .A1(G902), .A2(n598), .ZN(n459) );
  XNOR2_X1 U403 ( .A(n453), .B(n452), .ZN(n462) );
  XNOR2_X1 U404 ( .A(G119), .B(KEYINPUT3), .ZN(n452) );
  XOR2_X1 U405 ( .A(G101), .B(G113), .Z(n453) );
  XNOR2_X1 U406 ( .A(n486), .B(n479), .ZN(n359) );
  XNOR2_X1 U407 ( .A(n449), .B(n450), .ZN(n400) );
  NAND2_X1 U408 ( .A1(n648), .A2(n551), .ZN(n416) );
  NOR2_X1 U409 ( .A1(n629), .A2(n583), .ZN(n571) );
  INV_X1 U410 ( .A(n569), .ZN(n580) );
  INV_X2 U411 ( .A(G953), .ZN(n711) );
  INV_X1 U412 ( .A(n597), .ZN(n411) );
  XNOR2_X1 U413 ( .A(n457), .B(n427), .ZN(n675) );
  INV_X1 U414 ( .A(KEYINPUT46), .ZN(n364) );
  INV_X1 U415 ( .A(KEYINPUT64), .ZN(n391) );
  NAND2_X1 U416 ( .A1(n390), .A2(KEYINPUT64), .ZN(n389) );
  INV_X1 U417 ( .A(KEYINPUT44), .ZN(n390) );
  NAND2_X1 U418 ( .A1(n511), .A2(n651), .ZN(n367) );
  INV_X1 U419 ( .A(KEYINPUT66), .ZN(n397) );
  XNOR2_X1 U420 ( .A(n457), .B(n366), .ZN(n598) );
  XNOR2_X1 U421 ( .A(n363), .B(n456), .ZN(n366) );
  XNOR2_X1 U422 ( .A(n462), .B(n347), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n383), .B(n382), .ZN(n490) );
  INV_X1 U424 ( .A(KEYINPUT8), .ZN(n382) );
  NAND2_X1 U425 ( .A1(n711), .A2(G234), .ZN(n383) );
  INV_X1 U426 ( .A(KEYINPUT4), .ZN(n420) );
  INV_X1 U427 ( .A(KEYINPUT76), .ZN(n463) );
  NAND2_X1 U428 ( .A1(G234), .A2(G237), .ZN(n430) );
  NAND2_X1 U429 ( .A1(n580), .A2(n579), .ZN(n640) );
  OR2_X1 U430 ( .A1(G237), .A2(G902), .ZN(n497) );
  XNOR2_X1 U431 ( .A(G128), .B(G119), .ZN(n440) );
  XNOR2_X1 U432 ( .A(G110), .B(KEYINPUT24), .ZN(n441) );
  XNOR2_X1 U433 ( .A(KEYINPUT86), .B(G902), .ZN(n403) );
  XOR2_X1 U434 ( .A(G122), .B(G134), .Z(n492) );
  XOR2_X1 U435 ( .A(KEYINPUT94), .B(G140), .Z(n478) );
  XNOR2_X1 U436 ( .A(G143), .B(G113), .ZN(n477) );
  XNOR2_X1 U437 ( .A(KEYINPUT93), .B(KEYINPUT12), .ZN(n472) );
  INV_X1 U438 ( .A(n421), .ZN(n480) );
  XNOR2_X1 U439 ( .A(n692), .B(n393), .ZN(n468) );
  INV_X1 U440 ( .A(KEYINPUT70), .ZN(n393) );
  NAND2_X1 U441 ( .A1(n404), .A2(n406), .ZN(n379) );
  XNOR2_X1 U442 ( .A(n507), .B(n506), .ZN(n544) );
  AND2_X1 U443 ( .A1(n520), .A2(n505), .ZN(n507) );
  XNOR2_X1 U444 ( .A(n526), .B(KEYINPUT19), .ZN(n556) );
  XNOR2_X1 U445 ( .A(n396), .B(n395), .ZN(n394) );
  INV_X1 U446 ( .A(KEYINPUT28), .ZN(n395) );
  XNOR2_X1 U447 ( .A(n362), .B(n413), .ZN(n693) );
  INV_X1 U448 ( .A(n462), .ZN(n413) );
  XNOR2_X1 U449 ( .A(n359), .B(n461), .ZN(n362) );
  XNOR2_X1 U450 ( .A(n543), .B(KEYINPUT103), .ZN(n718) );
  XNOR2_X1 U451 ( .A(n508), .B(n401), .ZN(n719) );
  XNOR2_X1 U452 ( .A(KEYINPUT108), .B(KEYINPUT40), .ZN(n401) );
  AND2_X1 U453 ( .A1(n544), .A2(n530), .ZN(n508) );
  AND2_X1 U454 ( .A1(n376), .A2(n375), .ZN(n624) );
  INV_X1 U455 ( .A(n549), .ZN(n375) );
  NAND2_X1 U456 ( .A1(n576), .A2(n560), .ZN(n561) );
  NAND2_X1 U457 ( .A1(n360), .A2(n346), .ZN(n524) );
  XNOR2_X1 U458 ( .A(n522), .B(KEYINPUT105), .ZN(n360) );
  XNOR2_X1 U459 ( .A(n372), .B(KEYINPUT78), .ZN(n616) );
  NOR2_X1 U460 ( .A1(n527), .A2(n556), .ZN(n372) );
  NAND2_X1 U461 ( .A1(n565), .A2(n564), .ZN(n613) );
  AND2_X1 U462 ( .A1(n374), .A2(n639), .ZN(n609) );
  XNOR2_X1 U463 ( .A(n567), .B(KEYINPUT91), .ZN(n374) );
  XNOR2_X1 U464 ( .A(n675), .B(n351), .ZN(n676) );
  INV_X1 U465 ( .A(KEYINPUT56), .ZN(n368) );
  XOR2_X1 U466 ( .A(n669), .B(n354), .Z(n344) );
  AND2_X1 U467 ( .A1(n723), .A2(n613), .ZN(n345) );
  AND2_X1 U468 ( .A1(n523), .A2(n529), .ZN(n346) );
  AND2_X1 U469 ( .A1(n474), .A2(G210), .ZN(n347) );
  XOR2_X1 U470 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n348) );
  AND2_X1 U471 ( .A1(n613), .A2(KEYINPUT64), .ZN(n349) );
  XOR2_X1 U472 ( .A(KEYINPUT104), .B(KEYINPUT30), .Z(n350) );
  XOR2_X1 U473 ( .A(n674), .B(n673), .Z(n351) );
  XOR2_X1 U474 ( .A(KEYINPUT77), .B(KEYINPUT35), .Z(n352) );
  NAND2_X1 U475 ( .A1(n391), .A2(KEYINPUT44), .ZN(n353) );
  XNOR2_X1 U476 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n354) );
  XNOR2_X1 U477 ( .A(KEYINPUT123), .B(KEYINPUT59), .ZN(n355) );
  XOR2_X1 U478 ( .A(KEYINPUT62), .B(KEYINPUT109), .Z(n356) );
  NAND2_X1 U479 ( .A1(n723), .A2(n386), .ZN(n385) );
  XNOR2_X2 U480 ( .A(n561), .B(KEYINPUT32), .ZN(n723) );
  XNOR2_X1 U481 ( .A(n509), .B(n510), .ZN(n569) );
  XNOR2_X1 U482 ( .A(n429), .B(n428), .ZN(n509) );
  AND2_X2 U483 ( .A1(n534), .A2(n535), .ZN(n536) );
  NAND2_X1 U484 ( .A1(n358), .A2(n720), .ZN(n370) );
  NAND2_X1 U485 ( .A1(n531), .A2(KEYINPUT47), .ZN(n358) );
  XNOR2_X1 U486 ( .A(n538), .B(n539), .ZN(n540) );
  NAND2_X1 U487 ( .A1(n588), .A2(n361), .ZN(n589) );
  NAND2_X1 U488 ( .A1(n520), .A2(n566), .ZN(n521) );
  XNOR2_X1 U489 ( .A(n483), .B(n482), .ZN(n679) );
  XOR2_X1 U490 ( .A(KEYINPUT11), .B(KEYINPUT95), .Z(n473) );
  XNOR2_X2 U491 ( .A(n511), .B(n512), .ZN(n559) );
  XNOR2_X2 U492 ( .A(n459), .B(n458), .ZN(n511) );
  XNOR2_X2 U493 ( .A(n596), .B(n548), .ZN(n709) );
  OR2_X2 U494 ( .A1(n541), .A2(n521), .ZN(n522) );
  NAND2_X1 U495 ( .A1(n405), .A2(KEYINPUT2), .ZN(n404) );
  NAND2_X1 U496 ( .A1(n700), .A2(n596), .ZN(n405) );
  XNOR2_X1 U497 ( .A(n369), .B(n368), .ZN(G51) );
  NAND2_X1 U498 ( .A1(n672), .A2(n671), .ZN(n369) );
  XNOR2_X1 U499 ( .A(n370), .B(KEYINPUT79), .ZN(n533) );
  XNOR2_X1 U500 ( .A(n371), .B(n605), .ZN(G57) );
  NOR2_X2 U501 ( .A1(n603), .A2(n691), .ZN(n371) );
  INV_X1 U502 ( .A(n551), .ZN(n381) );
  XNOR2_X1 U503 ( .A(n373), .B(KEYINPUT122), .ZN(G54) );
  NOR2_X2 U504 ( .A1(n678), .A2(n691), .ZN(n373) );
  XNOR2_X1 U505 ( .A(n518), .B(KEYINPUT36), .ZN(n376) );
  XNOR2_X2 U506 ( .A(n485), .B(n484), .ZN(n529) );
  XNOR2_X1 U507 ( .A(n377), .B(KEYINPUT60), .ZN(G60) );
  NOR2_X2 U508 ( .A1(n682), .A2(n691), .ZN(n377) );
  XNOR2_X1 U509 ( .A(n475), .B(n418), .ZN(n476) );
  XNOR2_X1 U510 ( .A(n705), .B(n476), .ZN(n483) );
  XNOR2_X2 U511 ( .A(n378), .B(G146), .ZN(n467) );
  NOR2_X1 U512 ( .A1(n379), .A2(n628), .ZN(n666) );
  INV_X1 U513 ( .A(n562), .ZN(n633) );
  XNOR2_X2 U514 ( .A(n399), .B(n400), .ZN(n562) );
  NAND2_X1 U515 ( .A1(n385), .A2(n384), .ZN(n388) );
  NAND2_X1 U516 ( .A1(n388), .A2(n387), .ZN(n588) );
  NAND2_X1 U517 ( .A1(n723), .A2(n349), .ZN(n387) );
  XNOR2_X1 U518 ( .A(n468), .B(n392), .ZN(n469) );
  XNOR2_X1 U519 ( .A(n467), .B(n348), .ZN(n392) );
  XNOR2_X2 U520 ( .A(KEYINPUT74), .B(G110), .ZN(n692) );
  OR2_X2 U521 ( .A1(n583), .A2(n416), .ZN(n415) );
  NAND2_X1 U522 ( .A1(n394), .A2(n460), .ZN(n527) );
  NAND2_X1 U523 ( .A1(n513), .A2(n568), .ZN(n396) );
  XNOR2_X1 U524 ( .A(n451), .B(KEYINPUT68), .ZN(n513) );
  XNOR2_X2 U525 ( .A(n398), .B(n397), .ZN(n579) );
  NAND2_X1 U526 ( .A1(n562), .A2(n551), .ZN(n398) );
  NOR2_X1 U527 ( .A1(n689), .A2(G902), .ZN(n399) );
  NAND2_X1 U528 ( .A1(n407), .A2(n700), .ZN(n406) );
  XNOR2_X2 U529 ( .A(n595), .B(KEYINPUT45), .ZN(n700) );
  NOR2_X1 U530 ( .A1(n709), .A2(KEYINPUT2), .ZN(n407) );
  NAND2_X1 U531 ( .A1(n590), .A2(KEYINPUT44), .ZN(n585) );
  XNOR2_X2 U532 ( .A(n408), .B(n352), .ZN(n590) );
  NAND2_X1 U533 ( .A1(n409), .A2(n346), .ZN(n408) );
  XNOR2_X1 U534 ( .A(n584), .B(KEYINPUT34), .ZN(n409) );
  XNOR2_X2 U535 ( .A(n487), .B(n420), .ZN(n466) );
  XNOR2_X2 U536 ( .A(n419), .B(G128), .ZN(n487) );
  XNOR2_X2 U537 ( .A(n412), .B(n471), .ZN(n541) );
  NAND2_X1 U538 ( .A1(n669), .A2(n597), .ZN(n412) );
  XNOR2_X1 U539 ( .A(n693), .B(n414), .ZN(n669) );
  XNOR2_X1 U540 ( .A(n470), .B(n469), .ZN(n414) );
  NOR2_X2 U541 ( .A1(n563), .A2(n559), .ZN(n576) );
  XNOR2_X2 U542 ( .A(n415), .B(KEYINPUT22), .ZN(n563) );
  XNOR2_X1 U543 ( .A(n670), .B(n344), .ZN(n672) );
  XNOR2_X1 U544 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U545 ( .A(n681), .B(n680), .ZN(n682) );
  BUF_X1 U546 ( .A(n627), .Z(n656) );
  XOR2_X2 U547 ( .A(KEYINPUT10), .B(n467), .Z(n705) );
  XOR2_X1 U548 ( .A(n478), .B(n477), .Z(n417) );
  AND2_X1 U549 ( .A1(G214), .A2(n474), .ZN(n418) );
  XNOR2_X1 U550 ( .A(n464), .B(n463), .ZN(n465) );
  XNOR2_X1 U551 ( .A(n466), .B(n465), .ZN(n470) );
  INV_X1 U552 ( .A(n501), .ZN(n502) );
  XNOR2_X1 U553 ( .A(n417), .B(n481), .ZN(n482) );
  XNOR2_X1 U554 ( .A(n598), .B(n356), .ZN(n600) );
  XNOR2_X1 U555 ( .A(n600), .B(n599), .ZN(n601) );
  XNOR2_X1 U556 ( .A(n602), .B(n601), .ZN(n603) );
  XNOR2_X1 U557 ( .A(n446), .B(n447), .ZN(n689) );
  XNOR2_X1 U558 ( .A(KEYINPUT98), .B(n530), .ZN(n618) );
  XNOR2_X1 U559 ( .A(n604), .B(KEYINPUT85), .ZN(n605) );
  NOR2_X1 U560 ( .A1(G952), .A2(n711), .ZN(n691) );
  XOR2_X1 U561 ( .A(G107), .B(G104), .Z(n423) );
  NAND2_X1 U562 ( .A1(G227), .A2(n711), .ZN(n422) );
  XNOR2_X1 U563 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U564 ( .A(KEYINPUT88), .B(n438), .ZN(n706) );
  XOR2_X1 U565 ( .A(n424), .B(n706), .Z(n426) );
  XOR2_X1 U566 ( .A(G101), .B(n468), .Z(n425) );
  XNOR2_X1 U567 ( .A(n426), .B(n425), .ZN(n427) );
  NOR2_X1 U568 ( .A1(G902), .A2(n675), .ZN(n429) );
  XNOR2_X1 U569 ( .A(KEYINPUT69), .B(G469), .ZN(n428) );
  BUF_X1 U570 ( .A(n509), .Z(n566) );
  XOR2_X1 U571 ( .A(n566), .B(KEYINPUT107), .Z(n460) );
  XOR2_X1 U572 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n431) );
  XNOR2_X1 U573 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U574 ( .A1(G952), .A2(n432), .ZN(n662) );
  NOR2_X1 U575 ( .A1(G953), .A2(n662), .ZN(n554) );
  NAND2_X1 U576 ( .A1(G902), .A2(n432), .ZN(n552) );
  NOR2_X1 U577 ( .A1(G900), .A2(n552), .ZN(n433) );
  NAND2_X1 U578 ( .A1(G953), .A2(n433), .ZN(n434) );
  XNOR2_X1 U579 ( .A(KEYINPUT99), .B(n434), .ZN(n435) );
  NOR2_X1 U580 ( .A1(n554), .A2(n435), .ZN(n501) );
  XOR2_X1 U581 ( .A(KEYINPUT90), .B(KEYINPUT21), .Z(n437) );
  NAND2_X1 U582 ( .A1(G221), .A2(n448), .ZN(n436) );
  XNOR2_X1 U583 ( .A(n437), .B(n436), .ZN(n551) );
  INV_X1 U584 ( .A(n438), .ZN(n439) );
  XNOR2_X1 U585 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U586 ( .A(KEYINPUT23), .B(KEYINPUT89), .Z(n442) );
  XNOR2_X1 U587 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U588 ( .A(n444), .B(n443), .Z(n447) );
  NAND2_X1 U589 ( .A1(G221), .A2(n490), .ZN(n445) );
  XNOR2_X1 U590 ( .A(n705), .B(n445), .ZN(n446) );
  XOR2_X1 U591 ( .A(KEYINPUT25), .B(KEYINPUT75), .Z(n450) );
  NAND2_X1 U592 ( .A1(G217), .A2(n448), .ZN(n449) );
  XNOR2_X1 U593 ( .A(n455), .B(n454), .ZN(n456) );
  XNOR2_X1 U594 ( .A(G472), .B(KEYINPUT71), .ZN(n458) );
  INV_X1 U595 ( .A(n511), .ZN(n639) );
  NAND2_X1 U596 ( .A1(n497), .A2(G210), .ZN(n471) );
  XOR2_X1 U597 ( .A(KEYINPUT72), .B(KEYINPUT16), .Z(n461) );
  NAND2_X1 U598 ( .A1(G224), .A2(n711), .ZN(n464) );
  XNOR2_X1 U599 ( .A(KEYINPUT38), .B(n541), .ZN(n646) );
  XNOR2_X1 U600 ( .A(KEYINPUT13), .B(G475), .ZN(n485) );
  XNOR2_X1 U601 ( .A(n473), .B(n472), .ZN(n475) );
  XNOR2_X1 U602 ( .A(n479), .B(n480), .ZN(n481) );
  XOR2_X1 U603 ( .A(KEYINPUT7), .B(KEYINPUT9), .Z(n489) );
  XNOR2_X1 U604 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U605 ( .A(n489), .B(n488), .ZN(n494) );
  NAND2_X1 U606 ( .A1(G217), .A2(n490), .ZN(n491) );
  XNOR2_X1 U607 ( .A(n492), .B(n491), .ZN(n493) );
  XNOR2_X1 U608 ( .A(n494), .B(n493), .ZN(n683) );
  NOR2_X1 U609 ( .A1(G902), .A2(n683), .ZN(n496) );
  XNOR2_X1 U610 ( .A(KEYINPUT96), .B(G478), .ZN(n495) );
  XNOR2_X1 U611 ( .A(n496), .B(n495), .ZN(n528) );
  INV_X1 U612 ( .A(n528), .ZN(n523) );
  NOR2_X1 U613 ( .A1(n529), .A2(n523), .ZN(n648) );
  NAND2_X1 U614 ( .A1(n646), .A2(n648), .ZN(n654) );
  NAND2_X1 U615 ( .A1(n497), .A2(G214), .ZN(n498) );
  XNOR2_X1 U616 ( .A(n499), .B(KEYINPUT41), .ZN(n645) );
  NOR2_X1 U617 ( .A1(n527), .A2(n645), .ZN(n500) );
  XNOR2_X1 U618 ( .A(KEYINPUT42), .B(n500), .ZN(n722) );
  INV_X1 U619 ( .A(n525), .ZN(n651) );
  AND2_X1 U620 ( .A1(n579), .A2(n502), .ZN(n503) );
  AND2_X1 U621 ( .A1(n646), .A2(n566), .ZN(n505) );
  INV_X1 U622 ( .A(KEYINPUT39), .ZN(n506) );
  INV_X1 U623 ( .A(KEYINPUT1), .ZN(n510) );
  INV_X1 U624 ( .A(n580), .ZN(n630) );
  XNOR2_X1 U625 ( .A(n630), .B(KEYINPUT84), .ZN(n549) );
  INV_X1 U626 ( .A(KEYINPUT6), .ZN(n512) );
  INV_X1 U627 ( .A(n559), .ZN(n581) );
  NAND2_X1 U628 ( .A1(n513), .A2(n618), .ZN(n514) );
  XOR2_X1 U629 ( .A(KEYINPUT100), .B(n515), .Z(n516) );
  NOR2_X1 U630 ( .A1(n525), .A2(n516), .ZN(n537) );
  INV_X1 U631 ( .A(n537), .ZN(n517) );
  NOR2_X1 U632 ( .A1(n517), .A2(n541), .ZN(n518) );
  NOR2_X1 U633 ( .A1(n519), .A2(n624), .ZN(n535) );
  NOR2_X1 U634 ( .A1(n529), .A2(n528), .ZN(n621) );
  NOR2_X1 U635 ( .A1(n530), .A2(n621), .ZN(n574) );
  INV_X1 U636 ( .A(n574), .ZN(n647) );
  NAND2_X1 U637 ( .A1(n616), .A2(n647), .ZN(n531) );
  OR2_X1 U638 ( .A1(KEYINPUT47), .A2(n531), .ZN(n532) );
  XNOR2_X1 U639 ( .A(n536), .B(KEYINPUT48), .ZN(n547) );
  XOR2_X1 U640 ( .A(KEYINPUT43), .B(KEYINPUT101), .Z(n539) );
  NAND2_X1 U641 ( .A1(n537), .A2(n630), .ZN(n538) );
  XNOR2_X1 U642 ( .A(KEYINPUT102), .B(n540), .ZN(n542) );
  NAND2_X1 U643 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U644 ( .A1(n544), .A2(n621), .ZN(n626) );
  INV_X1 U645 ( .A(n626), .ZN(n545) );
  NOR2_X1 U646 ( .A1(n718), .A2(n545), .ZN(n546) );
  AND2_X2 U647 ( .A1(n547), .A2(n546), .ZN(n596) );
  INV_X1 U648 ( .A(KEYINPUT80), .ZN(n548) );
  OR2_X1 U649 ( .A1(n562), .A2(n549), .ZN(n550) );
  XNOR2_X1 U650 ( .A(KEYINPUT97), .B(n550), .ZN(n560) );
  INV_X1 U651 ( .A(G898), .ZN(n698) );
  NAND2_X1 U652 ( .A1(G953), .A2(n698), .ZN(n694) );
  NOR2_X1 U653 ( .A1(n552), .A2(n694), .ZN(n553) );
  NOR2_X1 U654 ( .A1(n554), .A2(n553), .ZN(n555) );
  NOR2_X1 U655 ( .A1(n556), .A2(n555), .ZN(n558) );
  INV_X1 U656 ( .A(KEYINPUT0), .ZN(n557) );
  XNOR2_X1 U657 ( .A(n558), .B(n557), .ZN(n583) );
  NOR2_X1 U658 ( .A1(n563), .A2(n562), .ZN(n565) );
  NOR2_X1 U659 ( .A1(n568), .A2(n580), .ZN(n564) );
  INV_X1 U660 ( .A(n579), .ZN(n629) );
  NAND2_X1 U661 ( .A1(n566), .A2(n571), .ZN(n567) );
  NOR2_X1 U662 ( .A1(n639), .A2(n630), .ZN(n570) );
  NAND2_X1 U663 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U664 ( .A(KEYINPUT31), .B(n572), .ZN(n622) );
  NOR2_X1 U665 ( .A1(n609), .A2(n622), .ZN(n573) );
  NOR2_X1 U666 ( .A1(n574), .A2(n573), .ZN(n578) );
  NOR2_X1 U667 ( .A1(n633), .A2(n580), .ZN(n575) );
  NAND2_X1 U668 ( .A1(n576), .A2(n575), .ZN(n606) );
  INV_X1 U669 ( .A(n606), .ZN(n577) );
  NOR2_X1 U670 ( .A1(n578), .A2(n577), .ZN(n587) );
  XNOR2_X1 U671 ( .A(n582), .B(KEYINPUT33), .ZN(n627) );
  NOR2_X1 U672 ( .A1(n583), .A2(n627), .ZN(n584) );
  XNOR2_X1 U673 ( .A(n585), .B(KEYINPUT82), .ZN(n586) );
  XNOR2_X1 U674 ( .A(n589), .B(KEYINPUT81), .ZN(n594) );
  NOR2_X1 U675 ( .A1(n590), .A2(KEYINPUT44), .ZN(n591) );
  XOR2_X1 U676 ( .A(KEYINPUT65), .B(n591), .Z(n592) );
  NAND2_X1 U677 ( .A1(n592), .A2(n345), .ZN(n593) );
  NAND2_X1 U678 ( .A1(n594), .A2(n593), .ZN(n595) );
  NAND2_X1 U679 ( .A1(n687), .A2(G472), .ZN(n602) );
  XOR2_X1 U680 ( .A(KEYINPUT110), .B(KEYINPUT83), .Z(n599) );
  XOR2_X1 U681 ( .A(KEYINPUT63), .B(KEYINPUT111), .Z(n604) );
  XNOR2_X1 U682 ( .A(G101), .B(KEYINPUT112), .ZN(n607) );
  XNOR2_X1 U683 ( .A(n607), .B(n606), .ZN(G3) );
  NAND2_X1 U684 ( .A1(n618), .A2(n609), .ZN(n608) );
  XNOR2_X1 U685 ( .A(n608), .B(G104), .ZN(G6) );
  XOR2_X1 U686 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n611) );
  NAND2_X1 U687 ( .A1(n609), .A2(n621), .ZN(n610) );
  XNOR2_X1 U688 ( .A(n611), .B(n610), .ZN(n612) );
  XNOR2_X1 U689 ( .A(G107), .B(n612), .ZN(G9) );
  XNOR2_X1 U690 ( .A(G110), .B(n613), .ZN(G12) );
  XOR2_X1 U691 ( .A(G128), .B(KEYINPUT29), .Z(n615) );
  NAND2_X1 U692 ( .A1(n621), .A2(n616), .ZN(n614) );
  XNOR2_X1 U693 ( .A(n615), .B(n614), .ZN(G30) );
  NAND2_X1 U694 ( .A1(n616), .A2(n618), .ZN(n617) );
  XNOR2_X1 U695 ( .A(n617), .B(G146), .ZN(G48) );
  NAND2_X1 U696 ( .A1(n618), .A2(n622), .ZN(n619) );
  XNOR2_X1 U697 ( .A(n619), .B(KEYINPUT114), .ZN(n620) );
  XNOR2_X1 U698 ( .A(G113), .B(n620), .ZN(G15) );
  NAND2_X1 U699 ( .A1(n622), .A2(n621), .ZN(n623) );
  XNOR2_X1 U700 ( .A(n623), .B(G116), .ZN(G18) );
  XNOR2_X1 U701 ( .A(n624), .B(G125), .ZN(n625) );
  XNOR2_X1 U702 ( .A(n625), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U703 ( .A(G134), .B(n626), .ZN(G36) );
  NOR2_X1 U704 ( .A1(n645), .A2(n656), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n630), .A2(n629), .ZN(n631) );
  XNOR2_X1 U706 ( .A(n631), .B(KEYINPUT50), .ZN(n632) );
  NAND2_X1 U707 ( .A1(n632), .A2(n639), .ZN(n638) );
  XOR2_X1 U708 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n635) );
  NAND2_X1 U709 ( .A1(n633), .A2(n381), .ZN(n634) );
  XNOR2_X1 U710 ( .A(n635), .B(n634), .ZN(n636) );
  XNOR2_X1 U711 ( .A(n636), .B(KEYINPUT115), .ZN(n637) );
  NOR2_X1 U712 ( .A1(n638), .A2(n637), .ZN(n642) );
  NOR2_X1 U713 ( .A1(n640), .A2(n639), .ZN(n641) );
  NOR2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U715 ( .A(KEYINPUT51), .B(n643), .Z(n644) );
  NOR2_X1 U716 ( .A1(n645), .A2(n644), .ZN(n659) );
  NAND2_X1 U717 ( .A1(n647), .A2(n646), .ZN(n650) );
  INV_X1 U718 ( .A(n648), .ZN(n649) );
  NAND2_X1 U719 ( .A1(n650), .A2(n649), .ZN(n652) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n654), .A2(n653), .ZN(n655) );
  XNOR2_X1 U722 ( .A(KEYINPUT117), .B(n655), .ZN(n657) );
  NOR2_X1 U723 ( .A1(n657), .A2(n656), .ZN(n658) );
  NOR2_X1 U724 ( .A1(n659), .A2(n658), .ZN(n661) );
  XNOR2_X1 U725 ( .A(KEYINPUT52), .B(KEYINPUT118), .ZN(n660) );
  XNOR2_X1 U726 ( .A(n661), .B(n660), .ZN(n663) );
  NOR2_X1 U727 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U728 ( .A(n664), .B(KEYINPUT119), .ZN(n665) );
  NAND2_X1 U729 ( .A1(n666), .A2(n665), .ZN(n667) );
  NOR2_X1 U730 ( .A1(n667), .A2(G953), .ZN(n668) );
  XNOR2_X1 U731 ( .A(n668), .B(KEYINPUT53), .ZN(G75) );
  NAND2_X1 U732 ( .A1(n687), .A2(G210), .ZN(n670) );
  INV_X1 U733 ( .A(n691), .ZN(n671) );
  NAND2_X1 U734 ( .A1(n687), .A2(G469), .ZN(n677) );
  XOR2_X1 U735 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n674) );
  XNOR2_X1 U736 ( .A(KEYINPUT58), .B(KEYINPUT57), .ZN(n673) );
  NAND2_X1 U737 ( .A1(n687), .A2(G475), .ZN(n681) );
  XNOR2_X1 U738 ( .A(n679), .B(n355), .ZN(n680) );
  XNOR2_X1 U739 ( .A(n683), .B(KEYINPUT124), .ZN(n685) );
  NAND2_X1 U740 ( .A1(G478), .A2(n687), .ZN(n684) );
  XNOR2_X1 U741 ( .A(n685), .B(n684), .ZN(n686) );
  NOR2_X1 U742 ( .A1(n691), .A2(n686), .ZN(G63) );
  NAND2_X1 U743 ( .A1(G217), .A2(n687), .ZN(n688) );
  XNOR2_X1 U744 ( .A(n689), .B(n688), .ZN(n690) );
  NOR2_X1 U745 ( .A1(n691), .A2(n690), .ZN(G66) );
  XNOR2_X1 U746 ( .A(n693), .B(n692), .ZN(n695) );
  NAND2_X1 U747 ( .A1(n695), .A2(n694), .ZN(n704) );
  NAND2_X1 U748 ( .A1(G953), .A2(G224), .ZN(n696) );
  XOR2_X1 U749 ( .A(KEYINPUT61), .B(n696), .Z(n697) );
  NOR2_X1 U750 ( .A1(n698), .A2(n697), .ZN(n699) );
  XNOR2_X1 U751 ( .A(n699), .B(KEYINPUT125), .ZN(n702) );
  NAND2_X1 U752 ( .A1(n700), .A2(n711), .ZN(n701) );
  NAND2_X1 U753 ( .A1(n702), .A2(n701), .ZN(n703) );
  XOR2_X1 U754 ( .A(n704), .B(n703), .Z(G69) );
  XNOR2_X1 U755 ( .A(n706), .B(n705), .ZN(n708) );
  XNOR2_X1 U756 ( .A(n708), .B(n707), .ZN(n713) );
  XNOR2_X1 U757 ( .A(KEYINPUT126), .B(n713), .ZN(n710) );
  XNOR2_X1 U758 ( .A(n710), .B(n709), .ZN(n712) );
  NAND2_X1 U759 ( .A1(n712), .A2(n711), .ZN(n717) );
  XNOR2_X1 U760 ( .A(G227), .B(n713), .ZN(n714) );
  NAND2_X1 U761 ( .A1(n714), .A2(G900), .ZN(n715) );
  NAND2_X1 U762 ( .A1(n715), .A2(G953), .ZN(n716) );
  NAND2_X1 U763 ( .A1(n717), .A2(n716), .ZN(G72) );
  XOR2_X1 U764 ( .A(G140), .B(n718), .Z(G42) );
  XOR2_X1 U765 ( .A(n719), .B(G131), .Z(G33) );
  XOR2_X1 U766 ( .A(n590), .B(G122), .Z(G24) );
  XOR2_X1 U767 ( .A(n720), .B(G143), .Z(n721) );
  XNOR2_X1 U768 ( .A(KEYINPUT113), .B(n721), .ZN(G45) );
  XOR2_X1 U769 ( .A(G137), .B(n722), .Z(G39) );
  XOR2_X1 U770 ( .A(n723), .B(G119), .Z(n724) );
  XNOR2_X1 U771 ( .A(KEYINPUT127), .B(n724), .ZN(G21) );
endmodule

