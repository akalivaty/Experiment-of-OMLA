

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582;

  XOR2_X1 U322 ( .A(G64GAT), .B(G92GAT), .Z(n290) );
  AND2_X1 U323 ( .A1(n394), .A2(n552), .ZN(n395) );
  INV_X1 U324 ( .A(KEYINPUT54), .ZN(n419) );
  XOR2_X1 U325 ( .A(n386), .B(n373), .Z(n573) );
  XNOR2_X1 U326 ( .A(n441), .B(KEYINPUT58), .ZN(n442) );
  XNOR2_X1 U327 ( .A(n443), .B(n442), .ZN(G1351GAT) );
  XOR2_X1 U328 ( .A(KEYINPUT11), .B(KEYINPUT72), .Z(n292) );
  XNOR2_X1 U329 ( .A(G92GAT), .B(KEYINPUT71), .ZN(n291) );
  XNOR2_X1 U330 ( .A(n292), .B(n291), .ZN(n297) );
  XOR2_X1 U331 ( .A(G36GAT), .B(G190GAT), .Z(n409) );
  XNOR2_X1 U332 ( .A(G50GAT), .B(KEYINPUT69), .ZN(n293) );
  XNOR2_X1 U333 ( .A(n293), .B(G162GAT), .ZN(n314) );
  XOR2_X1 U334 ( .A(n409), .B(n314), .Z(n295) );
  XNOR2_X1 U335 ( .A(G134GAT), .B(G218GAT), .ZN(n294) );
  XNOR2_X1 U336 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U337 ( .A(n297), .B(n296), .ZN(n308) );
  XOR2_X1 U338 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n299) );
  NAND2_X1 U339 ( .A1(G232GAT), .A2(G233GAT), .ZN(n298) );
  XNOR2_X1 U340 ( .A(n299), .B(n298), .ZN(n300) );
  XOR2_X1 U341 ( .A(n300), .B(KEYINPUT70), .Z(n306) );
  XOR2_X1 U342 ( .A(G29GAT), .B(G43GAT), .Z(n302) );
  XNOR2_X1 U343 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U344 ( .A(n302), .B(n301), .ZN(n350) );
  XOR2_X1 U345 ( .A(KEYINPUT67), .B(G85GAT), .Z(n304) );
  XNOR2_X1 U346 ( .A(G99GAT), .B(G106GAT), .ZN(n303) );
  XNOR2_X1 U347 ( .A(n304), .B(n303), .ZN(n363) );
  XNOR2_X1 U348 ( .A(n350), .B(n363), .ZN(n305) );
  XNOR2_X1 U349 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U350 ( .A(n308), .B(n307), .Z(n552) );
  XOR2_X1 U351 ( .A(KEYINPUT23), .B(KEYINPUT22), .Z(n310) );
  XNOR2_X1 U352 ( .A(G204GAT), .B(KEYINPUT83), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U354 ( .A(n311), .B(G106GAT), .Z(n313) );
  XOR2_X1 U355 ( .A(G148GAT), .B(G78GAT), .Z(n370) );
  XNOR2_X1 U356 ( .A(G22GAT), .B(n370), .ZN(n312) );
  XNOR2_X1 U357 ( .A(n313), .B(n312), .ZN(n318) );
  XOR2_X1 U358 ( .A(n314), .B(KEYINPUT24), .Z(n316) );
  NAND2_X1 U359 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U360 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U361 ( .A(n318), .B(n317), .Z(n327) );
  XOR2_X1 U362 ( .A(KEYINPUT86), .B(KEYINPUT3), .Z(n320) );
  XNOR2_X1 U363 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n319) );
  XNOR2_X1 U364 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U365 ( .A(G141GAT), .B(n321), .Z(n341) );
  XNOR2_X1 U366 ( .A(G211GAT), .B(KEYINPUT84), .ZN(n322) );
  XNOR2_X1 U367 ( .A(n322), .B(KEYINPUT21), .ZN(n323) );
  XOR2_X1 U368 ( .A(n323), .B(KEYINPUT85), .Z(n325) );
  XNOR2_X1 U369 ( .A(G197GAT), .B(G218GAT), .ZN(n324) );
  XNOR2_X1 U370 ( .A(n325), .B(n324), .ZN(n410) );
  XNOR2_X1 U371 ( .A(n341), .B(n410), .ZN(n326) );
  XNOR2_X1 U372 ( .A(n327), .B(n326), .ZN(n461) );
  XOR2_X1 U373 ( .A(KEYINPUT1), .B(KEYINPUT4), .Z(n329) );
  XNOR2_X1 U374 ( .A(KEYINPUT6), .B(KEYINPUT88), .ZN(n328) );
  XNOR2_X1 U375 ( .A(n329), .B(n328), .ZN(n345) );
  XOR2_X1 U376 ( .A(G85GAT), .B(G148GAT), .Z(n331) );
  XNOR2_X1 U377 ( .A(G29GAT), .B(G162GAT), .ZN(n330) );
  XNOR2_X1 U378 ( .A(n331), .B(n330), .ZN(n335) );
  XOR2_X1 U379 ( .A(G57GAT), .B(KEYINPUT87), .Z(n333) );
  XNOR2_X1 U380 ( .A(G113GAT), .B(G1GAT), .ZN(n332) );
  XNOR2_X1 U381 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U382 ( .A(n335), .B(n334), .Z(n343) );
  XOR2_X1 U383 ( .A(G120GAT), .B(G127GAT), .Z(n337) );
  XNOR2_X1 U384 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n336) );
  XNOR2_X1 U385 ( .A(n337), .B(n336), .ZN(n429) );
  XOR2_X1 U386 ( .A(n429), .B(KEYINPUT5), .Z(n339) );
  NAND2_X1 U387 ( .A1(G225GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U388 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U389 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U390 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U391 ( .A(n345), .B(n344), .ZN(n513) );
  INV_X1 U392 ( .A(n513), .ZN(n485) );
  XOR2_X1 U393 ( .A(G113GAT), .B(G15GAT), .Z(n426) );
  XNOR2_X1 U394 ( .A(G22GAT), .B(G1GAT), .ZN(n346) );
  XNOR2_X1 U395 ( .A(n346), .B(KEYINPUT66), .ZN(n387) );
  XOR2_X1 U396 ( .A(n426), .B(n387), .Z(n348) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U398 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U399 ( .A(n349), .B(KEYINPUT29), .Z(n352) );
  XNOR2_X1 U400 ( .A(n350), .B(KEYINPUT65), .ZN(n351) );
  XNOR2_X1 U401 ( .A(n352), .B(n351), .ZN(n360) );
  XOR2_X1 U402 ( .A(G197GAT), .B(G141GAT), .Z(n354) );
  XNOR2_X1 U403 ( .A(G50GAT), .B(G36GAT), .ZN(n353) );
  XNOR2_X1 U404 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U405 ( .A(KEYINPUT64), .B(KEYINPUT30), .Z(n356) );
  XNOR2_X1 U406 ( .A(G169GAT), .B(G8GAT), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U408 ( .A(n358), .B(n357), .Z(n359) );
  XOR2_X1 U409 ( .A(n360), .B(n359), .Z(n499) );
  INV_X1 U410 ( .A(n499), .ZN(n567) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G57GAT), .ZN(n361) );
  XOR2_X1 U412 ( .A(n361), .B(KEYINPUT13), .Z(n386) );
  XNOR2_X1 U413 ( .A(G176GAT), .B(G204GAT), .ZN(n362) );
  XNOR2_X1 U414 ( .A(n290), .B(n362), .ZN(n404) );
  XNOR2_X1 U415 ( .A(n363), .B(n404), .ZN(n368) );
  XOR2_X1 U416 ( .A(KEYINPUT31), .B(KEYINPUT33), .Z(n365) );
  NAND2_X1 U417 ( .A1(G230GAT), .A2(G233GAT), .ZN(n364) );
  XNOR2_X1 U418 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U419 ( .A(n366), .B(KEYINPUT68), .Z(n367) );
  XNOR2_X1 U420 ( .A(n368), .B(n367), .ZN(n369) );
  XOR2_X1 U421 ( .A(n369), .B(KEYINPUT32), .Z(n372) );
  XNOR2_X1 U422 ( .A(G120GAT), .B(n370), .ZN(n371) );
  XNOR2_X1 U423 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U424 ( .A(n573), .B(KEYINPUT41), .Z(n498) );
  NOR2_X1 U425 ( .A1(n567), .A2(n498), .ZN(n374) );
  XNOR2_X1 U426 ( .A(n374), .B(KEYINPUT46), .ZN(n392) );
  XOR2_X1 U427 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n376) );
  XNOR2_X1 U428 ( .A(G15GAT), .B(G64GAT), .ZN(n375) );
  XNOR2_X1 U429 ( .A(n376), .B(n375), .ZN(n391) );
  XOR2_X1 U430 ( .A(G8GAT), .B(G183GAT), .Z(n407) );
  XOR2_X1 U431 ( .A(G78GAT), .B(G211GAT), .Z(n378) );
  XNOR2_X1 U432 ( .A(G127GAT), .B(G155GAT), .ZN(n377) );
  XNOR2_X1 U433 ( .A(n378), .B(n377), .ZN(n379) );
  XOR2_X1 U434 ( .A(n407), .B(n379), .Z(n381) );
  NAND2_X1 U435 ( .A1(G231GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U436 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT73), .Z(n383) );
  XNOR2_X1 U438 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n382) );
  XNOR2_X1 U439 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U440 ( .A(n385), .B(n384), .Z(n389) );
  XOR2_X1 U441 ( .A(n387), .B(n386), .Z(n388) );
  XNOR2_X1 U442 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U443 ( .A(n391), .B(n390), .ZN(n565) );
  INV_X1 U444 ( .A(n565), .ZN(n478) );
  NOR2_X1 U445 ( .A1(n392), .A2(n478), .ZN(n393) );
  XNOR2_X1 U446 ( .A(n393), .B(KEYINPUT108), .ZN(n394) );
  INV_X1 U447 ( .A(n552), .ZN(n396) );
  XNOR2_X1 U448 ( .A(n395), .B(KEYINPUT47), .ZN(n401) );
  INV_X1 U449 ( .A(n573), .ZN(n451) );
  XOR2_X1 U450 ( .A(KEYINPUT36), .B(n396), .Z(n579) );
  NOR2_X1 U451 ( .A1(n579), .A2(n565), .ZN(n397) );
  XOR2_X1 U452 ( .A(KEYINPUT45), .B(n397), .Z(n398) );
  NOR2_X1 U453 ( .A1(n451), .A2(n398), .ZN(n399) );
  NAND2_X1 U454 ( .A1(n399), .A2(n567), .ZN(n400) );
  NAND2_X1 U455 ( .A1(n401), .A2(n400), .ZN(n403) );
  XNOR2_X1 U456 ( .A(KEYINPUT109), .B(KEYINPUT48), .ZN(n402) );
  XNOR2_X1 U457 ( .A(n403), .B(n402), .ZN(n527) );
  XOR2_X1 U458 ( .A(n404), .B(KEYINPUT89), .Z(n406) );
  NAND2_X1 U459 ( .A1(G226GAT), .A2(G233GAT), .ZN(n405) );
  XNOR2_X1 U460 ( .A(n406), .B(n405), .ZN(n408) );
  XOR2_X1 U461 ( .A(n408), .B(n407), .Z(n412) );
  XNOR2_X1 U462 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U463 ( .A(n412), .B(n411), .ZN(n417) );
  XNOR2_X1 U464 ( .A(KEYINPUT17), .B(KEYINPUT19), .ZN(n413) );
  XNOR2_X1 U465 ( .A(n413), .B(KEYINPUT79), .ZN(n414) );
  XOR2_X1 U466 ( .A(n414), .B(KEYINPUT80), .Z(n416) );
  XNOR2_X1 U467 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n415) );
  XOR2_X1 U468 ( .A(n416), .B(n415), .Z(n437) );
  XOR2_X1 U469 ( .A(n417), .B(n437), .Z(n489) );
  XNOR2_X1 U470 ( .A(KEYINPUT117), .B(n489), .ZN(n418) );
  NOR2_X1 U471 ( .A1(n527), .A2(n418), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n420), .B(n419), .ZN(n421) );
  NOR2_X1 U473 ( .A1(n485), .A2(n421), .ZN(n446) );
  NAND2_X1 U474 ( .A1(n461), .A2(n446), .ZN(n422) );
  XNOR2_X1 U475 ( .A(n422), .B(KEYINPUT55), .ZN(n440) );
  XOR2_X1 U476 ( .A(KEYINPUT82), .B(G71GAT), .Z(n424) );
  XNOR2_X1 U477 ( .A(G190GAT), .B(G176GAT), .ZN(n423) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U479 ( .A(n425), .B(G99GAT), .Z(n428) );
  XNOR2_X1 U480 ( .A(G43GAT), .B(n426), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n428), .B(n427), .ZN(n433) );
  XOR2_X1 U482 ( .A(G183GAT), .B(n429), .Z(n431) );
  NAND2_X1 U483 ( .A1(G227GAT), .A2(G233GAT), .ZN(n430) );
  XNOR2_X1 U484 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U485 ( .A(n433), .B(n432), .Z(n439) );
  XOR2_X1 U486 ( .A(KEYINPUT78), .B(KEYINPUT20), .Z(n435) );
  XNOR2_X1 U487 ( .A(KEYINPUT81), .B(KEYINPUT77), .ZN(n434) );
  XNOR2_X1 U488 ( .A(n435), .B(n434), .ZN(n436) );
  XOR2_X1 U489 ( .A(n437), .B(n436), .Z(n438) );
  XOR2_X1 U490 ( .A(n439), .B(n438), .Z(n519) );
  INV_X1 U491 ( .A(n519), .ZN(n528) );
  NAND2_X1 U492 ( .A1(n440), .A2(n528), .ZN(n564) );
  NOR2_X1 U493 ( .A1(n552), .A2(n564), .ZN(n443) );
  INV_X1 U494 ( .A(G190GAT), .ZN(n441) );
  XNOR2_X1 U495 ( .A(KEYINPUT26), .B(KEYINPUT90), .ZN(n445) );
  NOR2_X1 U496 ( .A1(n528), .A2(n461), .ZN(n444) );
  XNOR2_X1 U497 ( .A(n445), .B(n444), .ZN(n543) );
  NAND2_X1 U498 ( .A1(n543), .A2(n446), .ZN(n447) );
  XOR2_X1 U499 ( .A(n447), .B(KEYINPUT121), .Z(n578) );
  NOR2_X1 U500 ( .A1(n565), .A2(n578), .ZN(n448) );
  XNOR2_X1 U501 ( .A(n448), .B(KEYINPUT126), .ZN(n450) );
  INV_X1 U502 ( .A(G211GAT), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n450), .B(n449), .ZN(G1354GAT) );
  NOR2_X1 U504 ( .A1(n451), .A2(n567), .ZN(n482) );
  XOR2_X1 U505 ( .A(KEYINPUT16), .B(KEYINPUT76), .Z(n453) );
  NAND2_X1 U506 ( .A1(n478), .A2(n552), .ZN(n452) );
  XNOR2_X1 U507 ( .A(n453), .B(n452), .ZN(n465) );
  NAND2_X1 U508 ( .A1(n528), .A2(n489), .ZN(n454) );
  NAND2_X1 U509 ( .A1(n461), .A2(n454), .ZN(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT25), .B(n455), .Z(n457) );
  XNOR2_X1 U511 ( .A(n489), .B(KEYINPUT27), .ZN(n460) );
  NAND2_X1 U512 ( .A1(n543), .A2(n460), .ZN(n456) );
  NAND2_X1 U513 ( .A1(n457), .A2(n456), .ZN(n458) );
  NAND2_X1 U514 ( .A1(n513), .A2(n458), .ZN(n459) );
  XOR2_X1 U515 ( .A(KEYINPUT91), .B(n459), .Z(n464) );
  NAND2_X1 U516 ( .A1(n485), .A2(n460), .ZN(n526) );
  NOR2_X1 U517 ( .A1(n528), .A2(n526), .ZN(n462) );
  XOR2_X1 U518 ( .A(n461), .B(KEYINPUT28), .Z(n495) );
  INV_X1 U519 ( .A(n495), .ZN(n530) );
  NAND2_X1 U520 ( .A1(n462), .A2(n530), .ZN(n463) );
  NAND2_X1 U521 ( .A1(n464), .A2(n463), .ZN(n479) );
  AND2_X1 U522 ( .A1(n465), .A2(n479), .ZN(n500) );
  NAND2_X1 U523 ( .A1(n482), .A2(n500), .ZN(n475) );
  NOR2_X1 U524 ( .A1(n513), .A2(n475), .ZN(n467) );
  XNOR2_X1 U525 ( .A(KEYINPUT34), .B(KEYINPUT92), .ZN(n466) );
  XNOR2_X1 U526 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U527 ( .A(G1GAT), .B(n468), .Z(G1324GAT) );
  INV_X1 U528 ( .A(n489), .ZN(n516) );
  NOR2_X1 U529 ( .A1(n516), .A2(n475), .ZN(n470) );
  XNOR2_X1 U530 ( .A(G8GAT), .B(KEYINPUT93), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(G1325GAT) );
  NOR2_X1 U532 ( .A1(n475), .A2(n519), .ZN(n474) );
  XOR2_X1 U533 ( .A(KEYINPUT94), .B(KEYINPUT95), .Z(n472) );
  XNOR2_X1 U534 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n471) );
  XNOR2_X1 U535 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(G1326GAT) );
  NOR2_X1 U537 ( .A1(n530), .A2(n475), .ZN(n476) );
  XOR2_X1 U538 ( .A(KEYINPUT96), .B(n476), .Z(n477) );
  XNOR2_X1 U539 ( .A(G22GAT), .B(n477), .ZN(G1327GAT) );
  NOR2_X1 U540 ( .A1(n579), .A2(n478), .ZN(n480) );
  NAND2_X1 U541 ( .A1(n480), .A2(n479), .ZN(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT37), .B(n481), .ZN(n512) );
  NAND2_X1 U543 ( .A1(n512), .A2(n482), .ZN(n484) );
  XOR2_X1 U544 ( .A(KEYINPUT98), .B(KEYINPUT38), .Z(n483) );
  XNOR2_X1 U545 ( .A(n484), .B(n483), .ZN(n494) );
  NAND2_X1 U546 ( .A1(n494), .A2(n485), .ZN(n488) );
  XNOR2_X1 U547 ( .A(G29GAT), .B(KEYINPUT97), .ZN(n486) );
  XNOR2_X1 U548 ( .A(n486), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n488), .B(n487), .ZN(G1328GAT) );
  XOR2_X1 U550 ( .A(G36GAT), .B(KEYINPUT99), .Z(n491) );
  NAND2_X1 U551 ( .A1(n494), .A2(n489), .ZN(n490) );
  XNOR2_X1 U552 ( .A(n491), .B(n490), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n494), .A2(n528), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XNOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT100), .ZN(n497) );
  NAND2_X1 U557 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U558 ( .A(n497), .B(n496), .ZN(G1331GAT) );
  BUF_X1 U559 ( .A(n498), .Z(n561) );
  NOR2_X1 U560 ( .A1(n499), .A2(n561), .ZN(n511) );
  NAND2_X1 U561 ( .A1(n511), .A2(n500), .ZN(n507) );
  NOR2_X1 U562 ( .A1(n513), .A2(n507), .ZN(n502) );
  XNOR2_X1 U563 ( .A(KEYINPUT101), .B(KEYINPUT42), .ZN(n501) );
  XNOR2_X1 U564 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(n503), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n516), .A2(n507), .ZN(n504) );
  XOR2_X1 U567 ( .A(KEYINPUT102), .B(n504), .Z(n505) );
  XNOR2_X1 U568 ( .A(G64GAT), .B(n505), .ZN(G1333GAT) );
  NOR2_X1 U569 ( .A1(n519), .A2(n507), .ZN(n506) );
  XOR2_X1 U570 ( .A(G71GAT), .B(n506), .Z(G1334GAT) );
  NOR2_X1 U571 ( .A1(n530), .A2(n507), .ZN(n509) );
  XNOR2_X1 U572 ( .A(KEYINPUT43), .B(KEYINPUT103), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n509), .B(n508), .ZN(n510) );
  XOR2_X1 U574 ( .A(G78GAT), .B(n510), .Z(G1335GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n511), .ZN(n523) );
  NOR2_X1 U576 ( .A1(n513), .A2(n523), .ZN(n514) );
  XOR2_X1 U577 ( .A(G85GAT), .B(n514), .Z(n515) );
  XNOR2_X1 U578 ( .A(KEYINPUT104), .B(n515), .ZN(G1336GAT) );
  NOR2_X1 U579 ( .A1(n516), .A2(n523), .ZN(n518) );
  XNOR2_X1 U580 ( .A(G92GAT), .B(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U582 ( .A1(n519), .A2(n523), .ZN(n520) );
  XOR2_X1 U583 ( .A(G99GAT), .B(n520), .Z(G1338GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(KEYINPUT106), .Z(n522) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n522), .B(n521), .ZN(n525) );
  NOR2_X1 U587 ( .A1(n530), .A2(n523), .ZN(n524) );
  XOR2_X1 U588 ( .A(n525), .B(n524), .Z(G1339GAT) );
  NOR2_X1 U589 ( .A1(n527), .A2(n526), .ZN(n542) );
  NAND2_X1 U590 ( .A1(n528), .A2(n542), .ZN(n529) );
  XOR2_X1 U591 ( .A(KEYINPUT110), .B(n529), .Z(n531) );
  NAND2_X1 U592 ( .A1(n531), .A2(n530), .ZN(n539) );
  NOR2_X1 U593 ( .A1(n567), .A2(n539), .ZN(n533) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(KEYINPUT111), .ZN(n532) );
  XNOR2_X1 U595 ( .A(n533), .B(n532), .ZN(G1340GAT) );
  NOR2_X1 U596 ( .A1(n561), .A2(n539), .ZN(n535) );
  XNOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n534) );
  XNOR2_X1 U598 ( .A(n535), .B(n534), .ZN(G1341GAT) );
  NOR2_X1 U599 ( .A1(n565), .A2(n539), .ZN(n537) );
  XNOR2_X1 U600 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n536) );
  XNOR2_X1 U601 ( .A(n537), .B(n536), .ZN(n538) );
  XOR2_X1 U602 ( .A(G127GAT), .B(n538), .Z(G1342GAT) );
  NOR2_X1 U603 ( .A1(n552), .A2(n539), .ZN(n541) );
  XNOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n543), .A2(n542), .ZN(n551) );
  NOR2_X1 U607 ( .A1(n567), .A2(n551), .ZN(n544) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n544), .Z(G1344GAT) );
  NOR2_X1 U609 ( .A1(n551), .A2(n561), .ZN(n548) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n546) );
  XNOR2_X1 U611 ( .A(G148GAT), .B(KEYINPUT113), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n547) );
  XNOR2_X1 U613 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NOR2_X1 U614 ( .A1(n565), .A2(n551), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT114), .B(n549), .Z(n550) );
  XNOR2_X1 U616 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U617 ( .A1(n552), .A2(n551), .ZN(n554) );
  XNOR2_X1 U618 ( .A(KEYINPUT115), .B(KEYINPUT116), .ZN(n553) );
  XNOR2_X1 U619 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  XNOR2_X1 U621 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n558) );
  NOR2_X1 U622 ( .A1(n564), .A2(n567), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n556), .B(KEYINPUT119), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  XNOR2_X1 U626 ( .A(G176GAT), .B(KEYINPUT120), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n563) );
  NOR2_X1 U628 ( .A1(n564), .A2(n561), .ZN(n562) );
  XOR2_X1 U629 ( .A(n563), .B(n562), .Z(G1349GAT) );
  NOR2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n566) );
  XOR2_X1 U631 ( .A(G183GAT), .B(n566), .Z(G1350GAT) );
  NOR2_X1 U632 ( .A1(n567), .A2(n578), .ZN(n572) );
  XOR2_X1 U633 ( .A(KEYINPUT60), .B(KEYINPUT123), .Z(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U635 ( .A(n569), .B(n568), .ZN(n570) );
  XNOR2_X1 U636 ( .A(KEYINPUT122), .B(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  NOR2_X1 U638 ( .A1(n578), .A2(n573), .ZN(n577) );
  XOR2_X1 U639 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n575) );
  XNOR2_X1 U640 ( .A(G204GAT), .B(KEYINPUT125), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT127), .B(KEYINPUT62), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(n582), .B(G218GAT), .ZN(G1355GAT) );
endmodule

