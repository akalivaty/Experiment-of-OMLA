//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 1 1 0 0 0 0 0 0 0 0 0 1 1 0 1 1 1 1 1 1 1 1 0 1 1 0 0 1 1 0 1 1 1 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 0 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:24:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n713, new_n714,
    new_n715, new_n716, new_n717, new_n718, new_n719, new_n720, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n733, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n757, new_n758, new_n759,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n825, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984, new_n985, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1027, new_n1028, new_n1029,
    new_n1030, new_n1031, new_n1032, new_n1033, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1053, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064, new_n1065, new_n1066, new_n1067;
  INV_X1    g000(.A(KEYINPUT25), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT77), .ZN(new_n188));
  INV_X1    g002(.A(G125), .ZN(new_n189));
  OAI211_X1 g003(.A(new_n188), .B(G140), .C1(new_n189), .C2(KEYINPUT76), .ZN(new_n190));
  INV_X1    g004(.A(G140), .ZN(new_n191));
  OAI21_X1  g005(.A(KEYINPUT77), .B1(new_n191), .B2(G125), .ZN(new_n192));
  INV_X1    g006(.A(KEYINPUT76), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n193), .A2(new_n191), .A3(G125), .ZN(new_n194));
  NAND4_X1  g008(.A1(new_n190), .A2(new_n192), .A3(new_n194), .A4(KEYINPUT16), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n189), .A2(G140), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT16), .ZN(new_n197));
  AOI21_X1  g011(.A(KEYINPUT78), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  AND2_X1   g012(.A1(new_n195), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT78), .ZN(new_n200));
  NOR2_X1   g014(.A1(new_n195), .A2(new_n200), .ZN(new_n201));
  OAI21_X1  g015(.A(G146), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(KEYINPUT78), .A3(KEYINPUT16), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n195), .A2(new_n198), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n204), .A2(new_n205), .A3(new_n206), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g022(.A1(G119), .A2(G128), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT66), .A2(G119), .ZN(new_n211));
  INV_X1    g025(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT66), .A2(G119), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G128), .ZN(new_n215));
  OAI21_X1  g029(.A(new_n210), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT75), .ZN(new_n217));
  XNOR2_X1  g031(.A(KEYINPUT66), .B(G119), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n209), .B1(new_n218), .B2(G128), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT75), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g035(.A(KEYINPUT24), .B(G110), .Z(new_n222));
  NAND3_X1  g036(.A1(new_n217), .A2(new_n221), .A3(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT23), .ZN(new_n224));
  OAI21_X1  g038(.A(new_n224), .B1(new_n214), .B2(G128), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n225), .B1(new_n216), .B2(new_n224), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(G110), .ZN(new_n227));
  NAND3_X1  g041(.A1(new_n208), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n189), .A2(G140), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n191), .A2(G125), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n229), .A2(new_n230), .A3(new_n205), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n226), .A2(G110), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n222), .B1(new_n217), .B2(new_n221), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n202), .B(new_n232), .C1(new_n233), .C2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n228), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G953), .ZN(new_n237));
  NAND3_X1  g051(.A1(new_n237), .A2(G221), .A3(G234), .ZN(new_n238));
  XNOR2_X1  g052(.A(new_n238), .B(KEYINPUT79), .ZN(new_n239));
  XNOR2_X1  g053(.A(KEYINPUT22), .B(G137), .ZN(new_n240));
  XNOR2_X1  g054(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g055(.A(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n236), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n228), .A2(new_n235), .A3(new_n241), .ZN(new_n244));
  AOI21_X1  g058(.A(G902), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n187), .B1(new_n245), .B2(KEYINPUT80), .ZN(new_n246));
  INV_X1    g060(.A(G902), .ZN(new_n247));
  INV_X1    g061(.A(new_n244), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n241), .B1(new_n228), .B2(new_n235), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n247), .B1(new_n248), .B2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT80), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(KEYINPUT25), .ZN(new_n252));
  INV_X1    g066(.A(G217), .ZN(new_n253));
  AOI21_X1  g067(.A(new_n253), .B1(G234), .B2(new_n247), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n246), .A2(new_n252), .A3(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n243), .A2(new_n244), .ZN(new_n256));
  NOR2_X1   g070(.A1(new_n254), .A2(G902), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT74), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT11), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n261), .B1(new_n262), .B2(G137), .ZN(new_n263));
  INV_X1    g077(.A(G137), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n264), .A2(KEYINPUT11), .A3(G134), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n262), .A2(G137), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G131), .ZN(new_n268));
  INV_X1    g082(.A(G131), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n263), .A2(new_n265), .A3(new_n269), .A4(new_n266), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n205), .A2(G143), .ZN(new_n272));
  INV_X1    g086(.A(G143), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n273), .A2(G146), .ZN(new_n274));
  NOR2_X1   g088(.A1(KEYINPUT0), .A2(G128), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n272), .A2(new_n274), .B1(new_n275), .B2(KEYINPUT64), .ZN(new_n276));
  AND2_X1   g090(.A1(KEYINPUT0), .A2(G128), .ZN(new_n277));
  OR2_X1    g091(.A1(KEYINPUT0), .A2(G128), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT64), .ZN(new_n279));
  AOI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  XNOR2_X1  g094(.A(G143), .B(G146), .ZN(new_n281));
  AOI22_X1  g095(.A1(new_n276), .A2(new_n280), .B1(new_n277), .B2(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n271), .A2(new_n282), .ZN(new_n283));
  OR2_X1    g097(.A1(KEYINPUT66), .A2(G119), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(G116), .A3(new_n211), .ZN(new_n285));
  INV_X1    g099(.A(G116), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G119), .ZN(new_n287));
  INV_X1    g101(.A(G113), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(KEYINPUT2), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT2), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n290), .A2(G113), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n285), .A2(new_n287), .A3(new_n292), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n292), .B1(new_n285), .B2(new_n287), .ZN(new_n294));
  NOR2_X1   g108(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(new_n266), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n262), .A2(G137), .ZN(new_n297));
  OAI21_X1  g111(.A(G131), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(KEYINPUT1), .B1(new_n273), .B2(G146), .ZN(new_n299));
  NOR2_X1   g113(.A1(new_n273), .A2(G146), .ZN(new_n300));
  NOR2_X1   g114(.A1(new_n205), .A2(G143), .ZN(new_n301));
  OAI211_X1 g115(.A(G128), .B(new_n299), .C1(new_n300), .C2(new_n301), .ZN(new_n302));
  OAI211_X1 g116(.A(new_n272), .B(new_n274), .C1(KEYINPUT1), .C2(new_n215), .ZN(new_n303));
  NAND4_X1  g117(.A1(new_n298), .A2(new_n302), .A3(new_n270), .A4(new_n303), .ZN(new_n304));
  NAND3_X1  g118(.A1(new_n283), .A2(new_n295), .A3(new_n304), .ZN(new_n305));
  INV_X1    g119(.A(KEYINPUT28), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g121(.A(KEYINPUT70), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n305), .A2(KEYINPUT70), .A3(new_n306), .ZN(new_n310));
  AND2_X1   g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT69), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n283), .A2(new_n304), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n285), .A2(new_n287), .ZN(new_n314));
  INV_X1    g128(.A(new_n292), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n285), .A2(new_n287), .A3(new_n292), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n313), .A2(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(new_n305), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n312), .B1(new_n320), .B2(KEYINPUT28), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n283), .A2(new_n295), .A3(new_n304), .ZN(new_n322));
  AOI21_X1  g136(.A(new_n295), .B1(new_n283), .B2(new_n304), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n312), .B(KEYINPUT28), .C1(new_n322), .C2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(new_n324), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n311), .B1(new_n321), .B2(new_n325), .ZN(new_n326));
  XOR2_X1   g140(.A(KEYINPUT67), .B(KEYINPUT27), .Z(new_n327));
  NOR2_X1   g141(.A1(G237), .A2(G953), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G210), .ZN(new_n329));
  XNOR2_X1  g143(.A(new_n327), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g144(.A(KEYINPUT26), .B(G101), .ZN(new_n331));
  XNOR2_X1  g145(.A(new_n330), .B(new_n331), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT30), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n333), .A2(KEYINPUT65), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n333), .A2(KEYINPUT65), .ZN(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  AOI211_X1 g150(.A(new_n334), .B(new_n336), .C1(new_n283), .C2(new_n304), .ZN(new_n337));
  NAND4_X1  g151(.A1(new_n283), .A2(KEYINPUT65), .A3(new_n333), .A4(new_n304), .ZN(new_n338));
  INV_X1    g152(.A(new_n338), .ZN(new_n339));
  OAI21_X1  g153(.A(new_n318), .B1(new_n337), .B2(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n332), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n340), .A2(new_n305), .A3(new_n341), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n326), .A2(new_n332), .B1(KEYINPUT31), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT31), .ZN(new_n344));
  NAND4_X1  g158(.A1(new_n340), .A2(new_n344), .A3(new_n305), .A4(new_n341), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT68), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n334), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n313), .A2(new_n348), .A3(new_n335), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n338), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n322), .B1(new_n350), .B2(new_n318), .ZN(new_n351));
  NAND4_X1  g165(.A1(new_n351), .A2(KEYINPUT68), .A3(new_n344), .A4(new_n341), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n347), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g167(.A1(new_n343), .A2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(G472), .A2(G902), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n355), .A2(KEYINPUT32), .ZN(new_n356));
  INV_X1    g170(.A(new_n356), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n260), .B1(new_n354), .B2(new_n357), .ZN(new_n358));
  AOI211_X1 g172(.A(KEYINPUT74), .B(new_n356), .C1(new_n343), .C2(new_n353), .ZN(new_n359));
  INV_X1    g173(.A(G472), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n361), .B1(new_n351), .B2(new_n341), .ZN(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n363), .B1(new_n332), .B2(new_n326), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n320), .A2(KEYINPUT28), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n332), .A2(new_n361), .ZN(new_n366));
  NAND4_X1  g180(.A1(new_n365), .A2(new_n309), .A3(new_n310), .A4(new_n366), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT73), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND4_X1  g183(.A1(new_n311), .A2(KEYINPUT73), .A3(new_n365), .A4(new_n366), .ZN(new_n370));
  AND3_X1   g184(.A1(new_n369), .A2(new_n370), .A3(new_n247), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n360), .B1(new_n364), .B2(new_n371), .ZN(new_n372));
  NOR3_X1   g186(.A1(new_n358), .A2(new_n359), .A3(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n353), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n342), .A2(KEYINPUT31), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n309), .A2(new_n310), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n365), .A2(KEYINPUT69), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n376), .B1(new_n377), .B2(new_n324), .ZN(new_n378));
  OAI21_X1  g192(.A(new_n375), .B1(new_n378), .B2(new_n341), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n355), .B1(new_n374), .B2(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n381));
  XOR2_X1   g195(.A(KEYINPUT71), .B(KEYINPUT32), .Z(new_n382));
  INV_X1    g196(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n380), .A2(new_n381), .A3(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(new_n355), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n385), .B1(new_n343), .B2(new_n353), .ZN(new_n386));
  OAI21_X1  g200(.A(KEYINPUT72), .B1(new_n386), .B2(new_n382), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n384), .A2(new_n387), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n259), .B1(new_n373), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT90), .ZN(new_n390));
  OAI21_X1  g204(.A(G210), .B1(G237), .B2(G902), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n285), .A2(KEYINPUT5), .A3(new_n287), .ZN(new_n393));
  NOR3_X1   g207(.A1(new_n212), .A2(new_n213), .A3(new_n286), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT5), .ZN(new_n395));
  AOI21_X1  g209(.A(new_n288), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  AOI21_X1  g210(.A(new_n293), .B1(new_n393), .B2(new_n396), .ZN(new_n397));
  INV_X1    g211(.A(KEYINPUT3), .ZN(new_n398));
  INV_X1    g212(.A(G104), .ZN(new_n399));
  OAI21_X1  g213(.A(new_n398), .B1(new_n399), .B2(G107), .ZN(new_n400));
  INV_X1    g214(.A(G107), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT3), .A3(G104), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(G101), .ZN(new_n404));
  OAI21_X1  g218(.A(KEYINPUT81), .B1(new_n401), .B2(G104), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT81), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n406), .A2(new_n399), .A3(G107), .ZN(new_n407));
  NAND4_X1  g221(.A1(new_n403), .A2(new_n404), .A3(new_n405), .A4(new_n407), .ZN(new_n408));
  OAI21_X1  g222(.A(KEYINPUT82), .B1(new_n399), .B2(G107), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT82), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n410), .A2(new_n401), .A3(G104), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n399), .A2(G107), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n409), .A2(new_n411), .A3(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n413), .A2(G101), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n408), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT84), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT84), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n408), .A2(new_n414), .A3(new_n417), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n397), .A2(new_n416), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n405), .A2(new_n407), .ZN(new_n420));
  AOI21_X1  g234(.A(new_n404), .B1(new_n420), .B2(new_n403), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT4), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n408), .A2(KEYINPUT4), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(new_n318), .C1(new_n421), .C2(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n419), .A2(new_n425), .ZN(new_n426));
  XNOR2_X1  g240(.A(G110), .B(G122), .ZN(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n426), .A2(KEYINPUT89), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT6), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n427), .B1(new_n419), .B2(new_n425), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT6), .ZN(new_n432));
  NAND3_X1  g246(.A1(new_n431), .A2(KEYINPUT89), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n430), .A2(new_n433), .ZN(new_n434));
  NAND3_X1  g248(.A1(new_n419), .A2(new_n425), .A3(new_n427), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT88), .ZN(new_n436));
  INV_X1    g250(.A(new_n431), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT88), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n419), .A2(new_n425), .A3(new_n438), .A4(new_n427), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(G224), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n441), .A2(G953), .ZN(new_n442));
  NOR2_X1   g256(.A1(new_n282), .A2(new_n189), .ZN(new_n443));
  AOI21_X1  g257(.A(G125), .B1(new_n302), .B2(new_n303), .ZN(new_n444));
  OAI21_X1  g258(.A(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n276), .A2(new_n280), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n281), .A2(new_n277), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(G125), .ZN(new_n449));
  INV_X1    g263(.A(new_n442), .ZN(new_n450));
  INV_X1    g264(.A(new_n444), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  AOI22_X1  g266(.A1(new_n434), .A2(new_n440), .B1(new_n445), .B2(new_n452), .ZN(new_n453));
  XOR2_X1   g267(.A(new_n427), .B(KEYINPUT8), .Z(new_n454));
  INV_X1    g268(.A(new_n415), .ZN(new_n455));
  OR2_X1    g269(.A1(new_n397), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n454), .B1(new_n456), .B2(new_n419), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n442), .A2(KEYINPUT7), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n458), .B1(new_n445), .B2(new_n452), .ZN(new_n459));
  AOI211_X1 g273(.A(KEYINPUT7), .B(new_n442), .C1(new_n449), .C2(new_n451), .ZN(new_n460));
  NOR3_X1   g274(.A1(new_n457), .A2(new_n459), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n436), .A2(new_n439), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(new_n247), .ZN(new_n464));
  OAI21_X1  g278(.A(new_n392), .B1(new_n453), .B2(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(new_n433), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n432), .B1(new_n431), .B2(KEYINPUT89), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n440), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n445), .A2(new_n452), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  AOI21_X1  g284(.A(G902), .B1(new_n461), .B2(new_n462), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n470), .A2(new_n471), .A3(new_n391), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n465), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G214), .B1(G237), .B2(G902), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n390), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n474), .ZN(new_n476));
  AOI211_X1 g290(.A(KEYINPUT90), .B(new_n476), .C1(new_n465), .C2(new_n472), .ZN(new_n477));
  INV_X1    g291(.A(G475), .ZN(new_n478));
  INV_X1    g292(.A(G237), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n479), .A2(new_n237), .A3(G214), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n273), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n328), .A2(G143), .A3(G214), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G131), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT17), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n481), .A2(new_n269), .A3(new_n482), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n483), .A2(KEYINPUT17), .A3(G131), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n202), .A2(new_n207), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  XNOR2_X1  g303(.A(G113), .B(G122), .ZN(new_n490));
  XNOR2_X1  g304(.A(new_n490), .B(new_n399), .ZN(new_n491));
  OAI21_X1  g305(.A(new_n232), .B1(new_n203), .B2(new_n205), .ZN(new_n492));
  INV_X1    g306(.A(KEYINPUT91), .ZN(new_n493));
  NAND2_X1  g307(.A1(KEYINPUT18), .A2(G131), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n481), .A2(new_n482), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n494), .ZN(new_n496));
  AND4_X1   g310(.A1(G143), .A2(new_n479), .A3(new_n237), .A4(G214), .ZN(new_n497));
  AOI21_X1  g311(.A(G143), .B1(new_n328), .B2(G214), .ZN(new_n498));
  OAI21_X1  g312(.A(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND4_X1  g313(.A1(new_n492), .A2(new_n493), .A3(new_n495), .A4(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n499), .A2(new_n495), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n190), .A2(new_n192), .A3(new_n194), .ZN(new_n502));
  AOI21_X1  g316(.A(new_n231), .B1(G146), .B2(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(KEYINPUT91), .B1(new_n501), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n500), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n489), .A2(new_n491), .A3(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT93), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT93), .ZN(new_n508));
  NAND4_X1  g322(.A1(new_n489), .A2(new_n505), .A3(new_n508), .A4(new_n491), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AND2_X1   g324(.A1(new_n489), .A2(new_n505), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n491), .B2(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n478), .B1(new_n512), .B2(new_n247), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT94), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n484), .A2(new_n486), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT19), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n229), .A2(new_n230), .A3(new_n516), .ZN(new_n517));
  INV_X1    g331(.A(KEYINPUT92), .ZN(new_n518));
  OR2_X1    g332(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n518), .ZN(new_n520));
  OAI211_X1 g334(.A(new_n519), .B(new_n520), .C1(new_n516), .C2(new_n203), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n515), .B1(new_n521), .B2(G146), .ZN(new_n522));
  INV_X1    g336(.A(new_n202), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n505), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(new_n491), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n514), .B1(new_n510), .B2(new_n526), .ZN(new_n527));
  AOI22_X1  g341(.A1(new_n507), .A2(new_n509), .B1(new_n525), .B2(new_n524), .ZN(new_n528));
  NOR2_X1   g342(.A1(G475), .A2(G902), .ZN(new_n529));
  INV_X1    g343(.A(new_n529), .ZN(new_n530));
  OAI22_X1  g344(.A1(new_n527), .A2(KEYINPUT20), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n510), .A2(new_n526), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n532), .A2(new_n514), .A3(new_n533), .A4(new_n529), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n513), .B1(new_n531), .B2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(G478), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(KEYINPUT15), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT9), .B(G234), .ZN(new_n538));
  NOR3_X1   g352(.A1(new_n538), .A2(new_n253), .A3(G953), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  OAI21_X1  g354(.A(KEYINPUT95), .B1(new_n286), .B2(G122), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT95), .ZN(new_n542));
  INV_X1    g356(.A(G122), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n542), .A2(new_n543), .A3(G116), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  AOI21_X1  g359(.A(new_n401), .B1(new_n545), .B2(KEYINPUT14), .ZN(new_n546));
  AOI22_X1  g360(.A1(new_n541), .A2(new_n544), .B1(new_n286), .B2(G122), .ZN(new_n547));
  INV_X1    g361(.A(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n546), .A2(new_n548), .ZN(new_n549));
  OAI221_X1 g363(.A(new_n545), .B1(KEYINPUT14), .B2(new_n401), .C1(G116), .C2(new_n543), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(KEYINPUT96), .B1(new_n273), .B2(G128), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT96), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n215), .A3(G143), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT97), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n273), .A2(G128), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n556), .B1(new_n555), .B2(new_n557), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n262), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n560), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n562), .A2(G134), .A3(new_n558), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n551), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  AOI21_X1  g378(.A(G134), .B1(new_n562), .B2(new_n558), .ZN(new_n565));
  INV_X1    g379(.A(KEYINPUT13), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n557), .A2(new_n566), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n273), .A2(KEYINPUT13), .A3(G128), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n555), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(G134), .ZN(new_n570));
  AND2_X1   g384(.A1(new_n547), .A2(new_n401), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n547), .A2(new_n401), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n570), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n565), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g388(.A(new_n540), .B1(new_n564), .B2(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n549), .A2(new_n550), .ZN(new_n576));
  NOR3_X1   g390(.A1(new_n559), .A2(new_n262), .A3(new_n560), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n576), .B1(new_n565), .B2(new_n577), .ZN(new_n578));
  OAI211_X1 g392(.A(new_n561), .B(new_n570), .C1(new_n572), .C2(new_n571), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n578), .A2(new_n579), .A3(new_n539), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT98), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g396(.A(KEYINPUT98), .B(new_n540), .C1(new_n564), .C2(new_n574), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n582), .A2(new_n247), .A3(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n537), .B1(new_n584), .B2(KEYINPUT99), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(KEYINPUT99), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT99), .ZN(new_n587));
  NAND4_X1  g401(.A1(new_n582), .A2(new_n587), .A3(new_n247), .A4(new_n583), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n585), .B1(new_n589), .B2(new_n537), .ZN(new_n590));
  XNOR2_X1  g404(.A(KEYINPUT21), .B(G898), .ZN(new_n591));
  XNOR2_X1  g405(.A(new_n591), .B(KEYINPUT100), .ZN(new_n592));
  NAND2_X1  g406(.A1(G234), .A2(G237), .ZN(new_n593));
  AND3_X1   g407(.A1(new_n593), .A2(G902), .A3(G953), .ZN(new_n594));
  AND2_X1   g408(.A1(new_n592), .A2(new_n594), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n593), .A2(G952), .A3(new_n237), .ZN(new_n596));
  OR2_X1    g410(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  XOR2_X1   g411(.A(new_n597), .B(KEYINPUT101), .Z(new_n598));
  NAND3_X1  g412(.A1(new_n535), .A2(new_n590), .A3(new_n598), .ZN(new_n599));
  NOR3_X1   g413(.A1(new_n475), .A2(new_n477), .A3(new_n599), .ZN(new_n600));
  INV_X1    g414(.A(G469), .ZN(new_n601));
  XNOR2_X1  g415(.A(G110), .B(G140), .ZN(new_n602));
  INV_X1    g416(.A(G227), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G953), .ZN(new_n604));
  XNOR2_X1  g418(.A(new_n602), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n302), .A2(new_n303), .ZN(new_n606));
  OAI21_X1  g420(.A(KEYINPUT83), .B1(new_n415), .B2(new_n606), .ZN(new_n607));
  AND2_X1   g421(.A1(new_n302), .A2(new_n303), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT83), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n608), .A2(new_n609), .A3(new_n408), .A4(new_n414), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  AND3_X1   g425(.A1(new_n408), .A2(new_n414), .A3(new_n417), .ZN(new_n612));
  AOI21_X1  g426(.A(new_n417), .B1(new_n408), .B2(new_n414), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n606), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n611), .A2(new_n614), .ZN(new_n615));
  AOI21_X1  g429(.A(KEYINPUT12), .B1(new_n615), .B2(new_n271), .ZN(new_n616));
  INV_X1    g430(.A(KEYINPUT12), .ZN(new_n617));
  INV_X1    g431(.A(new_n271), .ZN(new_n618));
  AOI211_X1 g432(.A(new_n617), .B(new_n618), .C1(new_n611), .C2(new_n614), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g434(.A(KEYINPUT10), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n606), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n416), .A2(new_n418), .A3(new_n622), .ZN(new_n623));
  OAI211_X1 g437(.A(new_n423), .B(new_n282), .C1(new_n421), .C2(new_n424), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g439(.A(KEYINPUT10), .B1(new_n607), .B2(new_n610), .ZN(new_n626));
  NOR3_X1   g440(.A1(new_n625), .A2(new_n626), .A3(new_n271), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n605), .B1(new_n620), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n612), .A2(new_n613), .ZN(new_n629));
  OR2_X1    g443(.A1(new_n424), .A2(new_n421), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n448), .B1(new_n422), .B2(new_n421), .ZN(new_n631));
  AOI22_X1  g445(.A1(new_n629), .A2(new_n622), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n611), .A2(new_n621), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(new_n633), .A3(new_n618), .ZN(new_n634));
  INV_X1    g448(.A(new_n605), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(new_n618), .B1(new_n632), .B2(new_n633), .ZN(new_n637));
  OAI21_X1  g451(.A(new_n628), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n601), .B1(new_n638), .B2(new_n247), .ZN(new_n639));
  INV_X1    g453(.A(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(KEYINPUT86), .ZN(new_n641));
  OAI21_X1  g455(.A(new_n605), .B1(new_n637), .B2(new_n627), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n416), .A2(new_n418), .ZN(new_n643));
  AOI22_X1  g457(.A1(new_n643), .A2(new_n606), .B1(new_n607), .B2(new_n610), .ZN(new_n644));
  OAI21_X1  g458(.A(new_n617), .B1(new_n644), .B2(new_n618), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n615), .A2(KEYINPUT12), .A3(new_n271), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n625), .A2(new_n626), .ZN(new_n648));
  AOI21_X1  g462(.A(new_n605), .B1(new_n648), .B2(new_n618), .ZN(new_n649));
  AOI22_X1  g463(.A1(new_n642), .A2(KEYINPUT85), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n271), .B1(new_n625), .B2(new_n626), .ZN(new_n651));
  AOI21_X1  g465(.A(new_n635), .B1(new_n634), .B2(new_n651), .ZN(new_n652));
  INV_X1    g466(.A(KEYINPUT85), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  AOI21_X1  g468(.A(G902), .B1(new_n650), .B2(new_n654), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n641), .B1(new_n655), .B2(new_n601), .ZN(new_n656));
  OAI22_X1  g470(.A1(new_n652), .A2(new_n653), .B1(new_n620), .B2(new_n636), .ZN(new_n657));
  AOI211_X1 g471(.A(KEYINPUT85), .B(new_n635), .C1(new_n634), .C2(new_n651), .ZN(new_n658));
  OAI211_X1 g472(.A(new_n601), .B(new_n247), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  NOR2_X1   g473(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n640), .B1(new_n656), .B2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(KEYINPUT87), .ZN(new_n662));
  OAI21_X1  g476(.A(G221), .B1(new_n538), .B2(G902), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n661), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n659), .A2(KEYINPUT86), .ZN(new_n665));
  NAND2_X1  g479(.A1(new_n642), .A2(KEYINPUT85), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n647), .A2(new_n649), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n654), .A3(new_n667), .ZN(new_n668));
  NAND4_X1  g482(.A1(new_n668), .A2(new_n641), .A3(new_n601), .A4(new_n247), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n639), .B1(new_n665), .B2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n663), .ZN(new_n671));
  OAI21_X1  g485(.A(KEYINPUT87), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND4_X1  g486(.A1(new_n389), .A2(new_n600), .A3(new_n664), .A4(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G101), .ZN(G3));
  AOI21_X1  g488(.A(new_n662), .B1(new_n661), .B2(new_n663), .ZN(new_n675));
  NOR3_X1   g489(.A1(new_n670), .A2(KEYINPUT87), .A3(new_n671), .ZN(new_n676));
  NOR2_X1   g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI21_X1  g491(.A(G902), .B1(new_n343), .B2(new_n353), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n380), .B1(new_n360), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g493(.A1(new_n679), .A2(new_n259), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n476), .B1(new_n465), .B2(new_n472), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n681), .A2(new_n598), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n531), .A2(new_n534), .ZN(new_n683));
  INV_X1    g497(.A(new_n513), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(KEYINPUT33), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n582), .A2(new_n686), .A3(new_n583), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n575), .A2(new_n580), .A3(KEYINPUT33), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n687), .A2(new_n688), .A3(G478), .A4(new_n247), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n584), .A2(new_n536), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n685), .A2(KEYINPUT102), .A3(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT102), .ZN(new_n693));
  INV_X1    g507(.A(new_n691), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n693), .B1(new_n535), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n682), .B1(new_n692), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n677), .A2(new_n680), .A3(new_n696), .ZN(new_n697));
  XOR2_X1   g511(.A(KEYINPUT34), .B(G104), .Z(new_n698));
  XNOR2_X1  g512(.A(new_n697), .B(new_n698), .ZN(G6));
  NAND2_X1  g513(.A1(new_n589), .A2(new_n537), .ZN(new_n700));
  INV_X1    g514(.A(new_n585), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n532), .A2(new_n529), .ZN(new_n703));
  NOR2_X1   g517(.A1(KEYINPUT103), .A2(KEYINPUT20), .ZN(new_n704));
  AND2_X1   g518(.A1(KEYINPUT103), .A2(KEYINPUT20), .ZN(new_n705));
  OAI21_X1  g519(.A(new_n703), .B1(new_n704), .B2(new_n705), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n706), .B1(new_n703), .B2(new_n705), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n702), .A2(new_n707), .A3(new_n684), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n682), .A2(new_n708), .ZN(new_n709));
  NAND3_X1  g523(.A1(new_n677), .A2(new_n680), .A3(new_n709), .ZN(new_n710));
  XOR2_X1   g524(.A(KEYINPUT35), .B(G107), .Z(new_n711));
  XNOR2_X1  g525(.A(new_n710), .B(new_n711), .ZN(G9));
  NOR2_X1   g526(.A1(new_n241), .A2(KEYINPUT36), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n236), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n714), .A2(new_n257), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n255), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(new_n716), .ZN(new_n717));
  NOR2_X1   g531(.A1(new_n679), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n600), .A2(new_n664), .A3(new_n672), .A4(new_n718), .ZN(new_n719));
  XOR2_X1   g533(.A(KEYINPUT37), .B(G110), .Z(new_n720));
  XNOR2_X1  g534(.A(new_n719), .B(new_n720), .ZN(G12));
  NAND2_X1  g535(.A1(new_n664), .A2(new_n672), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n681), .A2(new_n716), .ZN(new_n723));
  INV_X1    g537(.A(new_n723), .ZN(new_n724));
  INV_X1    g538(.A(G900), .ZN(new_n725));
  AOI21_X1  g539(.A(new_n596), .B1(new_n594), .B2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n726), .ZN(new_n727));
  NAND4_X1  g541(.A1(new_n702), .A2(new_n707), .A3(new_n684), .A4(new_n727), .ZN(new_n728));
  INV_X1    g542(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n381), .B1(new_n380), .B2(new_n383), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n386), .A2(KEYINPUT72), .A3(new_n382), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n354), .A2(new_n357), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT74), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n354), .A2(new_n260), .A3(new_n357), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n362), .B1(new_n378), .B2(new_n341), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n369), .A2(new_n370), .A3(new_n247), .ZN(new_n737));
  OAI21_X1  g551(.A(G472), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n735), .A3(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n724), .B(new_n729), .C1(new_n732), .C2(new_n739), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n722), .A2(new_n740), .ZN(new_n741));
  XNOR2_X1  g555(.A(new_n741), .B(new_n215), .ZN(G30));
  XOR2_X1   g556(.A(KEYINPUT104), .B(KEYINPUT38), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n473), .B(new_n743), .ZN(new_n744));
  NOR3_X1   g558(.A1(new_n744), .A2(new_n476), .A3(new_n716), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n358), .A2(new_n359), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n351), .A2(new_n332), .ZN(new_n747));
  OAI21_X1  g561(.A(new_n247), .B1(new_n320), .B2(new_n341), .ZN(new_n748));
  OAI21_X1  g562(.A(G472), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n388), .A2(new_n746), .A3(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n745), .A2(new_n685), .A3(new_n702), .A4(new_n750), .ZN(new_n751));
  XOR2_X1   g565(.A(new_n726), .B(KEYINPUT39), .Z(new_n752));
  NAND2_X1  g566(.A1(new_n677), .A2(new_n752), .ZN(new_n753));
  AOI21_X1  g567(.A(new_n751), .B1(new_n753), .B2(KEYINPUT40), .ZN(new_n754));
  OAI21_X1  g568(.A(new_n754), .B1(KEYINPUT40), .B2(new_n753), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n755), .B(G143), .ZN(G45));
  AOI21_X1  g570(.A(new_n723), .B1(new_n373), .B2(new_n388), .ZN(new_n757));
  NOR3_X1   g571(.A1(new_n535), .A2(new_n694), .A3(new_n726), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n757), .A2(new_n664), .A3(new_n672), .A4(new_n758), .ZN(new_n759));
  XNOR2_X1  g573(.A(new_n759), .B(G146), .ZN(G48));
  AOI21_X1  g574(.A(new_n601), .B1(new_n668), .B2(new_n247), .ZN(new_n761));
  AOI211_X1 g575(.A(new_n671), .B(new_n761), .C1(new_n665), .C2(new_n669), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n389), .A2(new_n696), .A3(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT105), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g579(.A1(new_n389), .A2(KEYINPUT105), .A3(new_n696), .A4(new_n762), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XOR2_X1   g581(.A(KEYINPUT41), .B(G113), .Z(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(KEYINPUT106), .ZN(new_n769));
  XNOR2_X1  g583(.A(new_n767), .B(new_n769), .ZN(G15));
  NAND2_X1  g584(.A1(new_n373), .A2(new_n388), .ZN(new_n771));
  INV_X1    g585(.A(new_n259), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n771), .A2(new_n709), .A3(new_n772), .A4(new_n762), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT107), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n389), .A2(KEYINPUT107), .A3(new_n709), .A4(new_n762), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G116), .ZN(G18));
  NAND2_X1  g592(.A1(new_n771), .A2(new_n724), .ZN(new_n779));
  INV_X1    g593(.A(new_n599), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n762), .A2(new_n780), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n779), .A2(new_n781), .ZN(new_n782));
  XOR2_X1   g596(.A(new_n782), .B(G119), .Z(G21));
  NOR2_X1   g597(.A1(new_n678), .A2(new_n360), .ZN(new_n784));
  AOI21_X1  g598(.A(new_n341), .B1(new_n311), .B2(new_n365), .ZN(new_n785));
  AOI21_X1  g599(.A(new_n785), .B1(KEYINPUT31), .B2(new_n342), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n385), .B1(new_n786), .B2(new_n353), .ZN(new_n787));
  NOR3_X1   g601(.A1(new_n784), .A2(new_n259), .A3(new_n787), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n762), .A2(new_n598), .A3(new_n788), .ZN(new_n789));
  INV_X1    g603(.A(KEYINPUT108), .ZN(new_n790));
  NAND3_X1  g604(.A1(new_n685), .A2(new_n702), .A3(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(KEYINPUT108), .B1(new_n535), .B2(new_n590), .ZN(new_n792));
  NAND3_X1  g606(.A1(new_n791), .A2(new_n792), .A3(new_n681), .ZN(new_n793));
  NOR2_X1   g607(.A1(new_n789), .A2(new_n793), .ZN(new_n794));
  XNOR2_X1  g608(.A(new_n794), .B(new_n543), .ZN(G24));
  NOR2_X1   g609(.A1(new_n784), .A2(new_n787), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n796), .A2(new_n758), .A3(new_n716), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n761), .B1(new_n665), .B2(new_n669), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n798), .A2(new_n663), .A3(new_n681), .ZN(new_n799));
  NOR2_X1   g613(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(new_n189), .ZN(G27));
  NOR2_X1   g615(.A1(new_n535), .A2(new_n694), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n802), .A2(new_n727), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(KEYINPUT42), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT109), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n665), .A2(new_n669), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n671), .B1(new_n806), .B2(new_n640), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n465), .A2(new_n472), .A3(new_n474), .ZN(new_n808));
  INV_X1    g622(.A(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n805), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n670), .A2(KEYINPUT109), .A3(new_n671), .A4(new_n808), .ZN(new_n811));
  OAI211_X1 g625(.A(new_n389), .B(new_n804), .C1(new_n810), .C2(new_n811), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n733), .B(new_n738), .C1(KEYINPUT32), .C2(new_n386), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n813), .A2(new_n772), .ZN(new_n814));
  INV_X1    g628(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n815), .A2(new_n758), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n809), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(KEYINPUT109), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n807), .A2(new_n805), .A3(new_n809), .ZN(new_n819));
  AOI21_X1  g633(.A(new_n816), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT42), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n812), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XOR2_X1   g636(.A(KEYINPUT110), .B(G131), .Z(new_n823));
  XNOR2_X1  g637(.A(new_n822), .B(new_n823), .ZN(G33));
  OAI211_X1 g638(.A(new_n389), .B(new_n729), .C1(new_n810), .C2(new_n811), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(G134), .ZN(G36));
  INV_X1    g640(.A(KEYINPUT45), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n638), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n638), .A2(new_n827), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n828), .A2(G469), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(G469), .A2(G902), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT46), .ZN(new_n833));
  AOI22_X1  g647(.A1(new_n832), .A2(new_n833), .B1(new_n669), .B2(new_n665), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n834), .B1(new_n833), .B2(new_n832), .ZN(new_n835));
  NAND2_X1  g649(.A1(new_n835), .A2(new_n663), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n535), .A2(new_n691), .ZN(new_n838));
  OR2_X1    g652(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(KEYINPUT43), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n839), .A2(new_n679), .A3(new_n716), .A4(new_n840), .ZN(new_n841));
  INV_X1    g655(.A(KEYINPUT44), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n808), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  OR2_X1    g657(.A1(new_n841), .A2(new_n842), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n837), .A2(new_n752), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  XNOR2_X1  g659(.A(new_n845), .B(G137), .ZN(G39));
  NOR4_X1   g660(.A1(new_n771), .A2(new_n772), .A3(new_n803), .A4(new_n808), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n835), .A2(KEYINPUT47), .A3(new_n663), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT47), .B1(new_n835), .B2(new_n663), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  OR2_X1    g664(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n850), .A2(KEYINPUT111), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g667(.A(new_n853), .B(G140), .ZN(G42));
  XOR2_X1   g668(.A(new_n798), .B(KEYINPUT113), .Z(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT49), .Z(new_n856));
  AND4_X1   g670(.A1(new_n388), .A2(new_n744), .A3(new_n746), .A4(new_n749), .ZN(new_n857));
  NOR4_X1   g671(.A1(new_n838), .A2(new_n259), .A3(new_n671), .A4(new_n476), .ZN(new_n858));
  XNOR2_X1  g672(.A(new_n858), .B(KEYINPUT112), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n857), .A3(new_n859), .ZN(new_n860));
  AOI211_X1 g674(.A(new_n723), .B(new_n728), .C1(new_n373), .C2(new_n388), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n800), .B1(new_n677), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT52), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n791), .A2(new_n792), .A3(new_n681), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n716), .A2(new_n726), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n864), .A2(new_n750), .A3(new_n807), .A4(new_n865), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n862), .A2(new_n863), .A3(new_n759), .A4(new_n866), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n759), .A2(new_n866), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n786), .A2(new_n353), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n355), .ZN(new_n870));
  OAI211_X1 g684(.A(new_n870), .B(new_n716), .C1(new_n360), .C2(new_n678), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n803), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n872), .A2(new_n681), .A3(new_n762), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n873), .B1(new_n722), .B2(new_n740), .ZN(new_n874));
  OAI21_X1  g688(.A(KEYINPUT52), .B1(new_n868), .B2(new_n874), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n867), .A2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(KEYINPUT116), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT116), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n867), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(new_n389), .ZN(new_n881));
  AOI21_X1  g695(.A(new_n881), .B1(new_n818), .B2(new_n819), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n758), .B(new_n815), .C1(new_n810), .C2(new_n811), .ZN(new_n883));
  AOI22_X1  g697(.A1(new_n882), .A2(new_n804), .B1(new_n883), .B2(KEYINPUT42), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n872), .B1(new_n810), .B2(new_n811), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n707), .A2(new_n590), .A3(new_n684), .A4(new_n727), .ZN(new_n886));
  NOR3_X1   g700(.A1(new_n886), .A2(new_n717), .A3(new_n808), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n664), .A2(new_n672), .A3(new_n771), .A4(new_n887), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n825), .A2(new_n885), .A3(new_n888), .ZN(new_n889));
  OAI22_X1  g703(.A1(new_n779), .A2(new_n781), .B1(new_n789), .B2(new_n793), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n890), .B1(new_n765), .B2(new_n766), .ZN(new_n891));
  NAND4_X1  g705(.A1(new_n884), .A2(new_n889), .A3(new_n891), .A4(new_n777), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n473), .A2(new_n474), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(KEYINPUT90), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n685), .A2(new_n590), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n681), .A2(new_n390), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n894), .A2(new_n895), .A3(new_n896), .A4(new_n598), .ZN(new_n897));
  INV_X1    g711(.A(KEYINPUT114), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(new_n475), .A2(new_n477), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n900), .A2(KEYINPUT114), .A3(new_n598), .A4(new_n895), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n664), .A2(new_n680), .A3(new_n672), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n719), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT115), .ZN(new_n905));
  INV_X1    g719(.A(KEYINPUT115), .ZN(new_n906));
  OAI211_X1 g720(.A(new_n906), .B(new_n719), .C1(new_n902), .C2(new_n903), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n894), .A2(new_n896), .A3(new_n598), .A4(new_n802), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n908), .A2(new_n672), .A3(new_n664), .A4(new_n680), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n909), .A2(new_n673), .ZN(new_n910));
  INV_X1    g724(.A(new_n910), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n905), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  NOR2_X1   g726(.A1(new_n892), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n880), .A2(new_n913), .A3(KEYINPUT53), .ZN(new_n914));
  INV_X1    g728(.A(KEYINPUT53), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n825), .A2(new_n885), .A3(new_n888), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n822), .A2(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(new_n890), .ZN(new_n918));
  AND3_X1   g732(.A1(new_n767), .A2(new_n777), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g733(.A(new_n910), .B1(new_n904), .B2(KEYINPUT115), .ZN(new_n920));
  NAND4_X1  g734(.A1(new_n917), .A2(new_n919), .A3(new_n920), .A4(new_n907), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n915), .B1(new_n921), .B2(new_n876), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n914), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n923), .A2(KEYINPUT54), .ZN(new_n924));
  AND3_X1   g738(.A1(new_n867), .A2(new_n878), .A3(new_n875), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n878), .B1(new_n867), .B2(new_n875), .ZN(new_n926));
  NOR2_X1   g740(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n915), .B1(new_n927), .B2(new_n921), .ZN(new_n928));
  XOR2_X1   g742(.A(KEYINPUT117), .B(KEYINPUT54), .Z(new_n929));
  NAND4_X1  g743(.A1(new_n913), .A2(KEYINPUT53), .A3(new_n867), .A4(new_n875), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n924), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g746(.A1(new_n839), .A2(new_n596), .A3(new_n788), .A4(new_n840), .ZN(new_n933));
  NOR2_X1   g747(.A1(new_n933), .A2(new_n808), .ZN(new_n934));
  OR2_X1    g748(.A1(new_n848), .A2(new_n849), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n855), .A2(new_n663), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g751(.A1(new_n762), .A2(new_n744), .A3(new_n476), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n933), .A2(new_n938), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT50), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n839), .A2(new_n840), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n798), .A2(new_n663), .A3(new_n596), .A4(new_n809), .ZN(new_n942));
  OR2_X1    g756(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(new_n943), .A2(new_n871), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n750), .A2(new_n942), .A3(new_n259), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n685), .A2(new_n691), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND4_X1  g761(.A1(new_n937), .A2(KEYINPUT51), .A3(new_n940), .A4(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n933), .A2(new_n799), .ZN(new_n949));
  INV_X1    g763(.A(G952), .ZN(new_n950));
  NOR3_X1   g764(.A1(new_n949), .A2(new_n950), .A3(G953), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n692), .A2(new_n695), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n945), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g767(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OR2_X1    g768(.A1(new_n954), .A2(KEYINPUT119), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT48), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n943), .A2(new_n814), .ZN(new_n957));
  INV_X1    g771(.A(KEYINPUT120), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n956), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n958), .B2(new_n957), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n954), .A2(KEYINPUT119), .ZN(new_n961));
  OAI211_X1 g775(.A(KEYINPUT120), .B(new_n956), .C1(new_n943), .C2(new_n814), .ZN(new_n962));
  AND4_X1   g776(.A1(new_n955), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n947), .A2(new_n940), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n936), .B1(new_n935), .B2(KEYINPUT118), .ZN(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(KEYINPUT118), .B2(new_n935), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n964), .B1(new_n966), .B2(new_n934), .ZN(new_n967));
  OAI211_X1 g781(.A(new_n948), .B(new_n963), .C1(new_n967), .C2(KEYINPUT51), .ZN(new_n968));
  NOR2_X1   g782(.A1(new_n932), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g783(.A1(G952), .A2(G953), .ZN(new_n970));
  OAI21_X1  g784(.A(new_n860), .B1(new_n969), .B2(new_n970), .ZN(G75));
  INV_X1    g785(.A(KEYINPUT56), .ZN(new_n972));
  XNOR2_X1  g786(.A(new_n468), .B(new_n469), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n973), .B(KEYINPUT55), .ZN(new_n974));
  INV_X1    g788(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(KEYINPUT53), .B1(new_n880), .B2(new_n913), .ZN(new_n976));
  NOR3_X1   g790(.A1(new_n921), .A2(new_n915), .A3(new_n876), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g792(.A1(G210), .A2(G902), .ZN(new_n979));
  OAI211_X1 g793(.A(new_n972), .B(new_n975), .C1(new_n978), .C2(new_n979), .ZN(new_n980));
  NOR2_X1   g794(.A1(new_n237), .A2(G952), .ZN(new_n981));
  INV_X1    g795(.A(new_n981), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g797(.A(KEYINPUT121), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n928), .A2(new_n930), .ZN(new_n985));
  INV_X1    g799(.A(new_n979), .ZN(new_n986));
  AOI21_X1  g800(.A(KEYINPUT56), .B1(new_n985), .B2(new_n986), .ZN(new_n987));
  OAI21_X1  g801(.A(new_n984), .B1(new_n987), .B2(new_n975), .ZN(new_n988));
  OAI21_X1  g802(.A(new_n972), .B1(new_n978), .B2(new_n979), .ZN(new_n989));
  NAND3_X1  g803(.A1(new_n989), .A2(KEYINPUT121), .A3(new_n974), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n983), .B1(new_n988), .B2(new_n990), .ZN(G51));
  XOR2_X1   g805(.A(new_n831), .B(KEYINPUT57), .Z(new_n992));
  INV_X1    g806(.A(new_n929), .ZN(new_n993));
  NOR3_X1   g807(.A1(new_n976), .A2(new_n977), .A3(new_n993), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n929), .B1(new_n928), .B2(new_n930), .ZN(new_n995));
  OAI21_X1  g809(.A(new_n992), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(new_n668), .ZN(new_n997));
  OR3_X1    g811(.A1(new_n978), .A2(new_n247), .A3(new_n830), .ZN(new_n998));
  AOI21_X1  g812(.A(new_n981), .B1(new_n997), .B2(new_n998), .ZN(G54));
  AND2_X1   g813(.A1(KEYINPUT58), .A2(G475), .ZN(new_n1000));
  NAND3_X1  g814(.A1(new_n985), .A2(G902), .A3(new_n1000), .ZN(new_n1001));
  AND2_X1   g815(.A1(new_n1001), .A2(new_n528), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1001), .A2(new_n528), .ZN(new_n1003));
  NOR3_X1   g817(.A1(new_n1002), .A2(new_n1003), .A3(new_n981), .ZN(G60));
  NAND2_X1  g818(.A1(new_n687), .A2(new_n688), .ZN(new_n1005));
  XNOR2_X1  g819(.A(KEYINPUT122), .B(KEYINPUT59), .ZN(new_n1006));
  NOR2_X1   g820(.A1(new_n536), .A2(new_n247), .ZN(new_n1007));
  XOR2_X1   g821(.A(new_n1006), .B(new_n1007), .Z(new_n1008));
  NOR2_X1   g822(.A1(new_n1005), .A2(new_n1008), .ZN(new_n1009));
  OAI21_X1  g823(.A(new_n1009), .B1(new_n994), .B2(new_n995), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n1010), .A2(new_n982), .ZN(new_n1011));
  INV_X1    g825(.A(new_n1005), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1008), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1012), .B1(new_n932), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n1011), .A2(new_n1014), .ZN(G63));
  NAND2_X1  g829(.A1(G217), .A2(G902), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1016), .B(KEYINPUT60), .ZN(new_n1017));
  OAI211_X1 g831(.A(new_n244), .B(new_n243), .C1(new_n978), .C2(new_n1017), .ZN(new_n1018));
  INV_X1    g832(.A(new_n1017), .ZN(new_n1019));
  OAI211_X1 g833(.A(new_n714), .B(new_n1019), .C1(new_n976), .C2(new_n977), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n1018), .A2(KEYINPUT61), .A3(new_n982), .A4(new_n1020), .ZN(new_n1021));
  AOI21_X1  g835(.A(new_n1017), .B1(new_n928), .B2(new_n930), .ZN(new_n1022));
  OAI211_X1 g836(.A(new_n1020), .B(new_n982), .C1(new_n1022), .C2(new_n256), .ZN(new_n1023));
  INV_X1    g837(.A(KEYINPUT61), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n1021), .A2(new_n1025), .ZN(G66));
  OAI21_X1  g840(.A(G953), .B1(new_n592), .B2(new_n441), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n919), .A2(new_n907), .A3(new_n920), .ZN(new_n1028));
  INV_X1    g842(.A(new_n1028), .ZN(new_n1029));
  OAI21_X1  g843(.A(new_n1027), .B1(new_n1029), .B2(G953), .ZN(new_n1030));
  OAI211_X1 g844(.A(new_n434), .B(new_n440), .C1(G898), .C2(new_n237), .ZN(new_n1031));
  XNOR2_X1  g845(.A(new_n1031), .B(KEYINPUT123), .ZN(new_n1032));
  XNOR2_X1  g846(.A(new_n1032), .B(KEYINPUT124), .ZN(new_n1033));
  XNOR2_X1  g847(.A(new_n1030), .B(new_n1033), .ZN(G69));
  XOR2_X1   g848(.A(new_n350), .B(KEYINPUT125), .Z(new_n1035));
  XNOR2_X1  g849(.A(new_n1035), .B(new_n521), .ZN(new_n1036));
  NAND4_X1  g850(.A1(new_n837), .A2(new_n752), .A3(new_n864), .A4(new_n815), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n845), .A2(new_n1037), .A3(new_n825), .ZN(new_n1038));
  AND2_X1   g852(.A1(new_n862), .A2(new_n759), .ZN(new_n1039));
  NAND4_X1  g853(.A1(new_n853), .A2(new_n884), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n237), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n603), .A2(G900), .A3(G953), .ZN(new_n1042));
  AOI21_X1  g856(.A(new_n1036), .B1(new_n1041), .B2(new_n1042), .ZN(new_n1043));
  NAND3_X1  g857(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n1044));
  OAI211_X1 g858(.A(new_n389), .B(new_n809), .C1(new_n802), .C2(new_n895), .ZN(new_n1045));
  OAI21_X1  g859(.A(new_n845), .B1(new_n753), .B2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g860(.A(new_n1046), .B1(new_n851), .B2(new_n852), .ZN(new_n1047));
  AND2_X1   g861(.A1(new_n755), .A2(new_n1039), .ZN(new_n1048));
  INV_X1    g862(.A(KEYINPUT62), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1047), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g864(.A1(new_n1048), .A2(new_n1049), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n237), .ZN(new_n1052));
  OAI21_X1  g866(.A(new_n1044), .B1(new_n1050), .B2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1043), .B1(new_n1053), .B2(new_n1036), .ZN(G72));
  XNOR2_X1  g868(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n1055));
  NOR2_X1   g869(.A1(new_n360), .A2(new_n247), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1055), .B(new_n1056), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT127), .ZN(new_n1058));
  OAI21_X1  g872(.A(new_n1058), .B1(new_n1040), .B2(new_n1028), .ZN(new_n1059));
  NAND2_X1  g873(.A1(new_n351), .A2(new_n332), .ZN(new_n1060));
  INV_X1    g874(.A(new_n1060), .ZN(new_n1061));
  AOI21_X1  g875(.A(new_n981), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g876(.A1(new_n1051), .A2(new_n1029), .ZN(new_n1063));
  OAI21_X1  g877(.A(new_n1058), .B1(new_n1050), .B2(new_n1063), .ZN(new_n1064));
  NAND2_X1  g878(.A1(new_n1064), .A2(new_n747), .ZN(new_n1065));
  INV_X1    g879(.A(new_n747), .ZN(new_n1066));
  NAND4_X1  g880(.A1(new_n923), .A2(new_n1066), .A3(new_n1060), .A4(new_n1057), .ZN(new_n1067));
  AND3_X1   g881(.A1(new_n1062), .A2(new_n1065), .A3(new_n1067), .ZN(G57));
endmodule


