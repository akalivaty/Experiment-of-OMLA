

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587;

  XNOR2_X1 U325 ( .A(G29GAT), .B(KEYINPUT7), .ZN(n296) );
  XNOR2_X1 U326 ( .A(n306), .B(n305), .ZN(n308) );
  XNOR2_X1 U327 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U328 ( .A(KEYINPUT45), .B(n339), .Z(n293) );
  XOR2_X1 U329 ( .A(n309), .B(KEYINPUT67), .Z(n294) );
  XOR2_X1 U330 ( .A(G92GAT), .B(G85GAT), .Z(n295) );
  INV_X1 U331 ( .A(KEYINPUT96), .ZN(n453) );
  XNOR2_X1 U332 ( .A(n453), .B(KEYINPUT25), .ZN(n454) );
  XNOR2_X1 U333 ( .A(n455), .B(n454), .ZN(n459) );
  INV_X1 U334 ( .A(KEYINPUT18), .ZN(n373) );
  XNOR2_X1 U335 ( .A(n374), .B(n373), .ZN(n375) );
  XNOR2_X1 U336 ( .A(n376), .B(n375), .ZN(n445) );
  XNOR2_X1 U337 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U338 ( .A(n317), .B(n316), .ZN(n323) );
  XOR2_X1 U339 ( .A(KEYINPUT41), .B(n574), .Z(n542) );
  INV_X1 U340 ( .A(G106GAT), .ZN(n474) );
  XNOR2_X1 U341 ( .A(n384), .B(n383), .ZN(n516) );
  XNOR2_X1 U342 ( .A(n449), .B(KEYINPUT58), .ZN(n450) );
  XNOR2_X1 U343 ( .A(n474), .B(KEYINPUT44), .ZN(n475) );
  XNOR2_X1 U344 ( .A(n451), .B(n450), .ZN(G1351GAT) );
  XOR2_X1 U345 ( .A(G36GAT), .B(G190GAT), .Z(n382) );
  XNOR2_X1 U346 ( .A(n296), .B(KEYINPUT8), .ZN(n343) );
  XNOR2_X1 U347 ( .A(n382), .B(n343), .ZN(n298) );
  AND2_X1 U348 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U349 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U350 ( .A(KEYINPUT11), .B(n299), .Z(n306) );
  XNOR2_X1 U351 ( .A(G99GAT), .B(G106GAT), .ZN(n300) );
  XNOR2_X1 U352 ( .A(n295), .B(n300), .ZN(n309) );
  XNOR2_X1 U353 ( .A(n309), .B(KEYINPUT9), .ZN(n304) );
  XOR2_X1 U354 ( .A(KEYINPUT10), .B(KEYINPUT71), .Z(n302) );
  XNOR2_X1 U355 ( .A(G218GAT), .B(KEYINPUT72), .ZN(n301) );
  XOR2_X1 U356 ( .A(n302), .B(n301), .Z(n303) );
  XOR2_X1 U357 ( .A(G43GAT), .B(G134GAT), .Z(n430) );
  XOR2_X1 U358 ( .A(G50GAT), .B(G162GAT), .Z(n410) );
  XNOR2_X1 U359 ( .A(n430), .B(n410), .ZN(n307) );
  XNOR2_X1 U360 ( .A(n308), .B(n307), .ZN(n550) );
  NAND2_X1 U361 ( .A1(G230GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n294), .B(n310), .ZN(n311) );
  XNOR2_X1 U363 ( .A(n311), .B(KEYINPUT33), .ZN(n317) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G148GAT), .Z(n399) );
  XOR2_X1 U365 ( .A(n399), .B(KEYINPUT31), .Z(n315) );
  XOR2_X1 U366 ( .A(KEYINPUT32), .B(KEYINPUT70), .Z(n313) );
  XNOR2_X1 U367 ( .A(KEYINPUT66), .B(KEYINPUT68), .ZN(n312) );
  XOR2_X1 U368 ( .A(n313), .B(n312), .Z(n314) );
  XOR2_X1 U369 ( .A(G64GAT), .B(KEYINPUT69), .Z(n319) );
  XNOR2_X1 U370 ( .A(G176GAT), .B(G204GAT), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n369) );
  XOR2_X1 U372 ( .A(KEYINPUT13), .B(G57GAT), .Z(n321) );
  XNOR2_X1 U373 ( .A(G71GAT), .B(G78GAT), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n336) );
  XNOR2_X1 U375 ( .A(n369), .B(n336), .ZN(n322) );
  XNOR2_X1 U376 ( .A(n323), .B(n322), .ZN(n574) );
  XOR2_X1 U377 ( .A(G8GAT), .B(G183GAT), .Z(n367) );
  XOR2_X1 U378 ( .A(G22GAT), .B(G155GAT), .Z(n411) );
  XOR2_X1 U379 ( .A(n367), .B(n411), .Z(n325) );
  NAND2_X1 U380 ( .A1(G231GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U382 ( .A(KEYINPUT14), .B(KEYINPUT76), .Z(n327) );
  XNOR2_X1 U383 ( .A(KEYINPUT15), .B(KEYINPUT75), .ZN(n326) );
  XNOR2_X1 U384 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U385 ( .A(n329), .B(n328), .Z(n334) );
  XOR2_X1 U386 ( .A(G15GAT), .B(G1GAT), .Z(n344) );
  XOR2_X1 U387 ( .A(KEYINPUT73), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U388 ( .A(G127GAT), .B(G211GAT), .ZN(n330) );
  XNOR2_X1 U389 ( .A(n331), .B(n330), .ZN(n332) );
  XNOR2_X1 U390 ( .A(n344), .B(n332), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n335) );
  XOR2_X1 U392 ( .A(n335), .B(KEYINPUT12), .Z(n338) );
  XNOR2_X1 U393 ( .A(n336), .B(KEYINPUT74), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n338), .B(n337), .ZN(n577) );
  INV_X1 U395 ( .A(n577), .ZN(n470) );
  XNOR2_X1 U396 ( .A(n550), .B(KEYINPUT36), .ZN(n584) );
  NOR2_X1 U397 ( .A1(n470), .A2(n584), .ZN(n339) );
  NOR2_X1 U398 ( .A1(n574), .A2(n293), .ZN(n340) );
  XNOR2_X1 U399 ( .A(n340), .B(KEYINPUT111), .ZN(n358) );
  XOR2_X1 U400 ( .A(G197GAT), .B(G113GAT), .Z(n342) );
  XNOR2_X1 U401 ( .A(G169GAT), .B(G50GAT), .ZN(n341) );
  XNOR2_X1 U402 ( .A(n342), .B(n341), .ZN(n357) );
  XOR2_X1 U403 ( .A(n344), .B(n343), .Z(n346) );
  XNOR2_X1 U404 ( .A(G36GAT), .B(G43GAT), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n350) );
  XOR2_X1 U406 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n348) );
  NAND2_X1 U407 ( .A1(G229GAT), .A2(G233GAT), .ZN(n347) );
  XNOR2_X1 U408 ( .A(n348), .B(n347), .ZN(n349) );
  XOR2_X1 U409 ( .A(n350), .B(n349), .Z(n355) );
  XOR2_X1 U410 ( .A(KEYINPUT64), .B(G8GAT), .Z(n352) );
  XNOR2_X1 U411 ( .A(G141GAT), .B(G22GAT), .ZN(n351) );
  XNOR2_X1 U412 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n353), .B(KEYINPUT65), .ZN(n354) );
  XNOR2_X1 U414 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U415 ( .A(n357), .B(n356), .Z(n553) );
  INV_X1 U416 ( .A(n553), .ZN(n570) );
  NOR2_X1 U417 ( .A1(n358), .A2(n570), .ZN(n359) );
  XNOR2_X1 U418 ( .A(n359), .B(KEYINPUT112), .ZN(n365) );
  XNOR2_X1 U419 ( .A(KEYINPUT110), .B(n577), .ZN(n561) );
  NAND2_X1 U420 ( .A1(n542), .A2(n570), .ZN(n360) );
  XNOR2_X1 U421 ( .A(KEYINPUT46), .B(n360), .ZN(n361) );
  NAND2_X1 U422 ( .A1(n361), .A2(n550), .ZN(n362) );
  NOR2_X1 U423 ( .A1(n561), .A2(n362), .ZN(n363) );
  XOR2_X1 U424 ( .A(KEYINPUT47), .B(n363), .Z(n364) );
  NOR2_X1 U425 ( .A1(n365), .A2(n364), .ZN(n366) );
  XNOR2_X1 U426 ( .A(KEYINPUT48), .B(n366), .ZN(n522) );
  XNOR2_X1 U427 ( .A(G92GAT), .B(KEYINPUT92), .ZN(n368) );
  XNOR2_X1 U428 ( .A(n368), .B(n367), .ZN(n370) );
  XOR2_X1 U429 ( .A(n370), .B(n369), .Z(n380) );
  XOR2_X1 U430 ( .A(KEYINPUT79), .B(KEYINPUT19), .Z(n372) );
  XNOR2_X1 U431 ( .A(KEYINPUT81), .B(KEYINPUT17), .ZN(n371) );
  XNOR2_X1 U432 ( .A(n372), .B(n371), .ZN(n376) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(KEYINPUT80), .ZN(n374) );
  XOR2_X1 U434 ( .A(G211GAT), .B(KEYINPUT21), .Z(n378) );
  XNOR2_X1 U435 ( .A(G197GAT), .B(G218GAT), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n413) );
  XNOR2_X1 U437 ( .A(n445), .B(n413), .ZN(n379) );
  XOR2_X1 U438 ( .A(n380), .B(n379), .Z(n381) );
  XNOR2_X1 U439 ( .A(n382), .B(n381), .ZN(n384) );
  NAND2_X1 U440 ( .A1(G226GAT), .A2(G233GAT), .ZN(n383) );
  NOR2_X1 U441 ( .A1(n522), .A2(n516), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n385), .B(KEYINPUT54), .ZN(n566) );
  XOR2_X1 U443 ( .A(KEYINPUT5), .B(KEYINPUT6), .Z(n387) );
  XNOR2_X1 U444 ( .A(G57GAT), .B(KEYINPUT91), .ZN(n386) );
  XNOR2_X1 U445 ( .A(n387), .B(n386), .ZN(n391) );
  XOR2_X1 U446 ( .A(KEYINPUT1), .B(KEYINPUT87), .Z(n389) );
  XNOR2_X1 U447 ( .A(KEYINPUT86), .B(KEYINPUT4), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XOR2_X1 U449 ( .A(n391), .B(n390), .Z(n396) );
  XOR2_X1 U450 ( .A(KEYINPUT88), .B(KEYINPUT90), .Z(n393) );
  NAND2_X1 U451 ( .A1(G225GAT), .A2(G233GAT), .ZN(n392) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n394) );
  XNOR2_X1 U453 ( .A(KEYINPUT89), .B(n394), .ZN(n395) );
  XNOR2_X1 U454 ( .A(n396), .B(n395), .ZN(n404) );
  XOR2_X1 U455 ( .A(G85GAT), .B(G155GAT), .Z(n398) );
  XNOR2_X1 U456 ( .A(G1GAT), .B(G134GAT), .ZN(n397) );
  XNOR2_X1 U457 ( .A(n398), .B(n397), .ZN(n400) );
  XOR2_X1 U458 ( .A(n400), .B(n399), .Z(n402) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(G162GAT), .ZN(n401) );
  XNOR2_X1 U460 ( .A(n402), .B(n401), .ZN(n403) );
  XOR2_X1 U461 ( .A(n404), .B(n403), .Z(n408) );
  XNOR2_X1 U462 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n405) );
  XNOR2_X1 U463 ( .A(n405), .B(G127GAT), .ZN(n431) );
  XNOR2_X1 U464 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n406) );
  XNOR2_X1 U465 ( .A(n406), .B(KEYINPUT2), .ZN(n409) );
  XNOR2_X1 U466 ( .A(n431), .B(n409), .ZN(n407) );
  XNOR2_X1 U467 ( .A(n408), .B(n407), .ZN(n565) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n412) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n417) );
  XOR2_X1 U470 ( .A(G78GAT), .B(n413), .Z(n415) );
  NAND2_X1 U471 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U473 ( .A(n417), .B(n416), .Z(n425) );
  XOR2_X1 U474 ( .A(KEYINPUT23), .B(G148GAT), .Z(n419) );
  XNOR2_X1 U475 ( .A(G106GAT), .B(G204GAT), .ZN(n418) );
  XNOR2_X1 U476 ( .A(n419), .B(n418), .ZN(n423) );
  XOR2_X1 U477 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n421) );
  XNOR2_X1 U478 ( .A(KEYINPUT84), .B(KEYINPUT85), .ZN(n420) );
  XNOR2_X1 U479 ( .A(n421), .B(n420), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U481 ( .A(n425), .B(n424), .ZN(n456) );
  INV_X1 U482 ( .A(n456), .ZN(n426) );
  AND2_X1 U483 ( .A1(n565), .A2(n426), .ZN(n427) );
  AND2_X1 U484 ( .A1(n566), .A2(n427), .ZN(n429) );
  XNOR2_X1 U485 ( .A(KEYINPUT55), .B(KEYINPUT119), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n429), .B(n428), .ZN(n448) );
  XOR2_X1 U487 ( .A(n431), .B(n430), .Z(n433) );
  NAND2_X1 U488 ( .A1(G227GAT), .A2(G233GAT), .ZN(n432) );
  XNOR2_X1 U489 ( .A(n433), .B(n432), .ZN(n447) );
  XOR2_X1 U490 ( .A(KEYINPUT82), .B(KEYINPUT83), .Z(n435) );
  XNOR2_X1 U491 ( .A(G190GAT), .B(G99GAT), .ZN(n434) );
  XNOR2_X1 U492 ( .A(n435), .B(n434), .ZN(n443) );
  XOR2_X1 U493 ( .A(G120GAT), .B(G176GAT), .Z(n437) );
  XNOR2_X1 U494 ( .A(G15GAT), .B(KEYINPUT77), .ZN(n436) );
  XNOR2_X1 U495 ( .A(n437), .B(n436), .ZN(n441) );
  XOR2_X1 U496 ( .A(G71GAT), .B(G183GAT), .Z(n439) );
  XNOR2_X1 U497 ( .A(KEYINPUT78), .B(KEYINPUT20), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n439), .B(n438), .ZN(n440) );
  XOR2_X1 U499 ( .A(n441), .B(n440), .Z(n442) );
  XNOR2_X1 U500 ( .A(n443), .B(n442), .ZN(n444) );
  XOR2_X1 U501 ( .A(n445), .B(n444), .Z(n446) );
  XNOR2_X1 U502 ( .A(n447), .B(n446), .ZN(n524) );
  NAND2_X1 U503 ( .A1(n448), .A2(n524), .ZN(n560) );
  NOR2_X1 U504 ( .A1(n550), .A2(n560), .ZN(n451) );
  INV_X1 U505 ( .A(G190GAT), .ZN(n449) );
  XOR2_X1 U506 ( .A(n456), .B(KEYINPUT28), .Z(n511) );
  INV_X1 U507 ( .A(n524), .ZN(n519) );
  NOR2_X1 U508 ( .A1(n516), .A2(n519), .ZN(n452) );
  NOR2_X1 U509 ( .A1(n456), .A2(n452), .ZN(n455) );
  NAND2_X1 U510 ( .A1(n519), .A2(n456), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n457), .B(KEYINPUT26), .ZN(n567) );
  XNOR2_X1 U512 ( .A(n516), .B(KEYINPUT27), .ZN(n463) );
  NOR2_X1 U513 ( .A1(n567), .A2(n463), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n459), .A2(n458), .ZN(n460) );
  XNOR2_X1 U515 ( .A(n460), .B(KEYINPUT97), .ZN(n461) );
  NAND2_X1 U516 ( .A1(n461), .A2(n565), .ZN(n462) );
  XOR2_X1 U517 ( .A(KEYINPUT98), .B(n462), .Z(n469) );
  INV_X1 U518 ( .A(KEYINPUT95), .ZN(n467) );
  NOR2_X1 U519 ( .A1(n565), .A2(n463), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT93), .B(n464), .Z(n540) );
  NAND2_X1 U521 ( .A1(n540), .A2(n511), .ZN(n523) );
  XNOR2_X1 U522 ( .A(KEYINPUT94), .B(n523), .ZN(n465) );
  NOR2_X1 U523 ( .A1(n465), .A2(n524), .ZN(n466) );
  XNOR2_X1 U524 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n469), .A2(n468), .ZN(n479) );
  NOR2_X1 U526 ( .A1(n479), .A2(n584), .ZN(n471) );
  NAND2_X1 U527 ( .A1(n471), .A2(n470), .ZN(n472) );
  XNOR2_X1 U528 ( .A(n472), .B(KEYINPUT37), .ZN(n489) );
  XOR2_X1 U529 ( .A(n542), .B(KEYINPUT104), .Z(n555) );
  NOR2_X1 U530 ( .A1(n555), .A2(n570), .ZN(n503) );
  NAND2_X1 U531 ( .A1(n489), .A2(n503), .ZN(n473) );
  XNOR2_X1 U532 ( .A(n473), .B(KEYINPUT108), .ZN(n520) );
  NOR2_X1 U533 ( .A1(n511), .A2(n520), .ZN(n476) );
  XNOR2_X1 U534 ( .A(n476), .B(n475), .ZN(G1339GAT) );
  NOR2_X1 U535 ( .A1(n553), .A2(n574), .ZN(n490) );
  NAND2_X1 U536 ( .A1(n550), .A2(n577), .ZN(n477) );
  XNOR2_X1 U537 ( .A(KEYINPUT16), .B(n477), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n479), .A2(n478), .ZN(n502) );
  NAND2_X1 U539 ( .A1(n490), .A2(n502), .ZN(n485) );
  NOR2_X1 U540 ( .A1(n565), .A2(n485), .ZN(n480) );
  XOR2_X1 U541 ( .A(KEYINPUT34), .B(n480), .Z(n481) );
  XNOR2_X1 U542 ( .A(G1GAT), .B(n481), .ZN(G1324GAT) );
  NOR2_X1 U543 ( .A1(n516), .A2(n485), .ZN(n482) );
  XOR2_X1 U544 ( .A(G8GAT), .B(n482), .Z(G1325GAT) );
  NOR2_X1 U545 ( .A1(n519), .A2(n485), .ZN(n484) );
  XNOR2_X1 U546 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n483) );
  XNOR2_X1 U547 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NOR2_X1 U548 ( .A1(n511), .A2(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n486) );
  XNOR2_X1 U550 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U551 ( .A(G22GAT), .B(n488), .ZN(G1327GAT) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n494) );
  XOR2_X1 U553 ( .A(KEYINPUT38), .B(KEYINPUT101), .Z(n492) );
  NAND2_X1 U554 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U555 ( .A(n492), .B(n491), .ZN(n500) );
  NOR2_X1 U556 ( .A1(n565), .A2(n500), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NOR2_X1 U558 ( .A1(n516), .A2(n500), .ZN(n495) );
  XOR2_X1 U559 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT40), .B(KEYINPUT103), .Z(n497) );
  XNOR2_X1 U561 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(n499) );
  NOR2_X1 U563 ( .A1(n500), .A2(n519), .ZN(n498) );
  XOR2_X1 U564 ( .A(n499), .B(n498), .Z(G1330GAT) );
  NOR2_X1 U565 ( .A1(n511), .A2(n500), .ZN(n501) );
  XOR2_X1 U566 ( .A(G50GAT), .B(n501), .Z(G1331GAT) );
  NAND2_X1 U567 ( .A1(n503), .A2(n502), .ZN(n510) );
  NOR2_X1 U568 ( .A1(n565), .A2(n510), .ZN(n505) );
  XNOR2_X1 U569 ( .A(KEYINPUT105), .B(KEYINPUT42), .ZN(n504) );
  XNOR2_X1 U570 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(n506), .ZN(G1332GAT) );
  NOR2_X1 U572 ( .A1(n516), .A2(n510), .ZN(n507) );
  XOR2_X1 U573 ( .A(KEYINPUT106), .B(n507), .Z(n508) );
  XNOR2_X1 U574 ( .A(G64GAT), .B(n508), .ZN(G1333GAT) );
  NOR2_X1 U575 ( .A1(n519), .A2(n510), .ZN(n509) );
  XOR2_X1 U576 ( .A(G71GAT), .B(n509), .Z(G1334GAT) );
  NOR2_X1 U577 ( .A1(n511), .A2(n510), .ZN(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U580 ( .A(G78GAT), .B(n514), .Z(G1335GAT) );
  NOR2_X1 U581 ( .A1(n565), .A2(n520), .ZN(n515) );
  XOR2_X1 U582 ( .A(G85GAT), .B(n515), .Z(G1336GAT) );
  XNOR2_X1 U583 ( .A(G92GAT), .B(KEYINPUT109), .ZN(n518) );
  NOR2_X1 U584 ( .A1(n520), .A2(n516), .ZN(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n520), .A2(n519), .ZN(n521) );
  XOR2_X1 U587 ( .A(G99GAT), .B(n521), .Z(G1338GAT) );
  NOR2_X1 U588 ( .A1(n522), .A2(n523), .ZN(n525) );
  NAND2_X1 U589 ( .A1(n525), .A2(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n526), .B(KEYINPUT113), .ZN(n532) );
  NAND2_X1 U591 ( .A1(n570), .A2(n532), .ZN(n527) );
  XNOR2_X1 U592 ( .A(n527), .B(G113GAT), .ZN(G1340GAT) );
  INV_X1 U593 ( .A(n532), .ZN(n535) );
  NOR2_X1 U594 ( .A1(n535), .A2(n555), .ZN(n531) );
  XOR2_X1 U595 ( .A(KEYINPUT114), .B(KEYINPUT115), .Z(n529) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT49), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n561), .A2(n532), .ZN(n533) );
  XNOR2_X1 U600 ( .A(n533), .B(KEYINPUT50), .ZN(n534) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n534), .ZN(G1342GAT) );
  NOR2_X1 U602 ( .A1(n550), .A2(n535), .ZN(n537) );
  XNOR2_X1 U603 ( .A(KEYINPUT51), .B(KEYINPUT116), .ZN(n536) );
  XNOR2_X1 U604 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U605 ( .A(G134GAT), .B(n538), .ZN(G1343GAT) );
  NOR2_X1 U606 ( .A1(n567), .A2(n522), .ZN(n539) );
  NAND2_X1 U607 ( .A1(n540), .A2(n539), .ZN(n549) );
  NOR2_X1 U608 ( .A1(n553), .A2(n549), .ZN(n541) );
  XOR2_X1 U609 ( .A(G141GAT), .B(n541), .Z(G1344GAT) );
  XOR2_X1 U610 ( .A(G148GAT), .B(KEYINPUT117), .Z(n544) );
  INV_X1 U611 ( .A(n549), .ZN(n547) );
  NAND2_X1 U612 ( .A1(n547), .A2(n542), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n546) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  XNOR2_X1 U615 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NAND2_X1 U616 ( .A1(n547), .A2(n577), .ZN(n548) );
  XNOR2_X1 U617 ( .A(n548), .B(G155GAT), .ZN(G1346GAT) );
  NOR2_X1 U618 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U619 ( .A(KEYINPUT118), .B(n551), .Z(n552) );
  XNOR2_X1 U620 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  NOR2_X1 U621 ( .A1(n553), .A2(n560), .ZN(n554) );
  XOR2_X1 U622 ( .A(G169GAT), .B(n554), .Z(G1348GAT) );
  XNOR2_X1 U623 ( .A(KEYINPUT57), .B(KEYINPUT120), .ZN(n559) );
  NOR2_X1 U624 ( .A1(n555), .A2(n560), .ZN(n557) );
  XNOR2_X1 U625 ( .A(G176GAT), .B(KEYINPUT56), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n557), .B(n556), .ZN(n558) );
  XNOR2_X1 U627 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  XOR2_X1 U628 ( .A(G183GAT), .B(KEYINPUT121), .Z(n564) );
  INV_X1 U629 ( .A(n560), .ZN(n562) );
  NAND2_X1 U630 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1350GAT) );
  XOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n572) );
  NAND2_X1 U633 ( .A1(n566), .A2(n565), .ZN(n568) );
  NOR2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(KEYINPUT122), .ZN(n583) );
  NAND2_X1 U636 ( .A1(n583), .A2(n570), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  XOR2_X1 U639 ( .A(G204GAT), .B(KEYINPUT61), .Z(n576) );
  NAND2_X1 U640 ( .A1(n574), .A2(n583), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n579) );
  NAND2_X1 U643 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n582) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(n587) );
  INV_X1 U649 ( .A(n583), .ZN(n585) );
  NOR2_X1 U650 ( .A1(n585), .A2(n584), .ZN(n586) );
  XOR2_X1 U651 ( .A(n587), .B(n586), .Z(G1355GAT) );
endmodule

