

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586;

  AND2_X1 U320 ( .A1(G232GAT), .A2(G233GAT), .ZN(n288) );
  XNOR2_X1 U321 ( .A(n413), .B(n288), .ZN(n414) );
  INV_X1 U322 ( .A(KEYINPUT48), .ZN(n435) );
  XNOR2_X1 U323 ( .A(KEYINPUT54), .B(KEYINPUT124), .ZN(n452) );
  XNOR2_X1 U324 ( .A(n435), .B(KEYINPUT120), .ZN(n436) );
  XNOR2_X1 U325 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U326 ( .A(n437), .B(n436), .ZN(n534) );
  NOR2_X1 U327 ( .A1(n536), .A2(n456), .ZN(n568) );
  XOR2_X1 U328 ( .A(n469), .B(KEYINPUT28), .Z(n539) );
  XNOR2_X1 U329 ( .A(n457), .B(G176GAT), .ZN(n458) );
  XNOR2_X1 U330 ( .A(n459), .B(n458), .ZN(G1349GAT) );
  XOR2_X1 U331 ( .A(KEYINPUT86), .B(KEYINPUT88), .Z(n290) );
  XNOR2_X1 U332 ( .A(G169GAT), .B(KEYINPUT20), .ZN(n289) );
  XNOR2_X1 U333 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U334 ( .A(G120GAT), .B(G71GAT), .Z(n353) );
  XOR2_X1 U335 ( .A(G99GAT), .B(n353), .Z(n292) );
  XOR2_X1 U336 ( .A(G190GAT), .B(G134GAT), .Z(n413) );
  XNOR2_X1 U337 ( .A(G43GAT), .B(n413), .ZN(n291) );
  XNOR2_X1 U338 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U339 ( .A(n294), .B(n293), .Z(n296) );
  NAND2_X1 U340 ( .A1(G227GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U341 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U342 ( .A(n297), .B(G176GAT), .Z(n300) );
  XNOR2_X1 U343 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n298), .B(G127GAT), .ZN(n337) );
  XNOR2_X1 U345 ( .A(G15GAT), .B(n337), .ZN(n299) );
  XNOR2_X1 U346 ( .A(n300), .B(n299), .ZN(n304) );
  XOR2_X1 U347 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n302) );
  XNOR2_X1 U348 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n301) );
  XNOR2_X1 U349 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U350 ( .A(KEYINPUT17), .B(n303), .ZN(n450) );
  XNOR2_X1 U351 ( .A(n304), .B(n450), .ZN(n536) );
  XOR2_X1 U352 ( .A(KEYINPUT91), .B(G204GAT), .Z(n306) );
  XNOR2_X1 U353 ( .A(G197GAT), .B(G211GAT), .ZN(n305) );
  XNOR2_X1 U354 ( .A(n306), .B(n305), .ZN(n308) );
  XOR2_X1 U355 ( .A(KEYINPUT92), .B(KEYINPUT21), .Z(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n445) );
  XOR2_X1 U357 ( .A(KEYINPUT90), .B(KEYINPUT22), .Z(n310) );
  XNOR2_X1 U358 ( .A(G50GAT), .B(G106GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U360 ( .A(KEYINPUT23), .B(KEYINPUT94), .Z(n312) );
  XNOR2_X1 U361 ( .A(KEYINPUT89), .B(KEYINPUT24), .ZN(n311) );
  XNOR2_X1 U362 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U363 ( .A(n314), .B(n313), .Z(n319) );
  XOR2_X1 U364 ( .A(G141GAT), .B(G22GAT), .Z(n371) );
  XOR2_X1 U365 ( .A(G218GAT), .B(G162GAT), .Z(n417) );
  XOR2_X1 U366 ( .A(G148GAT), .B(G78GAT), .Z(n352) );
  XOR2_X1 U367 ( .A(n417), .B(n352), .Z(n316) );
  NAND2_X1 U368 ( .A1(G228GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U369 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n371), .B(n317), .ZN(n318) );
  XNOR2_X1 U371 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U372 ( .A(n320), .B(KEYINPUT96), .Z(n324) );
  XOR2_X1 U373 ( .A(G155GAT), .B(KEYINPUT3), .Z(n322) );
  XNOR2_X1 U374 ( .A(KEYINPUT2), .B(KEYINPUT93), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n326) );
  XNOR2_X1 U376 ( .A(n326), .B(KEYINPUT95), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n445), .B(n325), .ZN(n469) );
  XOR2_X1 U379 ( .A(n326), .B(KEYINPUT4), .Z(n328) );
  NAND2_X1 U380 ( .A1(G225GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U381 ( .A(n328), .B(n327), .ZN(n332) );
  XOR2_X1 U382 ( .A(G57GAT), .B(KEYINPUT6), .Z(n330) );
  XNOR2_X1 U383 ( .A(G1GAT), .B(KEYINPUT97), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U386 ( .A(KEYINPUT1), .B(G148GAT), .Z(n334) );
  XNOR2_X1 U387 ( .A(G141GAT), .B(G120GAT), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n341) );
  XOR2_X1 U390 ( .A(G85GAT), .B(G162GAT), .Z(n339) );
  XNOR2_X1 U391 ( .A(n337), .B(G134GAT), .ZN(n338) );
  XNOR2_X1 U392 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U393 ( .A(n341), .B(n340), .Z(n346) );
  XOR2_X1 U394 ( .A(KEYINPUT5), .B(KEYINPUT100), .Z(n343) );
  XNOR2_X1 U395 ( .A(KEYINPUT99), .B(KEYINPUT98), .ZN(n342) );
  XNOR2_X1 U396 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U397 ( .A(G29GAT), .B(n344), .ZN(n345) );
  XNOR2_X1 U398 ( .A(n346), .B(n345), .ZN(n532) );
  XOR2_X1 U399 ( .A(G92GAT), .B(G85GAT), .Z(n348) );
  XNOR2_X1 U400 ( .A(G99GAT), .B(G106GAT), .ZN(n347) );
  XNOR2_X1 U401 ( .A(n348), .B(n347), .ZN(n415) );
  XOR2_X1 U402 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n350) );
  XNOR2_X1 U403 ( .A(G204GAT), .B(KEYINPUT75), .ZN(n349) );
  XNOR2_X1 U404 ( .A(n350), .B(n349), .ZN(n351) );
  XOR2_X1 U405 ( .A(n415), .B(n351), .Z(n355) );
  XNOR2_X1 U406 ( .A(n353), .B(n352), .ZN(n354) );
  XNOR2_X1 U407 ( .A(n355), .B(n354), .ZN(n362) );
  XOR2_X1 U408 ( .A(KEYINPUT32), .B(KEYINPUT33), .Z(n357) );
  NAND2_X1 U409 ( .A1(G230GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U411 ( .A(n358), .B(KEYINPUT31), .Z(n360) );
  XOR2_X1 U412 ( .A(G176GAT), .B(G64GAT), .Z(n438) );
  XOR2_X1 U413 ( .A(G57GAT), .B(KEYINPUT13), .Z(n404) );
  XNOR2_X1 U414 ( .A(n438), .B(n404), .ZN(n359) );
  XNOR2_X1 U415 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n577) );
  XOR2_X1 U417 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n363) );
  XOR2_X1 U418 ( .A(n577), .B(n363), .Z(n554) );
  XOR2_X1 U419 ( .A(G43GAT), .B(G29GAT), .Z(n365) );
  XNOR2_X1 U420 ( .A(KEYINPUT7), .B(G50GAT), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n366) );
  XOR2_X1 U422 ( .A(n366), .B(KEYINPUT8), .Z(n368) );
  XNOR2_X1 U423 ( .A(G36GAT), .B(KEYINPUT70), .ZN(n367) );
  XNOR2_X1 U424 ( .A(n368), .B(n367), .ZN(n423) );
  XOR2_X1 U425 ( .A(KEYINPUT69), .B(KEYINPUT67), .Z(n370) );
  XNOR2_X1 U426 ( .A(KEYINPUT68), .B(KEYINPUT29), .ZN(n369) );
  XOR2_X1 U427 ( .A(n370), .B(n369), .Z(n377) );
  INV_X1 U428 ( .A(n377), .ZN(n375) );
  XOR2_X1 U429 ( .A(G113GAT), .B(G197GAT), .Z(n373) );
  XOR2_X1 U430 ( .A(G169GAT), .B(G8GAT), .Z(n447) );
  XNOR2_X1 U431 ( .A(n371), .B(n447), .ZN(n372) );
  XNOR2_X1 U432 ( .A(n373), .B(n372), .ZN(n376) );
  INV_X1 U433 ( .A(n376), .ZN(n374) );
  NAND2_X1 U434 ( .A1(n375), .A2(n374), .ZN(n379) );
  NAND2_X1 U435 ( .A1(n377), .A2(n376), .ZN(n378) );
  NAND2_X1 U436 ( .A1(n379), .A2(n378), .ZN(n381) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U438 ( .A(n381), .B(n380), .ZN(n383) );
  INV_X1 U439 ( .A(KEYINPUT66), .ZN(n382) );
  XNOR2_X1 U440 ( .A(n383), .B(n382), .ZN(n386) );
  XNOR2_X1 U441 ( .A(G15GAT), .B(G1GAT), .ZN(n384) );
  XNOR2_X1 U442 ( .A(n384), .B(KEYINPUT71), .ZN(n405) );
  XNOR2_X1 U443 ( .A(n405), .B(KEYINPUT30), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U445 ( .A(n423), .B(n387), .ZN(n431) );
  AND2_X1 U446 ( .A1(n554), .A2(n431), .ZN(n389) );
  INV_X1 U447 ( .A(KEYINPUT46), .ZN(n388) );
  XNOR2_X1 U448 ( .A(n389), .B(n388), .ZN(n390) );
  XNOR2_X1 U449 ( .A(n390), .B(KEYINPUT119), .ZN(n412) );
  XOR2_X1 U450 ( .A(G78GAT), .B(G211GAT), .Z(n392) );
  XNOR2_X1 U451 ( .A(G127GAT), .B(G71GAT), .ZN(n391) );
  XNOR2_X1 U452 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT82), .B(G64GAT), .Z(n394) );
  XNOR2_X1 U454 ( .A(G8GAT), .B(G183GAT), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U456 ( .A(n396), .B(n395), .Z(n401) );
  XOR2_X1 U457 ( .A(KEYINPUT84), .B(KEYINPUT81), .Z(n398) );
  NAND2_X1 U458 ( .A1(G231GAT), .A2(G233GAT), .ZN(n397) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U460 ( .A(KEYINPUT15), .B(n399), .ZN(n400) );
  XNOR2_X1 U461 ( .A(n401), .B(n400), .ZN(n411) );
  XOR2_X1 U462 ( .A(KEYINPUT83), .B(KEYINPUT80), .Z(n403) );
  XNOR2_X1 U463 ( .A(KEYINPUT12), .B(KEYINPUT14), .ZN(n402) );
  XNOR2_X1 U464 ( .A(n403), .B(n402), .ZN(n409) );
  XOR2_X1 U465 ( .A(n404), .B(G155GAT), .Z(n407) );
  XNOR2_X1 U466 ( .A(n405), .B(G22GAT), .ZN(n406) );
  XNOR2_X1 U467 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U468 ( .A(n409), .B(n408), .Z(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n581) );
  NOR2_X1 U470 ( .A1(n412), .A2(n581), .ZN(n426) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n416), .B(KEYINPUT65), .ZN(n419) );
  XOR2_X1 U473 ( .A(n417), .B(KEYINPUT77), .Z(n418) );
  XNOR2_X1 U474 ( .A(n419), .B(n418), .ZN(n425) );
  XOR2_X1 U475 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n421) );
  XNOR2_X1 U476 ( .A(KEYINPUT78), .B(KEYINPUT9), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U478 ( .A(n423), .B(n422), .Z(n424) );
  XNOR2_X1 U479 ( .A(n425), .B(n424), .ZN(n559) );
  NAND2_X1 U480 ( .A1(n426), .A2(n559), .ZN(n427) );
  XNOR2_X1 U481 ( .A(n427), .B(KEYINPUT47), .ZN(n434) );
  INV_X1 U482 ( .A(KEYINPUT79), .ZN(n428) );
  XNOR2_X1 U483 ( .A(n428), .B(n559), .ZN(n546) );
  XNOR2_X1 U484 ( .A(KEYINPUT36), .B(n546), .ZN(n584) );
  INV_X1 U485 ( .A(n581), .ZN(n492) );
  NOR2_X1 U486 ( .A1(n584), .A2(n492), .ZN(n429) );
  XNOR2_X1 U487 ( .A(n429), .B(KEYINPUT45), .ZN(n430) );
  NAND2_X1 U488 ( .A1(n430), .A2(n577), .ZN(n432) );
  INV_X1 U489 ( .A(n431), .ZN(n507) );
  XNOR2_X1 U490 ( .A(KEYINPUT72), .B(n431), .ZN(n563) );
  NOR2_X1 U491 ( .A1(n432), .A2(n563), .ZN(n433) );
  NOR2_X1 U492 ( .A1(n434), .A2(n433), .ZN(n437) );
  XOR2_X1 U493 ( .A(n438), .B(KEYINPUT101), .Z(n440) );
  NAND2_X1 U494 ( .A1(G226GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U495 ( .A(n440), .B(n439), .ZN(n444) );
  XOR2_X1 U496 ( .A(G92GAT), .B(G218GAT), .Z(n442) );
  XNOR2_X1 U497 ( .A(G36GAT), .B(G190GAT), .ZN(n441) );
  XNOR2_X1 U498 ( .A(n442), .B(n441), .ZN(n443) );
  XOR2_X1 U499 ( .A(n444), .B(n443), .Z(n449) );
  INV_X1 U500 ( .A(n445), .ZN(n446) );
  XNOR2_X1 U501 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U502 ( .A(n449), .B(n448), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n522) );
  NAND2_X1 U504 ( .A1(n534), .A2(n522), .ZN(n453) );
  NOR2_X1 U505 ( .A1(n532), .A2(n454), .ZN(n574) );
  AND2_X1 U506 ( .A1(n469), .A2(n574), .ZN(n455) );
  XNOR2_X1 U507 ( .A(n455), .B(KEYINPUT55), .ZN(n456) );
  NAND2_X1 U508 ( .A1(n568), .A2(n554), .ZN(n459) );
  XOR2_X1 U509 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n457) );
  XNOR2_X1 U510 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n481) );
  NAND2_X1 U511 ( .A1(n577), .A2(n563), .ZN(n460) );
  XNOR2_X1 U512 ( .A(n460), .B(KEYINPUT76), .ZN(n496) );
  XOR2_X1 U513 ( .A(KEYINPUT16), .B(KEYINPUT85), .Z(n462) );
  NAND2_X1 U514 ( .A1(n581), .A2(n546), .ZN(n461) );
  XNOR2_X1 U515 ( .A(n462), .B(n461), .ZN(n478) );
  XOR2_X1 U516 ( .A(n522), .B(KEYINPUT27), .Z(n468) );
  NOR2_X1 U517 ( .A1(n539), .A2(n468), .ZN(n463) );
  NAND2_X1 U518 ( .A1(n536), .A2(n463), .ZN(n464) );
  NAND2_X1 U519 ( .A1(n532), .A2(n464), .ZN(n477) );
  INV_X1 U520 ( .A(n536), .ZN(n524) );
  NAND2_X1 U521 ( .A1(n522), .A2(n524), .ZN(n465) );
  XNOR2_X1 U522 ( .A(KEYINPUT104), .B(n465), .ZN(n466) );
  NAND2_X1 U523 ( .A1(n466), .A2(n469), .ZN(n467) );
  XOR2_X1 U524 ( .A(KEYINPUT25), .B(n467), .Z(n475) );
  INV_X1 U525 ( .A(n468), .ZN(n533) );
  NOR2_X1 U526 ( .A1(n469), .A2(n524), .ZN(n471) );
  XNOR2_X1 U527 ( .A(KEYINPUT102), .B(KEYINPUT26), .ZN(n470) );
  XNOR2_X1 U528 ( .A(n471), .B(n470), .ZN(n573) );
  NAND2_X1 U529 ( .A1(n533), .A2(n573), .ZN(n472) );
  XNOR2_X1 U530 ( .A(n472), .B(KEYINPUT103), .ZN(n473) );
  NOR2_X1 U531 ( .A1(n473), .A2(n532), .ZN(n474) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n476) );
  NAND2_X1 U533 ( .A1(n477), .A2(n476), .ZN(n491) );
  OR2_X1 U534 ( .A1(n478), .A2(n491), .ZN(n508) );
  NOR2_X1 U535 ( .A1(n496), .A2(n508), .ZN(n479) );
  XOR2_X1 U536 ( .A(KEYINPUT105), .B(n479), .Z(n487) );
  NAND2_X1 U537 ( .A1(n532), .A2(n487), .ZN(n480) );
  XNOR2_X1 U538 ( .A(n481), .B(n480), .ZN(G1324GAT) );
  XOR2_X1 U539 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n483) );
  NAND2_X1 U540 ( .A1(n487), .A2(n522), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U542 ( .A(G8GAT), .B(n484), .ZN(G1325GAT) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U544 ( .A1(n487), .A2(n524), .ZN(n485) );
  XNOR2_X1 U545 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  NAND2_X1 U546 ( .A1(n487), .A2(n539), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT108), .B(KEYINPUT111), .Z(n490) );
  XNOR2_X1 U549 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n500) );
  NOR2_X1 U551 ( .A1(n584), .A2(n491), .ZN(n493) );
  NAND2_X1 U552 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(n494), .B(KEYINPUT109), .ZN(n495) );
  XNOR2_X1 U554 ( .A(KEYINPUT37), .B(n495), .ZN(n520) );
  NOR2_X1 U555 ( .A1(n496), .A2(n520), .ZN(n498) );
  XNOR2_X1 U556 ( .A(KEYINPUT110), .B(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U557 ( .A(n498), .B(n497), .ZN(n505) );
  NAND2_X1 U558 ( .A1(n505), .A2(n532), .ZN(n499) );
  XOR2_X1 U559 ( .A(n500), .B(n499), .Z(G1328GAT) );
  NAND2_X1 U560 ( .A1(n505), .A2(n522), .ZN(n501) );
  XNOR2_X1 U561 ( .A(n501), .B(KEYINPUT112), .ZN(n502) );
  XNOR2_X1 U562 ( .A(G36GAT), .B(n502), .ZN(G1329GAT) );
  NAND2_X1 U563 ( .A1(n524), .A2(n505), .ZN(n503) );
  XNOR2_X1 U564 ( .A(n503), .B(KEYINPUT40), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G43GAT), .B(n504), .ZN(G1330GAT) );
  NAND2_X1 U566 ( .A1(n505), .A2(n539), .ZN(n506) );
  XNOR2_X1 U567 ( .A(n506), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT113), .B(KEYINPUT42), .Z(n510) );
  NAND2_X1 U569 ( .A1(n507), .A2(n554), .ZN(n519) );
  NOR2_X1 U570 ( .A1(n508), .A2(n519), .ZN(n516) );
  NAND2_X1 U571 ( .A1(n516), .A2(n532), .ZN(n509) );
  XNOR2_X1 U572 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(n511), .ZN(G1332GAT) );
  NAND2_X1 U574 ( .A1(n516), .A2(n522), .ZN(n512) );
  XNOR2_X1 U575 ( .A(n512), .B(KEYINPUT114), .ZN(n513) );
  XNOR2_X1 U576 ( .A(G64GAT), .B(n513), .ZN(G1333GAT) );
  XOR2_X1 U577 ( .A(G71GAT), .B(KEYINPUT115), .Z(n515) );
  NAND2_X1 U578 ( .A1(n516), .A2(n524), .ZN(n514) );
  XNOR2_X1 U579 ( .A(n515), .B(n514), .ZN(G1334GAT) );
  XOR2_X1 U580 ( .A(G78GAT), .B(KEYINPUT43), .Z(n518) );
  NAND2_X1 U581 ( .A1(n516), .A2(n539), .ZN(n517) );
  XNOR2_X1 U582 ( .A(n518), .B(n517), .ZN(G1335GAT) );
  NOR2_X1 U583 ( .A1(n520), .A2(n519), .ZN(n527) );
  NAND2_X1 U584 ( .A1(n532), .A2(n527), .ZN(n521) );
  XNOR2_X1 U585 ( .A(G85GAT), .B(n521), .ZN(G1336GAT) );
  NAND2_X1 U586 ( .A1(n527), .A2(n522), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U588 ( .A1(n524), .A2(n527), .ZN(n525) );
  XNOR2_X1 U589 ( .A(n525), .B(KEYINPUT116), .ZN(n526) );
  XNOR2_X1 U590 ( .A(G99GAT), .B(n526), .ZN(G1338GAT) );
  XNOR2_X1 U591 ( .A(G106GAT), .B(KEYINPUT117), .ZN(n531) );
  XOR2_X1 U592 ( .A(KEYINPUT44), .B(KEYINPUT118), .Z(n529) );
  NAND2_X1 U593 ( .A1(n527), .A2(n539), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(n530) );
  XNOR2_X1 U595 ( .A(n531), .B(n530), .ZN(G1339GAT) );
  AND2_X1 U596 ( .A1(n533), .A2(n532), .ZN(n535) );
  NAND2_X1 U597 ( .A1(n535), .A2(n534), .ZN(n552) );
  NOR2_X1 U598 ( .A1(n536), .A2(n552), .ZN(n537) );
  XNOR2_X1 U599 ( .A(n537), .B(KEYINPUT121), .ZN(n538) );
  NOR2_X1 U600 ( .A1(n539), .A2(n538), .ZN(n547) );
  NAND2_X1 U601 ( .A1(n563), .A2(n547), .ZN(n540) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n540), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(KEYINPUT122), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U604 ( .A1(n547), .A2(n554), .ZN(n541) );
  XNOR2_X1 U605 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U606 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  NAND2_X1 U607 ( .A1(n581), .A2(n547), .ZN(n544) );
  XNOR2_X1 U608 ( .A(n544), .B(KEYINPUT50), .ZN(n545) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT123), .B(KEYINPUT51), .Z(n549) );
  INV_X1 U611 ( .A(n546), .ZN(n567) );
  NAND2_X1 U612 ( .A1(n547), .A2(n567), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n549), .B(n548), .ZN(n550) );
  XOR2_X1 U614 ( .A(G134GAT), .B(n550), .Z(G1343GAT) );
  INV_X1 U615 ( .A(n573), .ZN(n551) );
  NOR2_X1 U616 ( .A1(n552), .A2(n551), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n561), .A2(n431), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n556) );
  NAND2_X1 U620 ( .A1(n561), .A2(n554), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n556), .B(n555), .ZN(n557) );
  XNOR2_X1 U622 ( .A(G148GAT), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U623 ( .A1(n581), .A2(n561), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G155GAT), .ZN(G1346GAT) );
  INV_X1 U625 ( .A(n559), .ZN(n560) );
  NAND2_X1 U626 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U627 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n568), .A2(n563), .ZN(n564) );
  XNOR2_X1 U629 ( .A(n564), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U630 ( .A(G183GAT), .B(KEYINPUT125), .Z(n566) );
  NAND2_X1 U631 ( .A1(n568), .A2(n581), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n566), .B(n565), .ZN(G1350GAT) );
  NAND2_X1 U633 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(n569), .B(KEYINPUT58), .ZN(n570) );
  XNOR2_X1 U635 ( .A(G190GAT), .B(n570), .ZN(G1351GAT) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n571), .B(KEYINPUT60), .ZN(n572) );
  XOR2_X1 U638 ( .A(KEYINPUT126), .B(n572), .Z(n576) );
  NAND2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n583) );
  INV_X1 U640 ( .A(n583), .ZN(n580) );
  NAND2_X1 U641 ( .A1(n580), .A2(n431), .ZN(n575) );
  XNOR2_X1 U642 ( .A(n576), .B(n575), .ZN(G1352GAT) );
  XOR2_X1 U643 ( .A(G204GAT), .B(KEYINPUT61), .Z(n579) );
  OR2_X1 U644 ( .A1(n583), .A2(n577), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U649 ( .A(KEYINPUT62), .B(n585), .Z(n586) );
  XNOR2_X1 U650 ( .A(G218GAT), .B(n586), .ZN(G1355GAT) );
endmodule

