//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 0 1 0 1 1 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:00 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n652, new_n653, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n679, new_n680, new_n681, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n706, new_n707, new_n708,
    new_n709, new_n711, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n793, new_n794, new_n796, new_n797, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n847, new_n848, new_n850, new_n851, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n878,
    new_n879, new_n880, new_n881, new_n882, new_n883, new_n884, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n934, new_n935;
  XNOR2_X1  g000(.A(G15gat), .B(G43gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  XNOR2_X1  g003(.A(KEYINPUT27), .B(G183gat), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(KEYINPUT68), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND3_X1  g006(.A1(new_n206), .A2(KEYINPUT28), .A3(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT28), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT67), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n205), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G183gat), .ZN(new_n212));
  AND2_X1   g011(.A1(new_n212), .A2(KEYINPUT27), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n207), .B1(new_n213), .B2(KEYINPUT67), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n209), .B1(new_n211), .B2(new_n214), .ZN(new_n215));
  AOI22_X1  g014(.A1(new_n208), .A2(new_n215), .B1(G183gat), .B2(G190gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(G169gat), .A2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT66), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n217), .B(new_n218), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT26), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g020(.A(new_n221), .B(KEYINPUT69), .Z(new_n222));
  NAND2_X1  g021(.A1(G169gat), .A2(G176gat), .ZN(new_n223));
  XOR2_X1   g022(.A(new_n223), .B(KEYINPUT65), .Z(new_n224));
  OAI21_X1  g023(.A(new_n224), .B1(new_n220), .B2(new_n217), .ZN(new_n225));
  OAI21_X1  g024(.A(new_n216), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  XNOR2_X1  g025(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n228), .B1(G169gat), .B2(G176gat), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n217), .A2(KEYINPUT23), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n224), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g030(.A1(new_n212), .A2(new_n207), .A3(KEYINPUT24), .ZN(new_n232));
  INV_X1    g031(.A(new_n232), .ZN(new_n233));
  XNOR2_X1  g032(.A(G183gat), .B(G190gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT24), .ZN(new_n235));
  OAI21_X1  g034(.A(new_n233), .B1(new_n234), .B2(new_n235), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n227), .B1(new_n231), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n224), .A2(KEYINPUT25), .A3(new_n229), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n238), .A2(new_n236), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n219), .A2(KEYINPUT23), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n226), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(G113gat), .B(G120gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n243), .A2(KEYINPUT1), .ZN(new_n244));
  XNOR2_X1  g043(.A(G127gat), .B(G134gat), .ZN(new_n245));
  OR2_X1    g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT70), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n243), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n249));
  INV_X1    g048(.A(G120gat), .ZN(new_n250));
  OR3_X1    g049(.A1(new_n247), .A2(new_n250), .A3(G113gat), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n248), .A2(new_n249), .A3(new_n245), .A4(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n242), .A2(KEYINPUT71), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n226), .A2(new_n241), .ZN(new_n255));
  OR2_X1    g054(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n253), .A2(KEYINPUT71), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n256), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n254), .A2(G227gat), .A3(G233gat), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT33), .ZN(new_n260));
  AOI21_X1  g059(.A(new_n204), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n259), .A2(KEYINPUT32), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  OAI211_X1 g062(.A(new_n259), .B(KEYINPUT32), .C1(new_n260), .C2(new_n204), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT34), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n258), .ZN(new_n267));
  NAND2_X1  g066(.A1(G227gat), .A2(G233gat), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND3_X1   g068(.A1(new_n267), .A2(new_n266), .A3(new_n268), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n265), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n269), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n272), .A2(new_n263), .A3(new_n264), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n271), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g073(.A(G197gat), .B(G204gat), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT22), .ZN(new_n276));
  INV_X1    g075(.A(G211gat), .ZN(new_n277));
  INV_X1    g076(.A(G218gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  XNOR2_X1  g079(.A(G211gat), .B(G218gat), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  NOR2_X1   g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(new_n283), .B(KEYINPUT75), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(KEYINPUT73), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT73), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n281), .A2(new_n286), .ZN(new_n287));
  AND3_X1   g086(.A1(new_n285), .A2(new_n280), .A3(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AND2_X1   g089(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  OR2_X1    g090(.A1(new_n288), .A2(new_n289), .ZN(new_n292));
  AND2_X1   g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  XOR2_X1   g092(.A(KEYINPUT81), .B(G155gat), .Z(new_n294));
  NAND2_X1  g093(.A1(new_n294), .A2(G162gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT2), .ZN(new_n296));
  XOR2_X1   g095(.A(G141gat), .B(G148gat), .Z(new_n297));
  XNOR2_X1  g096(.A(G155gat), .B(G162gat), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n296), .A2(new_n297), .A3(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT2), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n298), .A2(KEYINPUT80), .ZN(new_n302));
  NOR2_X1   g101(.A1(G155gat), .A2(G162gat), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n301), .B(new_n302), .C1(KEYINPUT80), .C2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n299), .A2(new_n304), .ZN(new_n305));
  OR2_X1    g104(.A1(new_n305), .A2(KEYINPUT3), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT76), .B(KEYINPUT29), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n292), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  AOI21_X1  g110(.A(KEYINPUT3), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n305), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n309), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n314), .A2(G228gat), .A3(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(G228gat), .A2(G233gat), .ZN(new_n316));
  INV_X1    g115(.A(new_n280), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n284), .B1(new_n281), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(KEYINPUT3), .B1(new_n318), .B2(new_n307), .ZN(new_n319));
  OAI211_X1 g118(.A(new_n309), .B(new_n316), .C1(new_n313), .C2(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(KEYINPUT31), .B(G50gat), .ZN(new_n321));
  INV_X1    g120(.A(new_n321), .ZN(new_n322));
  AND3_X1   g121(.A1(new_n315), .A2(new_n320), .A3(new_n322), .ZN(new_n323));
  AOI21_X1  g122(.A(new_n322), .B1(new_n315), .B2(new_n320), .ZN(new_n324));
  XNOR2_X1  g123(.A(G78gat), .B(G106gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n325), .B(G22gat), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  OR3_X1    g126(.A1(new_n323), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n327), .B1(new_n323), .B2(new_n324), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n328), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n274), .A2(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G225gat), .A2(G233gat), .ZN(new_n332));
  INV_X1    g131(.A(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n253), .ZN(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n305), .B2(KEYINPUT3), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n333), .B1(new_n306), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n305), .A2(new_n253), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n337), .A2(KEYINPUT82), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT82), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n305), .B2(new_n253), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n339), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n336), .B(new_n338), .C1(new_n342), .C2(KEYINPUT4), .ZN(new_n343));
  OAI211_X1 g142(.A(new_n339), .B(new_n341), .C1(new_n334), .C2(new_n313), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n344), .A2(new_n333), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n343), .A2(KEYINPUT5), .A3(new_n345), .ZN(new_n346));
  NOR2_X1   g145(.A1(new_n337), .A2(KEYINPUT4), .ZN(new_n347));
  AOI21_X1  g146(.A(new_n347), .B1(new_n342), .B2(KEYINPUT4), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT5), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n348), .A2(new_n349), .A3(new_n336), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  XNOR2_X1  g151(.A(G1gat), .B(G29gat), .ZN(new_n353));
  XNOR2_X1  g152(.A(new_n353), .B(KEYINPUT0), .ZN(new_n354));
  XNOR2_X1  g153(.A(G57gat), .B(G85gat), .ZN(new_n355));
  XOR2_X1   g154(.A(new_n354), .B(new_n355), .Z(new_n356));
  NOR2_X1   g155(.A1(new_n352), .A2(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT83), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT6), .ZN(new_n359));
  INV_X1    g158(.A(new_n356), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n359), .B1(new_n351), .B2(new_n360), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n357), .B1(new_n358), .B2(new_n361), .ZN(new_n362));
  OR2_X1    g161(.A1(new_n361), .A2(new_n358), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n351), .A2(KEYINPUT6), .A3(new_n360), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(G226gat), .A2(G233gat), .ZN(new_n367));
  INV_X1    g166(.A(new_n307), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n367), .B1(new_n242), .B2(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n255), .A2(G226gat), .A3(G233gat), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n371), .A2(new_n293), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n367), .B1(new_n242), .B2(KEYINPUT29), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n373), .A2(new_n370), .A3(new_n310), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT77), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT77), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n372), .A2(new_n377), .A3(new_n374), .ZN(new_n378));
  XNOR2_X1  g177(.A(G8gat), .B(G36gat), .ZN(new_n379));
  XNOR2_X1  g178(.A(G64gat), .B(G92gat), .ZN(new_n380));
  XOR2_X1   g179(.A(new_n379), .B(new_n380), .Z(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(KEYINPUT78), .Z(new_n382));
  INV_X1    g181(.A(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n376), .A2(new_n378), .A3(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n372), .A2(new_n374), .A3(new_n381), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT30), .ZN(new_n386));
  OR2_X1    g185(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT79), .ZN(new_n388));
  AND3_X1   g187(.A1(new_n385), .A2(new_n388), .A3(new_n386), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n384), .B(new_n387), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  NAND3_X1  g191(.A1(new_n331), .A2(new_n366), .A3(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT35), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n330), .A2(KEYINPUT35), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT72), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n271), .A2(new_n396), .A3(new_n273), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n265), .B(KEYINPUT72), .C1(new_n269), .C2(new_n270), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n397), .A2(new_n398), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n365), .B1(new_n357), .B2(new_n361), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n395), .A2(new_n399), .A3(new_n392), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n394), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT86), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(new_n375), .B2(KEYINPUT37), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT37), .ZN(new_n405));
  NAND4_X1  g204(.A1(new_n372), .A2(KEYINPUT86), .A3(new_n405), .A4(new_n374), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n381), .B1(new_n404), .B2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n376), .A2(KEYINPUT37), .A3(new_n378), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT38), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n382), .A2(KEYINPUT38), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n373), .A2(new_n370), .A3(new_n293), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT37), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n293), .B1(new_n369), .B2(new_n370), .ZN(new_n414));
  OAI21_X1  g213(.A(new_n411), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n404), .B2(new_n406), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n365), .B(new_n385), .C1(new_n357), .C2(new_n361), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n330), .B1(new_n410), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT85), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n306), .A2(new_n335), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n348), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(new_n333), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n356), .B1(new_n423), .B2(KEYINPUT39), .ZN(new_n424));
  OAI21_X1  g223(.A(KEYINPUT39), .B1(new_n344), .B2(new_n333), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n425), .B1(new_n422), .B2(new_n333), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT84), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  OR2_X1    g226(.A1(new_n427), .A2(KEYINPUT40), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n357), .B1(new_n427), .B2(KEYINPUT40), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n420), .B1(new_n392), .B2(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n391), .A2(KEYINPUT85), .A3(new_n429), .A4(new_n428), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n419), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(KEYINPUT36), .B1(new_n397), .B2(new_n398), .ZN(new_n434));
  AND2_X1   g233(.A1(new_n274), .A2(KEYINPUT36), .ZN(new_n435));
  NOR2_X1   g234(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  AND2_X1   g235(.A1(new_n364), .A2(new_n365), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n330), .B1(new_n437), .B2(new_n391), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n402), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(G36gat), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n441), .A2(KEYINPUT89), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n441), .A2(KEYINPUT89), .ZN(new_n443));
  OAI21_X1  g242(.A(G29gat), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G29gat), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n445), .A2(new_n441), .A3(KEYINPUT88), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT88), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(G29gat), .B2(G36gat), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n446), .A2(new_n448), .A3(KEYINPUT14), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT14), .ZN(new_n450));
  OAI211_X1 g249(.A(new_n447), .B(new_n450), .C1(G29gat), .C2(G36gat), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n444), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(G50gat), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(G43gat), .ZN(new_n455));
  INV_X1    g254(.A(G43gat), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(G50gat), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n455), .A2(new_n457), .A3(KEYINPUT15), .ZN(new_n458));
  XNOR2_X1  g257(.A(KEYINPUT91), .B(KEYINPUT15), .ZN(new_n459));
  OR3_X1    g258(.A1(new_n454), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n457), .A2(KEYINPUT93), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  OR2_X1    g261(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(KEYINPUT92), .A2(G43gat), .ZN(new_n464));
  AOI21_X1  g263(.A(G50gat), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n459), .B1(new_n462), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n453), .A2(new_n458), .A3(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n458), .ZN(new_n468));
  AND3_X1   g267(.A1(new_n452), .A2(KEYINPUT90), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT90), .B1(new_n452), .B2(new_n468), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT17), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  OAI211_X1 g272(.A(new_n467), .B(KEYINPUT17), .C1(new_n469), .C2(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(G85gat), .A2(G92gat), .ZN(new_n475));
  XNOR2_X1  g274(.A(new_n475), .B(KEYINPUT7), .ZN(new_n476));
  NAND2_X1  g275(.A1(G99gat), .A2(G106gat), .ZN(new_n477));
  INV_X1    g276(.A(G85gat), .ZN(new_n478));
  INV_X1    g277(.A(G92gat), .ZN(new_n479));
  AOI22_X1  g278(.A1(KEYINPUT8), .A2(new_n477), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  XNOR2_X1  g280(.A(G99gat), .B(G106gat), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n481), .B(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n473), .A2(new_n474), .A3(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(G232gat), .A2(G233gat), .ZN(new_n486));
  AOI22_X1  g285(.A1(new_n471), .A2(new_n483), .B1(KEYINPUT41), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  XOR2_X1   g287(.A(G190gat), .B(G218gat), .Z(new_n489));
  XNOR2_X1  g288(.A(new_n489), .B(KEYINPUT104), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n488), .B(new_n491), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n486), .A2(KEYINPUT41), .ZN(new_n493));
  XNOR2_X1  g292(.A(G134gat), .B(G162gat), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n493), .B(new_n494), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n492), .B(new_n495), .ZN(new_n496));
  XOR2_X1   g295(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(G155gat), .ZN(new_n498));
  XNOR2_X1  g297(.A(G183gat), .B(G211gat), .ZN(new_n499));
  XOR2_X1   g298(.A(new_n498), .B(new_n499), .Z(new_n500));
  INV_X1    g299(.A(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(G71gat), .ZN(new_n502));
  INV_X1    g301(.A(G78gat), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(G71gat), .A2(G78gat), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT103), .ZN(new_n507));
  INV_X1    g306(.A(new_n505), .ZN(new_n508));
  OR2_X1    g307(.A1(new_n508), .A2(KEYINPUT9), .ZN(new_n509));
  NOR2_X1   g308(.A1(G57gat), .A2(G64gat), .ZN(new_n510));
  INV_X1    g309(.A(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(G57gat), .A2(G64gat), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n507), .A2(new_n509), .A3(new_n511), .A4(new_n512), .ZN(new_n513));
  NAND3_X1  g312(.A1(new_n511), .A2(KEYINPUT101), .A3(new_n512), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT101), .ZN(new_n515));
  INV_X1    g314(.A(new_n512), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n515), .B1(new_n516), .B2(new_n510), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n509), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT100), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n505), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(KEYINPUT100), .B1(G71gat), .B2(G78gat), .ZN(new_n522));
  OAI21_X1  g321(.A(new_n504), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g323(.A(KEYINPUT102), .B1(new_n519), .B2(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n508), .A2(KEYINPUT9), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n526), .B1(new_n514), .B2(new_n517), .ZN(new_n527));
  INV_X1    g326(.A(KEYINPUT102), .ZN(new_n528));
  NOR3_X1   g327(.A1(new_n527), .A2(new_n528), .A3(new_n523), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n513), .B1(new_n525), .B2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n531), .A2(KEYINPUT21), .ZN(new_n532));
  NAND2_X1  g331(.A1(G231gat), .A2(G233gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n534), .A2(G127gat), .ZN(new_n535));
  INV_X1    g334(.A(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(G15gat), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(G22gat), .ZN(new_n538));
  INV_X1    g337(.A(G22gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n539), .A2(G15gat), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(G1gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT16), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n543), .A2(G1gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n538), .A3(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(G8gat), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT95), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT95), .ZN(new_n549));
  AOI211_X1 g348(.A(new_n549), .B(G8gat), .C1(new_n542), .C2(new_n545), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(G1gat), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G22gat), .ZN(new_n553));
  OAI211_X1 g352(.A(new_n545), .B(G8gat), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT94), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n542), .A2(KEYINPUT94), .A3(G8gat), .A4(new_n545), .ZN(new_n557));
  AND2_X1   g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n560), .B1(new_n531), .B2(KEYINPUT21), .ZN(new_n561));
  INV_X1    g360(.A(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n534), .A2(G127gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n536), .A2(new_n562), .A3(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n562), .B1(new_n536), .B2(new_n563), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n501), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n566), .ZN(new_n568));
  NAND3_X1  g367(.A1(new_n568), .A2(new_n564), .A3(new_n500), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n496), .B1(new_n567), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  INV_X1    g370(.A(KEYINPUT96), .ZN(new_n572));
  OAI21_X1  g371(.A(new_n572), .B1(new_n551), .B2(new_n558), .ZN(new_n573));
  AND3_X1   g372(.A1(new_n544), .A2(new_n538), .A3(new_n540), .ZN(new_n574));
  AOI21_X1  g373(.A(new_n552), .B1(new_n538), .B2(new_n540), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n547), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(new_n549), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n546), .A2(KEYINPUT95), .A3(new_n547), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n556), .A2(new_n557), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(KEYINPUT96), .A3(new_n580), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n473), .A2(new_n573), .A3(new_n474), .A4(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT97), .ZN(new_n583));
  AND3_X1   g382(.A1(new_n579), .A2(KEYINPUT96), .A3(new_n580), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT96), .B1(new_n579), .B2(new_n580), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT97), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n586), .A2(new_n587), .A3(new_n474), .A4(new_n473), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n560), .A2(new_n471), .ZN(new_n590));
  NAND2_X1  g389(.A1(G229gat), .A2(G233gat), .ZN(new_n591));
  XOR2_X1   g390(.A(new_n591), .B(KEYINPUT98), .Z(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n590), .A2(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n589), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT18), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n596), .A2(KEYINPUT99), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT99), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n594), .B1(new_n583), .B2(new_n588), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n599), .B1(new_n600), .B2(KEYINPUT18), .ZN(new_n601));
  XOR2_X1   g400(.A(new_n592), .B(KEYINPUT13), .Z(new_n602));
  OR2_X1    g401(.A1(new_n560), .A2(new_n471), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n590), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n604), .B1(new_n600), .B2(KEYINPUT18), .ZN(new_n605));
  XNOR2_X1  g404(.A(G113gat), .B(G141gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT11), .B(G169gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  XNOR2_X1  g408(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n610));
  XOR2_X1   g409(.A(new_n609), .B(new_n610), .Z(new_n611));
  NAND4_X1  g410(.A1(new_n598), .A2(new_n601), .A3(new_n605), .A4(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(new_n611), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n589), .A2(KEYINPUT18), .A3(new_n595), .ZN(new_n614));
  INV_X1    g413(.A(new_n604), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n600), .A2(KEYINPUT18), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n613), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n612), .A2(new_n618), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G230gat), .ZN(new_n621));
  INV_X1    g420(.A(G233gat), .ZN(new_n622));
  NOR2_X1   g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n530), .A2(new_n484), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n519), .A2(new_n524), .A3(KEYINPUT102), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n528), .B1(new_n527), .B2(new_n523), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g427(.A1(new_n628), .A2(new_n513), .A3(new_n483), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n624), .A2(new_n625), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n531), .A2(KEYINPUT10), .A3(new_n483), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n623), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(new_n623), .ZN(new_n633));
  AOI21_X1  g432(.A(new_n633), .B1(new_n624), .B2(new_n629), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(G176gat), .B(G204gat), .ZN(new_n636));
  XOR2_X1   g435(.A(new_n635), .B(new_n636), .Z(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  OR3_X1    g437(.A1(new_n632), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n638), .B1(new_n632), .B2(new_n634), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR3_X1   g440(.A1(new_n571), .A2(new_n620), .A3(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n440), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n366), .ZN(new_n644));
  XNOR2_X1  g443(.A(new_n644), .B(new_n552), .ZN(G1324gat));
  INV_X1    g444(.A(new_n643), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n547), .B1(new_n646), .B2(new_n391), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT16), .B(G8gat), .ZN(new_n648));
  NOR3_X1   g447(.A1(new_n643), .A2(new_n392), .A3(new_n648), .ZN(new_n649));
  OAI21_X1  g448(.A(KEYINPUT42), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n650), .B1(KEYINPUT42), .B2(new_n649), .ZN(G1325gat));
  OAI21_X1  g450(.A(G15gat), .B1(new_n643), .B2(new_n436), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n399), .A2(new_n537), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n652), .B1(new_n643), .B2(new_n653), .ZN(G1326gat));
  INV_X1    g453(.A(new_n330), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n643), .A2(new_n655), .ZN(new_n656));
  XOR2_X1   g455(.A(KEYINPUT43), .B(G22gat), .Z(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(G1327gat));
  AOI21_X1  g457(.A(new_n655), .B1(new_n366), .B2(new_n392), .ZN(new_n659));
  NOR3_X1   g458(.A1(new_n659), .A2(new_n435), .A3(new_n434), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n419), .A2(new_n431), .A3(new_n432), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n660), .A2(new_n661), .B1(new_n394), .B2(new_n401), .ZN(new_n662));
  INV_X1    g461(.A(new_n496), .ZN(new_n663));
  NOR2_X1   g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n567), .A2(new_n569), .ZN(new_n665));
  NOR3_X1   g464(.A1(new_n665), .A2(new_n620), .A3(new_n641), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n664), .A2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n445), .A3(new_n437), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n669), .B(KEYINPUT45), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT44), .ZN(new_n671));
  OAI21_X1  g470(.A(new_n671), .B1(new_n662), .B2(new_n663), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n440), .A2(KEYINPUT44), .A3(new_n496), .ZN(new_n673));
  AND2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n666), .B(KEYINPUT105), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(G29gat), .B1(new_n676), .B2(new_n366), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n670), .A2(new_n677), .ZN(G1328gat));
  NOR4_X1   g477(.A1(new_n667), .A2(new_n392), .A3(new_n442), .A4(new_n443), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT46), .ZN(new_n680));
  OAI22_X1  g479(.A1(new_n676), .A2(new_n392), .B1(new_n442), .B2(new_n443), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(G1329gat));
  AND2_X1   g481(.A1(new_n463), .A2(new_n464), .ZN(new_n683));
  INV_X1    g482(.A(new_n399), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n667), .B2(new_n684), .ZN(new_n685));
  OR2_X1    g484(.A1(new_n436), .A2(new_n683), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n685), .B1(new_n676), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n687), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g487(.A1(new_n672), .A2(new_n673), .A3(new_n330), .A4(new_n675), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n689), .A2(G50gat), .ZN(new_n690));
  AOI21_X1  g489(.A(KEYINPUT48), .B1(new_n690), .B2(KEYINPUT106), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n668), .A2(new_n454), .A3(new_n330), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(new_n690), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n691), .B(new_n693), .ZN(G1331gat));
  NAND2_X1  g493(.A1(new_n620), .A2(new_n641), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n571), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n440), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n698), .A2(new_n437), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g499(.A1(new_n697), .A2(new_n392), .ZN(new_n701));
  NOR2_X1   g500(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n703));
  OAI21_X1  g502(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n704), .B1(new_n701), .B2(new_n702), .ZN(G1333gat));
  NOR3_X1   g504(.A1(new_n697), .A2(G71gat), .A3(new_n684), .ZN(new_n706));
  OR2_X1    g505(.A1(new_n434), .A2(new_n435), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n698), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g507(.A(new_n706), .B1(G71gat), .B2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g509(.A1(new_n697), .A2(new_n655), .ZN(new_n711));
  XNOR2_X1  g510(.A(new_n711), .B(new_n503), .ZN(G1335gat));
  NOR2_X1   g511(.A1(new_n665), .A2(new_n695), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n674), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(G85gat), .B1(new_n714), .B2(new_n366), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT107), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  AOI211_X1 g516(.A(new_n619), .B(new_n665), .C1(new_n716), .C2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n440), .A2(new_n496), .A3(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n717), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n720), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n440), .A2(new_n496), .A3(new_n722), .A4(new_n718), .ZN(new_n723));
  AND2_X1   g522(.A1(new_n721), .A2(new_n723), .ZN(new_n724));
  NAND4_X1  g523(.A1(new_n724), .A2(new_n478), .A3(new_n437), .A4(new_n641), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n715), .A2(new_n725), .ZN(G1336gat));
  NAND4_X1  g525(.A1(new_n672), .A2(new_n673), .A3(new_n391), .A4(new_n713), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n727), .A2(G92gat), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  AOI21_X1  g528(.A(KEYINPUT52), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n392), .A2(G92gat), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n721), .A2(new_n641), .A3(new_n723), .A4(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g533(.A(new_n728), .B(new_n732), .C1(new_n729), .C2(KEYINPUT52), .ZN(new_n735));
  AND2_X1   g534(.A1(new_n734), .A2(new_n735), .ZN(G1337gat));
  OAI21_X1  g535(.A(G99gat), .B1(new_n714), .B2(new_n436), .ZN(new_n737));
  INV_X1    g536(.A(new_n641), .ZN(new_n738));
  NOR3_X1   g537(.A1(new_n684), .A2(G99gat), .A3(new_n738), .ZN(new_n739));
  XOR2_X1   g538(.A(new_n739), .B(KEYINPUT109), .Z(new_n740));
  NAND2_X1  g539(.A1(new_n724), .A2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n737), .A2(new_n741), .ZN(G1338gat));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n655), .A2(G106gat), .ZN(new_n744));
  NAND4_X1  g543(.A1(new_n721), .A2(new_n641), .A3(new_n723), .A4(new_n744), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n743), .B1(new_n745), .B2(KEYINPUT110), .ZN(new_n746));
  NAND4_X1  g545(.A1(new_n672), .A2(new_n673), .A3(new_n330), .A4(new_n713), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(G106gat), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(new_n745), .ZN(new_n749));
  XNOR2_X1  g548(.A(new_n746), .B(new_n749), .ZN(G1339gat));
  NAND2_X1  g549(.A1(new_n630), .A2(new_n631), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(new_n633), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n630), .A2(new_n631), .A3(new_n623), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n752), .A2(KEYINPUT54), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT54), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n637), .B1(new_n632), .B2(new_n755), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n754), .A2(KEYINPUT55), .A3(new_n756), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n639), .ZN(new_n758));
  AOI21_X1  g557(.A(KEYINPUT55), .B1(new_n754), .B2(new_n756), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n760), .A2(new_n612), .A3(new_n496), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n603), .A2(new_n590), .A3(new_n602), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n593), .B1(new_n589), .B2(new_n590), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT111), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n762), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g564(.A(KEYINPUT111), .B(new_n593), .C1(new_n589), .C2(new_n590), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n609), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n761), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n619), .A2(new_n760), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n767), .A2(new_n612), .A3(new_n641), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n771), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n663), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n773), .B1(new_n771), .B2(new_n772), .ZN(new_n776));
  OAI21_X1  g575(.A(new_n770), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n665), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n777), .A2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n570), .A2(new_n620), .A3(new_n738), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n330), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n366), .A2(new_n391), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(new_n399), .A3(new_n782), .ZN(new_n783));
  OAI21_X1  g582(.A(G113gat), .B1(new_n783), .B2(new_n620), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT113), .ZN(new_n785));
  INV_X1    g584(.A(new_n780), .ZN(new_n786));
  AOI21_X1  g585(.A(new_n786), .B1(new_n777), .B2(new_n778), .ZN(new_n787));
  INV_X1    g586(.A(new_n782), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(new_n331), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n790), .A2(G113gat), .A3(new_n620), .ZN(new_n791));
  OR2_X1    g590(.A1(new_n785), .A2(new_n791), .ZN(G1340gat));
  NOR3_X1   g591(.A1(new_n783), .A2(new_n250), .A3(new_n738), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n331), .A3(new_n641), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n793), .B1(new_n250), .B2(new_n794), .ZN(G1341gat));
  OAI21_X1  g594(.A(G127gat), .B1(new_n783), .B2(new_n778), .ZN(new_n796));
  OR2_X1    g595(.A1(new_n778), .A2(G127gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n796), .B1(new_n790), .B2(new_n797), .ZN(G1342gat));
  OR2_X1    g597(.A1(new_n663), .A2(G134gat), .ZN(new_n799));
  OAI22_X1  g598(.A1(new_n790), .A2(new_n799), .B1(KEYINPUT115), .B2(KEYINPUT56), .ZN(new_n800));
  NAND2_X1  g599(.A1(KEYINPUT115), .A2(KEYINPUT56), .ZN(new_n801));
  XOR2_X1   g600(.A(new_n800), .B(new_n801), .Z(new_n802));
  OAI21_X1  g601(.A(G134gat), .B1(new_n783), .B2(new_n663), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n804));
  AND2_X1   g603(.A1(new_n803), .A2(KEYINPUT114), .ZN(new_n805));
  OAI21_X1  g604(.A(new_n802), .B1(new_n804), .B2(new_n805), .ZN(G1343gat));
  NAND2_X1  g605(.A1(new_n436), .A2(new_n330), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT117), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n789), .ZN(new_n809));
  OR3_X1    g608(.A1(new_n809), .A2(G141gat), .A3(new_n620), .ZN(new_n810));
  AOI21_X1  g609(.A(KEYINPUT99), .B1(new_n596), .B2(new_n597), .ZN(new_n811));
  NOR3_X1   g610(.A1(new_n600), .A2(new_n599), .A3(KEYINPUT18), .ZN(new_n812));
  NOR2_X1   g611(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n616), .A2(new_n613), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n738), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  AOI22_X1  g614(.A1(new_n815), .A2(new_n767), .B1(new_n619), .B2(new_n760), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n816), .A2(new_n496), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n778), .B1(new_n817), .B2(new_n769), .ZN(new_n818));
  OR2_X1    g617(.A1(new_n818), .A2(KEYINPUT116), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n786), .B1(new_n818), .B2(KEYINPUT116), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT57), .B1(new_n821), .B2(new_n655), .ZN(new_n822));
  NOR2_X1   g621(.A1(new_n787), .A2(new_n655), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT57), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n707), .A2(new_n788), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n822), .A2(new_n825), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(G141gat), .B1(new_n827), .B2(new_n620), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n810), .A2(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n829), .A2(KEYINPUT58), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT58), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n810), .A2(new_n828), .A3(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n830), .A2(new_n832), .ZN(G1344gat));
  INV_X1    g632(.A(new_n827), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT59), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n834), .A2(new_n835), .A3(new_n641), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n823), .A2(KEYINPUT57), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n655), .B1(new_n818), .B2(new_n780), .ZN(new_n838));
  OR3_X1    g637(.A1(new_n838), .A2(KEYINPUT118), .A3(KEYINPUT57), .ZN(new_n839));
  OAI21_X1  g638(.A(KEYINPUT118), .B1(new_n838), .B2(KEYINPUT57), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n837), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n841), .A2(new_n641), .A3(new_n826), .ZN(new_n842));
  NAND2_X1  g641(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n843));
  INV_X1    g642(.A(new_n809), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n835), .B1(new_n844), .B2(new_n641), .ZN(new_n845));
  OAI221_X1 g644(.A(new_n836), .B1(new_n842), .B2(new_n843), .C1(G148gat), .C2(new_n845), .ZN(G1345gat));
  OAI21_X1  g645(.A(new_n294), .B1(new_n827), .B2(new_n778), .ZN(new_n847));
  OR2_X1    g646(.A1(new_n778), .A2(new_n294), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n847), .B1(new_n809), .B2(new_n848), .ZN(G1346gat));
  AOI21_X1  g648(.A(G162gat), .B1(new_n844), .B2(new_n496), .ZN(new_n850));
  AND2_X1   g649(.A1(new_n496), .A2(G162gat), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n850), .B1(new_n834), .B2(new_n851), .ZN(G1347gat));
  NAND2_X1  g651(.A1(new_n366), .A2(new_n391), .ZN(new_n853));
  NOR2_X1   g652(.A1(new_n684), .A2(new_n853), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n781), .A2(new_n854), .ZN(new_n855));
  INV_X1    g654(.A(G169gat), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n855), .A2(new_n856), .A3(new_n620), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n331), .A2(new_n391), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT120), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n331), .A2(KEYINPUT120), .A3(new_n391), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g661(.A(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT119), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n787), .B2(new_n437), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n771), .A2(new_n772), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(KEYINPUT112), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n867), .A2(new_n663), .A3(new_n774), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n665), .B1(new_n868), .B2(new_n770), .ZN(new_n869));
  OAI211_X1 g668(.A(KEYINPUT119), .B(new_n366), .C1(new_n869), .C2(new_n786), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n863), .B1(new_n865), .B2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n871), .A2(new_n619), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n857), .B1(new_n872), .B2(new_n856), .ZN(G1348gat));
  OAI21_X1  g672(.A(G176gat), .B1(new_n855), .B2(new_n738), .ZN(new_n874));
  INV_X1    g673(.A(new_n871), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n738), .A2(G176gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(G1349gat));
  INV_X1    g676(.A(KEYINPUT124), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT122), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n496), .B1(new_n816), .B2(new_n773), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n769), .B1(new_n880), .B2(new_n867), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n780), .B1(new_n881), .B2(new_n665), .ZN(new_n882));
  NAND4_X1  g681(.A1(new_n882), .A2(new_n655), .A3(new_n665), .A4(new_n854), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(KEYINPUT121), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT121), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n781), .A2(new_n885), .A3(new_n665), .A4(new_n854), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n884), .A2(G183gat), .A3(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(KEYINPUT123), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n865), .A2(new_n870), .ZN(new_n889));
  AND2_X1   g688(.A1(new_n665), .A2(new_n206), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n889), .A2(new_n862), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n887), .A2(new_n888), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n212), .B1(new_n883), .B2(KEYINPUT121), .ZN(new_n893));
  AOI22_X1  g692(.A1(new_n886), .A2(new_n893), .B1(new_n871), .B2(new_n890), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n879), .A2(KEYINPUT60), .ZN(new_n895));
  AOI22_X1  g694(.A1(new_n879), .A2(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(KEYINPUT60), .B1(new_n894), .B2(new_n888), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n878), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  INV_X1    g697(.A(KEYINPUT60), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n892), .A2(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(KEYINPUT122), .B1(new_n894), .B2(new_n888), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n887), .A2(new_n891), .A3(new_n895), .ZN(new_n902));
  OAI211_X1 g701(.A(KEYINPUT124), .B(new_n900), .C1(new_n901), .C2(new_n902), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n898), .A2(new_n903), .ZN(G1350gat));
  NAND3_X1  g703(.A1(new_n871), .A2(new_n207), .A3(new_n496), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n781), .A2(new_n496), .A3(new_n854), .ZN(new_n906));
  INV_X1    g705(.A(KEYINPUT61), .ZN(new_n907));
  AND3_X1   g706(.A1(new_n906), .A2(new_n907), .A3(G190gat), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n906), .B2(G190gat), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n905), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  XOR2_X1   g709(.A(new_n910), .B(KEYINPUT125), .Z(G1351gat));
  NOR2_X1   g710(.A1(new_n707), .A2(new_n853), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n841), .A2(new_n912), .ZN(new_n913));
  INV_X1    g712(.A(G197gat), .ZN(new_n914));
  NOR3_X1   g713(.A1(new_n913), .A2(new_n914), .A3(new_n620), .ZN(new_n915));
  AOI211_X1 g714(.A(new_n392), .B(new_n807), .C1(new_n865), .C2(new_n870), .ZN(new_n916));
  AOI21_X1  g715(.A(G197gat), .B1(new_n916), .B2(new_n619), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n915), .A2(new_n917), .ZN(G1352gat));
  XNOR2_X1  g717(.A(KEYINPUT126), .B(G204gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n841), .A2(new_n641), .A3(new_n912), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n738), .A2(new_n919), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n916), .A2(new_n921), .ZN(new_n922));
  AOI22_X1  g721(.A1(new_n919), .A2(new_n920), .B1(new_n922), .B2(KEYINPUT62), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n922), .A2(KEYINPUT62), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT127), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  NOR3_X1   g725(.A1(new_n922), .A2(KEYINPUT127), .A3(KEYINPUT62), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n923), .B1(new_n926), .B2(new_n927), .ZN(G1353gat));
  NAND3_X1  g727(.A1(new_n916), .A2(new_n277), .A3(new_n665), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n841), .A2(new_n665), .A3(new_n912), .ZN(new_n930));
  AND3_X1   g729(.A1(new_n930), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n931));
  AOI21_X1  g730(.A(KEYINPUT63), .B1(new_n930), .B2(G211gat), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n929), .B1(new_n931), .B2(new_n932), .ZN(G1354gat));
  OAI21_X1  g732(.A(G218gat), .B1(new_n913), .B2(new_n663), .ZN(new_n934));
  NAND3_X1  g733(.A1(new_n916), .A2(new_n278), .A3(new_n496), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n934), .A2(new_n935), .ZN(G1355gat));
endmodule


