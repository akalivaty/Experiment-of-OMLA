//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 1 0 0 1 0 0 1 0 1 0 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:40:13 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1289, new_n1290, new_n1291;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0008(.A1(new_n206), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND3_X1  g0010(.A1(KEYINPUT66), .A2(G1), .A3(G13), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(KEYINPUT66), .B1(G1), .B2(G13), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n210), .A2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(KEYINPUT0), .ZN(new_n218));
  NAND2_X1  g0018(.A1(G1), .A2(G20), .ZN(new_n219));
  OR3_X1    g0019(.A1(new_n219), .A2(KEYINPUT65), .A3(G13), .ZN(new_n220));
  OAI21_X1  g0020(.A(KEYINPUT65), .B1(new_n219), .B2(G13), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI211_X1 g0022(.A(new_n222), .B(G250), .C1(G257), .C2(G264), .ZN(new_n223));
  OAI21_X1  g0023(.A(new_n217), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(new_n218), .B2(new_n223), .ZN(new_n225));
  XOR2_X1   g0025(.A(new_n225), .B(KEYINPUT67), .Z(new_n226));
  AOI22_X1  g0026(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n227));
  INV_X1    g0027(.A(G77), .ZN(new_n228));
  INV_X1    g0028(.A(G244), .ZN(new_n229));
  INV_X1    g0029(.A(G107), .ZN(new_n230));
  INV_X1    g0030(.A(G264), .ZN(new_n231));
  OAI221_X1 g0031(.A(new_n227), .B1(new_n228), .B2(new_n229), .C1(new_n230), .C2(new_n231), .ZN(new_n232));
  AOI22_X1  g0032(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n233));
  AOI22_X1  g0033(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n234));
  NAND2_X1  g0034(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  OAI21_X1  g0035(.A(new_n219), .B1(new_n232), .B2(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  NOR2_X1   g0038(.A1(new_n226), .A2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G238), .B(G244), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G232), .ZN(new_n241));
  XNOR2_X1  g0041(.A(KEYINPUT2), .B(G226), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XOR2_X1   g0043(.A(G264), .B(G270), .Z(new_n244));
  XNOR2_X1  g0044(.A(G250), .B(G257), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n243), .B(new_n246), .ZN(G358));
  XOR2_X1   g0047(.A(G87), .B(G97), .Z(new_n248));
  XNOR2_X1  g0048(.A(G107), .B(G116), .ZN(new_n249));
  XNOR2_X1  g0049(.A(new_n248), .B(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G50), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(G68), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n203), .A2(G50), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  XNOR2_X1  g0054(.A(G58), .B(G77), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n250), .B(new_n256), .ZN(G351));
  INV_X1    g0057(.A(new_n213), .ZN(new_n258));
  NAND3_X1  g0058(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(new_n211), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G1), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n251), .B1(new_n261), .B2(G20), .ZN(new_n265));
  AOI22_X1  g0065(.A1(new_n264), .A2(new_n265), .B1(new_n251), .B2(new_n263), .ZN(new_n266));
  OAI21_X1  g0066(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT8), .B(G58), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n215), .A2(G33), .ZN(new_n270));
  INV_X1    g0070(.A(new_n270), .ZN(new_n271));
  NOR2_X1   g0071(.A1(G20), .A2(G33), .ZN(new_n272));
  AOI22_X1  g0072(.A1(new_n269), .A2(new_n271), .B1(G150), .B2(new_n272), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n267), .A2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(new_n260), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n266), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g0076(.A(new_n276), .B(KEYINPUT9), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n278), .A2(KEYINPUT69), .ZN(new_n279));
  INV_X1    g0079(.A(KEYINPUT69), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n280), .A2(G33), .A3(G41), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  INV_X1    g0082(.A(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n279), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  AND2_X1   g0084(.A1(new_n284), .A2(G274), .ZN(new_n285));
  INV_X1    g0085(.A(G41), .ZN(new_n286));
  INV_X1    g0086(.A(G45), .ZN(new_n287));
  AOI21_X1  g0087(.A(G1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n282), .B1(KEYINPUT69), .B2(new_n278), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n288), .B1(new_n289), .B2(new_n281), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n285), .A2(new_n288), .B1(G226), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  INV_X1    g0092(.A(G1698), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n292), .A2(G222), .A3(new_n293), .ZN(new_n294));
  XNOR2_X1  g0094(.A(new_n294), .B(KEYINPUT70), .ZN(new_n295));
  INV_X1    g0095(.A(G33), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(KEYINPUT3), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT3), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G33), .ZN(new_n299));
  NAND2_X1  g0099(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  NOR2_X1   g0100(.A1(new_n300), .A2(new_n293), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G223), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n302), .B1(new_n228), .B2(new_n292), .ZN(new_n303));
  NOR2_X1   g0103(.A1(new_n295), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n278), .B1(new_n212), .B2(new_n213), .ZN(new_n305));
  OAI211_X1 g0105(.A(G190), .B(new_n291), .C1(new_n304), .C2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  INV_X1    g0107(.A(new_n291), .ZN(new_n308));
  OAI21_X1  g0108(.A(G200), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n277), .A2(new_n306), .A3(new_n309), .ZN(new_n310));
  XNOR2_X1  g0110(.A(new_n310), .B(KEYINPUT10), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n301), .A2(G238), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n292), .A2(G232), .A3(new_n293), .ZN(new_n313));
  OAI211_X1 g0113(.A(new_n312), .B(new_n313), .C1(new_n230), .C2(new_n292), .ZN(new_n314));
  INV_X1    g0114(.A(new_n305), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n284), .A2(G274), .A3(new_n288), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n290), .A2(G244), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G179), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n269), .A2(new_n272), .B1(G20), .B2(G77), .ZN(new_n323));
  XNOR2_X1  g0123(.A(KEYINPUT15), .B(G87), .ZN(new_n324));
  INV_X1    g0124(.A(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(new_n271), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n275), .B1(new_n323), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n327), .B1(new_n228), .B2(new_n263), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n261), .A2(G20), .ZN(new_n329));
  NAND3_X1  g0129(.A1(new_n264), .A2(G77), .A3(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n319), .A2(new_n332), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n322), .A2(new_n331), .A3(new_n333), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  AOI22_X1  g0135(.A1(new_n320), .A2(G190), .B1(new_n331), .B2(KEYINPUT72), .ZN(new_n336));
  INV_X1    g0136(.A(new_n331), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT72), .ZN(new_n338));
  AOI22_X1  g0138(.A1(new_n337), .A2(new_n338), .B1(G200), .B2(new_n319), .ZN(new_n339));
  AOI21_X1  g0139(.A(new_n335), .B1(new_n336), .B2(new_n339), .ZN(new_n340));
  AOI21_X1  g0140(.A(KEYINPUT74), .B1(new_n263), .B2(new_n203), .ZN(new_n341));
  XNOR2_X1  g0141(.A(new_n341), .B(KEYINPUT12), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n264), .A2(G68), .A3(new_n329), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT75), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n272), .A2(G50), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n347), .B1(new_n215), .B2(G68), .C1(new_n228), .C2(new_n270), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n260), .ZN(new_n349));
  XNOR2_X1  g0149(.A(new_n349), .B(KEYINPUT11), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n342), .A2(KEYINPUT75), .A3(new_n343), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n346), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  MUX2_X1   g0152(.A(G226), .B(G232), .S(G1698), .Z(new_n353));
  NAND2_X1  g0153(.A1(new_n353), .A2(new_n292), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G97), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n356), .A2(new_n315), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT13), .ZN(new_n358));
  INV_X1    g0158(.A(new_n288), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n284), .A2(G238), .A3(new_n359), .ZN(new_n360));
  NAND4_X1  g0160(.A1(new_n357), .A2(new_n358), .A3(new_n317), .A4(new_n360), .ZN(new_n361));
  AOI22_X1  g0161(.A1(new_n353), .A2(new_n292), .B1(G33), .B2(G97), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n317), .B(new_n360), .C1(new_n362), .C2(new_n305), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n363), .A2(KEYINPUT13), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n361), .A2(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(KEYINPUT14), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(new_n366), .A3(G169), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n367), .B1(new_n321), .B2(new_n365), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n366), .B1(new_n365), .B2(G169), .ZN(new_n369));
  OAI21_X1  g0169(.A(new_n352), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n352), .B1(G200), .B2(new_n365), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n361), .A2(new_n364), .A3(G190), .ZN(new_n372));
  XNOR2_X1  g0172(.A(new_n372), .B(KEYINPUT73), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n370), .A2(new_n374), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n307), .A2(new_n308), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT71), .B1(new_n376), .B2(G169), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n376), .A2(new_n321), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n376), .A2(KEYINPUT71), .A3(new_n321), .ZN(new_n380));
  NAND3_X1  g0180(.A1(new_n379), .A2(new_n276), .A3(new_n380), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n311), .A2(new_n340), .A3(new_n375), .A4(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT79), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n204), .A2(new_n205), .A3(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n272), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT76), .B1(new_n298), .B2(G33), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT76), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n389), .A2(new_n296), .A3(KEYINPUT3), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n388), .A2(new_n390), .A3(new_n299), .ZN(new_n391));
  INV_X1    g0191(.A(KEYINPUT7), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n391), .A2(new_n392), .A3(new_n215), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G68), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n392), .B1(new_n391), .B2(new_n215), .ZN(new_n395));
  OAI211_X1 g0195(.A(KEYINPUT16), .B(new_n387), .C1(new_n394), .C2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT16), .ZN(new_n397));
  OAI21_X1  g0197(.A(new_n392), .B1(new_n292), .B2(G20), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n300), .A2(KEYINPUT7), .A3(new_n215), .ZN(new_n399));
  AOI21_X1  g0199(.A(new_n203), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n386), .A2(G20), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n272), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  OAI21_X1  g0203(.A(new_n397), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  NAND3_X1  g0204(.A1(new_n396), .A2(new_n404), .A3(new_n260), .ZN(new_n405));
  INV_X1    g0205(.A(G200), .ZN(new_n406));
  NOR2_X1   g0206(.A1(G223), .A2(G1698), .ZN(new_n407));
  INV_X1    g0207(.A(G226), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n407), .B1(new_n408), .B2(G1698), .ZN(new_n409));
  NAND4_X1  g0209(.A1(new_n409), .A2(new_n299), .A3(new_n388), .A4(new_n390), .ZN(new_n410));
  NAND2_X1  g0210(.A1(G33), .A2(G87), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n305), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n284), .A2(G232), .A3(new_n359), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n317), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n406), .B1(new_n412), .B2(new_n414), .ZN(new_n415));
  NAND2_X1  g0215(.A1(new_n408), .A2(G1698), .ZN(new_n416));
  OAI21_X1  g0216(.A(new_n416), .B1(G223), .B2(G1698), .ZN(new_n417));
  OAI21_X1  g0217(.A(new_n411), .B1(new_n391), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(new_n315), .ZN(new_n419));
  INV_X1    g0219(.A(G190), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n419), .A2(new_n420), .A3(new_n317), .A4(new_n413), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n415), .A2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n268), .B1(new_n261), .B2(G20), .ZN(new_n423));
  AOI22_X1  g0223(.A1(new_n264), .A2(new_n423), .B1(new_n263), .B2(new_n268), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n405), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(KEYINPUT17), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  NAND4_X1  g0227(.A1(new_n405), .A2(new_n422), .A3(KEYINPUT17), .A4(new_n424), .ZN(new_n428));
  AND2_X1   g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g0229(.A1(new_n405), .A2(new_n424), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n332), .B1(new_n412), .B2(new_n414), .ZN(new_n431));
  AND2_X1   g0231(.A1(new_n317), .A2(new_n413), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(new_n321), .A3(new_n419), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT77), .ZN(new_n434));
  AND3_X1   g0234(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n434), .B1(new_n431), .B2(new_n433), .ZN(new_n436));
  OAI21_X1  g0236(.A(KEYINPUT78), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NOR3_X1   g0237(.A1(new_n412), .A2(new_n414), .A3(G179), .ZN(new_n438));
  AOI21_X1  g0238(.A(G169), .B1(new_n432), .B2(new_n419), .ZN(new_n439));
  OAI21_X1  g0239(.A(KEYINPUT77), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT78), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n431), .A2(new_n433), .A3(new_n434), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n430), .B1(new_n437), .B2(new_n443), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT18), .ZN(new_n445));
  OAI21_X1  g0245(.A(new_n429), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  AOI211_X1 g0246(.A(KEYINPUT18), .B(new_n430), .C1(new_n437), .C2(new_n443), .ZN(new_n447));
  NOR2_X1   g0247(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n383), .A2(new_n384), .A3(new_n448), .ZN(new_n449));
  INV_X1    g0249(.A(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(KEYINPUT79), .B1(new_n382), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n449), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT24), .ZN(new_n454));
  NAND4_X1  g0254(.A1(new_n388), .A2(new_n390), .A3(new_n215), .A4(new_n299), .ZN(new_n455));
  NAND2_X1  g0255(.A1(KEYINPUT22), .A2(G87), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G87), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n458), .A2(G20), .ZN(new_n459));
  AOI21_X1  g0259(.A(KEYINPUT22), .B1(new_n292), .B2(new_n459), .ZN(new_n460));
  OAI21_X1  g0260(.A(KEYINPUT87), .B1(new_n457), .B2(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(KEYINPUT22), .ZN(new_n462));
  INV_X1    g0262(.A(new_n459), .ZN(new_n463));
  OAI21_X1  g0263(.A(new_n462), .B1(new_n300), .B2(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT87), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n455), .C2(new_n456), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(G33), .A2(G116), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n468), .A2(G20), .ZN(new_n469));
  AOI21_X1  g0269(.A(KEYINPUT23), .B1(new_n230), .B2(G20), .ZN(new_n470));
  INV_X1    g0270(.A(new_n470), .ZN(new_n471));
  NAND3_X1  g0271(.A1(new_n230), .A2(KEYINPUT23), .A3(G20), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n469), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  AOI21_X1  g0273(.A(new_n454), .B1(new_n467), .B2(new_n473), .ZN(new_n474));
  INV_X1    g0274(.A(new_n473), .ZN(new_n475));
  AOI211_X1 g0275(.A(KEYINPUT24), .B(new_n475), .C1(new_n461), .C2(new_n466), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n260), .B1(new_n474), .B2(new_n476), .ZN(new_n477));
  OR2_X1    g0277(.A1(G250), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G257), .B2(new_n293), .ZN(new_n479));
  INV_X1    g0279(.A(G294), .ZN(new_n480));
  OAI22_X1  g0280(.A1(new_n391), .A2(new_n479), .B1(new_n296), .B2(new_n480), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n481), .A2(new_n315), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n261), .B(G45), .C1(new_n286), .C2(KEYINPUT5), .ZN(new_n483));
  INV_X1    g0283(.A(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT82), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT5), .ZN(new_n486));
  OAI21_X1  g0286(.A(new_n485), .B1(new_n486), .B2(G41), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n286), .A2(KEYINPUT82), .A3(KEYINPUT5), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI22_X1  g0289(.A1(new_n484), .A2(new_n489), .B1(new_n289), .B2(new_n281), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G264), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n483), .B1(new_n487), .B2(new_n488), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n285), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n482), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n420), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G200), .B2(new_n494), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n261), .A2(G33), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT80), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AOI21_X1  g0299(.A(KEYINPUT80), .B1(new_n261), .B2(G33), .ZN(new_n500));
  NOR4_X1   g0300(.A1(new_n260), .A2(new_n499), .A3(new_n263), .A4(new_n500), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT25), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n262), .B2(G107), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n263), .A2(KEYINPUT25), .A3(new_n230), .ZN(new_n504));
  AOI22_X1  g0304(.A1(new_n501), .A2(G107), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n477), .A2(new_n496), .A3(new_n505), .ZN(new_n506));
  INV_X1    g0306(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n494), .A2(new_n321), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n508), .B1(G169), .B2(new_n494), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n509), .B1(new_n477), .B2(new_n505), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  AND2_X1   g0312(.A1(KEYINPUT4), .A2(G244), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n297), .A2(new_n299), .A3(new_n513), .A4(new_n293), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n297), .A2(new_n299), .A3(G250), .A4(G1698), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G283), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT4), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n229), .A2(G1698), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n518), .B1(new_n391), .B2(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n315), .ZN(new_n523));
  AOI22_X1  g0323(.A1(new_n490), .A2(G257), .B1(new_n285), .B2(new_n492), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n272), .A2(G77), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT6), .ZN(new_n527));
  INV_X1    g0327(.A(G97), .ZN(new_n528));
  NOR3_X1   g0328(.A1(new_n527), .A2(new_n528), .A3(G107), .ZN(new_n529));
  XNOR2_X1  g0329(.A(G97), .B(G107), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n529), .B1(new_n527), .B2(new_n530), .ZN(new_n531));
  OAI21_X1  g0331(.A(new_n526), .B1(new_n531), .B2(new_n215), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n230), .B1(new_n398), .B2(new_n399), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n260), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n262), .A2(G97), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n535), .B1(new_n501), .B2(G97), .ZN(new_n536));
  AOI22_X1  g0336(.A1(new_n525), .A2(new_n332), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n305), .B1(new_n517), .B2(new_n521), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT81), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  AOI211_X1 g0340(.A(KEYINPUT81), .B(new_n305), .C1(new_n517), .C2(new_n521), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n321), .B(new_n524), .C1(new_n540), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  XNOR2_X1  g0343(.A(new_n538), .B(new_n539), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n406), .B1(new_n544), .B2(new_n524), .ZN(new_n545));
  OAI211_X1 g0345(.A(new_n534), .B(new_n536), .C1(new_n525), .C2(new_n420), .ZN(new_n546));
  OAI21_X1  g0346(.A(new_n543), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n229), .A2(G1698), .ZN(new_n548));
  OAI21_X1  g0348(.A(new_n548), .B1(G238), .B2(G1698), .ZN(new_n549));
  OAI21_X1  g0349(.A(new_n468), .B1(new_n391), .B2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n315), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n261), .A2(G45), .ZN(new_n552));
  MUX2_X1   g0352(.A(G274), .B(G250), .S(new_n552), .Z(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n284), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n406), .B1(new_n551), .B2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT19), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n458), .A2(new_n528), .A3(new_n230), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n355), .A2(new_n215), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR3_X1   g0360(.A1(new_n270), .A2(KEYINPUT19), .A3(new_n528), .ZN(new_n561));
  OAI22_X1  g0361(.A1(new_n203), .A2(new_n455), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  AOI22_X1  g0362(.A1(new_n562), .A2(new_n260), .B1(new_n263), .B2(new_n324), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n501), .A2(G87), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n556), .A2(KEYINPUT83), .A3(new_n563), .A4(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(KEYINPUT83), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n563), .A2(new_n564), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n566), .B1(new_n567), .B2(new_n555), .ZN(new_n568));
  AOI22_X1  g0368(.A1(new_n315), .A2(new_n550), .B1(new_n553), .B2(new_n284), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(G190), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n565), .A2(new_n568), .A3(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n501), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n563), .B1(new_n324), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n551), .A2(new_n554), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n574), .A2(new_n332), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n569), .A2(new_n321), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n573), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n571), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n512), .B1(new_n547), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n490), .A2(G270), .B1(new_n285), .B2(new_n492), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n300), .A2(G303), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n231), .A2(G1698), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(G257), .B2(G1698), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n581), .B1(new_n391), .B2(new_n583), .ZN(new_n584));
  INV_X1    g0384(.A(KEYINPUT85), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n315), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g0386(.A1(G257), .A2(G1698), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n587), .B1(new_n231), .B2(G1698), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n588), .A2(new_n299), .A3(new_n388), .A4(new_n390), .ZN(new_n589));
  AOI21_X1  g0389(.A(KEYINPUT85), .B1(new_n589), .B2(new_n581), .ZN(new_n590));
  OAI21_X1  g0390(.A(new_n580), .B1(new_n586), .B2(new_n590), .ZN(new_n591));
  AOI21_X1  g0391(.A(G20), .B1(G33), .B2(G283), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n296), .A2(G97), .ZN(new_n593));
  INV_X1    g0393(.A(G116), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n592), .A2(new_n593), .B1(G20), .B2(new_n594), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n260), .A2(new_n595), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n260), .A2(KEYINPUT20), .A3(new_n595), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NOR2_X1   g0400(.A1(new_n499), .A2(new_n500), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n264), .A2(G116), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n263), .A2(new_n594), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n600), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  NAND4_X1  g0404(.A1(new_n591), .A2(new_n604), .A3(KEYINPUT21), .A4(G169), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n584), .A2(new_n585), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n589), .A2(KEYINPUT85), .A3(new_n581), .ZN(new_n607));
  NAND3_X1  g0407(.A1(new_n606), .A2(new_n315), .A3(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n604), .A2(new_n608), .A3(G179), .A4(new_n580), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n604), .B1(new_n591), .B2(G200), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n611), .B1(new_n420), .B2(new_n591), .ZN(new_n612));
  AOI22_X1  g0412(.A1(new_n598), .A2(new_n599), .B1(new_n594), .B2(new_n263), .ZN(new_n613));
  AOI21_X1  g0413(.A(new_n332), .B1(new_n613), .B2(new_n602), .ZN(new_n614));
  AOI211_X1 g0414(.A(KEYINPUT86), .B(KEYINPUT21), .C1(new_n614), .C2(new_n591), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT86), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n591), .A2(G169), .A3(new_n604), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT21), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n616), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  OAI211_X1 g0419(.A(new_n610), .B(new_n612), .C1(new_n615), .C2(new_n619), .ZN(new_n620));
  INV_X1    g0420(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(new_n524), .B1(new_n540), .B2(new_n541), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n622), .A2(G200), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n534), .A2(new_n536), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n490), .A2(G257), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n625), .A2(new_n493), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n626), .A2(new_n538), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n624), .B1(new_n627), .B2(G190), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n623), .A2(new_n628), .B1(new_n542), .B2(new_n537), .ZN(new_n629));
  NAND4_X1  g0429(.A1(new_n629), .A2(KEYINPUT84), .A3(new_n577), .A4(new_n571), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n511), .A2(new_n579), .A3(new_n621), .A4(new_n630), .ZN(new_n631));
  NOR2_X1   g0431(.A1(new_n453), .A2(new_n631), .ZN(G372));
  INV_X1    g0432(.A(new_n381), .ZN(new_n633));
  AOI21_X1  g0433(.A(new_n334), .B1(new_n373), .B2(new_n371), .ZN(new_n634));
  INV_X1    g0434(.A(new_n370), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n429), .B1(new_n634), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n440), .A2(new_n442), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n405), .A2(new_n424), .ZN(new_n638));
  AND3_X1   g0438(.A1(new_n637), .A2(new_n445), .A3(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n445), .B1(new_n637), .B2(new_n638), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n636), .A2(new_n641), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n633), .B1(new_n642), .B2(new_n311), .ZN(new_n643));
  OAI21_X1  g0443(.A(KEYINPUT26), .B1(new_n578), .B2(new_n543), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n556), .A2(new_n563), .A3(new_n564), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n645), .A2(KEYINPUT88), .ZN(new_n646));
  OR3_X1    g0446(.A1(new_n567), .A2(new_n555), .A3(KEYINPUT88), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n646), .A2(new_n647), .A3(new_n570), .ZN(new_n648));
  INV_X1    g0448(.A(new_n543), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT26), .ZN(new_n650));
  NAND4_X1  g0450(.A1(new_n648), .A2(new_n649), .A3(new_n650), .A4(new_n577), .ZN(new_n651));
  XNOR2_X1  g0451(.A(new_n577), .B(KEYINPUT89), .ZN(new_n652));
  AND3_X1   g0452(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  NAND4_X1  g0453(.A1(new_n629), .A2(new_n648), .A3(new_n506), .A4(new_n577), .ZN(new_n654));
  INV_X1    g0454(.A(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n605), .A2(new_n609), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n617), .A2(new_n618), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n657), .A2(KEYINPUT86), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n617), .A2(new_n616), .A3(new_n618), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n656), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g0460(.A(new_n510), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n655), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n653), .A2(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n664), .ZN(new_n665));
  OAI21_X1  g0465(.A(new_n643), .B1(new_n453), .B2(new_n665), .ZN(G369));
  NAND3_X1  g0466(.A1(new_n261), .A2(new_n215), .A3(G13), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n667), .A2(KEYINPUT90), .A3(KEYINPUT27), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(KEYINPUT90), .B1(new_n667), .B2(KEYINPUT27), .ZN(new_n670));
  OAI221_X1 g0470(.A(G213), .B1(KEYINPUT27), .B2(new_n667), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(G343), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g0473(.A1(new_n604), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n621), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(new_n660), .B2(new_n674), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n676), .A2(G330), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  AND2_X1   g0478(.A1(new_n477), .A2(new_n505), .ZN(new_n679));
  INV_X1    g0479(.A(new_n673), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n511), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n681), .B1(new_n661), .B2(new_n680), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n678), .A2(new_n682), .ZN(new_n683));
  XNOR2_X1  g0483(.A(new_n683), .B(KEYINPUT91), .ZN(new_n684));
  NOR2_X1   g0484(.A1(new_n660), .A2(new_n673), .ZN(new_n685));
  AOI22_X1  g0485(.A1(new_n685), .A2(new_n511), .B1(new_n510), .B2(new_n680), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n684), .A2(new_n686), .ZN(G399));
  INV_X1    g0487(.A(new_n222), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  NOR2_X1   g0489(.A1(new_n558), .A2(G116), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR3_X1   g0491(.A1(new_n689), .A2(new_n261), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g0492(.A(new_n692), .B1(new_n210), .B2(new_n689), .ZN(new_n693));
  XNOR2_X1  g0493(.A(new_n693), .B(KEYINPUT92), .ZN(new_n694));
  XOR2_X1   g0494(.A(new_n694), .B(KEYINPUT28), .Z(new_n695));
  INV_X1    g0495(.A(G330), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n620), .A2(new_n507), .A3(new_n510), .ZN(new_n697));
  NAND4_X1  g0497(.A1(new_n697), .A2(new_n579), .A3(new_n630), .A4(new_n680), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n580), .A2(G179), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n482), .A2(new_n491), .ZN(new_n700));
  NOR3_X1   g0500(.A1(new_n699), .A2(new_n700), .A3(new_n574), .ZN(new_n701));
  NAND4_X1  g0501(.A1(new_n701), .A2(KEYINPUT30), .A3(new_n627), .A4(new_n608), .ZN(new_n702));
  INV_X1    g0502(.A(KEYINPUT30), .ZN(new_n703));
  INV_X1    g0503(.A(new_n700), .ZN(new_n704));
  NAND4_X1  g0504(.A1(new_n704), .A2(G179), .A3(new_n569), .A4(new_n580), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n627), .A2(new_n608), .ZN(new_n706));
  OAI21_X1  g0506(.A(new_n703), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NOR3_X1   g0507(.A1(new_n494), .A2(G179), .A3(new_n569), .ZN(new_n708));
  NAND3_X1  g0508(.A1(new_n708), .A2(new_n622), .A3(new_n591), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n702), .A2(new_n707), .A3(new_n709), .ZN(new_n710));
  AND3_X1   g0510(.A1(new_n710), .A2(KEYINPUT31), .A3(new_n673), .ZN(new_n711));
  AOI21_X1  g0511(.A(KEYINPUT31), .B1(new_n710), .B2(new_n673), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n696), .B1(new_n698), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n662), .A2(KEYINPUT94), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n610), .B1(new_n615), .B2(new_n619), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n716), .A2(new_n510), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT94), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  OAI21_X1  g0519(.A(new_n655), .B1(new_n715), .B2(new_n719), .ZN(new_n720));
  XNOR2_X1  g0520(.A(new_n652), .B(KEYINPUT93), .ZN(new_n721));
  NAND4_X1  g0521(.A1(new_n649), .A2(new_n650), .A3(new_n577), .A4(new_n571), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n648), .A2(new_n577), .ZN(new_n723));
  OAI21_X1  g0523(.A(KEYINPUT26), .B1(new_n723), .B2(new_n543), .ZN(new_n724));
  AND3_X1   g0524(.A1(new_n721), .A2(new_n722), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g0525(.A(new_n673), .B1(new_n720), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT29), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n673), .B1(new_n653), .B2(new_n663), .ZN(new_n728));
  OR2_X1    g0528(.A1(new_n728), .A2(KEYINPUT29), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n714), .B1(new_n727), .B2(new_n729), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n695), .B1(new_n730), .B2(G1), .ZN(G364));
  XOR2_X1   g0531(.A(new_n677), .B(KEYINPUT95), .Z(new_n732));
  INV_X1    g0532(.A(G13), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(G20), .ZN(new_n734));
  AOI21_X1  g0534(.A(new_n261), .B1(new_n734), .B2(G45), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n689), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OAI211_X1 g0538(.A(new_n732), .B(new_n738), .C1(G330), .C2(new_n676), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  XOR2_X1   g0542(.A(new_n742), .B(KEYINPUT97), .Z(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n332), .A2(KEYINPUT98), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n215), .B1(KEYINPUT98), .B2(new_n332), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n214), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n744), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n222), .A2(G355), .A3(new_n292), .ZN(new_n751));
  INV_X1    g0551(.A(new_n391), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n688), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g0553(.A(new_n753), .B1(G45), .B2(new_n209), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n256), .A2(new_n287), .ZN(new_n755));
  OAI221_X1 g0555(.A(new_n751), .B1(G116), .B2(new_n222), .C1(new_n754), .C2(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n750), .B1(new_n756), .B2(KEYINPUT96), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(KEYINPUT96), .B2(new_n756), .ZN(new_n758));
  NAND3_X1  g0558(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n759), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(new_n215), .A2(G179), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G190), .A3(G200), .ZN(new_n763));
  OAI22_X1  g0563(.A1(new_n761), .A2(new_n203), .B1(new_n763), .B2(new_n458), .ZN(new_n764));
  NAND3_X1  g0564(.A1(new_n762), .A2(new_n420), .A3(G200), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  AOI211_X1 g0566(.A(new_n300), .B(new_n764), .C1(G107), .C2(new_n766), .ZN(new_n767));
  NOR4_X1   g0567(.A1(new_n215), .A2(new_n321), .A3(new_n420), .A4(G200), .ZN(new_n768));
  INV_X1    g0568(.A(KEYINPUT99), .ZN(new_n769));
  AND2_X1   g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n768), .A2(new_n769), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR4_X1   g0572(.A1(new_n215), .A2(new_n321), .A3(G190), .A4(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n774));
  INV_X1    g0574(.A(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n773), .A2(KEYINPUT100), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI221_X1 g0577(.A(new_n767), .B1(new_n202), .B2(new_n772), .C1(new_n228), .C2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(G179), .A2(G200), .ZN(new_n779));
  NAND3_X1  g0579(.A1(new_n779), .A2(G20), .A3(new_n420), .ZN(new_n780));
  INV_X1    g0580(.A(G159), .ZN(new_n781));
  NOR2_X1   g0581(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT32), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n759), .A2(new_n420), .ZN(new_n784));
  INV_X1    g0584(.A(new_n784), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n215), .B1(new_n779), .B2(G190), .ZN(new_n786));
  OAI221_X1 g0586(.A(new_n783), .B1(new_n251), .B2(new_n785), .C1(new_n528), .C2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n773), .ZN(new_n788));
  INV_X1    g0588(.A(G311), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(new_n780), .ZN(new_n791));
  AOI211_X1 g0591(.A(new_n292), .B(new_n790), .C1(G329), .C2(new_n791), .ZN(new_n792));
  XNOR2_X1  g0592(.A(KEYINPUT33), .B(G317), .ZN(new_n793));
  OR2_X1    g0593(.A1(new_n793), .A2(KEYINPUT101), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n793), .A2(KEYINPUT101), .ZN(new_n795));
  NAND3_X1  g0595(.A1(new_n794), .A2(new_n760), .A3(new_n795), .ZN(new_n796));
  INV_X1    g0596(.A(G322), .ZN(new_n797));
  OAI211_X1 g0597(.A(new_n792), .B(new_n796), .C1(new_n797), .C2(new_n772), .ZN(new_n798));
  INV_X1    g0598(.A(new_n786), .ZN(new_n799));
  AOI22_X1  g0599(.A1(new_n799), .A2(G294), .B1(G326), .B2(new_n784), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  INV_X1    g0601(.A(G303), .ZN(new_n802));
  OAI221_X1 g0602(.A(new_n800), .B1(new_n801), .B2(new_n765), .C1(new_n802), .C2(new_n763), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n778), .A2(new_n787), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n738), .B1(new_n804), .B2(new_n748), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n758), .B(new_n805), .C1(new_n676), .C2(new_n743), .ZN(new_n806));
  XNOR2_X1  g0606(.A(new_n806), .B(KEYINPUT102), .ZN(new_n807));
  NAND2_X1  g0607(.A1(new_n739), .A2(new_n807), .ZN(G396));
  NAND2_X1  g0608(.A1(new_n335), .A2(new_n680), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n339), .A2(new_n336), .B1(new_n331), .B2(new_n673), .ZN(new_n810));
  OAI21_X1  g0610(.A(new_n809), .B1(new_n810), .B2(new_n335), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n665), .B2(new_n673), .ZN(new_n812));
  MUX2_X1   g0612(.A(new_n673), .B(new_n810), .S(new_n334), .Z(new_n813));
  NOR2_X1   g0613(.A1(new_n717), .A2(new_n654), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n644), .A2(new_n651), .A3(new_n652), .ZN(new_n815));
  OAI211_X1 g0615(.A(new_n813), .B(new_n680), .C1(new_n814), .C2(new_n815), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n714), .B1(new_n812), .B2(new_n816), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n817), .A2(new_n737), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n812), .A2(new_n714), .A3(new_n816), .ZN(new_n819));
  AND2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n748), .ZN(new_n821));
  NAND2_X1  g0621(.A1(new_n821), .A2(new_n741), .ZN(new_n822));
  OAI22_X1  g0622(.A1(new_n786), .A2(new_n528), .B1(new_n780), .B2(new_n789), .ZN(new_n823));
  INV_X1    g0623(.A(new_n777), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n823), .B1(new_n824), .B2(G116), .ZN(new_n825));
  OAI22_X1  g0625(.A1(new_n761), .A2(new_n801), .B1(new_n785), .B2(new_n802), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n826), .B1(G87), .B2(new_n766), .ZN(new_n827));
  OAI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(new_n480), .C2(new_n772), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n300), .B1(new_n763), .B2(new_n230), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT103), .Z(new_n830));
  NOR2_X1   g0630(.A1(new_n828), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n766), .A2(G68), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n251), .B2(new_n763), .C1(new_n202), .C2(new_n786), .ZN(new_n833));
  AOI211_X1 g0633(.A(new_n391), .B(new_n833), .C1(G132), .C2(new_n791), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT104), .Z(new_n835));
  AOI22_X1  g0635(.A1(G137), .A2(new_n784), .B1(new_n760), .B2(G150), .ZN(new_n836));
  INV_X1    g0636(.A(G143), .ZN(new_n837));
  OAI221_X1 g0637(.A(new_n836), .B1(new_n777), .B2(new_n781), .C1(new_n772), .C2(new_n837), .ZN(new_n838));
  XOR2_X1   g0638(.A(new_n838), .B(KEYINPUT34), .Z(new_n839));
  INV_X1    g0639(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n831), .B1(new_n835), .B2(new_n840), .ZN(new_n841));
  OAI221_X1 g0641(.A(new_n737), .B1(G77), .B2(new_n822), .C1(new_n841), .C2(new_n821), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n740), .B2(new_n811), .ZN(new_n843));
  NOR2_X1   g0643(.A1(new_n820), .A2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(G384));
  NOR2_X1   g0645(.A1(new_n734), .A2(new_n261), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n713), .B1(new_n631), .B2(new_n673), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT106), .ZN(new_n848));
  AND3_X1   g0648(.A1(new_n352), .A2(new_n848), .A3(new_n673), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n848), .B1(new_n352), .B2(new_n673), .ZN(new_n850));
  NOR2_X1   g0650(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n375), .A2(new_n851), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n370), .A2(new_n374), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n853), .B1(new_n850), .B2(new_n849), .ZN(new_n854));
  AOI21_X1  g0654(.A(new_n811), .B1(new_n852), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n847), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(KEYINPUT110), .ZN(new_n857));
  INV_X1    g0657(.A(KEYINPUT38), .ZN(new_n858));
  INV_X1    g0658(.A(new_n671), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n638), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n860), .A2(new_n425), .ZN(new_n861));
  NOR3_X1   g0661(.A1(new_n444), .A2(KEYINPUT37), .A3(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT107), .ZN(new_n863));
  OAI21_X1  g0663(.A(new_n387), .B1(new_n394), .B2(new_n395), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(new_n397), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n865), .A2(new_n260), .A3(new_n396), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n424), .A2(new_n866), .B1(new_n440), .B2(new_n442), .ZN(new_n867));
  AND3_X1   g0667(.A1(new_n405), .A2(new_n422), .A3(new_n424), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n863), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n866), .A2(new_n424), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n637), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(KEYINPUT107), .A3(new_n425), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n671), .B1(new_n866), .B2(new_n424), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n869), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g0675(.A(new_n862), .B1(new_n875), .B2(KEYINPUT37), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n427), .A2(new_n428), .ZN(new_n877));
  NOR3_X1   g0677(.A1(new_n435), .A2(new_n436), .A3(KEYINPUT78), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n441), .B1(new_n440), .B2(new_n442), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n638), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n877), .B1(new_n880), .B2(KEYINPUT18), .ZN(new_n881));
  INV_X1    g0681(.A(new_n447), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n874), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n858), .B1(new_n876), .B2(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n873), .B1(new_n446), .B2(new_n447), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT37), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n868), .B1(new_n637), .B2(new_n870), .ZN(new_n887));
  AOI21_X1  g0687(.A(new_n873), .B1(new_n887), .B2(KEYINPUT107), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n886), .B1(new_n888), .B2(new_n869), .ZN(new_n889));
  OAI211_X1 g0689(.A(new_n885), .B(KEYINPUT38), .C1(new_n889), .C2(new_n862), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n884), .A2(KEYINPUT108), .A3(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT108), .ZN(new_n892));
  OAI211_X1 g0692(.A(new_n892), .B(new_n858), .C1(new_n876), .C2(new_n883), .ZN(new_n893));
  INV_X1    g0693(.A(KEYINPUT110), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n847), .A2(new_n855), .A3(new_n894), .ZN(new_n895));
  NAND4_X1  g0695(.A1(new_n857), .A2(new_n891), .A3(new_n893), .A4(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT40), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n860), .A2(new_n425), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n637), .A2(new_n638), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n886), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n862), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n860), .B1(new_n641), .B2(new_n429), .ZN(new_n903));
  OAI21_X1  g0703(.A(new_n858), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n890), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(new_n905), .ZN(new_n906));
  NAND3_X1  g0706(.A1(new_n847), .A2(new_n855), .A3(KEYINPUT40), .ZN(new_n907));
  OAI21_X1  g0707(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  XOR2_X1   g0708(.A(new_n908), .B(KEYINPUT111), .Z(new_n909));
  AND2_X1   g0709(.A1(new_n452), .A2(new_n847), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n696), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n911), .B1(new_n909), .B2(new_n910), .ZN(new_n912));
  XOR2_X1   g0712(.A(new_n912), .B(KEYINPUT112), .Z(new_n913));
  INV_X1    g0713(.A(KEYINPUT39), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n890), .A2(new_n914), .A3(new_n904), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT109), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n890), .A2(new_n904), .A3(KEYINPUT109), .A4(new_n914), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g0719(.A1(new_n891), .A2(KEYINPUT39), .A3(new_n893), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n635), .A2(new_n680), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n852), .A2(new_n854), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n809), .B(KEYINPUT105), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n926), .B1(new_n816), .B2(new_n928), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(new_n891), .A3(new_n893), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n671), .B1(new_n639), .B2(new_n640), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n924), .A2(new_n933), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n727), .A2(new_n452), .A3(new_n729), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n643), .ZN(new_n936));
  XNOR2_X1  g0736(.A(new_n934), .B(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n846), .B1(new_n913), .B2(new_n937), .ZN(new_n938));
  OAI21_X1  g0738(.A(new_n938), .B1(new_n913), .B2(new_n937), .ZN(new_n939));
  INV_X1    g0739(.A(new_n531), .ZN(new_n940));
  OR2_X1    g0740(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n940), .A2(KEYINPUT35), .ZN(new_n942));
  NAND4_X1  g0742(.A1(new_n941), .A2(G116), .A3(new_n216), .A4(new_n942), .ZN(new_n943));
  XNOR2_X1  g0743(.A(new_n943), .B(KEYINPUT36), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n385), .A2(G77), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n252), .B1(new_n209), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n946), .A2(G1), .A3(new_n733), .ZN(new_n947));
  NAND3_X1  g0747(.A1(new_n939), .A2(new_n944), .A3(new_n947), .ZN(G367));
  NAND2_X1  g0748(.A1(new_n624), .A2(new_n673), .ZN(new_n949));
  AND2_X1   g0749(.A1(new_n629), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g0750(.A(new_n950), .B(KEYINPUT113), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n649), .A2(new_n673), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n953), .A2(new_n511), .A3(new_n685), .ZN(new_n954));
  OR2_X1    g0754(.A1(new_n954), .A2(KEYINPUT42), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n543), .B1(new_n951), .B2(new_n661), .ZN(new_n956));
  AOI22_X1  g0756(.A1(new_n954), .A2(KEYINPUT42), .B1(new_n680), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n567), .A2(new_n673), .ZN(new_n959));
  MUX2_X1   g0759(.A(new_n652), .B(new_n723), .S(new_n959), .Z(new_n960));
  INV_X1    g0760(.A(KEYINPUT43), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n960), .A2(new_n961), .ZN(new_n963));
  NAND3_X1  g0763(.A1(new_n958), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  NAND4_X1  g0764(.A1(new_n955), .A2(new_n957), .A3(new_n961), .A4(new_n960), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g0766(.A(new_n953), .ZN(new_n967));
  NOR2_X1   g0767(.A1(new_n684), .A2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n966), .B(new_n968), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n689), .B(KEYINPUT41), .Z(new_n970));
  NAND2_X1  g0770(.A1(new_n685), .A2(new_n511), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n682), .B2(new_n685), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n677), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n973), .B1(new_n732), .B2(new_n972), .ZN(new_n974));
  AND2_X1   g0774(.A1(new_n974), .A2(new_n730), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n953), .A2(new_n686), .ZN(new_n976));
  XNOR2_X1  g0776(.A(new_n976), .B(KEYINPUT44), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n953), .A2(new_n686), .ZN(new_n978));
  INV_X1    g0778(.A(KEYINPUT45), .ZN(new_n979));
  XNOR2_X1  g0779(.A(new_n978), .B(new_n979), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n684), .A2(new_n977), .A3(new_n980), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n977), .A2(new_n980), .ZN(new_n982));
  INV_X1    g0782(.A(KEYINPUT91), .ZN(new_n983));
  XNOR2_X1  g0783(.A(new_n683), .B(new_n983), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n982), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g0785(.A1(new_n975), .A2(new_n981), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n970), .B1(new_n986), .B2(new_n730), .ZN(new_n987));
  OAI21_X1  g0787(.A(new_n969), .B1(new_n987), .B2(new_n736), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n749), .B1(new_n222), .B2(new_n324), .ZN(new_n989));
  INV_X1    g0789(.A(new_n753), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n246), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n737), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n824), .A2(G50), .B1(G159), .B2(new_n760), .ZN(new_n993));
  OR2_X1    g0793(.A1(new_n993), .A2(KEYINPUT115), .ZN(new_n994));
  INV_X1    g0794(.A(G137), .ZN(new_n995));
  OAI22_X1  g0795(.A1(new_n763), .A2(new_n202), .B1(new_n995), .B2(new_n780), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n785), .A2(new_n837), .B1(new_n786), .B2(new_n203), .ZN(new_n997));
  INV_X1    g0797(.A(new_n772), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n996), .B(new_n997), .C1(new_n998), .C2(G150), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n292), .B1(new_n765), .B2(new_n228), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n1000), .B(KEYINPUT116), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n993), .A2(KEYINPUT115), .ZN(new_n1002));
  NAND4_X1  g0802(.A1(new_n994), .A2(new_n999), .A3(new_n1001), .A4(new_n1002), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(G303), .A2(new_n998), .B1(new_n824), .B2(G283), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n761), .A2(new_n480), .B1(new_n785), .B2(new_n789), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(G107), .B2(new_n799), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT46), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n1007), .B1(new_n763), .B2(new_n594), .ZN(new_n1008));
  OR3_X1    g0808(.A1(new_n763), .A2(new_n1007), .A3(new_n594), .ZN(new_n1009));
  NAND4_X1  g0809(.A1(new_n1004), .A2(new_n1006), .A3(new_n1008), .A4(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(G317), .ZN(new_n1011));
  OAI221_X1 g0811(.A(new_n391), .B1(new_n1011), .B2(new_n780), .C1(new_n765), .C2(new_n528), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT114), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n1003), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  XOR2_X1   g0814(.A(KEYINPUT117), .B(KEYINPUT47), .Z(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n992), .B1(new_n1016), .B2(new_n748), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n960), .A2(new_n744), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n988), .A2(new_n1019), .ZN(G387));
  NOR3_X1   g0820(.A1(new_n975), .A2(G41), .A3(new_n688), .ZN(new_n1021));
  OAI21_X1  g0821(.A(new_n1021), .B1(new_n730), .B2(new_n974), .ZN(new_n1022));
  OR2_X1    g0822(.A1(new_n682), .A2(new_n743), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n753), .B1(new_n243), .B2(new_n287), .ZN(new_n1024));
  NAND3_X1  g0824(.A1(new_n222), .A2(new_n691), .A3(new_n292), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OR3_X1    g0826(.A1(new_n268), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1027));
  OAI21_X1  g0827(.A(KEYINPUT50), .B1(new_n268), .B2(G50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(G45), .B1(G68), .B2(G77), .ZN(new_n1029));
  NAND4_X1  g0829(.A1(new_n1027), .A2(new_n690), .A3(new_n1028), .A4(new_n1029), .ZN(new_n1030));
  AOI22_X1  g0830(.A1(new_n1026), .A2(new_n1030), .B1(new_n230), .B2(new_n688), .ZN(new_n1031));
  OAI21_X1  g0831(.A(new_n737), .B1(new_n1031), .B2(new_n750), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n998), .A2(G50), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n785), .A2(new_n781), .B1(new_n763), .B2(new_n228), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1034), .B1(new_n269), .B2(new_n760), .ZN(new_n1035));
  INV_X1    g0835(.A(G150), .ZN(new_n1036));
  NOR2_X1   g0836(.A1(new_n780), .A2(new_n1036), .ZN(new_n1037));
  AOI211_X1 g0837(.A(new_n391), .B(new_n1037), .C1(G68), .C2(new_n773), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n766), .A2(G97), .B1(new_n799), .B2(new_n325), .ZN(new_n1039));
  NAND4_X1  g0839(.A1(new_n1033), .A2(new_n1035), .A3(new_n1038), .A4(new_n1039), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n752), .B1(G326), .B2(new_n791), .ZN(new_n1041));
  OAI22_X1  g0841(.A1(new_n763), .A2(new_n480), .B1(new_n786), .B2(new_n801), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G311), .A2(new_n760), .B1(new_n784), .B2(G322), .ZN(new_n1043));
  OAI221_X1 g0843(.A(new_n1043), .B1(new_n777), .B2(new_n802), .C1(new_n772), .C2(new_n1011), .ZN(new_n1044));
  INV_X1    g0844(.A(KEYINPUT48), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n1042), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(new_n1045), .B2(new_n1044), .ZN(new_n1047));
  INV_X1    g0847(.A(KEYINPUT49), .ZN(new_n1048));
  OAI221_X1 g0848(.A(new_n1041), .B1(new_n594), .B2(new_n765), .C1(new_n1047), .C2(new_n1048), .ZN(new_n1049));
  AND2_X1   g0849(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1040), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n1032), .B1(new_n1051), .B2(new_n748), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n974), .A2(new_n736), .B1(new_n1023), .B2(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1022), .A2(new_n1053), .ZN(G393));
  INV_X1    g0854(.A(KEYINPUT118), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n985), .A2(new_n981), .A3(new_n1055), .ZN(new_n1056));
  NAND3_X1  g0856(.A1(new_n982), .A2(KEYINPUT118), .A3(new_n984), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g0858(.A(new_n689), .B(new_n986), .C1(new_n1058), .C2(new_n975), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n967), .A2(new_n744), .ZN(new_n1060));
  OAI21_X1  g0860(.A(new_n749), .B1(new_n528), .B2(new_n222), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n990), .A2(new_n250), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n737), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n772), .A2(new_n789), .B1(new_n1011), .B2(new_n785), .ZN(new_n1064));
  XOR2_X1   g0864(.A(new_n1064), .B(KEYINPUT52), .Z(new_n1065));
  OAI221_X1 g0865(.A(new_n300), .B1(new_n797), .B2(new_n780), .C1(new_n788), .C2(new_n480), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n761), .A2(new_n802), .B1(new_n765), .B2(new_n230), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n763), .A2(new_n801), .B1(new_n786), .B2(new_n594), .ZN(new_n1068));
  NOR4_X1   g0868(.A1(new_n1065), .A2(new_n1066), .A3(new_n1067), .A4(new_n1068), .ZN(new_n1069));
  OAI22_X1  g0869(.A1(new_n772), .A2(new_n781), .B1(new_n1036), .B2(new_n785), .ZN(new_n1070));
  XOR2_X1   g0870(.A(new_n1070), .B(KEYINPUT51), .Z(new_n1071));
  AOI22_X1  g0871(.A1(new_n766), .A2(G87), .B1(new_n799), .B2(G77), .ZN(new_n1072));
  OAI221_X1 g0872(.A(new_n1072), .B1(new_n203), .B2(new_n763), .C1(new_n251), .C2(new_n761), .ZN(new_n1073));
  OAI221_X1 g0873(.A(new_n752), .B1(new_n837), .B2(new_n780), .C1(new_n777), .C2(new_n268), .ZN(new_n1074));
  NOR3_X1   g0874(.A1(new_n1071), .A2(new_n1073), .A3(new_n1074), .ZN(new_n1075));
  OR2_X1    g0875(.A1(new_n1069), .A2(new_n1075), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n1063), .B1(new_n1076), .B2(new_n748), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1058), .A2(new_n736), .B1(new_n1060), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1059), .A2(new_n1078), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1079), .A2(KEYINPUT119), .ZN(new_n1080));
  INV_X1    g0880(.A(KEYINPUT119), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1059), .A2(new_n1078), .A3(new_n1081), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1080), .A2(new_n1082), .ZN(G390));
  AOI21_X1  g0883(.A(new_n927), .B1(new_n726), .B2(new_n813), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n925), .B1(new_n714), .B2(new_n813), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n847), .A2(G330), .A3(new_n813), .A4(new_n925), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n1084), .A2(new_n1086), .A3(new_n1087), .ZN(new_n1088));
  INV_X1    g0888(.A(KEYINPUT120), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n714), .A2(KEYINPUT120), .A3(new_n813), .A4(new_n925), .ZN(new_n1091));
  AOI21_X1  g0891(.A(new_n1085), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n927), .B1(new_n728), .B2(new_n813), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1088), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n452), .A2(new_n714), .ZN(new_n1095));
  AND3_X1   g0895(.A1(new_n935), .A2(new_n1095), .A3(new_n643), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n922), .B1(new_n1093), .B2(new_n926), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n919), .A2(new_n920), .A3(new_n1098), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n906), .A2(new_n923), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n1100), .B1(new_n1084), .B2(new_n926), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1099), .A2(new_n1101), .A3(new_n1087), .ZN(new_n1102));
  INV_X1    g0902(.A(new_n1102), .ZN(new_n1103));
  NAND2_X1  g0903(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1104), .B1(new_n1099), .B2(new_n1101), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1097), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1099), .A2(new_n1101), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1104), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1107), .A2(new_n1108), .ZN(new_n1109));
  NAND4_X1  g0909(.A1(new_n1109), .A2(new_n1096), .A3(new_n1094), .A4(new_n1102), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n1106), .A2(new_n1110), .A3(new_n689), .ZN(new_n1111));
  NAND3_X1  g0911(.A1(new_n1109), .A2(new_n736), .A3(new_n1102), .ZN(new_n1112));
  INV_X1    g0912(.A(KEYINPUT123), .ZN(new_n1113));
  OAI21_X1  g0913(.A(new_n737), .B1(new_n269), .B2(new_n822), .ZN(new_n1114));
  INV_X1    g0914(.A(G125), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n292), .B1(new_n780), .B2(new_n1115), .C1(new_n765), .C2(new_n251), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1116), .B1(new_n998), .B2(G132), .ZN(new_n1117));
  INV_X1    g0917(.A(G128), .ZN(new_n1118));
  OAI22_X1  g0918(.A1(new_n785), .A2(new_n1118), .B1(new_n786), .B2(new_n781), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1119), .B1(G137), .B2(new_n760), .ZN(new_n1120));
  XNOR2_X1  g0920(.A(KEYINPUT54), .B(G143), .ZN(new_n1121));
  XOR2_X1   g0921(.A(new_n1121), .B(KEYINPUT121), .Z(new_n1122));
  NAND2_X1  g0922(.A1(new_n824), .A2(new_n1122), .ZN(new_n1123));
  NOR2_X1   g0923(.A1(new_n763), .A2(new_n1036), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(new_n1124), .B(KEYINPUT53), .ZN(new_n1125));
  NAND4_X1  g0925(.A1(new_n1117), .A2(new_n1120), .A3(new_n1123), .A4(new_n1125), .ZN(new_n1126));
  OAI221_X1 g0926(.A(new_n300), .B1(new_n780), .B2(new_n480), .C1(new_n763), .C2(new_n458), .ZN(new_n1127));
  OAI221_X1 g0927(.A(new_n832), .B1(new_n228), .B2(new_n786), .C1(new_n785), .C2(new_n801), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(G116), .C2(new_n998), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n824), .A2(G97), .B1(G107), .B2(new_n760), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(KEYINPUT122), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(KEYINPUT122), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g0934(.A(new_n1126), .B1(new_n1132), .B2(new_n1134), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1114), .B1(new_n1135), .B2(new_n748), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1136), .B1(new_n921), .B2(new_n741), .ZN(new_n1137));
  AND3_X1   g0937(.A1(new_n1112), .A2(new_n1113), .A3(new_n1137), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1113), .B1(new_n1112), .B2(new_n1137), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1111), .B1(new_n1138), .B2(new_n1139), .ZN(G378));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n276), .A2(new_n859), .ZN(new_n1143));
  NAND3_X1  g0943(.A1(new_n311), .A2(new_n381), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1143), .B1(new_n311), .B2(new_n381), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1142), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g0947(.A(new_n1146), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n1148), .A2(new_n1144), .A3(new_n1141), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n891), .A2(new_n893), .ZN(new_n1152));
  AND3_X1   g0952(.A1(new_n847), .A2(new_n894), .A3(new_n855), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n894), .B1(new_n847), .B2(new_n855), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n1153), .A2(new_n1154), .ZN(new_n1155));
  AOI21_X1  g0955(.A(KEYINPUT40), .B1(new_n1152), .B2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g0956(.A(G330), .B1(new_n906), .B2(new_n907), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1151), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n932), .B1(new_n921), .B2(new_n923), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1157), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n898), .A2(new_n1160), .A3(new_n1150), .ZN(new_n1161));
  AND3_X1   g0961(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1159), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1163));
  OAI21_X1  g0963(.A(KEYINPUT57), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1096), .ZN(new_n1165));
  NOR2_X1   g0965(.A1(new_n1103), .A2(new_n1105), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n1165), .B1(new_n1166), .B2(new_n1094), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n689), .B1(new_n1164), .B2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1110), .A2(new_n1096), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n1151), .B(new_n1157), .C1(new_n897), .C2(new_n896), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1150), .B1(new_n898), .B2(new_n1160), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n934), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g0972(.A1(new_n1158), .A2(new_n1159), .A3(new_n1161), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1172), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(KEYINPUT57), .B1(new_n1169), .B2(new_n1174), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1168), .A2(new_n1175), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n735), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1151), .A2(new_n740), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n737), .B1(G50), .B2(new_n822), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1122), .ZN(new_n1180));
  OAI22_X1  g0980(.A1(new_n1180), .A2(new_n763), .B1(new_n772), .B2(new_n1118), .ZN(new_n1181));
  OAI22_X1  g0981(.A1(new_n788), .A2(new_n995), .B1(new_n1036), .B2(new_n786), .ZN(new_n1182));
  INV_X1    g0982(.A(G132), .ZN(new_n1183));
  OAI22_X1  g0983(.A1(new_n761), .A2(new_n1183), .B1(new_n785), .B2(new_n1115), .ZN(new_n1184));
  NOR3_X1   g0984(.A1(new_n1181), .A2(new_n1182), .A3(new_n1184), .ZN(new_n1185));
  INV_X1    g0985(.A(new_n1185), .ZN(new_n1186));
  OR2_X1    g0986(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1186), .A2(KEYINPUT59), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n766), .A2(G159), .ZN(new_n1189));
  AOI211_X1 g0989(.A(G33), .B(G41), .C1(new_n791), .C2(G124), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1187), .A2(new_n1188), .A3(new_n1189), .A4(new_n1190), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n786), .A2(new_n203), .ZN(new_n1192));
  OAI22_X1  g0992(.A1(new_n788), .A2(new_n324), .B1(new_n801), .B2(new_n780), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1192), .B(new_n1193), .C1(new_n998), .C2(G107), .ZN(new_n1194));
  NOR2_X1   g0994(.A1(new_n765), .A2(new_n202), .ZN(new_n1195));
  OAI22_X1  g0995(.A1(new_n785), .A2(new_n594), .B1(new_n763), .B2(new_n228), .ZN(new_n1196));
  AOI211_X1 g0996(.A(new_n1195), .B(new_n1196), .C1(G97), .C2(new_n760), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1194), .A2(new_n286), .A3(new_n391), .A4(new_n1197), .ZN(new_n1198));
  INV_X1    g0998(.A(KEYINPUT58), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  OR2_X1    g1000(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1201));
  AOI21_X1  g1001(.A(G50), .B1(new_n296), .B2(new_n286), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1202), .B1(new_n752), .B2(G41), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n1191), .A2(new_n1200), .A3(new_n1201), .A4(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1179), .B1(new_n1204), .B2(new_n748), .ZN(new_n1205));
  AND2_X1   g1005(.A1(new_n1178), .A2(new_n1205), .ZN(new_n1206));
  NOR3_X1   g1006(.A1(new_n1176), .A2(new_n1177), .A3(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(G375));
  OR2_X1    g1008(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1209));
  INV_X1    g1009(.A(new_n970), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1209), .A2(new_n1210), .A3(new_n1097), .ZN(new_n1211));
  OAI22_X1  g1011(.A1(new_n788), .A2(new_n1036), .B1(new_n1118), .B2(new_n780), .ZN(new_n1212));
  AOI211_X1 g1012(.A(new_n391), .B(new_n1212), .C1(new_n998), .C2(G137), .ZN(new_n1213));
  OAI22_X1  g1013(.A1(new_n785), .A2(new_n1183), .B1(new_n763), .B2(new_n781), .ZN(new_n1214));
  AOI211_X1 g1014(.A(new_n1195), .B(new_n1214), .C1(G50), .C2(new_n799), .ZN(new_n1215));
  OAI211_X1 g1015(.A(new_n1213), .B(new_n1215), .C1(new_n761), .C2(new_n1180), .ZN(new_n1216));
  OAI22_X1  g1016(.A1(new_n777), .A2(new_n230), .B1(new_n594), .B2(new_n761), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT124), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n763), .A2(new_n528), .B1(new_n802), .B2(new_n780), .ZN(new_n1219));
  XOR2_X1   g1019(.A(new_n1219), .B(KEYINPUT126), .Z(new_n1220));
  NAND2_X1  g1020(.A1(new_n1218), .A2(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n998), .A2(G283), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n300), .B1(new_n765), .B2(new_n228), .ZN(new_n1223));
  OR2_X1    g1023(.A1(new_n1223), .A2(KEYINPUT125), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1223), .A2(KEYINPUT125), .ZN(new_n1225));
  AOI22_X1  g1025(.A1(new_n799), .A2(new_n325), .B1(G294), .B2(new_n784), .ZN(new_n1226));
  NAND4_X1  g1026(.A1(new_n1222), .A2(new_n1224), .A3(new_n1225), .A4(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1216), .B1(new_n1221), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1228), .A2(new_n748), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1229), .B(new_n737), .C1(G68), .C2(new_n822), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1230), .B1(new_n926), .B2(new_n740), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1094), .B2(new_n736), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1211), .A2(new_n1232), .ZN(G381));
  OR2_X1    g1033(.A1(G393), .A2(G396), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(G390), .A2(G384), .A3(new_n1234), .A4(G387), .ZN(new_n1235));
  INV_X1    g1035(.A(G381), .ZN(new_n1236));
  AND3_X1   g1036(.A1(new_n1111), .A2(new_n1112), .A3(new_n1137), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1235), .A2(new_n1207), .A3(new_n1236), .A4(new_n1237), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n672), .A2(G213), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1207), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(G407), .A2(G213), .A3(new_n1241), .ZN(G409));
  XNOR2_X1  g1042(.A(G393), .B(G396), .ZN(new_n1243));
  AND3_X1   g1043(.A1(new_n1080), .A2(G387), .A3(new_n1082), .ZN(new_n1244));
  AOI21_X1  g1044(.A(G387), .B1(new_n1080), .B2(new_n1082), .ZN(new_n1245));
  OAI21_X1  g1045(.A(new_n1243), .B1(new_n1244), .B2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(G387), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(G390), .A2(new_n1247), .ZN(new_n1248));
  INV_X1    g1048(.A(new_n1243), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1080), .A2(G387), .A3(new_n1082), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1248), .A2(new_n1249), .A3(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1246), .A2(new_n1251), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1206), .B1(new_n1174), .B2(new_n736), .ZN(new_n1253));
  OAI211_X1 g1053(.A(G378), .B(new_n1253), .C1(new_n1168), .C2(new_n1175), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1169), .A2(new_n1210), .A3(new_n1174), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1253), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n1237), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1240), .B1(new_n1254), .B2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1097), .A2(KEYINPUT60), .ZN(new_n1259));
  AND2_X1   g1059(.A1(new_n1259), .A2(new_n1209), .ZN(new_n1260));
  OAI21_X1  g1060(.A(new_n689), .B1(new_n1259), .B2(new_n1209), .ZN(new_n1261));
  OAI21_X1  g1061(.A(new_n1232), .B1(new_n1260), .B2(new_n1261), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1262), .A2(new_n844), .ZN(new_n1263));
  OAI211_X1 g1063(.A(G384), .B(new_n1232), .C1(new_n1260), .C2(new_n1261), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(new_n1264), .ZN(new_n1265));
  INV_X1    g1065(.A(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(KEYINPUT62), .B1(new_n1258), .B2(new_n1266), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n1254), .A2(new_n1257), .ZN(new_n1268));
  AOI21_X1  g1068(.A(KEYINPUT127), .B1(new_n1268), .B2(new_n1239), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT127), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1270), .B(new_n1240), .C1(new_n1254), .C2(new_n1257), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1269), .A2(new_n1271), .ZN(new_n1272));
  AND2_X1   g1072(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1267), .B1(new_n1272), .B2(new_n1273), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1240), .A2(G2897), .ZN(new_n1275));
  XNOR2_X1  g1075(.A(new_n1265), .B(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1276), .B1(new_n1269), .B2(new_n1271), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT61), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1277), .A2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1252), .B1(new_n1274), .B2(new_n1279), .ZN(new_n1280));
  NAND3_X1  g1080(.A1(new_n1272), .A2(KEYINPUT63), .A3(new_n1266), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1252), .A2(KEYINPUT61), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT63), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1258), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1283), .B1(new_n1284), .B2(new_n1265), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1276), .A2(new_n1284), .ZN(new_n1286));
  NAND4_X1  g1086(.A1(new_n1281), .A2(new_n1282), .A3(new_n1285), .A4(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1280), .A2(new_n1287), .ZN(G405));
  INV_X1    g1088(.A(new_n1237), .ZN(new_n1289));
  OAI21_X1  g1089(.A(new_n1254), .B1(new_n1207), .B2(new_n1289), .ZN(new_n1290));
  XNOR2_X1  g1090(.A(new_n1290), .B(new_n1266), .ZN(new_n1291));
  XNOR2_X1  g1091(.A(new_n1291), .B(new_n1252), .ZN(G402));
endmodule


