//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 1 0 0 0 0 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:18 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n532,
    new_n533, new_n534, new_n535, new_n536, new_n537, new_n538, new_n539,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n556,
    new_n558, new_n559, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n613, new_n614, new_n615, new_n618,
    new_n620, new_n621, new_n623, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1183, new_n1184;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XOR2_X1   g003(.A(KEYINPUT64), .B(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT65), .B(G44), .ZN(G218));
  XOR2_X1   g009(.A(KEYINPUT66), .B(G132), .Z(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n450));
  XNOR2_X1  g025(.A(KEYINPUT67), .B(KEYINPUT2), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n453), .A2(G567), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  OAI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(KEYINPUT68), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(KEYINPUT68), .B2(new_n457), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI211_X1 g037(.A(G137), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NAND3_X1  g038(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT70), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT70), .ZN(new_n467));
  NAND3_X1  g042(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  OAI21_X1  g044(.A(KEYINPUT69), .B1(new_n461), .B2(new_n462), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  INV_X1    g046(.A(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  INV_X1    g048(.A(KEYINPUT69), .ZN(new_n474));
  NAND2_X1  g049(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n475));
  NAND3_X1  g050(.A1(new_n473), .A2(new_n474), .A3(new_n475), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n470), .A2(new_n476), .A3(G125), .ZN(new_n477));
  NAND2_X1  g052(.A1(G113), .A2(G2104), .ZN(new_n478));
  AOI21_X1  g053(.A(new_n460), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n469), .A2(new_n479), .ZN(G160));
  AOI21_X1  g055(.A(G2105), .B1(new_n473), .B2(new_n475), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT71), .Z(new_n483));
  OR2_X1    g058(.A1(G100), .A2(G2105), .ZN(new_n484));
  OAI211_X1 g059(.A(new_n484), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n485));
  AND2_X1   g060(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  AOI21_X1  g061(.A(new_n460), .B1(new_n473), .B2(new_n475), .ZN(new_n487));
  XNOR2_X1  g062(.A(new_n487), .B(KEYINPUT72), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G124), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n486), .A2(new_n490), .ZN(new_n491));
  INV_X1    g066(.A(new_n491), .ZN(G162));
  OAI211_X1 g067(.A(G126), .B(G2105), .C1(new_n461), .C2(new_n462), .ZN(new_n493));
  OR2_X1    g068(.A1(G102), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G2105), .ZN(new_n496));
  NAND3_X1  g071(.A1(new_n494), .A2(new_n496), .A3(G2104), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n493), .A2(new_n497), .ZN(new_n498));
  INV_X1    g073(.A(G138), .ZN(new_n499));
  NOR3_X1   g074(.A1(new_n499), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n470), .A2(new_n476), .A3(new_n500), .ZN(new_n501));
  OAI211_X1 g076(.A(G138), .B(new_n460), .C1(new_n461), .C2(new_n462), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(KEYINPUT4), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n498), .B1(new_n501), .B2(new_n503), .ZN(G164));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  INV_X1    g080(.A(KEYINPUT73), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  OAI21_X1  g082(.A(new_n506), .B1(new_n507), .B2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND3_X1  g084(.A1(new_n509), .A2(KEYINPUT73), .A3(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n511), .A2(G62), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G75), .A2(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n505), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT6), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(new_n505), .ZN(new_n517));
  NAND2_X1  g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n511), .A2(G88), .A3(new_n512), .ZN(new_n521));
  NAND2_X1  g096(.A1(G50), .A2(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n515), .A2(new_n523), .ZN(G166));
  NAND2_X1  g099(.A1(new_n511), .A2(new_n512), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n520), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n526), .A2(G89), .ZN(new_n527));
  INV_X1    g102(.A(new_n518), .ZN(new_n528));
  NOR2_X1   g103(.A1(KEYINPUT6), .A2(G651), .ZN(new_n529));
  OAI21_X1  g104(.A(KEYINPUT74), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  INV_X1    g105(.A(KEYINPUT74), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(new_n531), .A3(new_n518), .ZN(new_n532));
  NAND3_X1  g107(.A1(new_n530), .A2(G543), .A3(new_n532), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G51), .ZN(new_n535));
  NAND3_X1  g110(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n536));
  XNOR2_X1  g111(.A(new_n536), .B(KEYINPUT7), .ZN(new_n537));
  AND2_X1   g112(.A1(new_n511), .A2(new_n512), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n538), .A2(G63), .A3(G651), .ZN(new_n539));
  AND4_X1   g114(.A1(new_n527), .A2(new_n535), .A3(new_n537), .A4(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n538), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n541));
  NOR2_X1   g116(.A1(new_n541), .A2(new_n505), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n538), .A2(new_n519), .ZN(new_n543));
  INV_X1    g118(.A(G90), .ZN(new_n544));
  INV_X1    g119(.A(G52), .ZN(new_n545));
  OAI22_X1  g120(.A1(new_n543), .A2(new_n544), .B1(new_n545), .B2(new_n533), .ZN(new_n546));
  NOR2_X1   g121(.A1(new_n542), .A2(new_n546), .ZN(G171));
  AOI22_X1  g122(.A1(G81), .A2(new_n526), .B1(new_n534), .B2(G43), .ZN(new_n548));
  NAND2_X1  g123(.A1(G68), .A2(G543), .ZN(new_n549));
  INV_X1    g124(.A(G56), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n549), .B1(new_n525), .B2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G651), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n548), .A2(new_n552), .ZN(new_n553));
  INV_X1    g128(.A(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G860), .ZN(G153));
  AND3_X1   g130(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n556), .A2(G36), .ZN(G176));
  NAND2_X1  g132(.A1(G1), .A2(G3), .ZN(new_n558));
  XNOR2_X1  g133(.A(new_n558), .B(KEYINPUT8), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n556), .A2(new_n559), .ZN(G188));
  NAND4_X1  g135(.A1(new_n530), .A2(new_n532), .A3(G53), .A4(G543), .ZN(new_n561));
  XOR2_X1   g136(.A(KEYINPUT76), .B(KEYINPUT9), .Z(new_n562));
  OAI21_X1  g137(.A(KEYINPUT77), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT77), .ZN(new_n564));
  INV_X1    g139(.A(new_n562), .ZN(new_n565));
  NAND4_X1  g140(.A1(new_n534), .A2(new_n564), .A3(G53), .A4(new_n565), .ZN(new_n566));
  NAND3_X1  g141(.A1(new_n561), .A2(KEYINPUT75), .A3(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(new_n568));
  AOI21_X1  g143(.A(KEYINPUT75), .B1(new_n561), .B2(KEYINPUT9), .ZN(new_n569));
  OAI211_X1 g144(.A(new_n563), .B(new_n566), .C1(new_n568), .C2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(G78), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G65), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n525), .B2(new_n572), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n573), .A2(G651), .B1(new_n526), .B2(G91), .ZN(new_n574));
  NAND2_X1  g149(.A1(new_n570), .A2(new_n574), .ZN(G299));
  INV_X1    g150(.A(G171), .ZN(G301));
  INV_X1    g151(.A(G168), .ZN(G286));
  INV_X1    g152(.A(G166), .ZN(G303));
  NAND4_X1  g153(.A1(new_n530), .A2(new_n532), .A3(G49), .A4(G543), .ZN(new_n579));
  NAND4_X1  g154(.A1(new_n511), .A2(G87), .A3(new_n512), .A4(new_n519), .ZN(new_n580));
  AOI21_X1  g155(.A(G74), .B1(new_n511), .B2(new_n512), .ZN(new_n581));
  OAI211_X1 g156(.A(new_n579), .B(new_n580), .C1(new_n581), .C2(new_n505), .ZN(G288));
  NAND3_X1  g157(.A1(new_n511), .A2(G61), .A3(new_n512), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(KEYINPUT78), .B1(G73), .B2(G543), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT78), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n538), .A2(new_n585), .A3(G61), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n505), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n538), .A2(G86), .ZN(new_n588));
  NAND2_X1  g163(.A1(G48), .A2(G543), .ZN(new_n589));
  AOI21_X1  g164(.A(new_n520), .B1(new_n588), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n538), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n505), .ZN(new_n594));
  AOI22_X1  g169(.A1(G85), .A2(new_n526), .B1(new_n534), .B2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n594), .A2(new_n595), .ZN(G290));
  NAND2_X1  g171(.A1(G301), .A2(G868), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n511), .A2(G66), .A3(new_n512), .ZN(new_n598));
  NAND2_X1  g173(.A1(G79), .A2(G543), .ZN(new_n599));
  AOI21_X1  g174(.A(new_n505), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G54), .ZN(new_n601));
  NOR2_X1   g176(.A1(new_n533), .A2(new_n601), .ZN(new_n602));
  OR3_X1    g177(.A1(new_n600), .A2(new_n602), .A3(KEYINPUT79), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT79), .B1(new_n600), .B2(new_n602), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n526), .A2(G92), .ZN(new_n606));
  INV_X1    g181(.A(KEYINPUT10), .ZN(new_n607));
  XNOR2_X1  g182(.A(new_n606), .B(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n597), .B1(new_n610), .B2(G868), .ZN(G284));
  OAI21_X1  g186(.A(new_n597), .B1(new_n610), .B2(G868), .ZN(G321));
  INV_X1    g187(.A(G868), .ZN(new_n613));
  NOR2_X1   g188(.A1(G286), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g189(.A(G299), .B(KEYINPUT80), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G297));
  AOI21_X1  g191(.A(new_n614), .B1(new_n615), .B2(new_n613), .ZN(G280));
  XNOR2_X1  g192(.A(KEYINPUT81), .B(G559), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n610), .B1(G860), .B2(new_n618), .ZN(G148));
  NAND2_X1  g194(.A1(new_n610), .A2(new_n618), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(G868), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(G868), .B2(new_n554), .ZN(G323));
  XNOR2_X1  g197(.A(KEYINPUT82), .B(KEYINPUT11), .ZN(new_n623));
  XNOR2_X1  g198(.A(G323), .B(new_n623), .ZN(G282));
  NAND2_X1  g199(.A1(new_n470), .A2(new_n476), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n460), .A2(G2104), .ZN(new_n626));
  NOR2_X1   g201(.A1(new_n625), .A2(new_n626), .ZN(new_n627));
  XOR2_X1   g202(.A(new_n627), .B(KEYINPUT12), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT83), .B(KEYINPUT13), .Z(new_n630));
  OR2_X1    g205(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n629), .A2(new_n630), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n481), .A2(G135), .ZN(new_n633));
  NOR2_X1   g208(.A1(new_n460), .A2(G111), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n635));
  INV_X1    g210(.A(G123), .ZN(new_n636));
  OAI221_X1 g211(.A(new_n633), .B1(new_n634), .B2(new_n635), .C1(new_n488), .C2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND3_X1  g213(.A1(new_n631), .A2(new_n632), .A3(new_n638), .ZN(G156));
  INV_X1    g214(.A(KEYINPUT14), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2427), .B(G2438), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2430), .ZN(new_n642));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  AOI21_X1  g218(.A(new_n640), .B1(new_n642), .B2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(new_n644), .B1(new_n643), .B2(new_n642), .ZN(new_n645));
  XNOR2_X1  g220(.A(G2451), .B(G2454), .ZN(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT16), .ZN(new_n647));
  XNOR2_X1  g222(.A(G1341), .B(G1348), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n645), .B(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2443), .B(G2446), .ZN(new_n651));
  NAND2_X1  g226(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n652), .A2(G14), .ZN(new_n653));
  NOR2_X1   g228(.A1(new_n650), .A2(new_n651), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n653), .A2(new_n654), .ZN(G401));
  XNOR2_X1  g230(.A(G2067), .B(G2678), .ZN(new_n656));
  XOR2_X1   g231(.A(G2072), .B(G2078), .Z(new_n657));
  XOR2_X1   g232(.A(new_n657), .B(KEYINPUT84), .Z(new_n658));
  AOI21_X1  g233(.A(new_n656), .B1(new_n658), .B2(KEYINPUT85), .ZN(new_n659));
  OAI21_X1  g234(.A(new_n659), .B1(KEYINPUT85), .B2(new_n658), .ZN(new_n660));
  XNOR2_X1  g235(.A(G2084), .B(G2090), .ZN(new_n661));
  XOR2_X1   g236(.A(new_n658), .B(KEYINPUT17), .Z(new_n662));
  INV_X1    g237(.A(new_n656), .ZN(new_n663));
  OAI211_X1 g238(.A(new_n660), .B(new_n661), .C1(new_n662), .C2(new_n663), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n661), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n658), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  NOR2_X1   g242(.A1(new_n656), .A2(new_n661), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n662), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n664), .A2(new_n667), .A3(new_n669), .ZN(new_n670));
  XOR2_X1   g245(.A(G2096), .B(G2100), .Z(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G227));
  XOR2_X1   g247(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n673));
  XNOR2_X1  g248(.A(G1971), .B(G1976), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n675), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT20), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n676), .A2(new_n677), .ZN(new_n681));
  NAND2_X1  g256(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n681), .A2(new_n678), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n682), .C1(new_n675), .C2(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n686), .B(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(G1981), .B(G1986), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n688), .B(new_n689), .ZN(G229));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G35), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G162), .B2(new_n691), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n693), .B(KEYINPUT29), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n694), .A2(G2090), .ZN(new_n695));
  NOR2_X1   g270(.A1(G29), .A2(G33), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n697));
  XOR2_X1   g272(.A(new_n697), .B(KEYINPUT25), .Z(new_n698));
  NAND2_X1  g273(.A1(new_n481), .A2(G139), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND2_X1  g275(.A1(G115), .A2(G2104), .ZN(new_n701));
  INV_X1    g276(.A(G127), .ZN(new_n702));
  OAI21_X1  g277(.A(new_n701), .B1(new_n625), .B2(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n700), .B1(new_n703), .B2(G2105), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n696), .B1(new_n704), .B2(G29), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G2072), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT91), .Z(new_n707));
  NAND2_X1  g282(.A1(new_n695), .A2(new_n707), .ZN(new_n708));
  INV_X1    g283(.A(G16), .ZN(new_n709));
  NOR2_X1   g284(.A1(G171), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(G5), .B2(new_n709), .ZN(new_n711));
  INV_X1    g286(.A(G1961), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  XOR2_X1   g288(.A(new_n713), .B(KEYINPUT97), .Z(new_n714));
  NOR2_X1   g289(.A1(new_n694), .A2(G2090), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n708), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n709), .A2(G21), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G168), .B2(new_n709), .ZN(new_n718));
  INV_X1    g293(.A(G1966), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(new_n705), .A2(G2072), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT90), .ZN(new_n722));
  XNOR2_X1  g297(.A(KEYINPUT31), .B(G11), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT30), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n691), .B1(new_n724), .B2(G28), .ZN(new_n725));
  AND2_X1   g300(.A1(new_n725), .A2(KEYINPUT96), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n724), .A2(G28), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n725), .B2(KEYINPUT96), .ZN(new_n728));
  OAI221_X1 g303(.A(new_n723), .B1(new_n726), .B2(new_n728), .C1(new_n637), .C2(new_n691), .ZN(new_n729));
  INV_X1    g304(.A(G2078), .ZN(new_n730));
  NOR2_X1   g305(.A1(G27), .A2(G29), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n731), .B1(G164), .B2(G29), .ZN(new_n732));
  INV_X1    g307(.A(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n729), .B1(new_n730), .B2(new_n733), .ZN(new_n734));
  AND2_X1   g309(.A1(new_n691), .A2(G32), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n489), .A2(G129), .ZN(new_n736));
  XNOR2_X1  g311(.A(new_n736), .B(KEYINPUT92), .ZN(new_n737));
  NAND3_X1  g312(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT94), .Z(new_n739));
  XOR2_X1   g314(.A(KEYINPUT93), .B(KEYINPUT26), .Z(new_n740));
  INV_X1    g315(.A(new_n740), .ZN(new_n741));
  AND2_X1   g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  NOR2_X1   g317(.A1(new_n739), .A2(new_n741), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n481), .A2(G141), .ZN(new_n744));
  INV_X1    g319(.A(G105), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n744), .B1(new_n745), .B2(new_n626), .ZN(new_n746));
  NOR3_X1   g321(.A1(new_n742), .A2(new_n743), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n737), .A2(new_n747), .ZN(new_n748));
  AOI21_X1  g323(.A(new_n735), .B1(new_n748), .B2(G29), .ZN(new_n749));
  XNOR2_X1  g324(.A(KEYINPUT27), .B(G1996), .ZN(new_n750));
  OAI221_X1 g325(.A(new_n734), .B1(new_n730), .B2(new_n733), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NAND2_X1  g326(.A1(new_n711), .A2(new_n712), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n691), .A2(G26), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT28), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n489), .A2(G128), .ZN(new_n755));
  OAI21_X1  g330(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n756));
  INV_X1    g331(.A(G116), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n756), .B1(new_n757), .B2(G2105), .ZN(new_n758));
  AOI21_X1  g333(.A(new_n758), .B1(new_n481), .B2(G140), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n755), .A2(new_n759), .ZN(new_n760));
  AOI21_X1  g335(.A(new_n754), .B1(new_n760), .B2(G29), .ZN(new_n761));
  XNOR2_X1  g336(.A(new_n761), .B(G2067), .ZN(new_n762));
  AND2_X1   g337(.A1(KEYINPUT24), .A2(G34), .ZN(new_n763));
  OAI21_X1  g338(.A(new_n691), .B1(KEYINPUT24), .B2(G34), .ZN(new_n764));
  OAI22_X1  g339(.A1(G160), .A2(new_n691), .B1(new_n763), .B2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n765), .A2(G2084), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(G2084), .ZN(new_n767));
  NAND4_X1  g342(.A1(new_n752), .A2(new_n762), .A3(new_n766), .A4(new_n767), .ZN(new_n768));
  NOR2_X1   g343(.A1(new_n751), .A2(new_n768), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n716), .A2(new_n720), .A3(new_n722), .A4(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n691), .A2(G25), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n481), .A2(G131), .ZN(new_n772));
  NOR2_X1   g347(.A1(new_n460), .A2(G107), .ZN(new_n773));
  OAI21_X1  g348(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n774));
  INV_X1    g349(.A(G119), .ZN(new_n775));
  OAI221_X1 g350(.A(new_n772), .B1(new_n773), .B2(new_n774), .C1(new_n488), .C2(new_n775), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n771), .B1(new_n776), .B2(G29), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT35), .B(G1991), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(KEYINPUT87), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n777), .B(new_n779), .ZN(new_n780));
  INV_X1    g355(.A(G290), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n781), .A2(G16), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n782), .B1(G16), .B2(G24), .ZN(new_n783));
  INV_X1    g358(.A(G1986), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n780), .B1(new_n783), .B2(new_n784), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(new_n784), .B2(new_n783), .ZN(new_n786));
  NAND2_X1  g361(.A1(new_n709), .A2(G6), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n787), .B1(new_n591), .B2(new_n709), .ZN(new_n788));
  XNOR2_X1  g363(.A(KEYINPUT32), .B(G1981), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(KEYINPUT88), .ZN(new_n790));
  OR2_X1    g365(.A1(new_n788), .A2(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n788), .A2(new_n790), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n709), .A2(G22), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G166), .B2(new_n709), .ZN(new_n794));
  INV_X1    g369(.A(G1971), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  MUX2_X1   g371(.A(G23), .B(G288), .S(G16), .Z(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT33), .B(G1976), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n797), .B(new_n798), .ZN(new_n799));
  NAND4_X1  g374(.A1(new_n791), .A2(new_n792), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  OR2_X1    g375(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n800), .A2(KEYINPUT34), .ZN(new_n802));
  NAND3_X1  g377(.A1(new_n786), .A2(new_n801), .A3(new_n802), .ZN(new_n803));
  XOR2_X1   g378(.A(new_n803), .B(KEYINPUT36), .Z(new_n804));
  NAND2_X1  g379(.A1(new_n749), .A2(new_n750), .ZN(new_n805));
  XOR2_X1   g380(.A(new_n805), .B(KEYINPUT95), .Z(new_n806));
  NOR2_X1   g381(.A1(new_n610), .A2(new_n709), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(G4), .B2(new_n709), .ZN(new_n808));
  INV_X1    g383(.A(G1348), .ZN(new_n809));
  OR2_X1    g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n808), .A2(new_n809), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n709), .A2(G19), .ZN(new_n812));
  OAI21_X1  g387(.A(new_n812), .B1(new_n554), .B2(new_n709), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT89), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(G1341), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n806), .A2(new_n810), .A3(new_n811), .A4(new_n815), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n709), .A2(G20), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT23), .Z(new_n818));
  AOI21_X1  g393(.A(new_n818), .B1(G299), .B2(G16), .ZN(new_n819));
  INV_X1    g394(.A(G1956), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  NOR4_X1   g396(.A1(new_n770), .A2(new_n804), .A3(new_n816), .A4(new_n821), .ZN(G311));
  INV_X1    g397(.A(G311), .ZN(G150));
  NAND2_X1  g398(.A1(new_n610), .A2(G559), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT38), .ZN(new_n825));
  AOI22_X1  g400(.A1(new_n538), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n826), .A2(new_n505), .ZN(new_n827));
  INV_X1    g402(.A(G93), .ZN(new_n828));
  INV_X1    g403(.A(G55), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n543), .A2(new_n828), .B1(new_n829), .B2(new_n533), .ZN(new_n830));
  OR2_X1    g405(.A1(new_n827), .A2(new_n830), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n831), .A2(new_n553), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n827), .A2(new_n830), .ZN(new_n833));
  NOR2_X1   g408(.A1(new_n554), .A2(new_n833), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n825), .B(new_n835), .ZN(new_n836));
  OR2_X1    g411(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n837));
  INV_X1    g412(.A(G860), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n836), .A2(KEYINPUT39), .ZN(new_n839));
  NAND3_X1  g414(.A1(new_n837), .A2(new_n838), .A3(new_n839), .ZN(new_n840));
  NOR2_X1   g415(.A1(new_n833), .A2(new_n838), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n841), .B(KEYINPUT37), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n840), .A2(new_n842), .ZN(G145));
  INV_X1    g418(.A(KEYINPUT98), .ZN(new_n844));
  OR2_X1    g419(.A1(new_n704), .A2(new_n844), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n748), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n501), .A2(new_n503), .ZN(new_n847));
  INV_X1    g422(.A(new_n498), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n760), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  OAI21_X1  g428(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n854));
  INV_X1    g429(.A(G118), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n854), .B1(new_n855), .B2(G2105), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n856), .B1(new_n481), .B2(G142), .ZN(new_n857));
  INV_X1    g432(.A(G130), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n857), .B1(new_n488), .B2(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(KEYINPUT100), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n859), .B(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(new_n776), .ZN(new_n862));
  XOR2_X1   g437(.A(new_n628), .B(KEYINPUT99), .Z(new_n863));
  INV_X1    g438(.A(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n862), .B(new_n864), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT101), .ZN(new_n866));
  NAND2_X1  g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n862), .B(new_n863), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT101), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n853), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  NAND4_X1  g445(.A1(new_n851), .A2(new_n865), .A3(new_n866), .A4(new_n852), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n491), .B(G160), .ZN(new_n873));
  XOR2_X1   g448(.A(new_n873), .B(new_n637), .Z(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(G37), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n870), .A2(new_n871), .A3(new_n874), .ZN(new_n878));
  NAND3_X1  g453(.A1(new_n876), .A2(new_n877), .A3(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g455(.A(G288), .B(KEYINPUT103), .ZN(new_n881));
  XOR2_X1   g456(.A(new_n881), .B(new_n591), .Z(new_n882));
  XNOR2_X1  g457(.A(G290), .B(G166), .ZN(new_n883));
  XOR2_X1   g458(.A(new_n882), .B(new_n883), .Z(new_n884));
  XOR2_X1   g459(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n885));
  XOR2_X1   g460(.A(new_n884), .B(new_n885), .Z(new_n886));
  OR2_X1    g461(.A1(G299), .A2(KEYINPUT102), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(new_n610), .ZN(new_n888));
  NAND2_X1  g463(.A1(G299), .A2(KEYINPUT102), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g466(.A1(new_n887), .A2(new_n610), .A3(new_n889), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g468(.A(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n620), .B(new_n835), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n893), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n891), .A2(KEYINPUT41), .A3(new_n892), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n901), .A2(new_n895), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n886), .A2(new_n897), .A3(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n886), .B1(new_n902), .B2(new_n897), .ZN(new_n904));
  OAI21_X1  g479(.A(G868), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(G868), .B2(new_n833), .ZN(G295));
  OAI21_X1  g481(.A(new_n905), .B1(G868), .B2(new_n833), .ZN(G331));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n908));
  OAI21_X1  g483(.A(G171), .B1(new_n832), .B2(new_n834), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n831), .A2(new_n553), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n554), .A2(new_n833), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(G301), .A3(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n909), .A2(G168), .A3(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(G168), .B1(new_n909), .B2(new_n912), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n899), .A2(new_n915), .A3(new_n900), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n894), .B1(new_n913), .B2(new_n914), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  AOI21_X1  g493(.A(G37), .B1(new_n918), .B2(new_n884), .ZN(new_n919));
  XNOR2_X1  g494(.A(KEYINPUT105), .B(KEYINPUT43), .ZN(new_n920));
  INV_X1    g495(.A(new_n884), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n916), .A2(new_n917), .A3(new_n921), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n920), .B1(new_n919), .B2(new_n922), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n908), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n919), .A2(new_n922), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT43), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n928), .A2(KEYINPUT44), .A3(new_n923), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n926), .A2(new_n929), .ZN(G397));
  XNOR2_X1  g505(.A(KEYINPUT106), .B(G1384), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n849), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n934));
  NOR2_X1   g509(.A1(G164), .A2(new_n931), .ZN(new_n935));
  INV_X1    g510(.A(KEYINPUT107), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n935), .A2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n938));
  INV_X1    g513(.A(G40), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n469), .A2(new_n479), .A3(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n934), .A2(new_n937), .A3(new_n938), .A4(new_n940), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT109), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n942), .A2(G1996), .A3(new_n748), .ZN(new_n943));
  XOR2_X1   g518(.A(new_n943), .B(KEYINPUT110), .Z(new_n944));
  NOR2_X1   g519(.A1(new_n941), .A2(G1996), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n737), .A3(new_n747), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n760), .A2(G2067), .ZN(new_n947));
  INV_X1    g522(.A(G2067), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n755), .A2(new_n948), .A3(new_n759), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n947), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n942), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g526(.A(new_n946), .B1(new_n951), .B2(KEYINPUT111), .ZN(new_n952));
  AOI21_X1  g527(.A(new_n952), .B1(KEYINPUT111), .B2(new_n951), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n776), .A2(new_n779), .ZN(new_n954));
  NOR2_X1   g529(.A1(new_n776), .A2(new_n779), .ZN(new_n955));
  OAI21_X1  g530(.A(new_n942), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(new_n941), .ZN(new_n957));
  NOR2_X1   g532(.A1(G290), .A2(G1986), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  XNOR2_X1  g534(.A(new_n959), .B(KEYINPUT48), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n944), .A2(new_n953), .A3(new_n956), .A4(new_n960), .ZN(new_n961));
  XNOR2_X1  g536(.A(new_n945), .B(KEYINPUT46), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n942), .B1(new_n748), .B2(new_n950), .ZN(new_n963));
  OR2_X1    g538(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(KEYINPUT127), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n962), .B1(new_n964), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT47), .ZN(new_n967));
  AND2_X1   g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n966), .A2(new_n967), .ZN(new_n969));
  OAI21_X1  g544(.A(new_n961), .B1(new_n968), .B2(new_n969), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n944), .A2(new_n953), .A3(new_n955), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n949), .ZN(new_n972));
  AOI21_X1  g547(.A(new_n970), .B1(new_n942), .B2(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(KEYINPUT126), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n781), .A2(new_n784), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n957), .B1(new_n975), .B2(new_n958), .ZN(new_n976));
  XOR2_X1   g551(.A(new_n976), .B(KEYINPUT108), .Z(new_n977));
  NAND4_X1  g552(.A1(new_n944), .A2(new_n953), .A3(new_n956), .A4(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(G651), .B1(new_n538), .B2(G74), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n979), .A2(G1976), .A3(new_n580), .A4(new_n579), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n477), .A2(new_n478), .ZN(new_n981));
  NAND2_X1  g556(.A1(new_n981), .A2(G2105), .ZN(new_n982));
  AND3_X1   g557(.A1(new_n463), .A2(new_n467), .A3(new_n464), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n467), .B1(new_n463), .B2(new_n464), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n982), .A2(new_n985), .A3(G40), .ZN(new_n986));
  INV_X1    g561(.A(G1384), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n849), .A2(new_n987), .ZN(new_n988));
  OAI211_X1 g563(.A(G8), .B(new_n980), .C1(new_n986), .C2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(KEYINPUT52), .ZN(new_n990));
  AOI21_X1  g565(.A(G1384), .B1(new_n847), .B2(new_n848), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n940), .A2(new_n991), .ZN(new_n992));
  XNOR2_X1  g567(.A(KEYINPUT115), .B(G1976), .ZN(new_n993));
  AOI21_X1  g568(.A(KEYINPUT52), .B1(G288), .B2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n992), .A2(G8), .A3(new_n980), .A4(new_n994), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n990), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n992), .A2(G8), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n588), .A2(new_n589), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n998), .A2(new_n519), .ZN(new_n999));
  INV_X1    g574(.A(G1981), .ZN(new_n1000));
  AND2_X1   g575(.A1(new_n584), .A2(new_n586), .ZN(new_n1001));
  OAI211_X1 g576(.A(new_n999), .B(new_n1000), .C1(new_n1001), .C2(new_n505), .ZN(new_n1002));
  OAI21_X1  g577(.A(G1981), .B1(new_n587), .B2(new_n590), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT49), .ZN(new_n1005));
  AOI21_X1  g580(.A(new_n997), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1002), .A2(KEYINPUT49), .A3(new_n1003), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n996), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT55), .B(G8), .C1(new_n515), .C2(new_n523), .ZN(new_n1009));
  XNOR2_X1  g584(.A(KEYINPUT113), .B(KEYINPUT114), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  INV_X1    g587(.A(KEYINPUT55), .ZN(new_n1013));
  INV_X1    g588(.A(G8), .ZN(new_n1014));
  OAI21_X1  g589(.A(new_n1013), .B1(G166), .B2(new_n1014), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n1011), .A2(new_n1012), .A3(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1018));
  INV_X1    g593(.A(KEYINPUT50), .ZN(new_n1019));
  NAND3_X1  g594(.A1(new_n849), .A2(new_n1019), .A3(new_n987), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n940), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(G2090), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n938), .B1(G164), .B2(G1384), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n932), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n940), .A2(new_n1023), .A3(new_n1024), .ZN(new_n1025));
  AOI22_X1  g600(.A1(new_n1021), .A2(new_n1022), .B1(new_n1025), .B2(new_n795), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1017), .B1(new_n1026), .B2(new_n1014), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n795), .ZN(new_n1028));
  OAI21_X1  g603(.A(KEYINPUT112), .B1(new_n991), .B2(new_n1019), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT112), .ZN(new_n1030));
  OAI211_X1 g605(.A(new_n1030), .B(KEYINPUT50), .C1(G164), .C2(G1384), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1029), .A2(new_n940), .A3(new_n1020), .A4(new_n1031), .ZN(new_n1032));
  OAI21_X1  g607(.A(new_n1028), .B1(new_n1032), .B2(G2090), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1033), .A2(G8), .A3(new_n1016), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G168), .A2(G8), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n986), .B1(new_n1019), .B2(new_n991), .ZN(new_n1036));
  INV_X1    g611(.A(G2084), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1036), .A2(new_n1037), .A3(new_n1029), .A4(new_n1031), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n849), .A2(KEYINPUT45), .A3(new_n987), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n940), .A2(new_n1023), .A3(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1040), .A2(new_n719), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1035), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n1008), .A2(new_n1027), .A3(new_n1034), .A4(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT63), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1043), .A2(new_n1044), .ZN(new_n1045));
  AND2_X1   g620(.A1(new_n1042), .A2(KEYINPUT63), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1033), .A2(G8), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(new_n1017), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1046), .A2(new_n1048), .A3(new_n1034), .A4(new_n1008), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1045), .A2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1051));
  INV_X1    g626(.A(new_n997), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1051), .A2(new_n1007), .A3(new_n1052), .ZN(new_n1053));
  NOR2_X1   g628(.A1(G288), .A2(G1976), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(new_n1002), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1034), .ZN(new_n1057));
  AOI22_X1  g632(.A1(new_n1056), .A2(new_n1052), .B1(new_n1057), .B2(new_n1008), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1050), .A2(new_n1058), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n940), .A2(new_n1031), .A3(new_n1020), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1030), .B1(new_n988), .B2(KEYINPUT50), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n712), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  NAND4_X1  g637(.A1(new_n940), .A2(new_n1024), .A3(new_n730), .A4(new_n1023), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT53), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(G2078), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n940), .A2(new_n1039), .A3(new_n1023), .A4(new_n1066), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1062), .A2(new_n1065), .A3(G301), .A4(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT125), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1032), .A2(new_n712), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1070));
  INV_X1    g645(.A(KEYINPUT125), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1070), .A2(new_n1071), .A3(G301), .A4(new_n1067), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1069), .A2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n1074));
  OAI21_X1  g649(.A(KEYINPUT123), .B1(new_n983), .B2(new_n984), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT123), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n466), .A2(new_n1076), .A3(new_n468), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1075), .A2(new_n1077), .A3(new_n982), .A4(G40), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT124), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  NOR2_X1   g655(.A1(new_n479), .A2(new_n939), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(new_n1075), .A3(new_n1077), .A4(KEYINPUT124), .ZN(new_n1082));
  AND2_X1   g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1066), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1084), .B1(new_n935), .B2(KEYINPUT45), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n938), .B1(new_n935), .B2(new_n936), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n933), .A2(KEYINPUT107), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1085), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n1062), .B(new_n1065), .C1(new_n1083), .C2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1074), .B1(new_n1089), .B2(G171), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1073), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n996), .ZN(new_n1092));
  AND4_X1   g667(.A1(new_n1027), .A2(new_n1034), .A3(new_n1053), .A4(new_n1092), .ZN(new_n1093));
  XOR2_X1   g668(.A(KEYINPUT122), .B(KEYINPUT54), .Z(new_n1094));
  NAND2_X1  g669(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n934), .A2(new_n937), .A3(new_n938), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1095), .A2(new_n1096), .A3(new_n1085), .ZN(new_n1097));
  AND3_X1   g672(.A1(new_n1070), .A2(new_n1097), .A3(G301), .ZN(new_n1098));
  AOI21_X1  g673(.A(G301), .B1(new_n1070), .B2(new_n1067), .ZN(new_n1099));
  OAI21_X1  g674(.A(new_n1094), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1091), .A2(new_n1093), .A3(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT57), .ZN(new_n1102));
  INV_X1    g677(.A(new_n574), .ZN(new_n1103));
  AND2_X1   g678(.A1(new_n566), .A2(new_n563), .ZN(new_n1104));
  INV_X1    g679(.A(new_n569), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n567), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1103), .B1(new_n1104), .B2(new_n1106), .ZN(new_n1107));
  OAI21_X1  g682(.A(new_n1102), .B1(new_n1107), .B2(KEYINPUT116), .ZN(new_n1108));
  INV_X1    g683(.A(KEYINPUT116), .ZN(new_n1109));
  NAND3_X1  g684(.A1(G299), .A2(new_n1109), .A3(KEYINPUT57), .ZN(new_n1110));
  NAND3_X1  g685(.A1(new_n940), .A2(new_n1018), .A3(new_n1020), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n820), .ZN(new_n1112));
  XNOR2_X1  g687(.A(KEYINPUT56), .B(G2072), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n940), .A2(new_n1024), .A3(new_n1023), .A4(new_n1113), .ZN(new_n1114));
  NAND4_X1  g689(.A1(new_n1108), .A2(new_n1110), .A3(new_n1112), .A4(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1116));
  AOI21_X1  g691(.A(KEYINPUT57), .B1(G299), .B2(new_n1109), .ZN(new_n1117));
  AOI211_X1 g692(.A(KEYINPUT116), .B(new_n1102), .C1(new_n570), .C2(new_n574), .ZN(new_n1118));
  OAI21_X1  g693(.A(new_n1116), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT117), .ZN(new_n1120));
  OAI21_X1  g695(.A(new_n1120), .B1(new_n992), .B2(G2067), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n986), .A2(new_n988), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1122), .A2(KEYINPUT117), .A3(new_n948), .ZN(new_n1123));
  AND2_X1   g698(.A1(new_n1121), .A2(new_n1123), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1032), .A2(new_n809), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n609), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n1119), .B1(new_n1126), .B2(KEYINPUT118), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1125), .A2(new_n1123), .A3(new_n1121), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1128), .A2(KEYINPUT118), .A3(new_n610), .ZN(new_n1129));
  INV_X1    g704(.A(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1115), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1131));
  AND4_X1   g706(.A1(new_n609), .A2(new_n1125), .A3(new_n1123), .A4(new_n1121), .ZN(new_n1132));
  OAI21_X1  g707(.A(KEYINPUT60), .B1(new_n1126), .B2(new_n1132), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT61), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1134), .A2(new_n1135), .ZN(new_n1136));
  XNOR2_X1  g711(.A(KEYINPUT58), .B(G1341), .ZN(new_n1137));
  OAI22_X1  g712(.A1(new_n1025), .A2(G1996), .B1(new_n1122), .B2(new_n1137), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT119), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n553), .B1(new_n1139), .B2(KEYINPUT59), .ZN(new_n1140));
  NAND2_X1  g715(.A1(new_n1138), .A2(new_n1140), .ZN(new_n1141));
  OR2_X1    g716(.A1(new_n1139), .A2(KEYINPUT59), .ZN(new_n1142));
  XOR2_X1   g717(.A(new_n1142), .B(KEYINPUT120), .Z(new_n1143));
  NAND2_X1  g718(.A1(new_n1141), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(KEYINPUT60), .ZN(new_n1145));
  AND3_X1   g720(.A1(new_n605), .A2(new_n1145), .A3(new_n608), .ZN(new_n1146));
  NAND4_X1  g721(.A1(new_n1146), .A2(new_n1125), .A3(new_n1123), .A4(new_n1121), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1143), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1138), .A2(new_n1140), .A3(new_n1148), .ZN(new_n1149));
  AND3_X1   g724(.A1(new_n1144), .A2(new_n1147), .A3(new_n1149), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1115), .A2(new_n1119), .A3(KEYINPUT61), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1133), .A2(new_n1136), .A3(new_n1150), .A4(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1101), .B1(new_n1131), .B2(new_n1152), .ZN(new_n1153));
  OAI211_X1 g728(.A(new_n1041), .B(G168), .C1(new_n1032), .C2(G2084), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1154), .A2(G8), .ZN(new_n1155));
  AOI21_X1  g730(.A(G168), .B1(new_n1038), .B2(new_n1041), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT51), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT121), .ZN(new_n1158));
  INV_X1    g733(.A(KEYINPUT51), .ZN(new_n1159));
  NAND3_X1  g734(.A1(new_n1154), .A2(new_n1159), .A3(G8), .ZN(new_n1160));
  AND3_X1   g735(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1158), .B1(new_n1157), .B2(new_n1160), .ZN(new_n1162));
  NOR2_X1   g737(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n1059), .B1(new_n1153), .B2(new_n1163), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT62), .ZN(new_n1165));
  OAI21_X1  g740(.A(new_n1165), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1157), .A2(new_n1160), .ZN(new_n1167));
  NAND2_X1  g742(.A1(new_n1167), .A2(KEYINPUT121), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1157), .A2(new_n1158), .A3(new_n1160), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1168), .A2(KEYINPUT62), .A3(new_n1169), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1093), .A2(new_n1099), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1166), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  AOI211_X1 g747(.A(new_n974), .B(new_n978), .C1(new_n1164), .C2(new_n1172), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1152), .A2(new_n1131), .ZN(new_n1174));
  INV_X1    g749(.A(new_n1101), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1174), .A2(new_n1163), .A3(new_n1175), .ZN(new_n1176));
  INV_X1    g751(.A(new_n1059), .ZN(new_n1177));
  NAND3_X1  g752(.A1(new_n1172), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(new_n978), .ZN(new_n1179));
  AOI21_X1  g754(.A(KEYINPUT126), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n973), .B1(new_n1173), .B2(new_n1180), .ZN(G329));
  assign    G231 = 1'b0;
  OAI21_X1  g756(.A(G319), .B1(new_n653), .B2(new_n654), .ZN(new_n1183));
  NOR3_X1   g757(.A1(G229), .A2(G227), .A3(new_n1183), .ZN(new_n1184));
  OAI211_X1 g758(.A(new_n879), .B(new_n1184), .C1(new_n924), .C2(new_n925), .ZN(G225));
  INV_X1    g759(.A(G225), .ZN(G308));
endmodule


