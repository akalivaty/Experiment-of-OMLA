//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 0 1 0 1 1 1 0 1 1 1 0 1 1 0 1 0 0 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:36 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n722, new_n723, new_n724,
    new_n725, new_n727, new_n728, new_n729, new_n730, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n842, new_n843, new_n844, new_n845, new_n847, new_n848, new_n849,
    new_n851, new_n852, new_n853, new_n854, new_n855, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n899, new_n900, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n971, new_n972;
  XOR2_X1   g000(.A(G141gat), .B(G148gat), .Z(new_n202));
  INV_X1    g001(.A(G155gat), .ZN(new_n203));
  INV_X1    g002(.A(G162gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G155gat), .A2(G162gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(KEYINPUT2), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n202), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  XNOR2_X1  g008(.A(G141gat), .B(G148gat), .ZN(new_n210));
  OAI211_X1 g009(.A(new_n206), .B(new_n205), .C1(new_n210), .C2(KEYINPUT2), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT3), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n209), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(KEYINPUT74), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT74), .ZN(new_n215));
  NAND4_X1  g014(.A1(new_n209), .A2(new_n211), .A3(new_n215), .A4(new_n212), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G127gat), .B(G134gat), .Z(new_n218));
  NOR2_X1   g017(.A1(new_n218), .A2(KEYINPUT1), .ZN(new_n219));
  INV_X1    g018(.A(G113gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n220), .A2(G120gat), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(KEYINPUT70), .ZN(new_n223));
  INV_X1    g022(.A(G120gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(G113gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n223), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n219), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n225), .A2(new_n221), .A3(KEYINPUT69), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT69), .B1(new_n225), .B2(new_n221), .ZN(new_n231));
  OAI21_X1  g030(.A(new_n218), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n227), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n209), .A2(new_n211), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(KEYINPUT3), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n217), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  INV_X1    g036(.A(new_n233), .ZN(new_n238));
  AND2_X1   g037(.A1(new_n209), .A2(new_n211), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n238), .A2(KEYINPUT4), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n232), .A3(new_n227), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  NAND4_X1  g042(.A1(new_n236), .A2(new_n237), .A3(new_n240), .A4(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(new_n237), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n233), .A2(new_n234), .ZN(new_n246));
  AOI22_X1  g045(.A1(new_n227), .A2(new_n232), .B1(new_n211), .B2(new_n209), .ZN(new_n247));
  OAI21_X1  g046(.A(new_n245), .B1(new_n246), .B2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT75), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  OAI211_X1 g049(.A(KEYINPUT75), .B(new_n245), .C1(new_n246), .C2(new_n247), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n244), .A2(new_n250), .A3(KEYINPUT5), .A4(new_n251), .ZN(new_n252));
  XNOR2_X1  g051(.A(G1gat), .B(G29gat), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n253), .B(KEYINPUT0), .ZN(new_n254));
  XNOR2_X1  g053(.A(G57gat), .B(G85gat), .ZN(new_n255));
  XOR2_X1   g054(.A(new_n254), .B(new_n255), .Z(new_n256));
  XNOR2_X1  g055(.A(new_n241), .B(KEYINPUT4), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT5), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n237), .A4(new_n236), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n252), .A2(new_n256), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT6), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n262), .A2(KEYINPUT76), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n252), .A2(new_n259), .ZN(new_n264));
  INV_X1    g063(.A(new_n256), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT76), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n260), .A2(new_n267), .A3(new_n261), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n263), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n256), .B1(new_n252), .B2(new_n259), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT6), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G8gat), .B(G36gat), .ZN(new_n273));
  XNOR2_X1  g072(.A(G64gat), .B(G92gat), .ZN(new_n274));
  XOR2_X1   g073(.A(new_n273), .B(new_n274), .Z(new_n275));
  INV_X1    g074(.A(new_n275), .ZN(new_n276));
  OR2_X1    g075(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n277));
  NAND2_X1  g076(.A1(KEYINPUT72), .A2(KEYINPUT22), .ZN(new_n278));
  INV_X1    g077(.A(G211gat), .ZN(new_n279));
  INV_X1    g078(.A(G218gat), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n278), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  XNOR2_X1  g080(.A(G211gat), .B(G218gat), .ZN(new_n282));
  XNOR2_X1  g081(.A(G197gat), .B(G204gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n281), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n282), .B1(new_n281), .B2(new_n283), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AND2_X1   g086(.A1(G226gat), .A2(G233gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT29), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT67), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT66), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT27), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G183gat), .ZN(new_n293));
  INV_X1    g092(.A(G183gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n291), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(G190gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n294), .A2(KEYINPUT27), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n292), .A2(G183gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n298), .A2(new_n299), .A3(KEYINPUT66), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n296), .A2(new_n297), .A3(new_n300), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n301), .A2(KEYINPUT28), .ZN(new_n302));
  NOR4_X1   g101(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT28), .A4(G190gat), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n290), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n303), .B1(new_n301), .B2(KEYINPUT28), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n305), .A2(KEYINPUT67), .ZN(new_n306));
  NAND2_X1  g105(.A1(G169gat), .A2(G176gat), .ZN(new_n307));
  OR2_X1    g106(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(KEYINPUT65), .ZN(new_n309));
  NOR2_X1   g108(.A1(G169gat), .A2(G176gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n311));
  AOI22_X1  g110(.A1(new_n308), .A2(new_n309), .B1(new_n311), .B2(KEYINPUT26), .ZN(new_n312));
  OR2_X1    g111(.A1(new_n311), .A2(KEYINPUT26), .ZN(new_n313));
  AOI22_X1  g112(.A1(new_n312), .A2(new_n313), .B1(G183gat), .B2(G190gat), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n304), .A2(new_n306), .A3(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n316), .A2(KEYINPUT64), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(KEYINPUT64), .ZN(new_n318));
  NAND3_X1  g117(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n319));
  OAI21_X1  g118(.A(new_n319), .B1(G183gat), .B2(G190gat), .ZN(new_n320));
  NOR3_X1   g119(.A1(new_n317), .A2(new_n318), .A3(new_n320), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT23), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n310), .B(new_n322), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n308), .A2(new_n309), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NOR2_X1   g124(.A1(new_n321), .A2(new_n325), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n320), .A2(new_n316), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n323), .A2(new_n324), .A3(KEYINPUT25), .ZN(new_n328));
  OAI22_X1  g127(.A1(new_n326), .A2(KEYINPUT25), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(KEYINPUT73), .B1(new_n315), .B2(new_n329), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n314), .B1(new_n305), .B2(KEYINPUT67), .ZN(new_n331));
  AOI211_X1 g130(.A(new_n290), .B(new_n303), .C1(new_n301), .C2(KEYINPUT28), .ZN(new_n332));
  OAI211_X1 g131(.A(new_n329), .B(KEYINPUT73), .C1(new_n331), .C2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  OAI21_X1  g133(.A(new_n289), .B1(new_n330), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n329), .B1(new_n331), .B2(new_n332), .ZN(new_n336));
  INV_X1    g135(.A(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n288), .ZN(new_n338));
  AOI21_X1  g137(.A(new_n287), .B1(new_n335), .B2(new_n338), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT73), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n336), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n341), .A2(new_n288), .A3(new_n333), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n336), .A2(new_n289), .ZN(new_n343));
  AND3_X1   g142(.A1(new_n342), .A2(new_n287), .A3(new_n343), .ZN(new_n344));
  OAI21_X1  g143(.A(new_n276), .B1(new_n339), .B2(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n342), .A2(new_n287), .A3(new_n343), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n341), .A2(new_n333), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n347), .A2(new_n289), .B1(new_n337), .B2(new_n288), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n346), .B(new_n275), .C1(new_n348), .C2(new_n287), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n345), .A2(KEYINPUT30), .A3(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n339), .A2(new_n344), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT30), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n351), .A2(new_n352), .A3(new_n275), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n350), .A2(new_n353), .ZN(new_n354));
  AND2_X1   g153(.A1(new_n272), .A2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(KEYINPUT82), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT29), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n217), .A2(new_n357), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT81), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n358), .A2(new_n359), .A3(new_n287), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n281), .A2(new_n283), .ZN(new_n361));
  INV_X1    g160(.A(new_n282), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(KEYINPUT29), .B1(new_n363), .B2(new_n284), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n212), .B1(new_n364), .B2(KEYINPUT80), .ZN(new_n365));
  OAI211_X1 g164(.A(KEYINPUT80), .B(new_n357), .C1(new_n285), .C2(new_n286), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g166(.A(new_n234), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT29), .B1(new_n214), .B2(new_n216), .ZN(new_n369));
  INV_X1    g168(.A(new_n287), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT81), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n360), .A2(new_n368), .A3(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G228gat), .A2(G233gat), .ZN(new_n373));
  INV_X1    g172(.A(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n364), .A2(KEYINPUT78), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n212), .B1(new_n364), .B2(KEYINPUT78), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n234), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n358), .A2(KEYINPUT79), .A3(new_n287), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT79), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n381), .B1(new_n369), .B2(new_n370), .ZN(new_n382));
  NAND4_X1  g181(.A1(new_n379), .A2(new_n380), .A3(new_n373), .A4(new_n382), .ZN(new_n383));
  AND3_X1   g182(.A1(new_n375), .A2(G22gat), .A3(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(G22gat), .B1(new_n375), .B2(new_n383), .ZN(new_n385));
  OAI21_X1  g184(.A(new_n356), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n375), .A2(new_n383), .ZN(new_n387));
  INV_X1    g186(.A(G22gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n375), .A2(G22gat), .A3(new_n383), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n389), .A2(KEYINPUT82), .A3(new_n390), .ZN(new_n391));
  XNOR2_X1  g190(.A(G78gat), .B(G106gat), .ZN(new_n392));
  INV_X1    g191(.A(G50gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  XOR2_X1   g193(.A(KEYINPUT77), .B(KEYINPUT31), .Z(new_n395));
  XNOR2_X1  g194(.A(new_n394), .B(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n386), .A2(new_n391), .A3(new_n397), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n389), .A2(KEYINPUT82), .A3(new_n390), .A4(new_n396), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT34), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n336), .A2(new_n238), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n329), .B(new_n233), .C1(new_n331), .C2(new_n332), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(G227gat), .A2(G233gat), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n401), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n404), .A2(new_n401), .A3(new_n405), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n406), .B1(KEYINPUT71), .B2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  NAND3_X1  g208(.A1(new_n402), .A2(new_n409), .A3(new_n403), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT32), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT33), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n410), .A2(new_n412), .ZN(new_n413));
  XOR2_X1   g212(.A(G15gat), .B(G43gat), .Z(new_n414));
  XNOR2_X1  g213(.A(G71gat), .B(G99gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n414), .B(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n411), .A2(new_n413), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(new_n416), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n410), .B(KEYINPUT32), .C1(new_n412), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT71), .ZN(new_n420));
  NAND4_X1  g219(.A1(new_n404), .A2(new_n420), .A3(new_n401), .A4(new_n405), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n408), .A2(new_n417), .A3(new_n419), .A4(new_n421), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n407), .A2(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n404), .A2(new_n405), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(KEYINPUT34), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n424), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n423), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n422), .A2(new_n428), .A3(KEYINPUT36), .ZN(new_n429));
  AOI21_X1  g228(.A(KEYINPUT36), .B1(new_n422), .B2(new_n428), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n355), .A2(new_n400), .B1(new_n429), .B2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n398), .A2(new_n399), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n237), .B1(new_n257), .B2(new_n236), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT39), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n265), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OR2_X1    g235(.A1(new_n246), .A2(new_n247), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT39), .B1(new_n437), .B2(new_n245), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n436), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(KEYINPUT40), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  OR3_X1    g240(.A1(new_n439), .A2(KEYINPUT83), .A3(new_n440), .ZN(new_n442));
  OAI21_X1  g241(.A(KEYINPUT83), .B1(new_n439), .B2(new_n440), .ZN(new_n443));
  AOI211_X1 g242(.A(new_n270), .B(new_n441), .C1(new_n442), .C2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(new_n354), .ZN(new_n445));
  AOI21_X1  g244(.A(new_n433), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT37), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n275), .B1(new_n351), .B2(new_n447), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n447), .B2(new_n351), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(KEYINPUT38), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n271), .B1(new_n262), .B2(new_n270), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n451), .B1(new_n275), .B2(new_n351), .ZN(new_n452));
  OR2_X1    g251(.A1(new_n348), .A2(new_n370), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n342), .A2(new_n370), .A3(new_n343), .ZN(new_n454));
  AND2_X1   g253(.A1(new_n454), .A2(KEYINPUT37), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT38), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n448), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT84), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT84), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n448), .A2(new_n456), .A3(new_n459), .ZN(new_n460));
  NAND4_X1  g259(.A1(new_n450), .A2(new_n452), .A3(new_n458), .A4(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n432), .A2(new_n462), .ZN(new_n463));
  AND3_X1   g262(.A1(new_n422), .A2(new_n428), .A3(KEYINPUT85), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT85), .B1(new_n422), .B2(new_n428), .ZN(new_n465));
  NOR2_X1   g264(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n266), .A2(new_n261), .A3(new_n260), .ZN(new_n467));
  AOI21_X1  g266(.A(KEYINPUT35), .B1(new_n467), .B2(new_n271), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n354), .A2(new_n399), .A3(new_n398), .A4(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(KEYINPUT86), .B1(new_n466), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT85), .ZN(new_n471));
  NOR2_X1   g270(.A1(new_n423), .A2(new_n427), .ZN(new_n472));
  AOI22_X1  g271(.A1(new_n408), .A2(new_n421), .B1(new_n417), .B2(new_n419), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n422), .A2(new_n428), .A3(KEYINPUT85), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(KEYINPUT35), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n451), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n478), .B1(new_n353), .B2(new_n350), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT86), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n476), .A2(new_n479), .A3(new_n480), .A4(new_n400), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n272), .A2(new_n354), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n398), .A2(new_n422), .A3(new_n428), .A4(new_n399), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT35), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n470), .A2(new_n481), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n463), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT100), .ZN(new_n487));
  XNOR2_X1  g286(.A(G190gat), .B(G218gat), .ZN(new_n488));
  INV_X1    g287(.A(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(G85gat), .A2(G92gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT7), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT101), .ZN(new_n492));
  NOR2_X1   g291(.A1(G85gat), .A2(G92gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(G99gat), .A2(G106gat), .ZN(new_n494));
  AOI211_X1 g293(.A(new_n492), .B(new_n493), .C1(KEYINPUT8), .C2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(G85gat), .ZN(new_n496));
  INV_X1    g295(.A(G92gat), .ZN(new_n497));
  AOI22_X1  g296(.A1(KEYINPUT8), .A2(new_n494), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NOR2_X1   g297(.A1(new_n498), .A2(KEYINPUT101), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n491), .B1(new_n495), .B2(new_n499), .ZN(new_n500));
  XOR2_X1   g299(.A(G99gat), .B(G106gat), .Z(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(new_n501), .ZN(new_n503));
  OAI211_X1 g302(.A(new_n503), .B(new_n491), .C1(new_n495), .C2(new_n499), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT102), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT102), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n504), .A3(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n393), .A2(G43gat), .ZN(new_n509));
  INV_X1    g308(.A(G43gat), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n510), .A2(G50gat), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n509), .A2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT15), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  INV_X1    g313(.A(G29gat), .ZN(new_n515));
  INV_X1    g314(.A(G36gat), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n515), .A2(new_n516), .A3(KEYINPUT14), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT14), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n518), .B1(G29gat), .B2(G36gat), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(KEYINPUT89), .B(G36gat), .ZN(new_n521));
  OAI211_X1 g320(.A(new_n514), .B(new_n520), .C1(new_n515), .C2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT91), .B1(new_n512), .B2(new_n513), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT91), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n509), .A2(new_n511), .A3(new_n524), .A4(KEYINPUT15), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n525), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n512), .A2(new_n513), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT88), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n517), .A2(new_n519), .A3(new_n529), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(new_n515), .B2(new_n521), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n529), .B1(new_n517), .B2(new_n519), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n528), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT90), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT90), .ZN(new_n535));
  OAI211_X1 g334(.A(new_n535), .B(new_n528), .C1(new_n531), .C2(new_n532), .ZN(new_n536));
  AOI21_X1  g335(.A(new_n527), .B1(new_n534), .B2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT17), .ZN(new_n538));
  NOR2_X1   g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  AOI211_X1 g338(.A(KEYINPUT17), .B(new_n527), .C1(new_n534), .C2(new_n536), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n506), .B(new_n508), .C1(new_n539), .C2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT41), .ZN(new_n542));
  NAND2_X1  g341(.A1(G232gat), .A2(G233gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n543), .B(KEYINPUT99), .ZN(new_n544));
  OAI22_X1  g343(.A1(new_n537), .A2(new_n505), .B1(new_n542), .B2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n545), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n489), .B1(new_n541), .B2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT103), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n487), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n506), .A2(new_n508), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n534), .A2(new_n536), .ZN(new_n551));
  INV_X1    g350(.A(new_n527), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT17), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n537), .A2(new_n538), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n550), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n488), .B1(new_n556), .B2(new_n545), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n489), .A3(new_n546), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(KEYINPUT103), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n542), .ZN(new_n560));
  XOR2_X1   g359(.A(G134gat), .B(G162gat), .Z(new_n561));
  XOR2_X1   g360(.A(new_n560), .B(new_n561), .Z(new_n562));
  AND3_X1   g361(.A1(new_n549), .A2(new_n559), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(new_n562), .B1(new_n549), .B2(new_n559), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(G8gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(G15gat), .B(G22gat), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n568), .A2(G1gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT16), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n568), .B1(new_n570), .B2(G1gat), .ZN(new_n571));
  AOI21_X1  g370(.A(new_n567), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n569), .A2(new_n567), .A3(new_n571), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(KEYINPUT92), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n573), .A2(KEYINPUT92), .A3(new_n574), .ZN(new_n578));
  NAND2_X1  g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(G57gat), .ZN(new_n580));
  INV_X1    g379(.A(G64gat), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G57gat), .A2(G64gat), .ZN(new_n583));
  AND2_X1   g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(KEYINPUT9), .ZN(new_n585));
  NOR2_X1   g384(.A1(G71gat), .A2(G78gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT95), .ZN(new_n587));
  NAND2_X1  g386(.A1(G71gat), .A2(G78gat), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI211_X1 g388(.A(new_n585), .B(new_n589), .C1(new_n587), .C2(new_n588), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT96), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n581), .B1(new_n591), .B2(new_n580), .ZN(new_n592));
  NAND3_X1  g391(.A1(KEYINPUT96), .A2(G57gat), .A3(G64gat), .ZN(new_n593));
  AND2_X1   g392(.A1(new_n586), .A2(KEYINPUT9), .ZN(new_n594));
  OAI211_X1 g393(.A(new_n592), .B(new_n593), .C1(new_n594), .C2(new_n584), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n590), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT98), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n590), .A2(KEYINPUT98), .A3(new_n595), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n598), .A2(KEYINPUT21), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n579), .A2(new_n600), .ZN(new_n601));
  AOI21_X1  g400(.A(KEYINPUT21), .B1(new_n590), .B2(new_n595), .ZN(new_n602));
  XOR2_X1   g401(.A(G127gat), .B(G155gat), .Z(new_n603));
  XNOR2_X1  g402(.A(new_n602), .B(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n601), .B(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G231gat), .A2(G233gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT97), .ZN(new_n607));
  XOR2_X1   g406(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G183gat), .B(G211gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n605), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n566), .A2(new_n613), .ZN(new_n614));
  OAI211_X1 g413(.A(new_n590), .B(new_n595), .C1(KEYINPUT104), .C2(new_n503), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n505), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT10), .ZN(new_n617));
  NOR2_X1   g416(.A1(new_n503), .A2(KEYINPUT104), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n596), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n619), .A2(new_n504), .A3(new_n502), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n616), .A2(new_n617), .A3(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(KEYINPUT105), .ZN(new_n622));
  AND2_X1   g421(.A1(new_n502), .A2(new_n504), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n623), .A2(KEYINPUT10), .A3(new_n598), .A4(new_n599), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n621), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n621), .B2(new_n624), .ZN(new_n626));
  NAND2_X1  g425(.A1(G230gat), .A2(G233gat), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  NOR3_X1   g427(.A1(new_n625), .A2(new_n626), .A3(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n616), .A2(new_n620), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n628), .ZN(new_n631));
  XOR2_X1   g430(.A(G120gat), .B(G148gat), .Z(new_n632));
  XNOR2_X1  g431(.A(new_n632), .B(KEYINPUT106), .ZN(new_n633));
  XNOR2_X1  g432(.A(G176gat), .B(G204gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NOR2_X1   g435(.A1(new_n629), .A2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n628), .B1(new_n621), .B2(new_n624), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n639), .B1(new_n630), .B2(new_n628), .ZN(new_n640));
  OR2_X1    g439(.A1(new_n640), .A2(new_n635), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n638), .A2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n614), .A2(new_n643), .ZN(new_n644));
  XNOR2_X1  g443(.A(G113gat), .B(G141gat), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(G197gat), .ZN(new_n646));
  XOR2_X1   g445(.A(KEYINPUT11), .B(G169gat), .Z(new_n647));
  XNOR2_X1  g446(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XOR2_X1   g447(.A(KEYINPUT87), .B(KEYINPUT12), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(KEYINPUT93), .ZN(new_n651));
  AOI21_X1  g450(.A(new_n575), .B1(new_n554), .B2(new_n555), .ZN(new_n652));
  AOI21_X1  g451(.A(KEYINPUT92), .B1(new_n573), .B2(new_n574), .ZN(new_n653));
  INV_X1    g452(.A(new_n574), .ZN(new_n654));
  NOR3_X1   g453(.A1(new_n654), .A2(new_n576), .A3(new_n572), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n553), .ZN(new_n657));
  NAND2_X1  g456(.A1(G229gat), .A2(G233gat), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n651), .B1(new_n652), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT18), .ZN(new_n661));
  INV_X1    g460(.A(new_n575), .ZN(new_n662));
  OAI21_X1  g461(.A(new_n662), .B1(new_n539), .B2(new_n540), .ZN(new_n663));
  AOI22_X1  g462(.A1(new_n656), .A2(new_n553), .B1(G229gat), .B2(G233gat), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n663), .A2(KEYINPUT93), .A3(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n660), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n663), .A2(KEYINPUT18), .A3(new_n664), .ZN(new_n667));
  XOR2_X1   g466(.A(new_n658), .B(KEYINPUT13), .Z(new_n668));
  NOR2_X1   g467(.A1(new_n579), .A2(new_n537), .ZN(new_n669));
  NOR2_X1   g468(.A1(new_n656), .A2(new_n553), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n668), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n650), .B1(new_n666), .B2(new_n672), .ZN(new_n673));
  AND3_X1   g472(.A1(new_n667), .A2(new_n671), .A3(new_n650), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n666), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(KEYINPUT94), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT94), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n666), .A2(new_n674), .A3(new_n677), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n673), .B1(new_n676), .B2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n644), .A2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n486), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n272), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g484(.A(KEYINPUT16), .B(G8gat), .Z(new_n686));
  AND3_X1   g485(.A1(new_n682), .A2(new_n445), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n567), .B1(new_n682), .B2(new_n445), .ZN(new_n688));
  OAI21_X1  g487(.A(KEYINPUT42), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT107), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n682), .A2(new_n445), .A3(new_n686), .ZN(new_n691));
  INV_X1    g490(.A(KEYINPUT42), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  AND3_X1   g492(.A1(new_n689), .A2(new_n690), .A3(new_n693), .ZN(new_n694));
  AOI21_X1  g493(.A(new_n690), .B1(new_n689), .B2(new_n693), .ZN(new_n695));
  NOR2_X1   g494(.A1(new_n694), .A2(new_n695), .ZN(G1325gat));
  OR3_X1    g495(.A1(new_n681), .A2(G15gat), .A3(new_n466), .ZN(new_n697));
  NOR2_X1   g496(.A1(new_n429), .A2(new_n430), .ZN(new_n698));
  INV_X1    g497(.A(new_n698), .ZN(new_n699));
  OAI21_X1  g498(.A(G15gat), .B1(new_n681), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n697), .A2(new_n700), .ZN(G1326gat));
  NOR2_X1   g500(.A1(new_n681), .A2(new_n400), .ZN(new_n702));
  XOR2_X1   g501(.A(KEYINPUT43), .B(G22gat), .Z(new_n703));
  XNOR2_X1  g502(.A(new_n702), .B(new_n703), .ZN(G1327gat));
  INV_X1    g503(.A(KEYINPUT44), .ZN(new_n705));
  AOI21_X1  g504(.A(new_n431), .B1(new_n461), .B2(new_n446), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n485), .A2(KEYINPUT108), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT108), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n470), .A2(new_n481), .A3(new_n708), .A4(new_n484), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n706), .B1(new_n707), .B2(new_n709), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n705), .B1(new_n710), .B2(new_n565), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n565), .B1(new_n463), .B2(new_n485), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n712), .A2(KEYINPUT44), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n711), .A2(new_n713), .ZN(new_n714));
  NOR3_X1   g513(.A1(new_n679), .A2(new_n612), .A3(new_n642), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(G29gat), .B1(new_n716), .B2(new_n272), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n712), .A2(new_n715), .ZN(new_n718));
  NOR3_X1   g517(.A1(new_n718), .A2(G29gat), .A3(new_n272), .ZN(new_n719));
  XOR2_X1   g518(.A(new_n719), .B(KEYINPUT45), .Z(new_n720));
  NAND2_X1  g519(.A1(new_n717), .A2(new_n720), .ZN(G1328gat));
  INV_X1    g520(.A(new_n521), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n722), .B1(new_n716), .B2(new_n354), .ZN(new_n723));
  NOR3_X1   g522(.A1(new_n718), .A2(new_n354), .A3(new_n722), .ZN(new_n724));
  XNOR2_X1  g523(.A(new_n724), .B(KEYINPUT46), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n723), .A2(new_n725), .ZN(G1329gat));
  NOR2_X1   g525(.A1(new_n699), .A2(new_n510), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n711), .A2(new_n713), .A3(new_n715), .A4(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(new_n510), .B1(new_n718), .B2(new_n466), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n728), .A2(new_n729), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(KEYINPUT47), .ZN(G1330gat));
  NOR2_X1   g530(.A1(new_n400), .A2(new_n393), .ZN(new_n732));
  NAND4_X1  g531(.A1(new_n711), .A2(new_n713), .A3(new_n715), .A4(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n393), .B1(new_n718), .B2(new_n400), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g534(.A(new_n735), .B(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g535(.A1(new_n614), .A2(new_n679), .A3(new_n642), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n710), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n738), .A2(new_n683), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g539(.A(new_n354), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n738), .A2(new_n741), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT109), .ZN(new_n743));
  OR2_X1    g542(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n744));
  XNOR2_X1  g543(.A(new_n743), .B(new_n744), .ZN(G1333gat));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n738), .A2(new_n746), .A3(new_n476), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n710), .A2(new_n699), .A3(new_n737), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n748), .B2(new_n746), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g549(.A1(new_n738), .A2(new_n433), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(G78gat), .ZN(G1335gat));
  INV_X1    g551(.A(new_n679), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n753), .A2(new_n612), .ZN(new_n754));
  INV_X1    g553(.A(new_n754), .ZN(new_n755));
  NOR2_X1   g554(.A1(new_n755), .A2(new_n643), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n711), .A2(new_n683), .A3(new_n713), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n496), .B1(new_n757), .B2(KEYINPUT110), .ZN(new_n758));
  OAI21_X1  g557(.A(new_n758), .B1(KEYINPUT110), .B2(new_n757), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n707), .A2(new_n709), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n565), .B1(new_n760), .B2(new_n463), .ZN(new_n761));
  AOI21_X1  g560(.A(KEYINPUT51), .B1(new_n761), .B2(new_n754), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  NOR4_X1   g562(.A1(new_n710), .A2(new_n763), .A3(new_n565), .A4(new_n755), .ZN(new_n764));
  OR2_X1    g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g564(.A1(new_n765), .A2(new_n496), .A3(new_n683), .A4(new_n642), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n759), .A2(new_n766), .ZN(G1336gat));
  NAND3_X1  g566(.A1(new_n445), .A2(new_n497), .A3(new_n642), .ZN(new_n768));
  XNOR2_X1  g567(.A(new_n768), .B(KEYINPUT111), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n762), .B2(new_n764), .ZN(new_n770));
  NAND4_X1  g569(.A1(new_n711), .A2(new_n445), .A3(new_n713), .A4(new_n756), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(G92gat), .ZN(new_n772));
  INV_X1    g571(.A(KEYINPUT112), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n770), .A2(new_n772), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(KEYINPUT52), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT52), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n770), .A2(new_n772), .A3(new_n773), .A4(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(G1337gat));
  NAND3_X1  g577(.A1(new_n714), .A2(new_n698), .A3(new_n756), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(G99gat), .ZN(new_n780));
  NOR3_X1   g579(.A1(new_n466), .A2(G99gat), .A3(new_n643), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1338gat));
  NOR3_X1   g582(.A1(new_n400), .A2(G106gat), .A3(new_n643), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(KEYINPUT114), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n785), .B1(new_n762), .B2(new_n764), .ZN(new_n786));
  NAND4_X1  g585(.A1(new_n711), .A2(new_n433), .A3(new_n713), .A4(new_n756), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n787), .A2(G106gat), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT113), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n789), .A2(new_n791), .A3(KEYINPUT53), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT53), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n786), .B(new_n788), .C1(new_n790), .C2(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n792), .A2(new_n794), .ZN(G1339gat));
  NAND3_X1  g594(.A1(new_n614), .A2(new_n679), .A3(new_n643), .ZN(new_n796));
  INV_X1    g595(.A(new_n796), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n658), .B1(new_n663), .B2(new_n657), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n669), .A2(new_n670), .A3(new_n668), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n648), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT115), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  OAI211_X1 g601(.A(KEYINPUT115), .B(new_n648), .C1(new_n798), .C2(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AND3_X1   g603(.A1(new_n666), .A2(new_n674), .A3(new_n677), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n677), .B1(new_n666), .B2(new_n674), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n642), .B(new_n804), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(KEYINPUT54), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n635), .B1(new_n639), .B2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n621), .A2(new_n624), .A3(new_n628), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(KEYINPUT54), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n629), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT55), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n637), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(KEYINPUT55), .B(new_n809), .C1(new_n629), .C2(new_n811), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n807), .B1(new_n679), .B2(new_n816), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n817), .A2(new_n565), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n814), .B(new_n815), .C1(new_n563), .C2(new_n564), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n804), .B1(new_n805), .B2(new_n806), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g620(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n818), .A2(new_n822), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT116), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n612), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  AOI21_X1  g624(.A(new_n821), .B1(new_n817), .B2(new_n565), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n826), .A2(KEYINPUT116), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n797), .B1(new_n825), .B2(new_n827), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n445), .A2(new_n272), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  NOR4_X1   g629(.A1(new_n828), .A2(new_n466), .A3(new_n433), .A4(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n831), .A2(new_n753), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n832), .A2(G113gat), .ZN(new_n833));
  NOR2_X1   g632(.A1(new_n828), .A2(new_n272), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n483), .A2(new_n445), .ZN(new_n835));
  NAND4_X1  g634(.A1(new_n834), .A2(new_n220), .A3(new_n753), .A4(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n837), .A2(KEYINPUT117), .ZN(new_n838));
  INV_X1    g637(.A(KEYINPUT117), .ZN(new_n839));
  NAND3_X1  g638(.A1(new_n833), .A2(new_n839), .A3(new_n836), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n838), .A2(new_n840), .ZN(G1340gat));
  NAND2_X1  g640(.A1(new_n834), .A2(new_n835), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  AOI21_X1  g642(.A(G120gat), .B1(new_n843), .B2(new_n642), .ZN(new_n844));
  NOR2_X1   g643(.A1(new_n643), .A2(new_n224), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n831), .B2(new_n845), .ZN(G1341gat));
  INV_X1    g645(.A(G127gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n843), .A2(new_n847), .A3(new_n612), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n831), .A2(new_n612), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n848), .B1(new_n847), .B2(new_n849), .ZN(G1342gat));
  OR4_X1    g649(.A1(KEYINPUT56), .A2(new_n842), .A3(G134gat), .A4(new_n565), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n831), .A2(new_n566), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n852), .A2(G134gat), .ZN(new_n853));
  OR2_X1    g652(.A1(new_n565), .A2(G134gat), .ZN(new_n854));
  OAI21_X1  g653(.A(KEYINPUT56), .B1(new_n842), .B2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n853), .A3(new_n855), .ZN(G1343gat));
  NOR2_X1   g655(.A1(new_n830), .A2(new_n698), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n613), .B1(new_n826), .B2(KEYINPUT116), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n824), .B(new_n821), .C1(new_n565), .C2(new_n817), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n796), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n860), .B2(new_n433), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n433), .A2(KEYINPUT57), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n823), .A2(new_n613), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n796), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n857), .B1(new_n861), .B2(new_n864), .ZN(new_n865));
  OAI21_X1  g664(.A(G141gat), .B1(new_n865), .B2(new_n679), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n698), .A2(new_n400), .ZN(new_n867));
  AND4_X1   g666(.A1(new_n683), .A2(new_n860), .A3(new_n354), .A4(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(G141gat), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n868), .A2(new_n869), .A3(new_n753), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n866), .A2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT58), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n872), .B1(new_n870), .B2(KEYINPUT118), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  OAI211_X1 g673(.A(new_n866), .B(new_n870), .C1(KEYINPUT118), .C2(new_n872), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1344gat));
  NAND2_X1  g675(.A1(new_n857), .A2(new_n642), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n797), .A2(KEYINPUT120), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT120), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n796), .A2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n863), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g680(.A(KEYINPUT57), .B1(new_n881), .B2(new_n433), .ZN(new_n882));
  INV_X1    g681(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n860), .A2(KEYINPUT57), .A3(new_n433), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n877), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(G148gat), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  OAI211_X1 g686(.A(new_n642), .B(new_n857), .C1(new_n861), .C2(new_n864), .ZN(new_n888));
  INV_X1    g687(.A(KEYINPUT119), .ZN(new_n889));
  NOR2_X1   g688(.A1(new_n886), .A2(KEYINPUT59), .ZN(new_n890));
  AND3_X1   g689(.A1(new_n888), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n888), .B2(new_n890), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n887), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n868), .A2(new_n886), .A3(new_n642), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(G1345gat));
  OAI21_X1  g694(.A(G155gat), .B1(new_n865), .B2(new_n613), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n868), .A2(new_n203), .A3(new_n612), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n896), .A2(new_n897), .ZN(G1346gat));
  OAI21_X1  g697(.A(G162gat), .B1(new_n865), .B2(new_n565), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n868), .A2(new_n204), .A3(new_n566), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(G1347gat));
  NOR2_X1   g700(.A1(new_n483), .A2(new_n354), .ZN(new_n902));
  INV_X1    g701(.A(new_n902), .ZN(new_n903));
  OAI21_X1  g702(.A(KEYINPUT121), .B1(new_n828), .B2(new_n683), .ZN(new_n904));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n860), .A2(new_n905), .A3(new_n272), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n903), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n679), .A2(G169gat), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  INV_X1    g708(.A(KEYINPUT123), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n828), .A2(new_n433), .ZN(new_n911));
  NAND3_X1  g710(.A1(new_n476), .A2(new_n272), .A3(new_n445), .ZN(new_n912));
  XOR2_X1   g711(.A(new_n912), .B(KEYINPUT122), .Z(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(new_n914));
  OAI21_X1  g713(.A(G169gat), .B1(new_n914), .B2(new_n679), .ZN(new_n915));
  AND3_X1   g714(.A1(new_n909), .A2(new_n910), .A3(new_n915), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n910), .B1(new_n909), .B2(new_n915), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(G1348gat));
  AOI21_X1  g717(.A(G176gat), .B1(new_n907), .B2(new_n642), .ZN(new_n919));
  INV_X1    g718(.A(G176gat), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n643), .A2(new_n920), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n860), .A2(new_n400), .A3(new_n913), .A4(new_n921), .ZN(new_n922));
  XNOR2_X1  g721(.A(new_n922), .B(KEYINPUT124), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OAI21_X1  g723(.A(KEYINPUT125), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n904), .A2(new_n906), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n642), .A3(new_n902), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n920), .ZN(new_n928));
  INV_X1    g727(.A(KEYINPUT125), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n928), .A2(new_n929), .A3(new_n923), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n925), .A2(new_n930), .ZN(G1349gat));
  AND3_X1   g730(.A1(new_n612), .A2(new_n296), .A3(new_n300), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n907), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G183gat), .B1(new_n914), .B2(new_n613), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n935), .A2(KEYINPUT60), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT60), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n933), .A2(new_n937), .A3(new_n934), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n936), .A2(new_n938), .ZN(G1350gat));
  NAND3_X1  g738(.A1(new_n907), .A2(new_n297), .A3(new_n566), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n911), .A2(new_n566), .A3(new_n913), .ZN(new_n941));
  NOR2_X1   g740(.A1(KEYINPUT126), .A2(KEYINPUT61), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n297), .B1(KEYINPUT126), .B2(KEYINPUT61), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n941), .A2(new_n942), .A3(new_n943), .ZN(new_n944));
  AOI21_X1  g743(.A(new_n942), .B1(new_n941), .B2(new_n943), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n940), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  NAND2_X1  g745(.A1(new_n883), .A2(new_n884), .ZN(new_n947));
  NOR3_X1   g746(.A1(new_n698), .A2(new_n683), .A3(new_n354), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  INV_X1    g749(.A(G197gat), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n679), .A2(new_n951), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n867), .A2(new_n445), .ZN(new_n953));
  INV_X1    g752(.A(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n926), .A2(new_n753), .A3(new_n954), .ZN(new_n955));
  AOI22_X1  g754(.A1(new_n950), .A2(new_n952), .B1(new_n955), .B2(new_n951), .ZN(G1352gat));
  XOR2_X1   g755(.A(KEYINPUT127), .B(G204gat), .Z(new_n957));
  NOR2_X1   g756(.A1(new_n643), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n926), .A2(new_n954), .A3(new_n958), .ZN(new_n959));
  OR2_X1    g758(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n960));
  OAI21_X1  g759(.A(new_n957), .B1(new_n949), .B2(new_n643), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n959), .A2(KEYINPUT62), .ZN(new_n962));
  NAND3_X1  g761(.A1(new_n960), .A2(new_n961), .A3(new_n962), .ZN(G1353gat));
  INV_X1    g762(.A(new_n884), .ZN(new_n964));
  OAI211_X1 g763(.A(new_n612), .B(new_n948), .C1(new_n964), .C2(new_n882), .ZN(new_n965));
  AND3_X1   g764(.A1(new_n965), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n966));
  AOI21_X1  g765(.A(KEYINPUT63), .B1(new_n965), .B2(G211gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n926), .A2(new_n954), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n612), .A2(new_n279), .ZN(new_n969));
  OAI22_X1  g768(.A1(new_n966), .A2(new_n967), .B1(new_n968), .B2(new_n969), .ZN(G1354gat));
  OAI21_X1  g769(.A(G218gat), .B1(new_n949), .B2(new_n565), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n566), .A2(new_n280), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n971), .B1(new_n968), .B2(new_n972), .ZN(G1355gat));
endmodule


