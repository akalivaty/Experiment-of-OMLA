

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591;

  XNOR2_X1 U326 ( .A(n506), .B(KEYINPUT113), .ZN(n507) );
  XNOR2_X1 U327 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U328 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U329 ( .A(n329), .B(n328), .ZN(n331) );
  NOR2_X1 U330 ( .A1(n560), .A2(n559), .ZN(n570) );
  XOR2_X1 U331 ( .A(KEYINPUT4), .B(KEYINPUT5), .Z(n295) );
  XNOR2_X1 U332 ( .A(G57GAT), .B(KEYINPUT1), .ZN(n294) );
  XNOR2_X1 U333 ( .A(n295), .B(n294), .ZN(n302) );
  XOR2_X1 U334 ( .A(G85GAT), .B(G162GAT), .Z(n297) );
  XNOR2_X1 U335 ( .A(G141GAT), .B(G148GAT), .ZN(n296) );
  XNOR2_X1 U336 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U337 ( .A(n298), .B(G127GAT), .Z(n300) );
  XOR2_X1 U338 ( .A(G113GAT), .B(G1GAT), .Z(n314) );
  XNOR2_X1 U339 ( .A(G29GAT), .B(n314), .ZN(n299) );
  XNOR2_X1 U340 ( .A(n300), .B(n299), .ZN(n301) );
  XNOR2_X1 U341 ( .A(n302), .B(n301), .ZN(n311) );
  XOR2_X1 U342 ( .A(KEYINPUT93), .B(KEYINPUT94), .Z(n304) );
  NAND2_X1 U343 ( .A1(G225GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U344 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U345 ( .A(n305), .B(KEYINPUT6), .Z(n309) );
  XNOR2_X1 U346 ( .A(G134GAT), .B(G120GAT), .ZN(n306) );
  XNOR2_X1 U347 ( .A(n306), .B(KEYINPUT0), .ZN(n416) );
  XNOR2_X1 U348 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n307) );
  XNOR2_X1 U349 ( .A(n307), .B(KEYINPUT2), .ZN(n427) );
  XNOR2_X1 U350 ( .A(n416), .B(n427), .ZN(n308) );
  XNOR2_X1 U351 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U352 ( .A(n311), .B(n310), .ZN(n553) );
  XOR2_X1 U353 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n313) );
  XNOR2_X1 U354 ( .A(G15GAT), .B(G197GAT), .ZN(n312) );
  XNOR2_X1 U355 ( .A(n313), .B(n312), .ZN(n337) );
  XOR2_X1 U356 ( .A(G36GAT), .B(G50GAT), .Z(n316) );
  XOR2_X1 U357 ( .A(G169GAT), .B(G8GAT), .Z(n406) );
  XNOR2_X1 U358 ( .A(n406), .B(n314), .ZN(n315) );
  XNOR2_X1 U359 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U360 ( .A(G141GAT), .B(G22GAT), .Z(n432) );
  XOR2_X1 U361 ( .A(n317), .B(n432), .Z(n330) );
  INV_X1 U362 ( .A(G29GAT), .ZN(n318) );
  NAND2_X1 U363 ( .A1(n318), .A2(G43GAT), .ZN(n321) );
  INV_X1 U364 ( .A(G43GAT), .ZN(n319) );
  NAND2_X1 U365 ( .A1(n319), .A2(G29GAT), .ZN(n320) );
  NAND2_X1 U366 ( .A1(n321), .A2(n320), .ZN(n323) );
  XNOR2_X1 U367 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n322) );
  XNOR2_X1 U368 ( .A(n323), .B(n322), .ZN(n386) );
  XOR2_X1 U369 ( .A(n386), .B(KEYINPUT70), .Z(n329) );
  XOR2_X1 U370 ( .A(KEYINPUT71), .B(KEYINPUT67), .Z(n325) );
  XNOR2_X1 U371 ( .A(KEYINPUT68), .B(KEYINPUT30), .ZN(n324) );
  XNOR2_X1 U372 ( .A(n325), .B(n324), .ZN(n327) );
  NAND2_X1 U373 ( .A1(G229GAT), .A2(G233GAT), .ZN(n326) );
  NAND2_X1 U374 ( .A1(n330), .A2(n331), .ZN(n335) );
  INV_X1 U375 ( .A(n330), .ZN(n333) );
  INV_X1 U376 ( .A(n331), .ZN(n332) );
  NAND2_X1 U377 ( .A1(n333), .A2(n332), .ZN(n334) );
  NAND2_X1 U378 ( .A1(n335), .A2(n334), .ZN(n336) );
  XOR2_X1 U379 ( .A(n337), .B(n336), .Z(n517) );
  XOR2_X1 U380 ( .A(KEYINPUT73), .B(KEYINPUT77), .Z(n339) );
  XNOR2_X1 U381 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n338) );
  XNOR2_X1 U382 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U383 ( .A(KEYINPUT32), .B(G120GAT), .Z(n341) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n340) );
  XNOR2_X1 U385 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U386 ( .A(n343), .B(n342), .Z(n349) );
  XOR2_X1 U387 ( .A(G64GAT), .B(KEYINPUT76), .Z(n345) );
  XNOR2_X1 U388 ( .A(G176GAT), .B(G204GAT), .ZN(n344) );
  XNOR2_X1 U389 ( .A(n345), .B(n344), .ZN(n403) );
  XOR2_X1 U390 ( .A(KEYINPUT72), .B(KEYINPUT13), .Z(n347) );
  XNOR2_X1 U391 ( .A(G71GAT), .B(G57GAT), .ZN(n346) );
  XNOR2_X1 U392 ( .A(n347), .B(n346), .ZN(n368) );
  XNOR2_X1 U393 ( .A(n403), .B(n368), .ZN(n348) );
  XNOR2_X1 U394 ( .A(n349), .B(n348), .ZN(n355) );
  XOR2_X1 U395 ( .A(G78GAT), .B(G148GAT), .Z(n351) );
  XNOR2_X1 U396 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n350) );
  XNOR2_X1 U397 ( .A(n351), .B(n350), .ZN(n428) );
  XOR2_X1 U398 ( .A(KEYINPUT75), .B(G92GAT), .Z(n353) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .ZN(n352) );
  XNOR2_X1 U400 ( .A(n353), .B(n352), .ZN(n385) );
  XOR2_X1 U401 ( .A(n428), .B(n385), .Z(n354) );
  XNOR2_X1 U402 ( .A(n355), .B(n354), .ZN(n580) );
  NAND2_X1 U403 ( .A1(n517), .A2(n580), .ZN(n471) );
  XOR2_X1 U404 ( .A(KEYINPUT84), .B(KEYINPUT16), .Z(n390) );
  XOR2_X1 U405 ( .A(G64GAT), .B(KEYINPUT81), .Z(n357) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(G211GAT), .ZN(n356) );
  XNOR2_X1 U407 ( .A(n357), .B(n356), .ZN(n361) );
  XOR2_X1 U408 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n359) );
  XNOR2_X1 U409 ( .A(G1GAT), .B(KEYINPUT15), .ZN(n358) );
  XNOR2_X1 U410 ( .A(n359), .B(n358), .ZN(n360) );
  XNOR2_X1 U411 ( .A(n361), .B(n360), .ZN(n372) );
  XOR2_X1 U412 ( .A(G15GAT), .B(G127GAT), .Z(n412) );
  XOR2_X1 U413 ( .A(G155GAT), .B(G78GAT), .Z(n363) );
  XNOR2_X1 U414 ( .A(G22GAT), .B(G183GAT), .ZN(n362) );
  XNOR2_X1 U415 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U416 ( .A(n412), .B(n364), .Z(n366) );
  NAND2_X1 U417 ( .A1(G231GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U418 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U419 ( .A(n367), .B(KEYINPUT83), .Z(n370) );
  XNOR2_X1 U420 ( .A(n368), .B(KEYINPUT82), .ZN(n369) );
  XNOR2_X1 U421 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U422 ( .A(n372), .B(n371), .ZN(n585) );
  XOR2_X1 U423 ( .A(KEYINPUT66), .B(KEYINPUT10), .Z(n374) );
  XNOR2_X1 U424 ( .A(G106GAT), .B(KEYINPUT79), .ZN(n373) );
  XNOR2_X1 U425 ( .A(n374), .B(n373), .ZN(n378) );
  XOR2_X1 U426 ( .A(G36GAT), .B(G190GAT), .Z(n405) );
  XOR2_X1 U427 ( .A(KEYINPUT11), .B(n405), .Z(n376) );
  XOR2_X1 U428 ( .A(G50GAT), .B(G162GAT), .Z(n431) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(n431), .ZN(n375) );
  XNOR2_X1 U430 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U431 ( .A(n378), .B(n377), .Z(n380) );
  NAND2_X1 U432 ( .A1(G232GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U433 ( .A(n380), .B(n379), .ZN(n384) );
  XOR2_X1 U434 ( .A(KEYINPUT78), .B(KEYINPUT80), .Z(n382) );
  XNOR2_X1 U435 ( .A(G134GAT), .B(KEYINPUT9), .ZN(n381) );
  XNOR2_X1 U436 ( .A(n382), .B(n381), .ZN(n383) );
  XOR2_X1 U437 ( .A(n384), .B(n383), .Z(n388) );
  XNOR2_X1 U438 ( .A(n386), .B(n385), .ZN(n387) );
  XNOR2_X1 U439 ( .A(n388), .B(n387), .ZN(n536) );
  NAND2_X1 U440 ( .A1(n585), .A2(n536), .ZN(n389) );
  XNOR2_X1 U441 ( .A(n390), .B(n389), .ZN(n456) );
  XOR2_X1 U442 ( .A(KEYINPUT95), .B(KEYINPUT81), .Z(n392) );
  NAND2_X1 U443 ( .A1(G226GAT), .A2(G233GAT), .ZN(n391) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XOR2_X1 U445 ( .A(n393), .B(G92GAT), .Z(n402) );
  XOR2_X1 U446 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n395) );
  XNOR2_X1 U447 ( .A(KEYINPUT87), .B(G183GAT), .ZN(n394) );
  XNOR2_X1 U448 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U449 ( .A(KEYINPUT18), .B(n396), .Z(n424) );
  XNOR2_X1 U450 ( .A(G211GAT), .B(KEYINPUT92), .ZN(n397) );
  XNOR2_X1 U451 ( .A(n397), .B(KEYINPUT91), .ZN(n398) );
  XOR2_X1 U452 ( .A(n398), .B(KEYINPUT21), .Z(n400) );
  XNOR2_X1 U453 ( .A(G197GAT), .B(G218GAT), .ZN(n399) );
  XNOR2_X1 U454 ( .A(n400), .B(n399), .ZN(n442) );
  XNOR2_X1 U455 ( .A(n424), .B(n442), .ZN(n401) );
  XNOR2_X1 U456 ( .A(n402), .B(n401), .ZN(n404) );
  XOR2_X1 U457 ( .A(n404), .B(n403), .Z(n408) );
  XNOR2_X1 U458 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U459 ( .A(n408), .B(n407), .ZN(n551) );
  XNOR2_X1 U460 ( .A(n551), .B(KEYINPUT27), .ZN(n446) );
  NOR2_X1 U461 ( .A1(n553), .A2(n446), .ZN(n409) );
  XOR2_X1 U462 ( .A(KEYINPUT96), .B(n409), .Z(n522) );
  XOR2_X1 U463 ( .A(KEYINPUT85), .B(G71GAT), .Z(n411) );
  XNOR2_X1 U464 ( .A(G190GAT), .B(G99GAT), .ZN(n410) );
  XNOR2_X1 U465 ( .A(n411), .B(n410), .ZN(n413) );
  XOR2_X1 U466 ( .A(n413), .B(n412), .Z(n415) );
  XNOR2_X1 U467 ( .A(G43GAT), .B(G113GAT), .ZN(n414) );
  XNOR2_X1 U468 ( .A(n415), .B(n414), .ZN(n420) );
  XOR2_X1 U469 ( .A(n416), .B(KEYINPUT86), .Z(n418) );
  NAND2_X1 U470 ( .A1(G227GAT), .A2(G233GAT), .ZN(n417) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U472 ( .A(n420), .B(n419), .Z(n426) );
  XOR2_X1 U473 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n422) );
  XNOR2_X1 U474 ( .A(G169GAT), .B(G176GAT), .ZN(n421) );
  XNOR2_X1 U475 ( .A(n422), .B(n421), .ZN(n423) );
  XNOR2_X1 U476 ( .A(n424), .B(n423), .ZN(n425) );
  XNOR2_X1 U477 ( .A(n426), .B(n425), .ZN(n560) );
  XNOR2_X1 U478 ( .A(n428), .B(n427), .ZN(n440) );
  XOR2_X1 U479 ( .A(KEYINPUT90), .B(KEYINPUT89), .Z(n430) );
  XNOR2_X1 U480 ( .A(G204GAT), .B(KEYINPUT24), .ZN(n429) );
  XNOR2_X1 U481 ( .A(n430), .B(n429), .ZN(n436) );
  XOR2_X1 U482 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n434) );
  XNOR2_X1 U483 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U484 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U485 ( .A(n436), .B(n435), .Z(n438) );
  NAND2_X1 U486 ( .A1(G228GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U487 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U488 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U489 ( .A(n442), .B(n441), .ZN(n556) );
  XNOR2_X1 U490 ( .A(KEYINPUT28), .B(n556), .ZN(n525) );
  NAND2_X1 U491 ( .A1(n560), .A2(n525), .ZN(n443) );
  NOR2_X1 U492 ( .A1(n522), .A2(n443), .ZN(n444) );
  XNOR2_X1 U493 ( .A(n444), .B(KEYINPUT97), .ZN(n455) );
  INV_X1 U494 ( .A(n560), .ZN(n523) );
  NOR2_X1 U495 ( .A1(n556), .A2(n523), .ZN(n445) );
  XNOR2_X1 U496 ( .A(n445), .B(KEYINPUT26), .ZN(n576) );
  INV_X1 U497 ( .A(n576), .ZN(n447) );
  NOR2_X1 U498 ( .A1(n447), .A2(n446), .ZN(n448) );
  XOR2_X1 U499 ( .A(KEYINPUT98), .B(n448), .Z(n452) );
  OR2_X1 U500 ( .A1(n560), .A2(n551), .ZN(n449) );
  NAND2_X1 U501 ( .A1(n556), .A2(n449), .ZN(n450) );
  XOR2_X1 U502 ( .A(KEYINPUT25), .B(n450), .Z(n451) );
  NAND2_X1 U503 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U504 ( .A1(n553), .A2(n453), .ZN(n454) );
  NAND2_X1 U505 ( .A1(n455), .A2(n454), .ZN(n467) );
  NAND2_X1 U506 ( .A1(n456), .A2(n467), .ZN(n482) );
  OR2_X1 U507 ( .A1(n471), .A2(n482), .ZN(n464) );
  NOR2_X1 U508 ( .A1(n553), .A2(n464), .ZN(n458) );
  XNOR2_X1 U509 ( .A(KEYINPUT99), .B(KEYINPUT34), .ZN(n457) );
  XNOR2_X1 U510 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U511 ( .A(G1GAT), .B(n459), .ZN(G1324GAT) );
  NOR2_X1 U512 ( .A1(n551), .A2(n464), .ZN(n460) );
  XOR2_X1 U513 ( .A(G8GAT), .B(n460), .Z(G1325GAT) );
  NOR2_X1 U514 ( .A1(n560), .A2(n464), .ZN(n462) );
  XNOR2_X1 U515 ( .A(KEYINPUT100), .B(KEYINPUT35), .ZN(n461) );
  XNOR2_X1 U516 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U517 ( .A(G15GAT), .B(n463), .ZN(G1326GAT) );
  NOR2_X1 U518 ( .A1(n525), .A2(n464), .ZN(n466) );
  XNOR2_X1 U519 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n465) );
  XNOR2_X1 U520 ( .A(n466), .B(n465), .ZN(G1327GAT) );
  XNOR2_X1 U521 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n474) );
  XNOR2_X1 U522 ( .A(KEYINPUT36), .B(n536), .ZN(n589) );
  INV_X1 U523 ( .A(n585), .ZN(n513) );
  NAND2_X1 U524 ( .A1(n513), .A2(n467), .ZN(n468) );
  NOR2_X1 U525 ( .A1(n589), .A2(n468), .ZN(n470) );
  XNOR2_X1 U526 ( .A(KEYINPUT102), .B(KEYINPUT37), .ZN(n469) );
  XNOR2_X1 U527 ( .A(n470), .B(n469), .ZN(n494) );
  NOR2_X1 U528 ( .A1(n494), .A2(n471), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT38), .B(n472), .Z(n479) );
  NOR2_X1 U530 ( .A1(n553), .A2(n479), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n474), .B(n473), .ZN(G1328GAT) );
  NOR2_X1 U532 ( .A1(n551), .A2(n479), .ZN(n475) );
  XOR2_X1 U533 ( .A(G36GAT), .B(n475), .Z(G1329GAT) );
  XNOR2_X1 U534 ( .A(KEYINPUT40), .B(KEYINPUT103), .ZN(n477) );
  NOR2_X1 U535 ( .A1(n560), .A2(n479), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(G43GAT), .B(n478), .ZN(G1330GAT) );
  NOR2_X1 U538 ( .A1(n525), .A2(n479), .ZN(n480) );
  XOR2_X1 U539 ( .A(G50GAT), .B(n480), .Z(G1331GAT) );
  XNOR2_X1 U540 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n481), .B(n580), .ZN(n543) );
  XNOR2_X1 U542 ( .A(KEYINPUT104), .B(n543), .ZN(n562) );
  INV_X1 U543 ( .A(n517), .ZN(n528) );
  NAND2_X1 U544 ( .A1(n562), .A2(n528), .ZN(n493) );
  OR2_X1 U545 ( .A1(n493), .A2(n482), .ZN(n489) );
  NOR2_X1 U546 ( .A1(n553), .A2(n489), .ZN(n483) );
  XOR2_X1 U547 ( .A(n483), .B(KEYINPUT42), .Z(n484) );
  XNOR2_X1 U548 ( .A(G57GAT), .B(n484), .ZN(G1332GAT) );
  NOR2_X1 U549 ( .A1(n551), .A2(n489), .ZN(n485) );
  XOR2_X1 U550 ( .A(G64GAT), .B(n485), .Z(G1333GAT) );
  NOR2_X1 U551 ( .A1(n560), .A2(n489), .ZN(n487) );
  XNOR2_X1 U552 ( .A(KEYINPUT105), .B(KEYINPUT106), .ZN(n486) );
  XNOR2_X1 U553 ( .A(n487), .B(n486), .ZN(n488) );
  XNOR2_X1 U554 ( .A(G71GAT), .B(n488), .ZN(G1334GAT) );
  NOR2_X1 U555 ( .A1(n525), .A2(n489), .ZN(n491) );
  XNOR2_X1 U556 ( .A(KEYINPUT107), .B(KEYINPUT43), .ZN(n490) );
  XNOR2_X1 U557 ( .A(n491), .B(n490), .ZN(n492) );
  XOR2_X1 U558 ( .A(G78GAT), .B(n492), .Z(G1335GAT) );
  XNOR2_X1 U559 ( .A(G85GAT), .B(KEYINPUT109), .ZN(n497) );
  NOR2_X1 U560 ( .A1(n494), .A2(n493), .ZN(n495) );
  XOR2_X1 U561 ( .A(KEYINPUT108), .B(n495), .Z(n503) );
  NOR2_X1 U562 ( .A1(n553), .A2(n503), .ZN(n496) );
  XNOR2_X1 U563 ( .A(n497), .B(n496), .ZN(G1336GAT) );
  NOR2_X1 U564 ( .A1(n551), .A2(n503), .ZN(n498) );
  XOR2_X1 U565 ( .A(KEYINPUT110), .B(n498), .Z(n499) );
  XNOR2_X1 U566 ( .A(G92GAT), .B(n499), .ZN(G1337GAT) );
  NOR2_X1 U567 ( .A1(n560), .A2(n503), .ZN(n500) );
  XOR2_X1 U568 ( .A(G99GAT), .B(n500), .Z(G1338GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT44), .B(KEYINPUT111), .Z(n502) );
  XNOR2_X1 U570 ( .A(G106GAT), .B(KEYINPUT112), .ZN(n501) );
  XNOR2_X1 U571 ( .A(n502), .B(n501), .ZN(n505) );
  NOR2_X1 U572 ( .A1(n525), .A2(n503), .ZN(n504) );
  XOR2_X1 U573 ( .A(n505), .B(n504), .Z(G1339GAT) );
  AND2_X1 U574 ( .A1(n543), .A2(n517), .ZN(n508) );
  INV_X1 U575 ( .A(KEYINPUT46), .ZN(n506) );
  NOR2_X1 U576 ( .A1(n585), .A2(n509), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n510), .B(KEYINPUT114), .ZN(n511) );
  NAND2_X1 U578 ( .A1(n511), .A2(n536), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n512), .B(KEYINPUT47), .ZN(n520) );
  NOR2_X1 U580 ( .A1(n589), .A2(n513), .ZN(n515) );
  XOR2_X1 U581 ( .A(KEYINPUT45), .B(KEYINPUT115), .Z(n514) );
  XNOR2_X1 U582 ( .A(n515), .B(n514), .ZN(n516) );
  NAND2_X1 U583 ( .A1(n580), .A2(n516), .ZN(n518) );
  NOR2_X1 U584 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U585 ( .A1(n520), .A2(n519), .ZN(n521) );
  XNOR2_X1 U586 ( .A(n521), .B(KEYINPUT48), .ZN(n550) );
  NOR2_X1 U587 ( .A1(n522), .A2(n550), .ZN(n540) );
  NAND2_X1 U588 ( .A1(n540), .A2(n523), .ZN(n524) );
  XOR2_X1 U589 ( .A(KEYINPUT116), .B(n524), .Z(n526) );
  NAND2_X1 U590 ( .A1(n526), .A2(n525), .ZN(n527) );
  XNOR2_X1 U591 ( .A(n527), .B(KEYINPUT117), .ZN(n537) );
  NAND2_X1 U592 ( .A1(n537), .A2(n517), .ZN(n529) );
  XNOR2_X1 U593 ( .A(n529), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT119), .B(KEYINPUT49), .Z(n531) );
  NAND2_X1 U595 ( .A1(n537), .A2(n562), .ZN(n530) );
  XNOR2_X1 U596 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U597 ( .A(G120GAT), .B(KEYINPUT118), .Z(n532) );
  XNOR2_X1 U598 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n585), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(G134GAT), .B(KEYINPUT51), .Z(n539) );
  INV_X1 U603 ( .A(n536), .ZN(n569) );
  NAND2_X1 U604 ( .A1(n537), .A2(n569), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n576), .A2(n540), .ZN(n541) );
  XOR2_X1 U607 ( .A(KEYINPUT120), .B(n541), .Z(n548) );
  NAND2_X1 U608 ( .A1(n517), .A2(n548), .ZN(n542) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n542), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n545) );
  NAND2_X1 U611 ( .A1(n548), .A2(n543), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U613 ( .A(G148GAT), .B(n546), .ZN(G1345GAT) );
  NAND2_X1 U614 ( .A1(n548), .A2(n585), .ZN(n547) );
  XNOR2_X1 U615 ( .A(n547), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U616 ( .A1(n548), .A2(n569), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U618 ( .A1(n551), .A2(n550), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT54), .ZN(n554) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(n555), .B(KEYINPUT65), .ZN(n577) );
  NAND2_X1 U622 ( .A1(n556), .A2(n577), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(KEYINPUT55), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(KEYINPUT121), .ZN(n559) );
  NAND2_X1 U625 ( .A1(n570), .A2(n517), .ZN(n561) );
  XNOR2_X1 U626 ( .A(n561), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n570), .ZN(n567) );
  XOR2_X1 U628 ( .A(KEYINPUT57), .B(KEYINPUT123), .Z(n564) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XOR2_X1 U631 ( .A(KEYINPUT56), .B(n565), .Z(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(G1349GAT) );
  NAND2_X1 U633 ( .A1(n570), .A2(n585), .ZN(n568) );
  XNOR2_X1 U634 ( .A(n568), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U635 ( .A1(n570), .A2(n569), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1351GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT124), .B(KEYINPUT125), .Z(n574) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT60), .B(n575), .Z(n579) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n588) );
  INV_X1 U643 ( .A(n588), .ZN(n586) );
  NAND2_X1 U644 ( .A1(n586), .A2(n517), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U646 ( .A1(n588), .A2(n580), .ZN(n584) );
  XOR2_X1 U647 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n582) );
  XNOR2_X1 U648 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n581) );
  XNOR2_X1 U649 ( .A(n582), .B(n581), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(G1353GAT) );
  NAND2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n587), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U653 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U654 ( .A(KEYINPUT62), .B(n590), .Z(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

