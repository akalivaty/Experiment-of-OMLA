//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 0 1 1 1 0 1 0 0 1 1 0 1 1 0 0 0 1 1 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:04 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n445, new_n447, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n548, new_n549, new_n550,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n570, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162, new_n1163;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT64), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  NAND2_X1  g019(.A1(G94), .A2(G452), .ZN(new_n445));
  XNOR2_X1  g020(.A(new_n445), .B(KEYINPUT66), .ZN(G173));
  XNOR2_X1  g021(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n447));
  AND2_X1   g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n447), .B(new_n448), .ZN(G223));
  NAND2_X1  g024(.A1(new_n448), .A2(G567), .ZN(G234));
  NAND2_X1  g025(.A1(new_n448), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NAND4_X1  g028(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n453), .A2(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(G325), .B(KEYINPUT68), .Z(G261));
  NAND2_X1  g031(.A1(new_n453), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  XNOR2_X1  g033(.A(new_n458), .B(KEYINPUT69), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n457), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G113), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  OR3_X1    g038(.A1(new_n462), .A2(new_n463), .A3(KEYINPUT70), .ZN(new_n464));
  OAI21_X1  g039(.A(KEYINPUT70), .B1(new_n462), .B2(new_n463), .ZN(new_n465));
  INV_X1    g040(.A(G125), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  OAI211_X1 g044(.A(new_n464), .B(new_n465), .C1(new_n466), .C2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n469), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n463), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n471), .A2(new_n474), .ZN(G160));
  INV_X1    g050(.A(G2105), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n469), .A2(new_n476), .ZN(new_n477));
  MUX2_X1   g052(.A(G100), .B(G112), .S(G2105), .Z(new_n478));
  AOI22_X1  g053(.A1(new_n477), .A2(G124), .B1(G2104), .B2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(G136), .ZN(new_n480));
  INV_X1    g055(.A(new_n472), .ZN(new_n481));
  OAI21_X1  g056(.A(new_n479), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  XNOR2_X1  g057(.A(new_n482), .B(KEYINPUT71), .ZN(G162));
  NAND2_X1  g058(.A1(new_n472), .A2(G138), .ZN(new_n484));
  INV_X1    g059(.A(KEYINPUT4), .ZN(new_n485));
  NAND2_X1  g060(.A1(G102), .A2(G2104), .ZN(new_n486));
  NAND2_X1  g061(.A1(KEYINPUT4), .A2(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(new_n486), .B1(new_n469), .B2(new_n487), .ZN(new_n488));
  AOI22_X1  g063(.A1(new_n484), .A2(new_n485), .B1(new_n476), .B2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(G114), .A2(G2104), .ZN(new_n490));
  INV_X1    g065(.A(G126), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n469), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n492), .A2(G2105), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n489), .A2(new_n493), .ZN(new_n494));
  INV_X1    g069(.A(new_n494), .ZN(G164));
  INV_X1    g070(.A(KEYINPUT5), .ZN(new_n496));
  INV_X1    g071(.A(G543), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  INV_X1    g078(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(new_n502), .ZN(new_n505));
  NAND2_X1  g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  AOI21_X1  g081(.A(new_n497), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G50), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n500), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  OAI21_X1  g086(.A(new_n508), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NOR2_X1   g087(.A1(new_n503), .A2(new_n512), .ZN(G166));
  NAND2_X1  g088(.A1(new_n507), .A2(G51), .ZN(new_n514));
  NAND3_X1  g089(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n515));
  XNOR2_X1  g090(.A(new_n515), .B(KEYINPUT7), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  AND2_X1   g092(.A1(KEYINPUT5), .A2(G543), .ZN(new_n518));
  NOR2_X1   g093(.A1(KEYINPUT5), .A2(G543), .ZN(new_n519));
  NOR2_X1   g094(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n509), .A2(G89), .ZN(new_n521));
  NAND2_X1  g096(.A1(G63), .A2(G651), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NOR2_X1   g098(.A1(new_n517), .A2(new_n523), .ZN(G168));
  AOI22_X1  g099(.A1(new_n500), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n525), .A2(new_n502), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n507), .A2(G52), .ZN(new_n527));
  INV_X1    g102(.A(G90), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n510), .B2(new_n528), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n526), .A2(new_n529), .ZN(G171));
  INV_X1    g105(.A(G56), .ZN(new_n531));
  AOI21_X1  g106(.A(new_n531), .B1(new_n498), .B2(new_n499), .ZN(new_n532));
  NAND2_X1  g107(.A1(G68), .A2(G543), .ZN(new_n533));
  INV_X1    g108(.A(new_n533), .ZN(new_n534));
  OAI21_X1  g109(.A(KEYINPUT72), .B1(new_n532), .B2(new_n534), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n536));
  OAI211_X1 g111(.A(new_n536), .B(new_n533), .C1(new_n520), .C2(new_n531), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n535), .A2(G651), .A3(new_n537), .ZN(new_n538));
  INV_X1    g113(.A(KEYINPUT73), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n498), .A2(new_n499), .B1(new_n505), .B2(new_n506), .ZN(new_n540));
  AOI22_X1  g115(.A1(new_n540), .A2(G81), .B1(new_n507), .B2(G43), .ZN(new_n541));
  AND3_X1   g116(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g117(.A(new_n539), .B1(new_n538), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g118(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  XOR2_X1   g122(.A(KEYINPUT74), .B(KEYINPUT8), .Z(new_n548));
  NAND2_X1  g123(.A1(G1), .A2(G3), .ZN(new_n549));
  XNOR2_X1  g124(.A(new_n548), .B(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n546), .A2(new_n550), .ZN(G188));
  NAND2_X1  g126(.A1(new_n507), .A2(G53), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT9), .ZN(new_n553));
  INV_X1    g128(.A(G65), .ZN(new_n554));
  INV_X1    g129(.A(G78), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n520), .A2(new_n554), .B1(new_n555), .B2(new_n497), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT76), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  OAI221_X1 g133(.A(KEYINPUT76), .B1(new_n555), .B2(new_n497), .C1(new_n520), .C2(new_n554), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n558), .A2(G651), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n510), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n540), .A2(KEYINPUT75), .ZN(new_n563));
  NAND3_X1  g138(.A1(new_n562), .A2(new_n563), .A3(G91), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n553), .A2(new_n560), .A3(new_n564), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n565), .B(KEYINPUT77), .ZN(G299));
  INV_X1    g141(.A(G171), .ZN(G301));
  INV_X1    g142(.A(G168), .ZN(G286));
  INV_X1    g143(.A(G166), .ZN(G303));
  AND2_X1   g144(.A1(new_n562), .A2(new_n563), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G87), .ZN(new_n571));
  OR2_X1    g146(.A1(new_n500), .A2(G74), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n572), .A2(G651), .B1(new_n507), .B2(G49), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n571), .A2(new_n573), .ZN(G288));
  AOI22_X1  g149(.A1(new_n500), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n575), .A2(new_n502), .ZN(new_n576));
  XNOR2_X1  g151(.A(new_n576), .B(KEYINPUT78), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n507), .A2(G48), .ZN(new_n578));
  INV_X1    g153(.A(new_n578), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n579), .B1(new_n570), .B2(G86), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n577), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n502), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n507), .A2(G47), .ZN(new_n584));
  INV_X1    g159(.A(G85), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n510), .B2(new_n585), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  INV_X1    g162(.A(new_n587), .ZN(G290));
  NAND2_X1  g163(.A1(G301), .A2(G868), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n562), .A2(new_n563), .A3(G92), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT10), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(G79), .A2(G543), .ZN(new_n593));
  INV_X1    g168(.A(G66), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n520), .B2(new_n594), .ZN(new_n595));
  AOI22_X1  g170(.A1(new_n595), .A2(G651), .B1(G54), .B2(new_n507), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT79), .ZN(new_n598));
  XNOR2_X1  g173(.A(new_n597), .B(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n589), .B1(new_n599), .B2(G868), .ZN(G321));
  NAND2_X1  g176(.A1(G286), .A2(G868), .ZN(new_n602));
  INV_X1    g177(.A(KEYINPUT77), .ZN(new_n603));
  XNOR2_X1  g178(.A(new_n565), .B(new_n603), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n602), .B1(new_n604), .B2(G868), .ZN(G297));
  OAI21_X1  g180(.A(new_n602), .B1(new_n604), .B2(G868), .ZN(G280));
  AND2_X1   g181(.A1(new_n592), .A2(new_n596), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(new_n598), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n597), .A2(KEYINPUT79), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  INV_X1    g185(.A(G860), .ZN(new_n611));
  AOI21_X1  g186(.A(new_n610), .B1(G559), .B2(new_n611), .ZN(new_n612));
  XNOR2_X1  g187(.A(new_n612), .B(KEYINPUT80), .ZN(G148));
  INV_X1    g188(.A(G868), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  INV_X1    g190(.A(G559), .ZN(new_n616));
  NAND3_X1  g191(.A1(new_n599), .A2(new_n615), .A3(new_n616), .ZN(new_n617));
  NAND3_X1  g192(.A1(new_n608), .A2(new_n616), .A3(new_n609), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n614), .B1(new_n617), .B2(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n620), .A2(KEYINPUT82), .ZN(new_n621));
  INV_X1    g196(.A(KEYINPUT82), .ZN(new_n622));
  INV_X1    g197(.A(new_n544), .ZN(new_n623));
  AOI21_X1  g198(.A(new_n622), .B1(new_n623), .B2(new_n614), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n621), .B1(new_n620), .B2(new_n624), .ZN(new_n625));
  INV_X1    g200(.A(KEYINPUT83), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n625), .B(new_n626), .ZN(G323));
  XNOR2_X1  g202(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g203(.A1(new_n472), .A2(G2104), .ZN(new_n629));
  XNOR2_X1  g204(.A(new_n629), .B(KEYINPUT12), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT13), .ZN(new_n631));
  INV_X1    g206(.A(G2100), .ZN(new_n632));
  OR2_X1    g207(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g208(.A1(new_n631), .A2(new_n632), .ZN(new_n634));
  NAND2_X1  g209(.A1(new_n472), .A2(G135), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n477), .A2(G123), .ZN(new_n636));
  OR3_X1    g211(.A1(new_n476), .A2(KEYINPUT84), .A3(G111), .ZN(new_n637));
  OAI21_X1  g212(.A(KEYINPUT84), .B1(new_n476), .B2(G111), .ZN(new_n638));
  OR2_X1    g213(.A1(G99), .A2(G2105), .ZN(new_n639));
  NAND4_X1  g214(.A1(new_n637), .A2(G2104), .A3(new_n638), .A4(new_n639), .ZN(new_n640));
  AND3_X1   g215(.A1(new_n635), .A2(new_n636), .A3(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(G2096), .ZN(new_n642));
  NAND3_X1  g217(.A1(new_n633), .A2(new_n634), .A3(new_n642), .ZN(G156));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(G2438), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(G2427), .ZN(new_n646));
  INV_X1    g221(.A(G2430), .ZN(new_n647));
  OR2_X1    g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n646), .A2(new_n647), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(KEYINPUT14), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2443), .B(G2446), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n650), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(G1341), .B(G1348), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g232(.A1(new_n657), .A2(G14), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n655), .A2(new_n656), .ZN(new_n659));
  OR2_X1    g234(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(KEYINPUT85), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n658), .B1(new_n660), .B2(new_n661), .ZN(G401));
  XOR2_X1   g237(.A(G2084), .B(G2090), .Z(new_n663));
  XNOR2_X1  g238(.A(G2072), .B(G2078), .ZN(new_n664));
  XNOR2_X1  g239(.A(G2067), .B(G2678), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g241(.A(new_n666), .B(KEYINPUT18), .Z(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NAND2_X1  g243(.A1(new_n664), .A2(KEYINPUT17), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g245(.A1(new_n670), .A2(new_n665), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n671), .B1(new_n668), .B2(new_n669), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n663), .A2(new_n665), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n664), .B1(new_n673), .B2(KEYINPUT17), .ZN(new_n674));
  OAI21_X1  g249(.A(new_n667), .B1(new_n672), .B2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT86), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT87), .Z(new_n677));
  XNOR2_X1  g252(.A(G2096), .B(G2100), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n679), .ZN(G227));
  XNOR2_X1  g255(.A(G1971), .B(G1976), .ZN(new_n681));
  XNOR2_X1  g256(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  XOR2_X1   g258(.A(G1956), .B(G2474), .Z(new_n684));
  XOR2_X1   g259(.A(G1961), .B(G1966), .Z(new_n685));
  NAND2_X1  g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(KEYINPUT89), .B(KEYINPUT20), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  OR2_X1    g264(.A1(new_n684), .A2(new_n685), .ZN(new_n690));
  NAND3_X1  g265(.A1(new_n683), .A2(new_n686), .A3(new_n690), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n689), .B(new_n691), .C1(new_n683), .C2(new_n690), .ZN(new_n692));
  XOR2_X1   g267(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  XOR2_X1   g269(.A(G1991), .B(G1996), .Z(new_n695));
  XNOR2_X1  g270(.A(G1981), .B(G1986), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n694), .B(new_n697), .ZN(G229));
  NOR2_X1   g273(.A1(G16), .A2(G23), .ZN(new_n699));
  XNOR2_X1  g274(.A(G288), .B(KEYINPUT93), .ZN(new_n700));
  AOI21_X1  g275(.A(new_n699), .B1(new_n700), .B2(G16), .ZN(new_n701));
  XNOR2_X1  g276(.A(KEYINPUT33), .B(G1976), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT94), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n701), .A2(new_n703), .ZN(new_n704));
  NOR2_X1   g279(.A1(new_n701), .A2(new_n703), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  OR2_X1    g281(.A1(G6), .A2(G16), .ZN(new_n707));
  INV_X1    g282(.A(G16), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n707), .B1(G305), .B2(new_n708), .ZN(new_n709));
  XOR2_X1   g284(.A(KEYINPUT32), .B(G1981), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  NOR2_X1   g286(.A1(G16), .A2(G22), .ZN(new_n712));
  AOI21_X1  g287(.A(new_n712), .B1(G166), .B2(G16), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1971), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  OAI21_X1  g291(.A(KEYINPUT34), .B1(new_n706), .B2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(KEYINPUT34), .ZN(new_n718));
  OAI211_X1 g293(.A(new_n715), .B(new_n718), .C1(new_n705), .C2(new_n704), .ZN(new_n719));
  INV_X1    g294(.A(G29), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n720), .A2(G25), .ZN(new_n721));
  MUX2_X1   g296(.A(G95), .B(G107), .S(G2105), .Z(new_n722));
  AOI22_X1  g297(.A1(new_n477), .A2(G119), .B1(G2104), .B2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(G131), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n723), .B1(new_n724), .B2(new_n481), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n725), .B(KEYINPUT90), .ZN(new_n726));
  INV_X1    g301(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n721), .B1(new_n727), .B2(new_n720), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT91), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n728), .B(new_n730), .Z(new_n731));
  INV_X1    g306(.A(G24), .ZN(new_n732));
  OAI21_X1  g307(.A(KEYINPUT92), .B1(new_n732), .B2(G16), .ZN(new_n733));
  OR3_X1    g308(.A1(new_n732), .A2(KEYINPUT92), .A3(G16), .ZN(new_n734));
  OAI211_X1 g309(.A(new_n733), .B(new_n734), .C1(new_n587), .C2(new_n708), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n735), .B(G1986), .ZN(new_n736));
  NOR2_X1   g311(.A1(new_n731), .A2(new_n736), .ZN(new_n737));
  NAND3_X1  g312(.A1(new_n717), .A2(new_n719), .A3(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(KEYINPUT95), .B(KEYINPUT36), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g315(.A(KEYINPUT102), .B(KEYINPUT23), .Z(new_n741));
  NAND2_X1  g316(.A1(new_n708), .A2(G20), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n743), .B1(new_n604), .B2(new_n708), .ZN(new_n744));
  XNOR2_X1  g319(.A(new_n744), .B(KEYINPUT103), .ZN(new_n745));
  INV_X1    g320(.A(G1956), .ZN(new_n746));
  OR2_X1    g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n745), .A2(new_n746), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n708), .A2(G4), .ZN(new_n749));
  AOI21_X1  g324(.A(new_n749), .B1(new_n610), .B2(G16), .ZN(new_n750));
  AND2_X1   g325(.A1(new_n750), .A2(G1348), .ZN(new_n751));
  NOR2_X1   g326(.A1(new_n750), .A2(G1348), .ZN(new_n752));
  OAI211_X1 g327(.A(new_n747), .B(new_n748), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n641), .A2(G29), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT99), .Z(new_n756));
  XNOR2_X1  g331(.A(KEYINPUT31), .B(G11), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT30), .B(G28), .Z(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n758), .B2(G29), .ZN(new_n759));
  NOR2_X1   g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G168), .A2(new_n708), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(new_n708), .B2(G21), .ZN(new_n762));
  INV_X1    g337(.A(G1966), .ZN(new_n763));
  NAND2_X1  g338(.A1(new_n708), .A2(G5), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G171), .B2(new_n708), .ZN(new_n765));
  AOI22_X1  g340(.A1(new_n762), .A2(new_n763), .B1(G1961), .B2(new_n765), .ZN(new_n766));
  OR2_X1    g341(.A1(new_n762), .A2(new_n763), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n760), .A2(new_n766), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n720), .A2(G32), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n477), .A2(G129), .ZN(new_n772));
  XOR2_X1   g347(.A(new_n772), .B(KEYINPUT97), .Z(new_n773));
  AND2_X1   g348(.A1(new_n473), .A2(G105), .ZN(new_n774));
  NAND3_X1  g349(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT26), .ZN(new_n776));
  AOI211_X1 g351(.A(new_n774), .B(new_n776), .C1(G141), .C2(new_n472), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n771), .B1(new_n778), .B2(G29), .ZN(new_n779));
  XOR2_X1   g354(.A(KEYINPUT27), .B(G1996), .Z(new_n780));
  XNOR2_X1  g355(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  XNOR2_X1  g356(.A(new_n779), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n473), .A2(G103), .ZN(new_n783));
  INV_X1    g358(.A(KEYINPUT25), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n473), .A2(KEYINPUT25), .A3(G103), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n472), .A2(G139), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  INV_X1    g362(.A(new_n469), .ZN(new_n788));
  AOI22_X1  g363(.A1(new_n788), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n787), .B1(new_n476), .B2(new_n789), .ZN(new_n790));
  MUX2_X1   g365(.A(G33), .B(new_n790), .S(G29), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G2072), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g368(.A1(new_n760), .A2(new_n766), .A3(KEYINPUT100), .A4(new_n767), .ZN(new_n794));
  NOR2_X1   g369(.A1(G27), .A2(G29), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G164), .B2(G29), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G2078), .ZN(new_n797));
  AND2_X1   g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NOR2_X1   g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n720), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n471), .A2(new_n474), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n800), .B1(new_n801), .B2(new_n720), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n802), .B(G2084), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G1961), .B2(new_n765), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n797), .A2(new_n804), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n770), .A2(new_n793), .A3(new_n794), .A4(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n806), .A2(KEYINPUT101), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n782), .A2(new_n797), .A3(new_n804), .A4(new_n792), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT101), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n808), .A2(new_n809), .A3(new_n770), .A4(new_n794), .ZN(new_n810));
  INV_X1    g385(.A(G2090), .ZN(new_n811));
  NOR2_X1   g386(.A1(G29), .A2(G35), .ZN(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G162), .B2(G29), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n813), .A2(KEYINPUT29), .ZN(new_n814));
  INV_X1    g389(.A(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(G162), .A2(G29), .ZN(new_n816));
  INV_X1    g391(.A(new_n812), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(KEYINPUT29), .A3(new_n817), .ZN(new_n818));
  AOI21_X1  g393(.A(new_n811), .B1(new_n815), .B2(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n818), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n820), .A2(new_n814), .A3(G2090), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n708), .A2(G19), .ZN(new_n822));
  OAI21_X1  g397(.A(new_n822), .B1(new_n544), .B2(new_n708), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n823), .B(G1341), .ZN(new_n824));
  MUX2_X1   g399(.A(G104), .B(G116), .S(G2105), .Z(new_n825));
  AOI22_X1  g400(.A1(new_n477), .A2(G128), .B1(G2104), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G140), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(new_n481), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n828), .A2(G29), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n720), .A2(G26), .ZN(new_n830));
  XNOR2_X1  g405(.A(new_n830), .B(KEYINPUT96), .ZN(new_n831));
  XNOR2_X1  g406(.A(new_n831), .B(KEYINPUT28), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n829), .A2(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(G2067), .ZN(new_n834));
  NOR4_X1   g409(.A1(new_n819), .A2(new_n821), .A3(new_n824), .A4(new_n834), .ZN(new_n835));
  AND3_X1   g410(.A1(new_n807), .A2(new_n810), .A3(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(new_n739), .ZN(new_n837));
  NAND4_X1  g412(.A1(new_n717), .A2(new_n719), .A3(new_n737), .A4(new_n837), .ZN(new_n838));
  NAND4_X1  g413(.A1(new_n740), .A2(new_n754), .A3(new_n836), .A4(new_n838), .ZN(G150));
  XNOR2_X1  g414(.A(G150), .B(KEYINPUT104), .ZN(G311));
  AOI22_X1  g415(.A1(new_n500), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n841), .A2(new_n502), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n507), .A2(G55), .ZN(new_n843));
  INV_X1    g418(.A(G93), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n510), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n842), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n611), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(KEYINPUT37), .ZN(new_n848));
  INV_X1    g423(.A(KEYINPUT105), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n538), .A2(new_n541), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n850), .A2(KEYINPUT73), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n538), .A2(new_n539), .A3(new_n541), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n846), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n846), .A2(new_n538), .A3(new_n541), .ZN(new_n854));
  INV_X1    g429(.A(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n849), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n846), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n857), .B1(new_n542), .B2(new_n543), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n858), .A2(KEYINPUT105), .A3(new_n854), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(KEYINPUT38), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n599), .A2(G559), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  OR2_X1    g438(.A1(new_n863), .A2(KEYINPUT39), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT106), .ZN(new_n865));
  AND2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  AOI21_X1  g441(.A(G860), .B1(new_n863), .B2(KEYINPUT39), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n867), .B1(new_n864), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n848), .B1(new_n866), .B2(new_n868), .ZN(G145));
  XNOR2_X1  g444(.A(G162), .B(new_n801), .ZN(new_n870));
  XNOR2_X1  g445(.A(new_n870), .B(new_n641), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT107), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n494), .A2(new_n872), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n489), .A2(KEYINPUT107), .A3(new_n493), .ZN(new_n874));
  AND2_X1   g449(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n875), .B(new_n828), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n630), .B(new_n725), .ZN(new_n877));
  MUX2_X1   g452(.A(G106), .B(G118), .S(G2105), .Z(new_n878));
  AOI22_X1  g453(.A1(new_n477), .A2(G130), .B1(G2104), .B2(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G142), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n879), .B1(new_n880), .B2(new_n481), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n877), .B(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n876), .B(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n778), .B(new_n790), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  NOR2_X1   g461(.A1(new_n883), .A2(new_n884), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n871), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n887), .ZN(new_n889));
  INV_X1    g464(.A(new_n871), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(new_n890), .A3(new_n885), .ZN(new_n891));
  INV_X1    g466(.A(G37), .ZN(new_n892));
  NAND3_X1  g467(.A1(new_n888), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n893), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g469(.A1(new_n857), .A2(G868), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n700), .B(new_n587), .ZN(new_n896));
  XNOR2_X1  g471(.A(G305), .B(G166), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n896), .A2(new_n898), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n700), .B(G290), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n900), .A2(new_n897), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(new_n615), .B1(new_n599), .B2(new_n616), .ZN(new_n903));
  NOR2_X1   g478(.A1(new_n618), .A2(KEYINPUT81), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n860), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n604), .A2(new_n607), .ZN(new_n906));
  NAND2_X1  g481(.A1(G299), .A2(new_n597), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(new_n908), .ZN(new_n909));
  NAND4_X1  g484(.A1(new_n617), .A2(new_n619), .A3(new_n859), .A4(new_n856), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n905), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n911), .ZN(new_n912));
  AND3_X1   g487(.A1(new_n906), .A2(new_n907), .A3(KEYINPUT41), .ZN(new_n913));
  AOI21_X1  g488(.A(KEYINPUT41), .B1(new_n906), .B2(new_n907), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  AOI21_X1  g491(.A(new_n916), .B1(new_n905), .B2(new_n910), .ZN(new_n917));
  NOR3_X1   g492(.A1(new_n912), .A2(new_n917), .A3(KEYINPUT42), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT42), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n905), .A2(new_n910), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n920), .A2(new_n915), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n919), .B1(new_n921), .B2(new_n911), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n902), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g498(.A(KEYINPUT42), .B1(new_n912), .B2(new_n917), .ZN(new_n924));
  INV_X1    g499(.A(new_n902), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n921), .A2(new_n911), .A3(new_n919), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n923), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n895), .B1(new_n928), .B2(G868), .ZN(G295));
  AOI21_X1  g504(.A(new_n895), .B1(new_n928), .B2(G868), .ZN(G331));
  INV_X1    g505(.A(KEYINPUT43), .ZN(new_n931));
  XNOR2_X1  g506(.A(G171), .B(G168), .ZN(new_n932));
  INV_X1    g507(.A(new_n932), .ZN(new_n933));
  AND3_X1   g508(.A1(new_n858), .A2(KEYINPUT105), .A3(new_n854), .ZN(new_n934));
  AOI21_X1  g509(.A(KEYINPUT105), .B1(new_n858), .B2(new_n854), .ZN(new_n935));
  OAI21_X1  g510(.A(new_n933), .B1(new_n934), .B2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT109), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n860), .A2(KEYINPUT109), .A3(new_n933), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n856), .A2(new_n859), .A3(new_n932), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(KEYINPUT108), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT108), .ZN(new_n942));
  NAND4_X1  g517(.A1(new_n856), .A2(new_n942), .A3(new_n859), .A4(new_n932), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n938), .A2(new_n939), .A3(new_n941), .A4(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT111), .B1(new_n944), .B2(new_n908), .ZN(new_n945));
  AND2_X1   g520(.A1(new_n941), .A2(new_n943), .ZN(new_n946));
  AOI21_X1  g521(.A(KEYINPUT109), .B1(new_n860), .B2(new_n933), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n937), .B(new_n932), .C1(new_n856), .C2(new_n859), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT111), .ZN(new_n950));
  NAND4_X1  g525(.A1(new_n946), .A2(new_n949), .A3(new_n950), .A4(new_n909), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n860), .A2(KEYINPUT110), .A3(new_n933), .ZN(new_n952));
  INV_X1    g527(.A(KEYINPUT110), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n936), .A2(new_n953), .A3(new_n940), .ZN(new_n954));
  NAND3_X1  g529(.A1(new_n915), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  NAND3_X1  g530(.A1(new_n945), .A2(new_n951), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(new_n925), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n954), .A2(new_n952), .ZN(new_n958));
  AOI22_X1  g533(.A1(new_n915), .A2(new_n944), .B1(new_n958), .B2(new_n909), .ZN(new_n959));
  AOI21_X1  g534(.A(G37), .B1(new_n959), .B2(new_n902), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n931), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n944), .A2(new_n915), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n958), .A2(new_n909), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n962), .A2(new_n902), .A3(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n964), .A2(new_n892), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n902), .B1(new_n962), .B2(new_n963), .ZN(new_n966));
  NOR3_X1   g541(.A1(new_n965), .A2(KEYINPUT43), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(KEYINPUT44), .B1(new_n961), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT44), .ZN(new_n969));
  AOI21_X1  g544(.A(KEYINPUT43), .B1(new_n957), .B2(new_n960), .ZN(new_n970));
  NOR3_X1   g545(.A1(new_n965), .A2(new_n931), .A3(new_n966), .ZN(new_n971));
  OAI21_X1  g546(.A(new_n969), .B1(new_n970), .B2(new_n971), .ZN(new_n972));
  AND2_X1   g547(.A1(new_n968), .A2(new_n972), .ZN(G397));
  INV_X1    g548(.A(G1384), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n875), .A2(new_n974), .ZN(new_n975));
  INV_X1    g550(.A(KEYINPUT45), .ZN(new_n976));
  AND3_X1   g551(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n977));
  NAND3_X1  g552(.A1(new_n975), .A2(new_n976), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(new_n978), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n828), .B(G2067), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT112), .ZN(new_n982));
  XOR2_X1   g557(.A(new_n778), .B(G1996), .Z(new_n983));
  OAI22_X1  g558(.A1(new_n981), .A2(new_n982), .B1(new_n978), .B2(new_n983), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n981), .A2(new_n982), .ZN(new_n986));
  XOR2_X1   g561(.A(new_n725), .B(new_n730), .Z(new_n987));
  NAND2_X1  g562(.A1(new_n979), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n985), .A2(new_n986), .A3(new_n988), .ZN(new_n989));
  XOR2_X1   g564(.A(new_n587), .B(G1986), .Z(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n979), .B2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n489), .B2(new_n493), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(new_n977), .ZN(new_n993));
  AND3_X1   g568(.A1(new_n993), .A2(KEYINPUT115), .A3(G8), .ZN(new_n994));
  AOI21_X1  g569(.A(KEYINPUT115), .B1(new_n993), .B2(G8), .ZN(new_n995));
  NOR2_X1   g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1981), .ZN(new_n997));
  AOI21_X1  g572(.A(new_n579), .B1(G86), .B2(new_n540), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n997), .B1(new_n577), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n1000), .B(KEYINPUT49), .C1(G1981), .C2(G305), .ZN(new_n1001));
  INV_X1    g576(.A(KEYINPUT49), .ZN(new_n1002));
  NOR2_X1   g577(.A1(G305), .A2(G1981), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1002), .B1(new_n1003), .B2(new_n999), .ZN(new_n1004));
  OAI211_X1 g579(.A(new_n1001), .B(new_n1004), .C1(new_n994), .C2(new_n995), .ZN(new_n1005));
  INV_X1    g580(.A(G1976), .ZN(new_n1006));
  INV_X1    g581(.A(G288), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  XOR2_X1   g583(.A(new_n1003), .B(KEYINPUT116), .Z(new_n1009));
  AOI21_X1  g584(.A(new_n996), .B1(new_n1008), .B2(new_n1009), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT114), .ZN(new_n1011));
  OAI211_X1 g586(.A(G303), .B(G8), .C1(new_n1011), .C2(KEYINPUT55), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(KEYINPUT55), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1012), .B(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n977), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n494), .A2(new_n974), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT50), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1019));
  AOI21_X1  g594(.A(new_n1015), .B1(new_n1018), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1020), .A2(new_n811), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n977), .B1(new_n992), .B2(KEYINPUT45), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND4_X1  g598(.A1(new_n873), .A2(KEYINPUT45), .A3(new_n974), .A4(new_n874), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1971), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  OAI21_X1  g600(.A(new_n1021), .B1(new_n1025), .B2(KEYINPUT113), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1025), .A2(KEYINPUT113), .ZN(new_n1027));
  OAI211_X1 g602(.A(G8), .B(new_n1014), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1028), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1007), .A2(KEYINPUT93), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT93), .ZN(new_n1031));
  NAND2_X1  g606(.A1(G288), .A2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1030), .A2(G1976), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1033), .B1(new_n994), .B2(new_n995), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT52), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT52), .B1(G288), .B2(new_n1006), .ZN(new_n1036));
  OAI211_X1 g611(.A(new_n1033), .B(new_n1036), .C1(new_n994), .C2(new_n995), .ZN(new_n1037));
  AND3_X1   g612(.A1(new_n1035), .A2(new_n1005), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(new_n1010), .B1(new_n1029), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1019), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n992), .A2(KEYINPUT50), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n977), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  XNOR2_X1  g617(.A(KEYINPUT117), .B(G1956), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  XNOR2_X1  g619(.A(KEYINPUT56), .B(G2072), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1023), .A2(new_n1024), .A3(new_n1045), .ZN(new_n1046));
  XOR2_X1   g621(.A(new_n565), .B(KEYINPUT57), .Z(new_n1047));
  AND3_X1   g622(.A1(new_n1044), .A2(new_n1046), .A3(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1047), .B1(new_n1044), .B2(new_n1046), .ZN(new_n1049));
  OAI22_X1  g624(.A1(new_n1020), .A2(G1348), .B1(G2067), .B2(new_n993), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n607), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1049), .B1(KEYINPUT118), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1051), .A2(KEYINPUT118), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1048), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  NAND2_X1  g629(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1055));
  INV_X1    g630(.A(new_n993), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT58), .B(G1341), .ZN(new_n1057));
  OAI22_X1  g632(.A1(new_n1055), .A2(G1996), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1058), .A2(new_n544), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1059), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1060), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1058), .A2(new_n544), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1061), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n993), .A2(G2067), .ZN(new_n1065));
  INV_X1    g640(.A(G1348), .ZN(new_n1066));
  AOI21_X1  g641(.A(new_n1065), .B1(new_n1042), .B2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1067), .A2(KEYINPUT60), .A3(new_n597), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n1069));
  NAND2_X1  g644(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n1067), .A2(KEYINPUT121), .A3(KEYINPUT60), .A4(new_n597), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT60), .ZN(new_n1072));
  OAI21_X1  g647(.A(new_n607), .B1(new_n1050), .B2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1070), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1050), .A2(new_n1072), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1064), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT120), .B1(new_n1048), .B2(new_n1049), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT61), .ZN(new_n1078));
  NAND2_X1  g653(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g654(.A(KEYINPUT120), .B(KEYINPUT61), .C1(new_n1048), .C2(new_n1049), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1079), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1054), .B1(new_n1076), .B2(new_n1081), .ZN(new_n1082));
  XOR2_X1   g657(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1083));
  INV_X1    g658(.A(G8), .ZN(new_n1084));
  INV_X1    g659(.A(G2084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1085), .B(new_n977), .C1(new_n1040), .C2(new_n1041), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1016), .A2(new_n976), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n763), .B1(new_n1087), .B2(new_n1022), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n1084), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  NOR2_X1   g664(.A1(G168), .A2(new_n1084), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1083), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT123), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1093));
  OR3_X1    g668(.A1(new_n1089), .A2(KEYINPUT51), .A3(new_n1090), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT123), .B(new_n1083), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1089), .A2(G286), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1021), .ZN(new_n1099));
  OAI21_X1  g674(.A(G8), .B1(new_n1099), .B2(new_n1025), .ZN(new_n1100));
  INV_X1    g675(.A(new_n1014), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1038), .A2(new_n1102), .A3(new_n1028), .ZN(new_n1103));
  XNOR2_X1  g678(.A(G171), .B(KEYINPUT54), .ZN(new_n1104));
  INV_X1    g679(.A(G1961), .ZN(new_n1105));
  NOR2_X1   g680(.A1(new_n1087), .A2(new_n1022), .ZN(new_n1106));
  INV_X1    g681(.A(KEYINPUT53), .ZN(new_n1107));
  NOR2_X1   g682(.A1(new_n1107), .A2(G2078), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1042), .A2(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  OAI21_X1  g684(.A(new_n1107), .B1(new_n1055), .B2(G2078), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1104), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n975), .A2(new_n976), .ZN(new_n1112));
  NAND4_X1  g687(.A1(new_n1112), .A2(new_n977), .A3(new_n1024), .A4(new_n1108), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1042), .A2(new_n1105), .ZN(new_n1114));
  AND3_X1   g689(.A1(new_n1113), .A2(new_n1114), .A3(new_n1104), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1111), .B1(new_n1115), .B2(new_n1110), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1098), .A2(new_n1103), .A3(new_n1116), .ZN(new_n1117));
  OAI21_X1  g692(.A(new_n1039), .B1(new_n1082), .B2(new_n1117), .ZN(new_n1118));
  AND2_X1   g693(.A1(new_n1089), .A2(G168), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n1038), .A2(new_n1028), .A3(new_n1102), .A4(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT63), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  AND2_X1   g697(.A1(new_n1119), .A2(KEYINPUT63), .ZN(new_n1123));
  OAI21_X1  g698(.A(G8), .B1(new_n1026), .B2(new_n1027), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1124), .A2(new_n1101), .ZN(new_n1125));
  NAND4_X1  g700(.A1(new_n1123), .A2(new_n1125), .A3(new_n1028), .A4(new_n1038), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n1122), .A2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1096), .A2(new_n1128), .A3(new_n1097), .ZN(new_n1129));
  AOI21_X1  g704(.A(G301), .B1(new_n1109), .B2(new_n1110), .ZN(new_n1130));
  AND4_X1   g705(.A1(new_n1102), .A2(new_n1038), .A3(new_n1028), .A4(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1129), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1128), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1133));
  OAI21_X1  g708(.A(new_n1127), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(new_n991), .B1(new_n1118), .B2(new_n1134), .ZN(new_n1135));
  NOR2_X1   g710(.A1(new_n978), .A2(G1996), .ZN(new_n1136));
  XOR2_X1   g711(.A(new_n1136), .B(KEYINPUT46), .Z(new_n1137));
  OAI21_X1  g712(.A(new_n979), .B1(new_n778), .B2(new_n980), .ZN(new_n1138));
  OR2_X1    g713(.A1(new_n1138), .A2(KEYINPUT125), .ZN(new_n1139));
  NAND2_X1  g714(.A1(new_n1138), .A2(KEYINPUT125), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1137), .A2(new_n1139), .A3(new_n1140), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(KEYINPUT47), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT47), .ZN(new_n1143));
  NAND4_X1  g718(.A1(new_n1137), .A2(new_n1139), .A3(new_n1143), .A4(new_n1140), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT126), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n989), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n985), .A2(KEYINPUT126), .A3(new_n986), .A4(new_n988), .ZN(new_n1148));
  NOR3_X1   g723(.A1(new_n978), .A2(G1986), .A3(G290), .ZN(new_n1149));
  XNOR2_X1  g724(.A(KEYINPUT127), .B(KEYINPUT48), .ZN(new_n1150));
  XNOR2_X1  g725(.A(new_n1149), .B(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1147), .A2(new_n1148), .A3(new_n1151), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n727), .A2(new_n730), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT124), .ZN(new_n1154));
  AND3_X1   g729(.A1(new_n985), .A2(new_n986), .A3(new_n1154), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n828), .A2(G2067), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n979), .B1(new_n1155), .B2(new_n1156), .ZN(new_n1157));
  AND3_X1   g732(.A1(new_n1145), .A2(new_n1152), .A3(new_n1157), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1135), .A2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g734(.A1(G229), .A2(new_n460), .ZN(new_n1161));
  NOR3_X1   g735(.A1(G401), .A2(G227), .A3(new_n1161), .ZN(new_n1162));
  NAND2_X1  g736(.A1(new_n893), .A2(new_n1162), .ZN(new_n1163));
  NOR3_X1   g737(.A1(new_n1163), .A2(new_n970), .A3(new_n971), .ZN(G308));
  OR3_X1    g738(.A1(new_n1163), .A2(new_n970), .A3(new_n971), .ZN(G225));
endmodule


