

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XOR2_X1 U321 ( .A(n298), .B(n297), .Z(n289) );
  XNOR2_X1 U322 ( .A(KEYINPUT54), .B(KEYINPUT125), .ZN(n290) );
  AND2_X1 U323 ( .A1(G232GAT), .A2(G233GAT), .ZN(n291) );
  INV_X1 U324 ( .A(KEYINPUT45), .ZN(n503) );
  XNOR2_X1 U325 ( .A(n504), .B(n503), .ZN(n506) );
  XNOR2_X1 U326 ( .A(n367), .B(n291), .ZN(n293) );
  XNOR2_X1 U327 ( .A(n543), .B(n290), .ZN(n563) );
  XNOR2_X1 U328 ( .A(n299), .B(n289), .ZN(n300) );
  XNOR2_X1 U329 ( .A(n301), .B(n300), .ZN(n303) );
  XOR2_X1 U330 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n444) );
  XOR2_X1 U331 ( .A(G134GAT), .B(KEYINPUT79), .Z(n367) );
  XNOR2_X1 U332 ( .A(G99GAT), .B(G85GAT), .ZN(n292) );
  XNOR2_X1 U333 ( .A(n292), .B(KEYINPUT75), .ZN(n413) );
  XNOR2_X1 U334 ( .A(n293), .B(n413), .ZN(n294) );
  XOR2_X1 U335 ( .A(n294), .B(KEYINPUT9), .Z(n301) );
  XOR2_X1 U336 ( .A(G29GAT), .B(G43GAT), .Z(n296) );
  XNOR2_X1 U337 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n295) );
  XNOR2_X1 U338 ( .A(n296), .B(n295), .ZN(n432) );
  XNOR2_X1 U339 ( .A(n432), .B(KEYINPUT11), .ZN(n299) );
  XOR2_X1 U340 ( .A(KEYINPUT10), .B(G92GAT), .Z(n298) );
  XNOR2_X1 U341 ( .A(G218GAT), .B(G106GAT), .ZN(n297) );
  XOR2_X1 U342 ( .A(G50GAT), .B(G162GAT), .Z(n386) );
  XOR2_X1 U343 ( .A(G36GAT), .B(G190GAT), .Z(n341) );
  XNOR2_X1 U344 ( .A(n386), .B(n341), .ZN(n302) );
  XNOR2_X1 U345 ( .A(n303), .B(n302), .ZN(n557) );
  XOR2_X1 U346 ( .A(KEYINPUT80), .B(G78GAT), .Z(n305) );
  XNOR2_X1 U347 ( .A(G183GAT), .B(G211GAT), .ZN(n304) );
  XNOR2_X1 U348 ( .A(n305), .B(n304), .ZN(n309) );
  XOR2_X1 U349 ( .A(KEYINPUT81), .B(KEYINPUT15), .Z(n307) );
  XNOR2_X1 U350 ( .A(G64GAT), .B(KEYINPUT14), .ZN(n306) );
  XNOR2_X1 U351 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U352 ( .A(n309), .B(n308), .ZN(n319) );
  XOR2_X1 U353 ( .A(G57GAT), .B(KEYINPUT71), .Z(n311) );
  XNOR2_X1 U354 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n310) );
  XNOR2_X1 U355 ( .A(n311), .B(n310), .ZN(n419) );
  XOR2_X1 U356 ( .A(n419), .B(KEYINPUT12), .Z(n313) );
  NAND2_X1 U357 ( .A1(G231GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U358 ( .A(n313), .B(n312), .ZN(n314) );
  XOR2_X1 U359 ( .A(G22GAT), .B(G155GAT), .Z(n385) );
  XOR2_X1 U360 ( .A(n314), .B(n385), .Z(n317) );
  XNOR2_X1 U361 ( .A(G1GAT), .B(KEYINPUT68), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n315), .B(G8GAT), .ZN(n431) );
  XOR2_X1 U363 ( .A(G15GAT), .B(G127GAT), .Z(n324) );
  XNOR2_X1 U364 ( .A(n431), .B(n324), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n317), .B(n316), .ZN(n318) );
  XOR2_X1 U366 ( .A(n319), .B(n318), .Z(n573) );
  NOR2_X1 U367 ( .A1(n557), .A2(n573), .ZN(n321) );
  XNOR2_X1 U368 ( .A(KEYINPUT16), .B(KEYINPUT82), .ZN(n320) );
  XNOR2_X1 U369 ( .A(n321), .B(n320), .ZN(n406) );
  XOR2_X1 U370 ( .A(G120GAT), .B(KEYINPUT83), .Z(n323) );
  XNOR2_X1 U371 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n322) );
  XNOR2_X1 U372 ( .A(n323), .B(n322), .ZN(n364) );
  XOR2_X1 U373 ( .A(n324), .B(n364), .Z(n326) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G134GAT), .ZN(n325) );
  XNOR2_X1 U375 ( .A(n326), .B(n325), .ZN(n330) );
  XOR2_X1 U376 ( .A(G176GAT), .B(G71GAT), .Z(n328) );
  NAND2_X1 U377 ( .A1(G227GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U378 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U379 ( .A(n330), .B(n329), .Z(n335) );
  XOR2_X1 U380 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n332) );
  XNOR2_X1 U381 ( .A(G190GAT), .B(G99GAT), .ZN(n331) );
  XNOR2_X1 U382 ( .A(n332), .B(n331), .ZN(n333) );
  XNOR2_X1 U383 ( .A(n333), .B(KEYINPUT86), .ZN(n334) );
  XNOR2_X1 U384 ( .A(n335), .B(n334), .ZN(n340) );
  XOR2_X1 U385 ( .A(KEYINPUT18), .B(G183GAT), .Z(n337) );
  XNOR2_X1 U386 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n336) );
  XNOR2_X1 U387 ( .A(n337), .B(n336), .ZN(n339) );
  XOR2_X1 U388 ( .A(KEYINPUT85), .B(KEYINPUT19), .Z(n338) );
  XOR2_X1 U389 ( .A(n339), .B(n338), .Z(n347) );
  XOR2_X1 U390 ( .A(n340), .B(n347), .Z(n547) );
  XOR2_X1 U391 ( .A(n341), .B(G8GAT), .Z(n343) );
  NAND2_X1 U392 ( .A1(G226GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U393 ( .A(n343), .B(n342), .ZN(n346) );
  XOR2_X1 U394 ( .A(KEYINPUT77), .B(G64GAT), .Z(n345) );
  XNOR2_X1 U395 ( .A(G176GAT), .B(G92GAT), .ZN(n344) );
  XNOR2_X1 U396 ( .A(n345), .B(n344), .ZN(n409) );
  XOR2_X1 U397 ( .A(n346), .B(n409), .Z(n354) );
  INV_X1 U398 ( .A(n347), .ZN(n352) );
  XNOR2_X1 U399 ( .A(G211GAT), .B(G218GAT), .ZN(n348) );
  XNOR2_X1 U400 ( .A(n348), .B(KEYINPUT21), .ZN(n349) );
  XOR2_X1 U401 ( .A(n349), .B(KEYINPUT88), .Z(n351) );
  XNOR2_X1 U402 ( .A(G197GAT), .B(G204GAT), .ZN(n350) );
  XNOR2_X1 U403 ( .A(n351), .B(n350), .ZN(n393) );
  XOR2_X1 U404 ( .A(n352), .B(n393), .Z(n353) );
  XNOR2_X1 U405 ( .A(n354), .B(n353), .ZN(n541) );
  XNOR2_X1 U406 ( .A(n541), .B(KEYINPUT94), .ZN(n355) );
  XNOR2_X1 U407 ( .A(n355), .B(KEYINPUT27), .ZN(n397) );
  XOR2_X1 U408 ( .A(KEYINPUT4), .B(KEYINPUT91), .Z(n357) );
  XNOR2_X1 U409 ( .A(KEYINPUT6), .B(KEYINPUT1), .ZN(n356) );
  XNOR2_X1 U410 ( .A(n357), .B(n356), .ZN(n377) );
  XOR2_X1 U411 ( .A(G85GAT), .B(G148GAT), .Z(n359) );
  XNOR2_X1 U412 ( .A(G127GAT), .B(G155GAT), .ZN(n358) );
  XNOR2_X1 U413 ( .A(n359), .B(n358), .ZN(n363) );
  XOR2_X1 U414 ( .A(KEYINPUT92), .B(KEYINPUT5), .Z(n361) );
  XNOR2_X1 U415 ( .A(G1GAT), .B(G57GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U417 ( .A(n363), .B(n362), .Z(n375) );
  XOR2_X1 U418 ( .A(n364), .B(KEYINPUT93), .Z(n366) );
  NAND2_X1 U419 ( .A1(G225GAT), .A2(G233GAT), .ZN(n365) );
  XNOR2_X1 U420 ( .A(n366), .B(n365), .ZN(n373) );
  XOR2_X1 U421 ( .A(n367), .B(G162GAT), .Z(n371) );
  XOR2_X1 U422 ( .A(KEYINPUT2), .B(KEYINPUT89), .Z(n369) );
  XNOR2_X1 U423 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n368) );
  XNOR2_X1 U424 ( .A(n369), .B(n368), .ZN(n380) );
  XNOR2_X1 U425 ( .A(G29GAT), .B(n380), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n371), .B(n370), .ZN(n372) );
  XNOR2_X1 U427 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U428 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U429 ( .A(n377), .B(n376), .Z(n562) );
  INV_X1 U430 ( .A(n562), .ZN(n486) );
  NAND2_X1 U431 ( .A1(n397), .A2(n486), .ZN(n526) );
  XOR2_X1 U432 ( .A(KEYINPUT24), .B(KEYINPUT87), .Z(n379) );
  XNOR2_X1 U433 ( .A(KEYINPUT23), .B(KEYINPUT90), .ZN(n378) );
  XNOR2_X1 U434 ( .A(n379), .B(n378), .ZN(n384) );
  XOR2_X1 U435 ( .A(n380), .B(KEYINPUT22), .Z(n382) );
  NAND2_X1 U436 ( .A1(G228GAT), .A2(G233GAT), .ZN(n381) );
  XNOR2_X1 U437 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U438 ( .A(n384), .B(n383), .ZN(n391) );
  XNOR2_X1 U439 ( .A(n386), .B(n385), .ZN(n389) );
  XOR2_X1 U440 ( .A(G78GAT), .B(G148GAT), .Z(n388) );
  XNOR2_X1 U441 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n420) );
  XNOR2_X1 U443 ( .A(n389), .B(n420), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U445 ( .A(n393), .B(n392), .ZN(n540) );
  XOR2_X1 U446 ( .A(KEYINPUT28), .B(n540), .Z(n493) );
  NOR2_X1 U447 ( .A1(n526), .A2(n493), .ZN(n512) );
  NAND2_X1 U448 ( .A1(n547), .A2(n512), .ZN(n405) );
  INV_X1 U449 ( .A(n547), .ZN(n491) );
  NOR2_X1 U450 ( .A1(n491), .A2(n540), .ZN(n395) );
  XNOR2_X1 U451 ( .A(KEYINPUT96), .B(KEYINPUT26), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n396) );
  XOR2_X1 U453 ( .A(KEYINPUT95), .B(n396), .Z(n564) );
  NAND2_X1 U454 ( .A1(n397), .A2(n564), .ZN(n402) );
  NAND2_X1 U455 ( .A1(n541), .A2(n491), .ZN(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT97), .B(n398), .Z(n399) );
  NAND2_X1 U457 ( .A1(n399), .A2(n540), .ZN(n400) );
  XOR2_X1 U458 ( .A(KEYINPUT25), .B(n400), .Z(n401) );
  NAND2_X1 U459 ( .A1(n402), .A2(n401), .ZN(n403) );
  NAND2_X1 U460 ( .A1(n403), .A2(n562), .ZN(n404) );
  NAND2_X1 U461 ( .A1(n405), .A2(n404), .ZN(n452) );
  NAND2_X1 U462 ( .A1(n406), .A2(n452), .ZN(n473) );
  XOR2_X1 U463 ( .A(G204GAT), .B(G120GAT), .Z(n408) );
  NAND2_X1 U464 ( .A1(G230GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n410) );
  XOR2_X1 U466 ( .A(n410), .B(n409), .Z(n418) );
  XOR2_X1 U467 ( .A(KEYINPUT73), .B(KEYINPUT32), .Z(n412) );
  XNOR2_X1 U468 ( .A(KEYINPUT31), .B(KEYINPUT72), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n416) );
  XNOR2_X1 U470 ( .A(n413), .B(KEYINPUT33), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n414), .B(KEYINPUT76), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n418), .B(n417), .ZN(n422) );
  XOR2_X1 U474 ( .A(n420), .B(n419), .Z(n421) );
  XOR2_X1 U475 ( .A(n422), .B(n421), .Z(n505) );
  INV_X1 U476 ( .A(n505), .ZN(n570) );
  XOR2_X1 U477 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n424) );
  XNOR2_X1 U478 ( .A(G141GAT), .B(G197GAT), .ZN(n423) );
  XNOR2_X1 U479 ( .A(n424), .B(n423), .ZN(n440) );
  XOR2_X1 U480 ( .A(G22GAT), .B(G15GAT), .Z(n426) );
  XNOR2_X1 U481 ( .A(G169GAT), .B(G113GAT), .ZN(n425) );
  XNOR2_X1 U482 ( .A(n426), .B(n425), .ZN(n428) );
  XOR2_X1 U483 ( .A(G36GAT), .B(G50GAT), .Z(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n436) );
  XNOR2_X1 U485 ( .A(KEYINPUT66), .B(KEYINPUT70), .ZN(n429) );
  XNOR2_X1 U486 ( .A(n429), .B(KEYINPUT69), .ZN(n430) );
  XOR2_X1 U487 ( .A(n430), .B(KEYINPUT29), .Z(n434) );
  XNOR2_X1 U488 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U489 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U490 ( .A(n436), .B(n435), .ZN(n438) );
  NAND2_X1 U491 ( .A1(G229GAT), .A2(G233GAT), .ZN(n437) );
  XNOR2_X1 U492 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n548) );
  NAND2_X1 U494 ( .A1(n570), .A2(n548), .ZN(n441) );
  XNOR2_X1 U495 ( .A(n441), .B(KEYINPUT78), .ZN(n456) );
  NOR2_X1 U496 ( .A1(n473), .A2(n456), .ZN(n442) );
  XNOR2_X1 U497 ( .A(n442), .B(KEYINPUT98), .ZN(n450) );
  NAND2_X1 U498 ( .A1(n450), .A2(n486), .ZN(n443) );
  XNOR2_X1 U499 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U500 ( .A(G1GAT), .B(n445), .ZN(G1324GAT) );
  NAND2_X1 U501 ( .A1(n450), .A2(n541), .ZN(n446) );
  XNOR2_X1 U502 ( .A(n446), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U503 ( .A(KEYINPUT35), .B(KEYINPUT100), .Z(n448) );
  NAND2_X1 U504 ( .A1(n450), .A2(n491), .ZN(n447) );
  XNOR2_X1 U505 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U506 ( .A(G15GAT), .B(n449), .ZN(G1326GAT) );
  NAND2_X1 U507 ( .A1(n450), .A2(n493), .ZN(n451) );
  XNOR2_X1 U508 ( .A(n451), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U509 ( .A(G29GAT), .B(KEYINPUT39), .Z(n460) );
  XOR2_X1 U510 ( .A(KEYINPUT36), .B(n557), .Z(n576) );
  NAND2_X1 U511 ( .A1(n573), .A2(n452), .ZN(n453) );
  NOR2_X1 U512 ( .A1(n576), .A2(n453), .ZN(n455) );
  XOR2_X1 U513 ( .A(KEYINPUT101), .B(KEYINPUT37), .Z(n454) );
  XNOR2_X1 U514 ( .A(n455), .B(n454), .ZN(n483) );
  NOR2_X1 U515 ( .A1(n456), .A2(n483), .ZN(n458) );
  XNOR2_X1 U516 ( .A(KEYINPUT102), .B(KEYINPUT38), .ZN(n457) );
  XNOR2_X1 U517 ( .A(n458), .B(n457), .ZN(n468) );
  NAND2_X1 U518 ( .A1(n468), .A2(n486), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n460), .B(n459), .ZN(G1328GAT) );
  XOR2_X1 U520 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n462) );
  NAND2_X1 U521 ( .A1(n468), .A2(n541), .ZN(n461) );
  XNOR2_X1 U522 ( .A(n462), .B(n461), .ZN(n463) );
  XNOR2_X1 U523 ( .A(G36GAT), .B(n463), .ZN(G1329GAT) );
  XNOR2_X1 U524 ( .A(G43GAT), .B(KEYINPUT105), .ZN(n467) );
  XOR2_X1 U525 ( .A(KEYINPUT40), .B(KEYINPUT106), .Z(n465) );
  NAND2_X1 U526 ( .A1(n468), .A2(n491), .ZN(n464) );
  XNOR2_X1 U527 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U528 ( .A(n467), .B(n466), .ZN(G1330GAT) );
  XOR2_X1 U529 ( .A(G50GAT), .B(KEYINPUT107), .Z(n470) );
  NAND2_X1 U530 ( .A1(n468), .A2(n493), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(G1331GAT) );
  XNOR2_X1 U532 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n475) );
  XNOR2_X1 U533 ( .A(KEYINPUT41), .B(KEYINPUT65), .ZN(n471) );
  XNOR2_X1 U534 ( .A(n471), .B(n505), .ZN(n551) );
  INV_X1 U535 ( .A(n548), .ZN(n566) );
  NAND2_X1 U536 ( .A1(n551), .A2(n566), .ZN(n472) );
  XNOR2_X1 U537 ( .A(n472), .B(KEYINPUT108), .ZN(n484) );
  NOR2_X1 U538 ( .A1(n484), .A2(n473), .ZN(n479) );
  NAND2_X1 U539 ( .A1(n479), .A2(n486), .ZN(n474) );
  XNOR2_X1 U540 ( .A(n475), .B(n474), .ZN(G1332GAT) );
  XOR2_X1 U541 ( .A(G64GAT), .B(KEYINPUT109), .Z(n477) );
  NAND2_X1 U542 ( .A1(n479), .A2(n541), .ZN(n476) );
  XNOR2_X1 U543 ( .A(n477), .B(n476), .ZN(G1333GAT) );
  NAND2_X1 U544 ( .A1(n491), .A2(n479), .ZN(n478) );
  XNOR2_X1 U545 ( .A(n478), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U546 ( .A(KEYINPUT110), .B(KEYINPUT43), .Z(n481) );
  NAND2_X1 U547 ( .A1(n479), .A2(n493), .ZN(n480) );
  XNOR2_X1 U548 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U549 ( .A(G78GAT), .B(n482), .ZN(G1335GAT) );
  NOR2_X1 U550 ( .A1(n484), .A2(n483), .ZN(n485) );
  XOR2_X1 U551 ( .A(KEYINPUT111), .B(n485), .Z(n494) );
  NAND2_X1 U552 ( .A1(n486), .A2(n494), .ZN(n487) );
  XNOR2_X1 U553 ( .A(n487), .B(KEYINPUT112), .ZN(n488) );
  XNOR2_X1 U554 ( .A(G85GAT), .B(n488), .ZN(G1336GAT) );
  XOR2_X1 U555 ( .A(G92GAT), .B(KEYINPUT113), .Z(n490) );
  NAND2_X1 U556 ( .A1(n494), .A2(n541), .ZN(n489) );
  XNOR2_X1 U557 ( .A(n490), .B(n489), .ZN(G1337GAT) );
  NAND2_X1 U558 ( .A1(n491), .A2(n494), .ZN(n492) );
  XNOR2_X1 U559 ( .A(n492), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U560 ( .A(KEYINPUT44), .B(KEYINPUT114), .Z(n496) );
  NAND2_X1 U561 ( .A1(n494), .A2(n493), .ZN(n495) );
  XNOR2_X1 U562 ( .A(n496), .B(n495), .ZN(n497) );
  XOR2_X1 U563 ( .A(G106GAT), .B(n497), .Z(G1339GAT) );
  XNOR2_X1 U564 ( .A(KEYINPUT48), .B(KEYINPUT64), .ZN(n511) );
  INV_X1 U565 ( .A(n573), .ZN(n555) );
  AND2_X1 U566 ( .A1(n548), .A2(n551), .ZN(n498) );
  XNOR2_X1 U567 ( .A(n498), .B(KEYINPUT46), .ZN(n499) );
  NOR2_X1 U568 ( .A1(n555), .A2(n499), .ZN(n500) );
  XNOR2_X1 U569 ( .A(n500), .B(KEYINPUT115), .ZN(n501) );
  NOR2_X1 U570 ( .A1(n557), .A2(n501), .ZN(n502) );
  XNOR2_X1 U571 ( .A(n502), .B(KEYINPUT47), .ZN(n509) );
  NOR2_X1 U572 ( .A1(n576), .A2(n573), .ZN(n504) );
  NOR2_X1 U573 ( .A1(n506), .A2(n505), .ZN(n507) );
  NAND2_X1 U574 ( .A1(n507), .A2(n566), .ZN(n508) );
  NAND2_X1 U575 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n542) );
  NAND2_X1 U577 ( .A1(n512), .A2(n542), .ZN(n513) );
  NOR2_X1 U578 ( .A1(n547), .A2(n513), .ZN(n522) );
  NAND2_X1 U579 ( .A1(n548), .A2(n522), .ZN(n514) );
  XNOR2_X1 U580 ( .A(n514), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U581 ( .A(KEYINPUT49), .B(KEYINPUT117), .Z(n516) );
  NAND2_X1 U582 ( .A1(n522), .A2(n551), .ZN(n515) );
  XNOR2_X1 U583 ( .A(n516), .B(n515), .ZN(n518) );
  XOR2_X1 U584 ( .A(G120GAT), .B(KEYINPUT116), .Z(n517) );
  XNOR2_X1 U585 ( .A(n518), .B(n517), .ZN(G1341GAT) );
  XOR2_X1 U586 ( .A(KEYINPUT50), .B(KEYINPUT118), .Z(n520) );
  NAND2_X1 U587 ( .A1(n522), .A2(n555), .ZN(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(n521) );
  XOR2_X1 U589 ( .A(G127GAT), .B(n521), .Z(G1342GAT) );
  XOR2_X1 U590 ( .A(G134GAT), .B(KEYINPUT51), .Z(n524) );
  NAND2_X1 U591 ( .A1(n522), .A2(n557), .ZN(n523) );
  XNOR2_X1 U592 ( .A(n524), .B(n523), .ZN(G1343GAT) );
  NAND2_X1 U593 ( .A1(n564), .A2(n542), .ZN(n525) );
  NOR2_X1 U594 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U595 ( .A(KEYINPUT119), .B(n527), .Z(n537) );
  NAND2_X1 U596 ( .A1(n548), .A2(n537), .ZN(n528) );
  XNOR2_X1 U597 ( .A(n528), .B(KEYINPUT120), .ZN(n529) );
  XNOR2_X1 U598 ( .A(G141GAT), .B(n529), .ZN(G1344GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT53), .B(KEYINPUT122), .Z(n531) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n530) );
  XNOR2_X1 U601 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U602 ( .A(KEYINPUT121), .B(n532), .Z(n534) );
  NAND2_X1 U603 ( .A1(n537), .A2(n551), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  XOR2_X1 U605 ( .A(G155GAT), .B(KEYINPUT123), .Z(n536) );
  NAND2_X1 U606 ( .A1(n537), .A2(n555), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(G1346GAT) );
  NAND2_X1 U608 ( .A1(n537), .A2(n557), .ZN(n538) );
  XNOR2_X1 U609 ( .A(n538), .B(KEYINPUT124), .ZN(n539) );
  XNOR2_X1 U610 ( .A(G162GAT), .B(n539), .ZN(G1347GAT) );
  AND2_X1 U611 ( .A1(n540), .A2(n562), .ZN(n544) );
  NAND2_X1 U612 ( .A1(n542), .A2(n541), .ZN(n543) );
  NAND2_X1 U613 ( .A1(n544), .A2(n563), .ZN(n545) );
  XOR2_X1 U614 ( .A(KEYINPUT55), .B(n545), .Z(n546) );
  NOR2_X2 U615 ( .A1(n547), .A2(n546), .ZN(n558) );
  NAND2_X1 U616 ( .A1(n548), .A2(n558), .ZN(n549) );
  XNOR2_X1 U617 ( .A(n549), .B(KEYINPUT126), .ZN(n550) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n550), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n553) );
  NAND2_X1 U620 ( .A1(n558), .A2(n551), .ZN(n552) );
  XNOR2_X1 U621 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U622 ( .A(G176GAT), .B(n554), .ZN(G1349GAT) );
  NAND2_X1 U623 ( .A1(n558), .A2(n555), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n556), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U625 ( .A(KEYINPUT58), .B(KEYINPUT127), .Z(n560) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U628 ( .A(G190GAT), .B(n561), .ZN(G1351GAT) );
  AND2_X1 U629 ( .A1(n563), .A2(n562), .ZN(n565) );
  NAND2_X1 U630 ( .A1(n565), .A2(n564), .ZN(n575) );
  NOR2_X1 U631 ( .A1(n566), .A2(n575), .ZN(n568) );
  XNOR2_X1 U632 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U634 ( .A(G197GAT), .B(n569), .ZN(G1352GAT) );
  NOR2_X1 U635 ( .A1(n570), .A2(n575), .ZN(n572) );
  XNOR2_X1 U636 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1353GAT) );
  NOR2_X1 U638 ( .A1(n573), .A2(n575), .ZN(n574) );
  XOR2_X1 U639 ( .A(G211GAT), .B(n574), .Z(G1354GAT) );
  NOR2_X1 U640 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U641 ( .A(KEYINPUT62), .B(n577), .Z(n578) );
  XNOR2_X1 U642 ( .A(G218GAT), .B(n578), .ZN(G1355GAT) );
endmodule

