

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n660, n661, n662, n663, n664, n665, n666, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778;

  INV_X1 U371 ( .A(n751), .ZN(n348) );
  INV_X1 U372 ( .A(n751), .ZN(n352) );
  XNOR2_X1 U373 ( .A(n601), .B(KEYINPUT39), .ZN(n602) );
  BUF_X1 U374 ( .A(n714), .Z(n358) );
  XNOR2_X1 U375 ( .A(n599), .B(KEYINPUT79), .ZN(n630) );
  OR2_X1 U376 ( .A1(n747), .A2(G902), .ZN(n393) );
  XNOR2_X1 U377 ( .A(n391), .B(n468), .ZN(n380) );
  XNOR2_X1 U378 ( .A(G146), .B(G125), .ZN(n509) );
  INV_X1 U379 ( .A(n347), .ZN(n660) );
  NAND2_X1 U380 ( .A1(n349), .A2(n348), .ZN(n347) );
  XNOR2_X2 U381 ( .A(n658), .B(n350), .ZN(n349) );
  INV_X1 U382 ( .A(n371), .ZN(n350) );
  INV_X1 U383 ( .A(n351), .ZN(n669) );
  NAND2_X1 U384 ( .A1(n353), .A2(n352), .ZN(n351) );
  XNOR2_X2 U385 ( .A(n666), .B(n354), .ZN(n353) );
  INV_X1 U386 ( .A(n665), .ZN(n354) );
  XNOR2_X1 U387 ( .A(n509), .B(KEYINPUT10), .ZN(n765) );
  BUF_X1 U388 ( .A(n596), .Z(n360) );
  XNOR2_X2 U389 ( .A(n603), .B(KEYINPUT40), .ZN(n662) );
  OR2_X2 U390 ( .A1(n741), .A2(G902), .ZN(n378) );
  INV_X2 U391 ( .A(n412), .ZN(n616) );
  NAND2_X2 U392 ( .A1(n413), .A2(n526), .ZN(n476) );
  NOR2_X2 U393 ( .A1(n576), .A2(n722), .ZN(n578) );
  AND2_X2 U394 ( .A1(n402), .A2(n626), .ZN(n584) );
  NAND2_X2 U395 ( .A1(n475), .A2(n709), .ZN(n611) );
  XNOR2_X1 U396 ( .A(n587), .B(n586), .ZN(n698) );
  AND2_X1 U397 ( .A1(n570), .A2(n585), .ZN(n477) );
  OR2_X1 U398 ( .A1(n424), .A2(KEYINPUT106), .ZN(n388) );
  NOR2_X1 U399 ( .A1(n441), .A2(n440), .ZN(n439) );
  XNOR2_X1 U400 ( .A(n470), .B(n469), .ZN(n404) );
  NOR2_X1 U401 ( .A1(n637), .A2(n634), .ZN(n625) );
  XNOR2_X1 U402 ( .A(n392), .B(KEYINPUT72), .ZN(n624) );
  XNOR2_X1 U403 ( .A(n502), .B(G478), .ZN(n571) );
  XNOR2_X1 U404 ( .A(n378), .B(G469), .ZN(n609) );
  NOR2_X1 U405 ( .A1(G953), .A2(G237), .ZN(n544) );
  XNOR2_X1 U406 ( .A(n409), .B(n410), .ZN(n596) );
  BUF_X1 U407 ( .A(n402), .Z(n355) );
  XNOR2_X1 U408 ( .A(n556), .B(n394), .ZN(n402) );
  BUF_X1 U409 ( .A(n747), .Z(n356) );
  BUF_X1 U410 ( .A(n607), .Z(n357) );
  XNOR2_X1 U411 ( .A(n514), .B(n406), .ZN(n768) );
  XNOR2_X2 U412 ( .A(n359), .B(KEYINPUT6), .ZN(n623) );
  BUF_X1 U413 ( .A(n596), .Z(n359) );
  NAND2_X2 U414 ( .A1(n418), .A2(n525), .ZN(n453) );
  XNOR2_X2 U415 ( .A(n454), .B(KEYINPUT19), .ZN(n418) );
  BUF_X1 U416 ( .A(n663), .Z(n745) );
  AND2_X1 U417 ( .A1(n620), .A2(n404), .ZN(n385) );
  NAND2_X1 U418 ( .A1(n704), .A2(n422), .ZN(n421) );
  NOR2_X1 U419 ( .A1(n382), .A2(n384), .ZN(n430) );
  XNOR2_X1 U420 ( .A(n385), .B(n621), .ZN(n384) );
  XNOR2_X1 U421 ( .A(n552), .B(n370), .ZN(n732) );
  NOR2_X1 U422 ( .A1(n575), .A2(n560), .ZN(n552) );
  NOR2_X1 U423 ( .A1(n559), .A2(n623), .ZN(n403) );
  XNOR2_X1 U424 ( .A(n491), .B(n435), .ZN(n572) );
  XNOR2_X1 U425 ( .A(n492), .B(n493), .ZN(n435) );
  XNOR2_X1 U426 ( .A(n463), .B(KEYINPUT105), .ZN(n704) );
  XOR2_X1 U427 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n516) );
  INV_X1 U428 ( .A(G119), .ZN(n505) );
  XNOR2_X1 U429 ( .A(n377), .B(G140), .ZN(n538) );
  INV_X1 U430 ( .A(G137), .ZN(n377) );
  INV_X1 U431 ( .A(KEYINPUT8), .ZN(n468) );
  XOR2_X1 U432 ( .A(KEYINPUT12), .B(KEYINPUT99), .Z(n482) );
  XNOR2_X1 U433 ( .A(KEYINPUT78), .B(G110), .ZN(n503) );
  XNOR2_X1 U434 ( .A(n538), .B(n376), .ZN(n766) );
  INV_X1 U435 ( .A(KEYINPUT94), .ZN(n376) );
  XNOR2_X1 U436 ( .A(n631), .B(KEYINPUT48), .ZN(n632) );
  XOR2_X1 U437 ( .A(KEYINPUT23), .B(G110), .Z(n530) );
  XNOR2_X1 U438 ( .A(G119), .B(G128), .ZN(n529) );
  XNOR2_X1 U439 ( .A(n765), .B(n474), .ZN(n389) );
  XNOR2_X1 U440 ( .A(n532), .B(KEYINPUT24), .ZN(n474) );
  XNOR2_X1 U441 ( .A(n537), .B(KEYINPUT4), .ZN(n406) );
  XNOR2_X1 U442 ( .A(G134), .B(G131), .ZN(n537) );
  XOR2_X1 U443 ( .A(KEYINPUT81), .B(G101), .Z(n541) );
  INV_X1 U444 ( .A(n576), .ZN(n579) );
  INV_X1 U445 ( .A(KEYINPUT34), .ZN(n479) );
  INV_X1 U446 ( .A(KEYINPUT22), .ZN(n394) );
  AND2_X1 U447 ( .A1(n709), .A2(n553), .ZN(n554) );
  XNOR2_X1 U448 ( .A(n578), .B(n577), .ZN(n688) );
  XNOR2_X1 U449 ( .A(n471), .B(n608), .ZN(n619) );
  NOR2_X1 U450 ( .A1(n624), .A2(n360), .ZN(n471) );
  XNOR2_X1 U451 ( .A(n535), .B(n397), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n536), .B(n398), .ZN(n397) );
  NAND2_X1 U453 ( .A1(n602), .A2(n685), .ZN(n603) );
  INV_X1 U454 ( .A(n682), .ZN(n462) );
  XNOR2_X1 U455 ( .A(G113), .B(G101), .ZN(n506) );
  AND2_X1 U456 ( .A1(n424), .A2(n368), .ZN(n419) );
  XNOR2_X1 U457 ( .A(KEYINPUT90), .B(KEYINPUT92), .ZN(n515) );
  NOR2_X1 U458 ( .A1(n639), .A2(KEYINPUT85), .ZN(n441) );
  INV_X1 U459 ( .A(n661), .ZN(n440) );
  INV_X1 U460 ( .A(KEYINPUT85), .ZN(n444) );
  NAND2_X1 U461 ( .A1(G234), .A2(G237), .ZN(n520) );
  NOR2_X1 U462 ( .A1(n571), .A2(n572), .ZN(n709) );
  OR2_X1 U463 ( .A1(n575), .A2(n360), .ZN(n722) );
  OR2_X1 U464 ( .A1(G237), .A2(G902), .ZN(n480) );
  XNOR2_X1 U465 ( .A(KEYINPUT89), .B(KEYINPUT15), .ZN(n400) );
  NAND2_X1 U466 ( .A1(n595), .A2(n450), .ZN(n448) );
  NAND2_X1 U467 ( .A1(n607), .A2(n606), .ZN(n392) );
  INV_X1 U468 ( .A(KEYINPUT25), .ZN(n398) );
  XNOR2_X1 U469 ( .A(n550), .B(n405), .ZN(n648) );
  XNOR2_X1 U470 ( .A(n768), .B(G146), .ZN(n405) );
  XNOR2_X1 U471 ( .A(n457), .B(n549), .ZN(n758) );
  XNOR2_X1 U472 ( .A(n539), .B(n458), .ZN(n457) );
  XNOR2_X1 U473 ( .A(n459), .B(KEYINPUT16), .ZN(n458) );
  XOR2_X1 U474 ( .A(KEYINPUT7), .B(KEYINPUT103), .Z(n498) );
  XNOR2_X1 U475 ( .A(KEYINPUT9), .B(KEYINPUT102), .ZN(n497) );
  XNOR2_X1 U476 ( .A(G116), .B(G134), .ZN(n495) );
  XOR2_X1 U477 ( .A(G107), .B(G122), .Z(n496) );
  XNOR2_X1 U478 ( .A(n489), .B(n434), .ZN(n664) );
  XNOR2_X1 U479 ( .A(n490), .B(n765), .ZN(n434) );
  NAND2_X1 U480 ( .A1(n465), .A2(n571), .ZN(n464) );
  NOR2_X1 U481 ( .A1(n607), .A2(n716), .ZN(n714) );
  XNOR2_X1 U482 ( .A(n531), .B(n533), .ZN(n472) );
  XOR2_X1 U483 ( .A(KEYINPUT59), .B(n664), .Z(n665) );
  XNOR2_X1 U484 ( .A(n542), .B(n361), .ZN(n379) );
  OR2_X1 U485 ( .A1(n627), .A2(n626), .ZN(n437) );
  INV_X1 U486 ( .A(KEYINPUT35), .ZN(n372) );
  XNOR2_X1 U487 ( .A(n375), .B(n479), .ZN(n374) );
  XNOR2_X1 U488 ( .A(n401), .B(n461), .ZN(n778) );
  XNOR2_X1 U489 ( .A(n561), .B(KEYINPUT32), .ZN(n461) );
  INV_X1 U490 ( .A(KEYINPUT82), .ZN(n469) );
  NAND2_X1 U491 ( .A1(n619), .A2(n618), .ZN(n470) );
  INV_X1 U492 ( .A(n571), .ZN(n573) );
  XNOR2_X1 U493 ( .A(n616), .B(G137), .ZN(G39) );
  XOR2_X1 U494 ( .A(n541), .B(n540), .Z(n361) );
  XOR2_X1 U495 ( .A(n516), .B(n515), .Z(n362) );
  AND2_X1 U496 ( .A1(n623), .A2(n685), .ZN(n363) );
  INV_X1 U497 ( .A(n704), .ZN(n423) );
  AND2_X1 U498 ( .A1(n572), .A2(n571), .ZN(n364) );
  AND2_X1 U499 ( .A1(n404), .A2(n622), .ZN(n365) );
  INV_X1 U500 ( .A(n526), .ZN(n641) );
  XNOR2_X1 U501 ( .A(n400), .B(n399), .ZN(n526) );
  BUF_X1 U502 ( .A(n557), .Z(n713) );
  INV_X1 U503 ( .A(G902), .ZN(n399) );
  AND2_X1 U504 ( .A1(n670), .A2(n421), .ZN(n366) );
  AND2_X1 U505 ( .A1(n647), .A2(n652), .ZN(G63) );
  AND2_X1 U506 ( .A1(n423), .A2(KEYINPUT106), .ZN(n368) );
  XNOR2_X1 U507 ( .A(n464), .B(KEYINPUT104), .ZN(n673) );
  INV_X1 U508 ( .A(n673), .ZN(n395) );
  XNOR2_X1 U509 ( .A(KEYINPUT87), .B(KEYINPUT0), .ZN(n369) );
  INV_X1 U510 ( .A(KEYINPUT106), .ZN(n422) );
  XOR2_X1 U511 ( .A(KEYINPUT88), .B(KEYINPUT33), .Z(n370) );
  XNOR2_X1 U512 ( .A(n411), .B(n379), .ZN(n741) );
  XOR2_X1 U513 ( .A(n657), .B(n656), .Z(n371) );
  INV_X1 U514 ( .A(G953), .ZN(n753) );
  XNOR2_X2 U515 ( .A(n373), .B(n372), .ZN(n777) );
  NAND2_X1 U516 ( .A1(n374), .A2(n364), .ZN(n373) );
  NAND2_X1 U517 ( .A1(n732), .A2(n579), .ZN(n375) );
  NAND2_X1 U518 ( .A1(n380), .A2(G217), .ZN(n467) );
  NAND2_X1 U519 ( .A1(n380), .A2(G221), .ZN(n390) );
  NOR2_X1 U520 ( .A1(n381), .A2(n365), .ZN(n383) );
  NAND2_X1 U521 ( .A1(n437), .A2(n462), .ZN(n381) );
  NAND2_X1 U522 ( .A1(n383), .A2(n432), .ZN(n382) );
  XNOR2_X1 U523 ( .A(n514), .B(KEYINPUT4), .ZN(n387) );
  XNOR2_X2 U524 ( .A(n386), .B(n494), .ZN(n514) );
  XNOR2_X2 U525 ( .A(G143), .B(KEYINPUT66), .ZN(n386) );
  XNOR2_X1 U526 ( .A(n387), .B(n362), .ZN(n460) );
  NAND2_X1 U527 ( .A1(n388), .A2(n366), .ZN(n420) );
  XNOR2_X1 U528 ( .A(n582), .B(n425), .ZN(n424) );
  XNOR2_X1 U529 ( .A(n390), .B(n389), .ZN(n473) );
  NAND2_X1 U530 ( .A1(n511), .A2(G234), .ZN(n391) );
  XNOR2_X2 U531 ( .A(n393), .B(n396), .ZN(n607) );
  NAND2_X1 U532 ( .A1(n602), .A2(n395), .ZN(n661) );
  XNOR2_X1 U533 ( .A(n473), .B(n472), .ZN(n747) );
  NAND2_X1 U534 ( .A1(n403), .A2(n355), .ZN(n401) );
  NAND2_X1 U535 ( .A1(n404), .A2(n395), .ZN(n680) );
  NAND2_X1 U536 ( .A1(n404), .A2(n685), .ZN(n683) );
  NAND2_X1 U537 ( .A1(n584), .A2(n583), .ZN(n670) );
  BUF_X1 U538 ( .A(n688), .Z(n407) );
  BUF_X1 U539 ( .A(n706), .Z(n408) );
  NOR2_X1 U540 ( .A1(n648), .A2(G902), .ZN(n409) );
  XOR2_X1 U541 ( .A(n551), .B(G472), .Z(n410) );
  NAND2_X1 U542 ( .A1(n429), .A2(n617), .ZN(n428) );
  XNOR2_X1 U543 ( .A(n768), .B(G146), .ZN(n411) );
  XNOR2_X2 U544 ( .A(n615), .B(n614), .ZN(n412) );
  XNOR2_X2 U545 ( .A(n455), .B(n758), .ZN(n413) );
  NAND2_X1 U546 ( .A1(n460), .A2(n456), .ZN(n415) );
  NAND2_X1 U547 ( .A1(n414), .A2(n517), .ZN(n416) );
  NAND2_X1 U548 ( .A1(n416), .A2(n415), .ZN(n455) );
  INV_X1 U549 ( .A(n460), .ZN(n414) );
  BUF_X1 U550 ( .A(n696), .Z(n417) );
  AND2_X1 U551 ( .A1(n418), .A2(n609), .ZN(n618) );
  NOR2_X1 U552 ( .A1(n420), .A2(n419), .ZN(n585) );
  INV_X1 U553 ( .A(KEYINPUT98), .ZN(n425) );
  NAND2_X1 U554 ( .A1(n426), .A2(n612), .ZN(n615) );
  NAND2_X1 U555 ( .A1(n426), .A2(n732), .ZN(n733) );
  NAND2_X1 U556 ( .A1(n725), .A2(n426), .ZN(n726) );
  XNOR2_X2 U557 ( .A(n611), .B(KEYINPUT41), .ZN(n426) );
  NAND2_X1 U558 ( .A1(n428), .A2(n427), .ZN(n431) );
  NAND2_X1 U559 ( .A1(n436), .A2(n662), .ZN(n427) );
  INV_X1 U560 ( .A(n662), .ZN(n429) );
  NAND2_X1 U561 ( .A1(n431), .A2(n430), .ZN(n633) );
  NAND2_X1 U562 ( .A1(n412), .A2(KEYINPUT46), .ZN(n432) );
  NAND2_X1 U563 ( .A1(n442), .A2(n439), .ZN(n438) );
  NOR2_X1 U564 ( .A1(n688), .A2(n674), .ZN(n582) );
  NAND2_X1 U565 ( .A1(n534), .A2(G217), .ZN(n535) );
  XNOR2_X1 U566 ( .A(n527), .B(KEYINPUT20), .ZN(n534) );
  NOR2_X2 U567 ( .A1(n438), .A2(n445), .ZN(n770) );
  NAND2_X1 U568 ( .A1(n698), .A2(n770), .ZN(n696) );
  INV_X1 U569 ( .A(n555), .ZN(n576) );
  AND2_X1 U570 ( .A1(n555), .A2(n358), .ZN(n580) );
  XNOR2_X2 U571 ( .A(n453), .B(n369), .ZN(n555) );
  NOR2_X1 U572 ( .A1(n694), .A2(n444), .ZN(n443) );
  NAND2_X1 U573 ( .A1(n363), .A2(n433), .ZN(n634) );
  NOR2_X1 U574 ( .A1(n624), .A2(n595), .ZN(n433) );
  INV_X1 U575 ( .A(n437), .ZN(n691) );
  NAND2_X1 U576 ( .A1(n616), .A2(n617), .ZN(n436) );
  NAND2_X1 U577 ( .A1(n640), .A2(n443), .ZN(n442) );
  NOR2_X1 U578 ( .A1(n640), .A2(KEYINPUT85), .ZN(n445) );
  NAND2_X1 U579 ( .A1(n446), .A2(n598), .ZN(n599) );
  NOR2_X1 U580 ( .A1(n451), .A2(n447), .ZN(n446) );
  NAND2_X1 U581 ( .A1(n449), .A2(n448), .ZN(n447) );
  NAND2_X1 U582 ( .A1(n360), .A2(n450), .ZN(n449) );
  INV_X1 U583 ( .A(n597), .ZN(n450) );
  NOR2_X1 U584 ( .A1(n360), .A2(n452), .ZN(n451) );
  NAND2_X1 U585 ( .A1(n705), .A2(n597), .ZN(n452) );
  NAND2_X1 U586 ( .A1(n628), .A2(n705), .ZN(n454) );
  INV_X1 U587 ( .A(n413), .ZN(n655) );
  INV_X1 U588 ( .A(n517), .ZN(n456) );
  INV_X1 U589 ( .A(G122), .ZN(n459) );
  NAND2_X1 U590 ( .A1(n568), .A2(n777), .ZN(n565) );
  NOR2_X1 U591 ( .A1(n679), .A2(n778), .ZN(n568) );
  NOR2_X2 U592 ( .A1(n581), .A2(n593), .ZN(n674) );
  NAND2_X1 U593 ( .A1(n574), .A2(n673), .ZN(n463) );
  INV_X1 U594 ( .A(n572), .ZN(n465) );
  XNOR2_X1 U595 ( .A(n501), .B(n466), .ZN(n644) );
  XNOR2_X1 U596 ( .A(n514), .B(n467), .ZN(n466) );
  NAND2_X1 U597 ( .A1(n423), .A2(n475), .ZN(n711) );
  XNOR2_X2 U598 ( .A(n610), .B(KEYINPUT111), .ZN(n475) );
  XNOR2_X1 U599 ( .A(n628), .B(n600), .ZN(n706) );
  XNOR2_X2 U600 ( .A(n476), .B(n519), .ZN(n628) );
  NAND2_X1 U601 ( .A1(n477), .A2(n478), .ZN(n587) );
  NAND2_X1 U602 ( .A1(n569), .A2(n568), .ZN(n478) );
  XNOR2_X1 U603 ( .A(n645), .B(n644), .ZN(n647) );
  INV_X1 U604 ( .A(n626), .ZN(n557) );
  XNOR2_X1 U605 ( .A(n609), .B(n543), .ZN(n626) );
  BUF_X1 U606 ( .A(n698), .Z(n752) );
  INV_X1 U607 ( .A(KEYINPUT95), .ZN(n532) );
  INV_X1 U608 ( .A(n716), .ZN(n553) );
  INV_X1 U609 ( .A(KEYINPUT123), .ZN(n746) );
  INV_X1 U610 ( .A(KEYINPUT108), .ZN(n562) );
  INV_X1 U611 ( .A(n751), .ZN(n652) );
  XNOR2_X1 U612 ( .A(n356), .B(n746), .ZN(n748) );
  XNOR2_X1 U613 ( .A(n749), .B(n748), .ZN(n750) );
  XNOR2_X1 U614 ( .A(KEYINPUT101), .B(KEYINPUT13), .ZN(n492) );
  NAND2_X1 U615 ( .A1(G214), .A2(n544), .ZN(n481) );
  XNOR2_X1 U616 ( .A(n482), .B(n481), .ZN(n490) );
  XOR2_X1 U617 ( .A(G104), .B(G122), .Z(n484) );
  XNOR2_X1 U618 ( .A(G113), .B(G131), .ZN(n483) );
  XNOR2_X1 U619 ( .A(n484), .B(n483), .ZN(n488) );
  XOR2_X1 U620 ( .A(KEYINPUT11), .B(KEYINPUT100), .Z(n486) );
  XNOR2_X1 U621 ( .A(G143), .B(G140), .ZN(n485) );
  XNOR2_X1 U622 ( .A(n486), .B(n485), .ZN(n487) );
  XOR2_X1 U623 ( .A(n488), .B(n487), .Z(n489) );
  NOR2_X1 U624 ( .A1(G902), .A2(n664), .ZN(n491) );
  INV_X1 U625 ( .A(G475), .ZN(n493) );
  INV_X1 U626 ( .A(G128), .ZN(n494) );
  XNOR2_X1 U627 ( .A(n496), .B(n495), .ZN(n500) );
  XNOR2_X1 U628 ( .A(n498), .B(n497), .ZN(n499) );
  XOR2_X1 U629 ( .A(n500), .B(n499), .Z(n501) );
  XNOR2_X2 U630 ( .A(G953), .B(KEYINPUT64), .ZN(n588) );
  INV_X1 U631 ( .A(n588), .ZN(n511) );
  NAND2_X1 U632 ( .A1(n644), .A2(n399), .ZN(n502) );
  XNOR2_X1 U633 ( .A(KEYINPUT76), .B(n480), .ZN(n518) );
  NAND2_X1 U634 ( .A1(n518), .A2(G214), .ZN(n705) );
  XOR2_X1 U635 ( .A(G104), .B(G107), .Z(n504) );
  XNOR2_X1 U636 ( .A(n504), .B(n503), .ZN(n539) );
  XNOR2_X1 U637 ( .A(n506), .B(n505), .ZN(n508) );
  XOR2_X1 U638 ( .A(KEYINPUT3), .B(G116), .Z(n507) );
  XNOR2_X1 U639 ( .A(n508), .B(n507), .ZN(n549) );
  INV_X1 U640 ( .A(n509), .ZN(n510) );
  XOR2_X1 U641 ( .A(KEYINPUT91), .B(n510), .Z(n513) );
  NAND2_X1 U642 ( .A1(G224), .A2(n511), .ZN(n512) );
  XNOR2_X1 U643 ( .A(n513), .B(n512), .ZN(n517) );
  AND2_X1 U644 ( .A1(n518), .A2(G210), .ZN(n519) );
  NOR2_X1 U645 ( .A1(G898), .A2(n753), .ZN(n760) );
  XNOR2_X1 U646 ( .A(n520), .B(KEYINPUT14), .ZN(n522) );
  NAND2_X1 U647 ( .A1(n522), .A2(G902), .ZN(n521) );
  XNOR2_X1 U648 ( .A(n521), .B(KEYINPUT93), .ZN(n589) );
  NAND2_X1 U649 ( .A1(n760), .A2(n589), .ZN(n524) );
  NAND2_X1 U650 ( .A1(G952), .A2(n522), .ZN(n730) );
  NOR2_X1 U651 ( .A1(G953), .A2(n730), .ZN(n591) );
  INV_X1 U652 ( .A(n591), .ZN(n523) );
  NAND2_X1 U653 ( .A1(n524), .A2(n523), .ZN(n525) );
  NAND2_X1 U654 ( .A1(G234), .A2(n526), .ZN(n527) );
  NAND2_X1 U655 ( .A1(G221), .A2(n534), .ZN(n528) );
  XNOR2_X1 U656 ( .A(n528), .B(KEYINPUT21), .ZN(n716) );
  XNOR2_X1 U657 ( .A(n530), .B(n529), .ZN(n533) );
  XOR2_X1 U658 ( .A(n538), .B(KEYINPUT73), .Z(n531) );
  XOR2_X1 U659 ( .A(KEYINPUT96), .B(KEYINPUT80), .Z(n536) );
  XNOR2_X1 U660 ( .A(n539), .B(n766), .ZN(n542) );
  NAND2_X1 U661 ( .A1(G227), .A2(n511), .ZN(n540) );
  XNOR2_X1 U662 ( .A(KEYINPUT1), .B(KEYINPUT69), .ZN(n543) );
  NAND2_X1 U663 ( .A1(n358), .A2(n557), .ZN(n575) );
  NAND2_X1 U664 ( .A1(n544), .A2(G210), .ZN(n545) );
  XNOR2_X1 U665 ( .A(n545), .B(G137), .ZN(n547) );
  XNOR2_X1 U666 ( .A(KEYINPUT77), .B(KEYINPUT5), .ZN(n546) );
  XNOR2_X1 U667 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U668 ( .A(n549), .B(n548), .ZN(n550) );
  INV_X1 U669 ( .A(KEYINPUT74), .ZN(n551) );
  INV_X1 U670 ( .A(n623), .ZN(n560) );
  INV_X1 U671 ( .A(KEYINPUT68), .ZN(n561) );
  NAND2_X1 U672 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U673 ( .A1(n607), .A2(n713), .ZN(n558) );
  XOR2_X1 U674 ( .A(KEYINPUT107), .B(n558), .Z(n559) );
  XNOR2_X1 U675 ( .A(n584), .B(n562), .ZN(n564) );
  INV_X1 U676 ( .A(n360), .ZN(n718) );
  NAND2_X1 U677 ( .A1(n357), .A2(n360), .ZN(n563) );
  NOR2_X1 U678 ( .A1(n564), .A2(n563), .ZN(n679) );
  NAND2_X1 U679 ( .A1(n565), .A2(KEYINPUT44), .ZN(n570) );
  INV_X1 U680 ( .A(KEYINPUT44), .ZN(n566) );
  NAND2_X1 U681 ( .A1(n777), .A2(n566), .ZN(n567) );
  XNOR2_X1 U682 ( .A(n567), .B(KEYINPUT71), .ZN(n569) );
  AND2_X1 U683 ( .A1(n573), .A2(n572), .ZN(n685) );
  INV_X1 U684 ( .A(n685), .ZN(n574) );
  XNOR2_X1 U685 ( .A(KEYINPUT97), .B(KEYINPUT31), .ZN(n577) );
  NAND2_X1 U686 ( .A1(n580), .A2(n360), .ZN(n581) );
  INV_X1 U687 ( .A(n609), .ZN(n593) );
  NOR2_X1 U688 ( .A1(n357), .A2(n623), .ZN(n583) );
  XOR2_X1 U689 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n586) );
  NAND2_X1 U690 ( .A1(n588), .A2(n589), .ZN(n590) );
  NOR2_X1 U691 ( .A1(G900), .A2(n590), .ZN(n592) );
  OR2_X1 U692 ( .A1(n592), .A2(n591), .ZN(n604) );
  NAND2_X1 U693 ( .A1(n714), .A2(n604), .ZN(n594) );
  NOR2_X1 U694 ( .A1(n594), .A2(n593), .ZN(n598) );
  INV_X1 U695 ( .A(n705), .ZN(n595) );
  XNOR2_X1 U696 ( .A(KEYINPUT109), .B(KEYINPUT30), .ZN(n597) );
  INV_X1 U697 ( .A(KEYINPUT38), .ZN(n600) );
  NAND2_X1 U698 ( .A1(n630), .A2(n408), .ZN(n601) );
  INV_X1 U699 ( .A(n604), .ZN(n605) );
  NOR2_X1 U700 ( .A1(n716), .A2(n605), .ZN(n606) );
  XNOR2_X1 U701 ( .A(KEYINPUT28), .B(KEYINPUT110), .ZN(n608) );
  AND2_X1 U702 ( .A1(n619), .A2(n609), .ZN(n612) );
  NAND2_X1 U703 ( .A1(n706), .A2(n705), .ZN(n610) );
  INV_X1 U704 ( .A(KEYINPUT112), .ZN(n613) );
  XNOR2_X1 U705 ( .A(n613), .B(KEYINPUT42), .ZN(n614) );
  INV_X1 U706 ( .A(KEYINPUT46), .ZN(n617) );
  NOR2_X1 U707 ( .A1(KEYINPUT75), .A2(n704), .ZN(n620) );
  INV_X1 U708 ( .A(KEYINPUT47), .ZN(n621) );
  AND2_X1 U709 ( .A1(KEYINPUT75), .A2(n704), .ZN(n622) );
  INV_X1 U710 ( .A(n628), .ZN(n637) );
  XOR2_X1 U711 ( .A(KEYINPUT36), .B(n625), .Z(n627) );
  AND2_X1 U712 ( .A1(n628), .A2(n364), .ZN(n629) );
  AND2_X1 U713 ( .A1(n630), .A2(n629), .ZN(n682) );
  INV_X1 U714 ( .A(KEYINPUT86), .ZN(n631) );
  XNOR2_X1 U715 ( .A(n633), .B(n632), .ZN(n640) );
  NOR2_X1 U716 ( .A1(n713), .A2(n634), .ZN(n636) );
  INV_X1 U717 ( .A(KEYINPUT43), .ZN(n635) );
  XNOR2_X1 U718 ( .A(n636), .B(n635), .ZN(n638) );
  AND2_X1 U719 ( .A1(n638), .A2(n637), .ZN(n694) );
  INV_X1 U720 ( .A(n694), .ZN(n639) );
  XNOR2_X1 U721 ( .A(n696), .B(KEYINPUT2), .ZN(n642) );
  NAND2_X1 U722 ( .A1(n642), .A2(n641), .ZN(n643) );
  XNOR2_X2 U723 ( .A(n643), .B(KEYINPUT67), .ZN(n663) );
  NAND2_X1 U724 ( .A1(n745), .A2(G478), .ZN(n645) );
  INV_X1 U725 ( .A(G952), .ZN(n646) );
  AND2_X1 U726 ( .A1(n588), .A2(n646), .ZN(n751) );
  NAND2_X1 U727 ( .A1(n663), .A2(G472), .ZN(n650) );
  XNOR2_X1 U728 ( .A(n648), .B(KEYINPUT62), .ZN(n649) );
  XNOR2_X1 U729 ( .A(n650), .B(n649), .ZN(n651) );
  INV_X1 U730 ( .A(n651), .ZN(n653) );
  NAND2_X1 U731 ( .A1(n653), .A2(n652), .ZN(n654) );
  XNOR2_X1 U732 ( .A(n654), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U733 ( .A1(n663), .A2(G210), .ZN(n658) );
  XOR2_X1 U734 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n657) );
  XNOR2_X1 U735 ( .A(n655), .B(KEYINPUT83), .ZN(n656) );
  XNOR2_X1 U736 ( .A(n660), .B(KEYINPUT56), .ZN(G51) );
  XNOR2_X1 U737 ( .A(n661), .B(G134), .ZN(G36) );
  XNOR2_X1 U738 ( .A(n662), .B(G131), .ZN(G33) );
  NAND2_X1 U739 ( .A1(n663), .A2(G475), .ZN(n666) );
  XNOR2_X1 U740 ( .A(KEYINPUT70), .B(KEYINPUT60), .ZN(n668) );
  XNOR2_X1 U741 ( .A(n669), .B(n668), .ZN(G60) );
  XNOR2_X1 U742 ( .A(G101), .B(n670), .ZN(G3) );
  XOR2_X1 U743 ( .A(G104), .B(KEYINPUT113), .Z(n672) );
  NAND2_X1 U744 ( .A1(n674), .A2(n685), .ZN(n671) );
  XNOR2_X1 U745 ( .A(n672), .B(n671), .ZN(G6) );
  XNOR2_X1 U746 ( .A(G107), .B(KEYINPUT114), .ZN(n678) );
  XOR2_X1 U747 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n676) );
  NAND2_X1 U748 ( .A1(n674), .A2(n395), .ZN(n675) );
  XNOR2_X1 U749 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U750 ( .A(n678), .B(n677), .ZN(G9) );
  XOR2_X1 U751 ( .A(G110), .B(n679), .Z(G12) );
  XOR2_X1 U752 ( .A(G128), .B(KEYINPUT29), .Z(n681) );
  XNOR2_X1 U753 ( .A(n681), .B(n680), .ZN(G30) );
  XOR2_X1 U754 ( .A(G143), .B(n682), .Z(G45) );
  XOR2_X1 U755 ( .A(G146), .B(KEYINPUT115), .Z(n684) );
  XNOR2_X1 U756 ( .A(n684), .B(n683), .ZN(G48) );
  NAND2_X1 U757 ( .A1(n407), .A2(n685), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n686), .B(KEYINPUT116), .ZN(n687) );
  XNOR2_X1 U759 ( .A(G113), .B(n687), .ZN(G15) );
  XOR2_X1 U760 ( .A(G116), .B(KEYINPUT117), .Z(n690) );
  NAND2_X1 U761 ( .A1(n407), .A2(n395), .ZN(n689) );
  XNOR2_X1 U762 ( .A(n690), .B(n689), .ZN(G18) );
  XNOR2_X1 U763 ( .A(n691), .B(KEYINPUT37), .ZN(n692) );
  XNOR2_X1 U764 ( .A(n692), .B(KEYINPUT118), .ZN(n693) );
  XNOR2_X1 U765 ( .A(G125), .B(n693), .ZN(G27) );
  XNOR2_X1 U766 ( .A(G140), .B(n694), .ZN(n695) );
  XNOR2_X1 U767 ( .A(n695), .B(KEYINPUT119), .ZN(G42) );
  NAND2_X1 U768 ( .A1(n417), .A2(KEYINPUT84), .ZN(n697) );
  XOR2_X1 U769 ( .A(KEYINPUT2), .B(n697), .Z(n703) );
  INV_X1 U770 ( .A(n770), .ZN(n699) );
  NAND2_X1 U771 ( .A1(n752), .A2(n699), .ZN(n701) );
  INV_X1 U772 ( .A(KEYINPUT84), .ZN(n700) );
  NAND2_X1 U773 ( .A1(n701), .A2(n700), .ZN(n702) );
  NAND2_X1 U774 ( .A1(n703), .A2(n702), .ZN(n737) );
  NOR2_X1 U775 ( .A1(n408), .A2(n705), .ZN(n707) );
  XOR2_X1 U776 ( .A(KEYINPUT120), .B(n707), .Z(n708) );
  NAND2_X1 U777 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U778 ( .A1(n711), .A2(n710), .ZN(n712) );
  NAND2_X1 U779 ( .A1(n712), .A2(n732), .ZN(n727) );
  NOR2_X1 U780 ( .A1(n358), .A2(n713), .ZN(n715) );
  XOR2_X1 U781 ( .A(KEYINPUT50), .B(n715), .Z(n721) );
  NAND2_X1 U782 ( .A1(n357), .A2(n716), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(KEYINPUT49), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U785 ( .A1(n721), .A2(n720), .ZN(n723) );
  NAND2_X1 U786 ( .A1(n723), .A2(n722), .ZN(n724) );
  XOR2_X1 U787 ( .A(KEYINPUT51), .B(n724), .Z(n725) );
  NAND2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U789 ( .A(KEYINPUT52), .B(n728), .Z(n729) );
  NOR2_X1 U790 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U791 ( .A(n731), .B(KEYINPUT121), .ZN(n734) );
  NAND2_X1 U792 ( .A1(n734), .A2(n733), .ZN(n735) );
  NOR2_X1 U793 ( .A1(G953), .A2(n735), .ZN(n736) );
  NAND2_X1 U794 ( .A1(n737), .A2(n736), .ZN(n738) );
  XOR2_X1 U795 ( .A(KEYINPUT53), .B(n738), .Z(G75) );
  NAND2_X1 U796 ( .A1(n745), .A2(G469), .ZN(n743) );
  XNOR2_X1 U797 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n739) );
  XOR2_X1 U798 ( .A(n739), .B(KEYINPUT57), .Z(n740) );
  XNOR2_X1 U799 ( .A(n741), .B(n740), .ZN(n742) );
  XNOR2_X1 U800 ( .A(n743), .B(n742), .ZN(n744) );
  NOR2_X1 U801 ( .A1(n751), .A2(n744), .ZN(G54) );
  NAND2_X1 U802 ( .A1(n745), .A2(G217), .ZN(n749) );
  NOR2_X1 U803 ( .A1(n751), .A2(n750), .ZN(G66) );
  NAND2_X1 U804 ( .A1(n753), .A2(n752), .ZN(n757) );
  NAND2_X1 U805 ( .A1(G953), .A2(G224), .ZN(n754) );
  XNOR2_X1 U806 ( .A(KEYINPUT61), .B(n754), .ZN(n755) );
  NAND2_X1 U807 ( .A1(n755), .A2(G898), .ZN(n756) );
  NAND2_X1 U808 ( .A1(n757), .A2(n756), .ZN(n763) );
  XOR2_X1 U809 ( .A(n758), .B(KEYINPUT125), .Z(n759) );
  NOR2_X1 U810 ( .A1(n760), .A2(n759), .ZN(n761) );
  XOR2_X1 U811 ( .A(KEYINPUT124), .B(n761), .Z(n762) );
  XNOR2_X1 U812 ( .A(n763), .B(n762), .ZN(n764) );
  XOR2_X1 U813 ( .A(KEYINPUT126), .B(n764), .Z(G69) );
  XOR2_X1 U814 ( .A(n765), .B(n766), .Z(n767) );
  XOR2_X1 U815 ( .A(n768), .B(n767), .Z(n772) );
  XNOR2_X1 U816 ( .A(n772), .B(KEYINPUT127), .ZN(n769) );
  XNOR2_X1 U817 ( .A(n770), .B(n769), .ZN(n771) );
  NAND2_X1 U818 ( .A1(n771), .A2(n511), .ZN(n776) );
  XNOR2_X1 U819 ( .A(n772), .B(G227), .ZN(n773) );
  NAND2_X1 U820 ( .A1(n773), .A2(G900), .ZN(n774) );
  NAND2_X1 U821 ( .A1(n774), .A2(G953), .ZN(n775) );
  NAND2_X1 U822 ( .A1(n776), .A2(n775), .ZN(G72) );
  XNOR2_X1 U823 ( .A(n777), .B(G122), .ZN(G24) );
  XOR2_X1 U824 ( .A(n778), .B(G119), .Z(G21) );
endmodule

