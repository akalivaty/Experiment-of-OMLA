//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 0 1 0 1 1 0 0 0 0 0 0 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 0 0 1 1 1 0 1 1 0 0 1 1 0 1 1 0 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n634, new_n635, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n803, new_n804, new_n806, new_n807,
    new_n808, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n860,
    new_n861, new_n863, new_n864, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n879, new_n880, new_n881, new_n883, new_n884, new_n885, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920;
  XOR2_X1   g000(.A(G113gat), .B(G120gat), .Z(new_n202));
  INV_X1    g001(.A(KEYINPUT1), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G134gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G127gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n206), .A2(KEYINPUT72), .ZN(new_n207));
  OAI21_X1  g006(.A(KEYINPUT73), .B1(new_n205), .B2(G127gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT72), .ZN(new_n209));
  NAND3_X1  g008(.A1(new_n209), .A2(new_n205), .A3(G127gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT73), .ZN(new_n211));
  INV_X1    g010(.A(G127gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n211), .A2(new_n212), .A3(G134gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n207), .A2(new_n208), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n204), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT74), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XOR2_X1   g016(.A(G141gat), .B(G148gat), .Z(new_n218));
  INV_X1    g017(.A(G155gat), .ZN(new_n219));
  INV_X1    g018(.A(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(KEYINPUT2), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n218), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g021(.A(G155gat), .B(G162gat), .ZN(new_n223));
  XNOR2_X1  g022(.A(new_n222), .B(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n212), .A2(G134gat), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n202), .A2(new_n203), .A3(new_n206), .A4(new_n225), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n217), .A2(new_n224), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT4), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT4), .ZN(new_n229));
  NAND4_X1  g028(.A1(new_n217), .A2(new_n229), .A3(new_n224), .A4(new_n226), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(KEYINPUT84), .A3(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n224), .B(KEYINPUT3), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n217), .A2(new_n226), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT84), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n227), .A2(new_n235), .A3(KEYINPUT4), .ZN(new_n236));
  NAND2_X1  g035(.A1(G225gat), .A2(G233gat), .ZN(new_n237));
  XOR2_X1   g036(.A(new_n237), .B(KEYINPUT83), .Z(new_n238));
  NOR2_X1   g037(.A1(new_n238), .A2(KEYINPUT5), .ZN(new_n239));
  NAND4_X1  g038(.A1(new_n231), .A2(new_n234), .A3(new_n236), .A4(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n233), .B(new_n224), .ZN(new_n241));
  INV_X1    g040(.A(new_n238), .ZN(new_n242));
  OAI21_X1  g041(.A(KEYINPUT5), .B1(new_n241), .B2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n228), .A2(new_n230), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n238), .B1(new_n232), .B2(new_n233), .ZN(new_n245));
  AND2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n240), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(G1gat), .B(G29gat), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n248), .B(KEYINPUT0), .ZN(new_n249));
  XNOR2_X1  g048(.A(G57gat), .B(G85gat), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n249), .B(new_n250), .Z(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n247), .A2(KEYINPUT6), .A3(new_n252), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT85), .ZN(new_n254));
  XNOR2_X1  g053(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT6), .ZN(new_n256));
  OAI21_X1  g055(.A(new_n256), .B1(new_n247), .B2(new_n252), .ZN(new_n257));
  INV_X1    g056(.A(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n247), .A2(new_n252), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XOR2_X1   g059(.A(G8gat), .B(G36gat), .Z(new_n261));
  XNOR2_X1  g060(.A(new_n261), .B(KEYINPUT82), .ZN(new_n262));
  XNOR2_X1  g061(.A(G64gat), .B(G92gat), .ZN(new_n263));
  XOR2_X1   g062(.A(new_n262), .B(new_n263), .Z(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(G197gat), .B(G204gat), .ZN(new_n266));
  INV_X1    g065(.A(G211gat), .ZN(new_n267));
  INV_X1    g066(.A(G218gat), .ZN(new_n268));
  OAI22_X1  g067(.A1(new_n267), .A2(new_n268), .B1(KEYINPUT79), .B2(KEYINPUT22), .ZN(new_n269));
  AND2_X1   g068(.A1(KEYINPUT79), .A2(KEYINPUT22), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  XOR2_X1   g070(.A(G211gat), .B(G218gat), .Z(new_n272));
  XNOR2_X1  g071(.A(new_n271), .B(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  XOR2_X1   g073(.A(KEYINPUT27), .B(G183gat), .Z(new_n275));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n276));
  NOR3_X1   g075(.A1(new_n275), .A2(new_n276), .A3(G190gat), .ZN(new_n277));
  INV_X1    g076(.A(G190gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT27), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  OAI21_X1  g080(.A(G183gat), .B1(KEYINPUT69), .B2(KEYINPUT27), .ZN(new_n282));
  XOR2_X1   g081(.A(KEYINPUT68), .B(G183gat), .Z(new_n283));
  OAI221_X1 g082(.A(new_n278), .B1(new_n281), .B2(new_n282), .C1(new_n283), .C2(new_n280), .ZN(new_n284));
  AOI21_X1  g083(.A(new_n277), .B1(new_n284), .B2(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(G169gat), .A2(G176gat), .ZN(new_n286));
  INV_X1    g085(.A(new_n286), .ZN(new_n287));
  NOR2_X1   g086(.A1(G169gat), .A2(G176gat), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT70), .ZN(new_n289));
  AOI21_X1  g088(.A(new_n287), .B1(new_n289), .B2(KEYINPUT26), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n290), .B1(KEYINPUT26), .B2(new_n289), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT71), .ZN(new_n292));
  NAND2_X1  g091(.A1(G183gat), .A2(G190gat), .ZN(new_n293));
  AND3_X1   g092(.A1(new_n291), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n292), .B1(new_n291), .B2(new_n293), .ZN(new_n295));
  OR3_X1    g094(.A1(new_n285), .A2(new_n294), .A3(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT23), .ZN(new_n297));
  XNOR2_X1  g096(.A(new_n288), .B(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n286), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n299), .A2(KEYINPUT65), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT65), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n298), .A2(new_n301), .A3(new_n286), .ZN(new_n302));
  NAND3_X1  g101(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT64), .ZN(new_n304));
  OR2_X1    g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n303), .A2(new_n304), .ZN(new_n306));
  OR2_X1    g105(.A1(G183gat), .A2(G190gat), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT24), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n293), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g108(.A1(new_n305), .A2(new_n306), .A3(new_n307), .A4(new_n309), .ZN(new_n310));
  NAND3_X1  g109(.A1(new_n300), .A2(new_n302), .A3(new_n310), .ZN(new_n311));
  INV_X1    g110(.A(KEYINPUT25), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT66), .ZN(new_n314));
  OAI21_X1  g113(.A(KEYINPUT25), .B1(new_n286), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n314), .B2(new_n286), .ZN(new_n316));
  AND2_X1   g115(.A1(new_n316), .A2(new_n298), .ZN(new_n317));
  XNOR2_X1  g116(.A(new_n303), .B(KEYINPUT67), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n318), .B(new_n309), .C1(G190gat), .C2(new_n283), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n313), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n296), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(G226gat), .A2(G233gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n323), .B(KEYINPUT80), .ZN(new_n324));
  AOI21_X1  g123(.A(KEYINPUT81), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  NOR3_X1   g124(.A1(new_n285), .A2(new_n294), .A3(new_n295), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n311), .A2(new_n312), .B1(new_n317), .B2(new_n319), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT29), .B1(new_n296), .B2(new_n321), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n328), .B1(new_n329), .B2(new_n324), .ZN(new_n330));
  AOI211_X1 g129(.A(new_n274), .B(new_n325), .C1(new_n330), .C2(KEYINPUT81), .ZN(new_n331));
  INV_X1    g130(.A(new_n328), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT29), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n322), .A2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(new_n324), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n332), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n336), .A2(new_n273), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n265), .B1(new_n331), .B2(new_n337), .ZN(new_n338));
  INV_X1    g137(.A(new_n337), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n325), .B1(new_n330), .B2(KEYINPUT81), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n273), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n339), .A2(new_n341), .A3(new_n264), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n338), .A2(new_n342), .A3(KEYINPUT30), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n337), .B1(new_n273), .B2(new_n340), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT30), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n345), .A3(new_n264), .ZN(new_n346));
  AOI22_X1  g145(.A1(new_n255), .A2(new_n260), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(new_n224), .ZN(new_n348));
  OAI21_X1  g147(.A(new_n333), .B1(new_n348), .B2(KEYINPUT3), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n349), .A2(new_n274), .ZN(new_n350));
  OR2_X1    g149(.A1(new_n273), .A2(KEYINPUT86), .ZN(new_n351));
  AND2_X1   g150(.A1(new_n271), .A2(new_n272), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT29), .B1(new_n352), .B2(KEYINPUT86), .ZN(new_n353));
  AOI21_X1  g152(.A(KEYINPUT3), .B1(new_n351), .B2(new_n353), .ZN(new_n354));
  OAI21_X1  g153(.A(new_n350), .B1(new_n354), .B2(new_n224), .ZN(new_n355));
  NAND2_X1  g154(.A1(G228gat), .A2(G233gat), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n356), .B1(new_n349), .B2(new_n274), .ZN(new_n357));
  NOR2_X1   g156(.A1(new_n274), .A2(KEYINPUT29), .ZN(new_n358));
  OAI21_X1  g157(.A(new_n348), .B1(new_n358), .B2(KEYINPUT3), .ZN(new_n359));
  AOI22_X1  g158(.A1(new_n355), .A2(new_n356), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g159(.A(G22gat), .ZN(new_n361));
  OR2_X1    g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n360), .A2(new_n361), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT87), .ZN(new_n365));
  AOI21_X1  g164(.A(new_n365), .B1(new_n360), .B2(new_n361), .ZN(new_n366));
  XOR2_X1   g165(.A(G78gat), .B(G106gat), .Z(new_n367));
  XNOR2_X1  g166(.A(KEYINPUT31), .B(G50gat), .ZN(new_n368));
  XNOR2_X1  g167(.A(new_n367), .B(new_n368), .ZN(new_n369));
  OAI21_X1  g168(.A(KEYINPUT88), .B1(new_n366), .B2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n366), .A2(KEYINPUT88), .A3(new_n369), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n364), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n369), .B1(new_n363), .B2(KEYINPUT87), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  NAND4_X1  g175(.A1(new_n376), .A2(new_n363), .A3(new_n362), .A4(new_n370), .ZN(new_n377));
  AND2_X1   g176(.A1(new_n373), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g177(.A(new_n217), .B(new_n226), .C1(new_n326), .C2(new_n327), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n296), .A2(new_n233), .A3(new_n321), .ZN(new_n380));
  NAND4_X1  g179(.A1(new_n379), .A2(new_n380), .A3(G227gat), .A4(G233gat), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT33), .ZN(new_n382));
  XOR2_X1   g181(.A(G15gat), .B(G43gat), .Z(new_n383));
  XNOR2_X1  g182(.A(G71gat), .B(G99gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n383), .B(new_n384), .ZN(new_n385));
  XNOR2_X1  g184(.A(KEYINPUT75), .B(KEYINPUT76), .ZN(new_n386));
  XNOR2_X1  g185(.A(new_n385), .B(new_n386), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n381), .B(KEYINPUT32), .C1(new_n382), .C2(new_n387), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n387), .B1(new_n381), .B2(KEYINPUT32), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT77), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n381), .A2(new_n382), .ZN(new_n391));
  AND3_X1   g190(.A1(new_n389), .A2(new_n390), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n390), .B1(new_n389), .B2(new_n391), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n388), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT34), .ZN(new_n395));
  AND2_X1   g194(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n396));
  NOR2_X1   g195(.A1(new_n395), .A2(KEYINPUT78), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n379), .A2(new_n380), .ZN(new_n398));
  NAND2_X1  g197(.A1(G227gat), .A2(G233gat), .ZN(new_n399));
  AOI211_X1 g198(.A(new_n396), .B(new_n397), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n398), .A2(new_n399), .A3(new_n397), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n394), .A2(new_n402), .ZN(new_n403));
  OAI221_X1 g202(.A(new_n388), .B1(new_n400), .B2(new_n401), .C1(new_n392), .C2(new_n393), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n347), .A2(new_n378), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(KEYINPUT35), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n373), .A2(new_n403), .A3(new_n377), .A4(new_n404), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n343), .A2(new_n346), .ZN(new_n409));
  OR3_X1    g208(.A1(new_n408), .A2(KEYINPUT35), .A3(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n255), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n251), .B1(new_n247), .B2(KEYINPUT91), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT92), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT91), .ZN(new_n414));
  OAI211_X1 g213(.A(new_n414), .B(new_n240), .C1(new_n243), .C2(new_n246), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n412), .A2(new_n413), .A3(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n412), .B2(new_n415), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n258), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT93), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n247), .A2(KEYINPUT91), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n421), .A2(new_n252), .A3(new_n415), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n422), .A2(KEYINPUT92), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(new_n416), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT93), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n424), .A2(new_n425), .A3(new_n258), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n411), .B1(new_n420), .B2(new_n426), .ZN(new_n427));
  OAI21_X1  g226(.A(new_n407), .B1(new_n410), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n231), .A2(new_n234), .A3(new_n236), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n238), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n241), .A2(new_n242), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT39), .A3(new_n431), .ZN(new_n432));
  XNOR2_X1  g231(.A(KEYINPUT89), .B(KEYINPUT39), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n238), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n251), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g234(.A1(KEYINPUT90), .A2(KEYINPUT40), .ZN(new_n436));
  INV_X1    g235(.A(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(new_n435), .B(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n438), .A2(new_n424), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n343), .A2(new_n346), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n378), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n339), .A2(new_n341), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n265), .B1(new_n442), .B2(KEYINPUT37), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT38), .ZN(new_n444));
  AND2_X1   g243(.A1(new_n340), .A2(new_n274), .ZN(new_n445));
  OAI21_X1  g244(.A(KEYINPUT37), .B1(new_n336), .B2(new_n274), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n444), .B1(new_n445), .B2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n342), .B1(new_n443), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT37), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n264), .B1(new_n344), .B2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n442), .A2(KEYINPUT37), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n444), .B1(new_n450), .B2(new_n451), .ZN(new_n452));
  NOR2_X1   g251(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n441), .B1(new_n427), .B2(new_n453), .ZN(new_n454));
  AND3_X1   g253(.A1(new_n403), .A2(new_n404), .A3(KEYINPUT36), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT36), .B1(new_n403), .B2(new_n404), .ZN(new_n456));
  OAI22_X1  g255(.A1(new_n455), .A2(new_n456), .B1(new_n347), .B2(new_n378), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n428), .B1(new_n454), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT98), .ZN(new_n459));
  AND2_X1   g258(.A1(G43gat), .A2(G50gat), .ZN(new_n460));
  NOR2_X1   g259(.A1(G43gat), .A2(G50gat), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT15), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  NOR3_X1   g261(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n463));
  OAI21_X1  g262(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n464));
  AOI21_X1  g263(.A(new_n463), .B1(KEYINPUT94), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n465), .B1(KEYINPUT94), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g265(.A1(G29gat), .A2(G36gat), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n462), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n464), .ZN(new_n469));
  OAI211_X1 g268(.A(new_n462), .B(new_n467), .C1(new_n469), .C2(new_n463), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT15), .ZN(new_n471));
  XOR2_X1   g270(.A(KEYINPUT95), .B(G43gat), .Z(new_n472));
  XNOR2_X1  g271(.A(KEYINPUT96), .B(G50gat), .ZN(new_n473));
  OAI22_X1  g272(.A1(new_n472), .A2(G50gat), .B1(new_n473), .B2(G43gat), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n470), .B1(new_n471), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g274(.A1(new_n468), .A2(new_n475), .ZN(new_n476));
  INV_X1    g275(.A(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(G15gat), .B(G22gat), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT16), .ZN(new_n479));
  OAI21_X1  g278(.A(new_n478), .B1(new_n479), .B2(G1gat), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n480), .B1(G1gat), .B2(new_n478), .ZN(new_n481));
  XNOR2_X1  g280(.A(new_n481), .B(G8gat), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n459), .B1(new_n477), .B2(new_n482), .ZN(new_n483));
  INV_X1    g282(.A(new_n482), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n484), .A2(KEYINPUT98), .A3(new_n476), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n477), .A2(new_n482), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n483), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(G229gat), .A2(G233gat), .ZN(new_n488));
  XOR2_X1   g287(.A(new_n488), .B(KEYINPUT13), .Z(new_n489));
  NAND2_X1  g288(.A1(new_n487), .A2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT99), .ZN(new_n491));
  XNOR2_X1  g290(.A(new_n490), .B(new_n491), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n482), .B(KEYINPUT97), .ZN(new_n493));
  INV_X1    g292(.A(KEYINPUT17), .ZN(new_n494));
  NOR2_X1   g293(.A1(new_n476), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n477), .A2(KEYINPUT17), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NAND3_X1  g296(.A1(new_n497), .A2(new_n488), .A3(new_n486), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT18), .ZN(new_n499));
  OR2_X1    g298(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n498), .A2(new_n499), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n492), .A2(new_n500), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G113gat), .B(G141gat), .ZN(new_n503));
  XNOR2_X1  g302(.A(new_n503), .B(G197gat), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT11), .B(G169gat), .Z(new_n505));
  XNOR2_X1  g304(.A(new_n504), .B(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(new_n506), .B(KEYINPUT12), .Z(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(new_n507), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n492), .A2(new_n500), .A3(new_n509), .A4(new_n501), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  AND3_X1   g310(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n512));
  INV_X1    g311(.A(G92gat), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT101), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT101), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(G92gat), .ZN(new_n516));
  INV_X1    g315(.A(G85gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n514), .A2(new_n516), .A3(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G85gat), .A2(G92gat), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(KEYINPUT7), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT7), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n521), .A2(G85gat), .A3(G92gat), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(G99gat), .ZN(new_n524));
  INV_X1    g323(.A(G106gat), .ZN(new_n525));
  OAI21_X1  g324(.A(KEYINPUT8), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n518), .A2(new_n523), .A3(new_n526), .ZN(new_n527));
  XNOR2_X1  g326(.A(G99gat), .B(G106gat), .ZN(new_n528));
  INV_X1    g327(.A(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(new_n529), .ZN(new_n530));
  NAND4_X1  g329(.A1(new_n518), .A2(new_n523), .A3(new_n528), .A4(new_n526), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n530), .A2(KEYINPUT102), .A3(new_n531), .ZN(new_n532));
  OR3_X1    g331(.A1(new_n527), .A2(KEYINPUT102), .A3(new_n529), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n512), .B1(new_n477), .B2(new_n534), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n496), .A2(new_n495), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n535), .B1(new_n536), .B2(new_n534), .ZN(new_n537));
  XOR2_X1   g336(.A(G190gat), .B(G218gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(new_n538), .B(new_n535), .C1(new_n536), .C2(new_n534), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT103), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT104), .ZN(new_n544));
  XNOR2_X1  g343(.A(G134gat), .B(G162gat), .ZN(new_n545));
  AOI21_X1  g344(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n543), .A2(new_n544), .A3(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n544), .B1(new_n543), .B2(new_n547), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n540), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n550), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n552), .A2(new_n539), .A3(new_n548), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  XNOR2_X1  g353(.A(G57gat), .B(G64gat), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OR2_X1    g355(.A1(G71gat), .A2(G78gat), .ZN(new_n557));
  NAND2_X1  g356(.A1(G71gat), .A2(G78gat), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n558), .A2(new_n560), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n559), .A3(new_n561), .ZN(new_n562));
  OAI211_X1 g361(.A(new_n558), .B(new_n557), .C1(new_n555), .C2(new_n560), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(KEYINPUT100), .B(KEYINPUT21), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(G231gat), .A2(G233gat), .ZN(new_n567));
  XNOR2_X1  g366(.A(new_n566), .B(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G127gat), .ZN(new_n569));
  INV_X1    g368(.A(new_n564), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n482), .B1(KEYINPUT21), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g370(.A(new_n569), .B(new_n571), .Z(new_n572));
  XNOR2_X1  g371(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(new_n219), .ZN(new_n574));
  XOR2_X1   g373(.A(G183gat), .B(G211gat), .Z(new_n575));
  XNOR2_X1  g374(.A(new_n574), .B(new_n575), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n572), .B(new_n576), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n554), .A2(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G120gat), .B(G148gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G176gat), .B(G204gat), .ZN(new_n580));
  XOR2_X1   g379(.A(new_n579), .B(new_n580), .Z(new_n581));
  INV_X1    g380(.A(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT10), .ZN(new_n583));
  AOI21_X1  g382(.A(new_n570), .B1(new_n532), .B2(new_n533), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT105), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n531), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(new_n530), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n527), .A2(new_n585), .A3(new_n529), .ZN(new_n588));
  AOI21_X1  g387(.A(new_n564), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n583), .B1(new_n584), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n564), .A2(new_n583), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n534), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n590), .A2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(G230gat), .A2(G233gat), .ZN(new_n594));
  AOI21_X1  g393(.A(KEYINPUT106), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT106), .ZN(new_n596));
  INV_X1    g395(.A(new_n594), .ZN(new_n597));
  AOI211_X1 g396(.A(new_n596), .B(new_n597), .C1(new_n590), .C2(new_n592), .ZN(new_n598));
  NOR2_X1   g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n534), .A2(new_n564), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n587), .A2(new_n588), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n601), .A2(new_n570), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n600), .A2(new_n602), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n603), .A2(new_n594), .ZN(new_n604));
  OAI21_X1  g403(.A(new_n582), .B1(new_n599), .B2(new_n604), .ZN(new_n605));
  AOI21_X1  g404(.A(KEYINPUT10), .B1(new_n600), .B2(new_n602), .ZN(new_n606));
  INV_X1    g405(.A(new_n592), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n594), .B1(new_n606), .B2(new_n607), .ZN(new_n608));
  OAI211_X1 g407(.A(new_n608), .B(new_n581), .C1(new_n594), .C2(new_n603), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n605), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n578), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT107), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n615), .A2(KEYINPUT107), .ZN(new_n616));
  NAND4_X1  g415(.A1(new_n458), .A2(new_n511), .A3(new_n614), .A4(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n255), .A2(new_n260), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n619), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g419(.A1(new_n617), .A2(new_n440), .ZN(new_n621));
  XNOR2_X1  g420(.A(KEYINPUT108), .B(KEYINPUT16), .ZN(new_n622));
  INV_X1    g421(.A(G8gat), .ZN(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n625), .B1(new_n623), .B2(new_n621), .ZN(new_n626));
  MUX2_X1   g425(.A(new_n625), .B(new_n626), .S(KEYINPUT42), .Z(G1325gat));
  NOR2_X1   g426(.A1(new_n455), .A2(new_n456), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  OAI21_X1  g428(.A(G15gat), .B1(new_n617), .B2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n403), .A2(new_n404), .ZN(new_n631));
  OR2_X1    g430(.A1(new_n631), .A2(G15gat), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n617), .B2(new_n632), .ZN(G1326gat));
  NOR2_X1   g432(.A1(new_n617), .A2(new_n378), .ZN(new_n634));
  XOR2_X1   g433(.A(KEYINPUT43), .B(G22gat), .Z(new_n635));
  XNOR2_X1  g434(.A(new_n634), .B(new_n635), .ZN(G1327gat));
  AOI21_X1  g435(.A(new_n425), .B1(new_n424), .B2(new_n258), .ZN(new_n637));
  AOI211_X1 g436(.A(KEYINPUT93), .B(new_n257), .C1(new_n423), .C2(new_n416), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n453), .B(new_n255), .C1(new_n637), .C2(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n441), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n457), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(new_n255), .B1(new_n637), .B2(new_n638), .ZN(new_n642));
  NOR3_X1   g441(.A1(new_n408), .A2(KEYINPUT35), .A3(new_n409), .ZN(new_n643));
  AOI22_X1  g442(.A1(new_n642), .A2(new_n643), .B1(new_n406), .B2(KEYINPUT35), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n554), .B1(new_n641), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n511), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n577), .A2(new_n611), .ZN(new_n648));
  NOR2_X1   g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n650), .A2(G29gat), .A3(new_n618), .ZN(new_n651));
  XOR2_X1   g450(.A(new_n651), .B(KEYINPUT45), .Z(new_n652));
  INV_X1    g451(.A(KEYINPUT44), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n645), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT44), .B(new_n554), .C1(new_n641), .C2(new_n644), .ZN(new_n655));
  AND2_X1   g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n656), .A2(new_n649), .ZN(new_n657));
  OAI21_X1  g456(.A(G29gat), .B1(new_n657), .B2(new_n618), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n652), .A2(new_n658), .ZN(G1328gat));
  OAI21_X1  g458(.A(G36gat), .B1(new_n657), .B2(new_n440), .ZN(new_n660));
  INV_X1    g459(.A(new_n554), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT46), .ZN(new_n662));
  NOR2_X1   g461(.A1(new_n662), .A2(KEYINPUT109), .ZN(new_n663));
  NOR4_X1   g462(.A1(new_n661), .A2(G36gat), .A3(new_n648), .A4(new_n663), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n458), .A2(new_n409), .A3(new_n511), .A4(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n662), .A2(KEYINPUT109), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n665), .B(new_n666), .Z(new_n667));
  NAND2_X1  g466(.A1(new_n660), .A2(new_n667), .ZN(G1329gat));
  NAND4_X1  g467(.A1(new_n654), .A2(new_n628), .A3(new_n649), .A4(new_n655), .ZN(new_n669));
  INV_X1    g468(.A(new_n472), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n631), .A2(new_n670), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n646), .A2(new_n649), .A3(new_n672), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n671), .A2(KEYINPUT47), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g473(.A1(new_n671), .A2(KEYINPUT111), .ZN(new_n675));
  INV_X1    g474(.A(KEYINPUT112), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g476(.A1(new_n646), .A2(KEYINPUT112), .A3(new_n649), .A4(new_n672), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT111), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n669), .B2(new_n670), .ZN(new_n681));
  NOR3_X1   g480(.A1(new_n675), .A2(new_n679), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g481(.A(KEYINPUT110), .B(KEYINPUT47), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n674), .B1(new_n682), .B2(new_n683), .ZN(G1330gat));
  OAI21_X1  g483(.A(new_n473), .B1(new_n650), .B2(new_n378), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n378), .A2(new_n473), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(new_n685), .B1(new_n657), .B2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n688), .B(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g488(.A1(new_n458), .A2(new_n647), .A3(new_n578), .A4(new_n610), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(new_n618), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g493(.A(new_n440), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT113), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n691), .A2(new_n696), .ZN(new_n697));
  OR2_X1    g496(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n698));
  NOR2_X1   g497(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(KEYINPUT114), .ZN(new_n700));
  AND3_X1   g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  AOI21_X1  g500(.A(new_n699), .B1(new_n698), .B2(new_n700), .ZN(new_n702));
  NOR2_X1   g501(.A1(new_n701), .A2(new_n702), .ZN(G1333gat));
  OR3_X1    g502(.A1(new_n690), .A2(G71gat), .A3(new_n631), .ZN(new_n704));
  OAI21_X1  g503(.A(G71gat), .B1(new_n690), .B2(new_n629), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  XOR2_X1   g505(.A(new_n706), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g506(.A1(new_n373), .A2(new_n377), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n691), .A2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(new_n709), .B(G78gat), .ZN(G1335gat));
  INV_X1    g509(.A(new_n577), .ZN(new_n711));
  NOR3_X1   g510(.A1(new_n711), .A2(new_n511), .A3(new_n611), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n656), .A2(new_n712), .ZN(new_n713));
  OAI21_X1  g512(.A(G85gat), .B1(new_n713), .B2(new_n618), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n711), .A2(new_n511), .ZN(new_n715));
  OAI211_X1 g514(.A(new_n554), .B(new_n715), .C1(new_n641), .C2(new_n644), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT51), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n458), .A2(KEYINPUT51), .A3(new_n554), .A4(new_n715), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n692), .A2(new_n517), .A3(new_n610), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n714), .B1(new_n721), .B2(new_n722), .ZN(G1336gat));
  NAND4_X1  g522(.A1(new_n654), .A2(new_n409), .A3(new_n655), .A4(new_n712), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n514), .A2(new_n516), .ZN(new_n725));
  NAND2_X1  g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n440), .A2(new_n611), .A3(G92gat), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n720), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT115), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n716), .A2(new_n731), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n732), .A2(new_n717), .ZN(new_n733));
  NAND3_X1  g532(.A1(new_n716), .A2(new_n731), .A3(KEYINPUT51), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n733), .A2(new_n734), .A3(new_n727), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n729), .B1(new_n735), .B2(new_n726), .ZN(new_n736));
  OAI21_X1  g535(.A(KEYINPUT116), .B1(new_n730), .B2(new_n736), .ZN(new_n737));
  INV_X1    g536(.A(KEYINPUT116), .ZN(new_n738));
  NAND3_X1  g537(.A1(new_n726), .A2(new_n728), .A3(new_n729), .ZN(new_n739));
  AND3_X1   g538(.A1(new_n716), .A2(new_n731), .A3(KEYINPUT51), .ZN(new_n740));
  AOI21_X1  g539(.A(KEYINPUT51), .B1(new_n716), .B2(new_n731), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  AOI22_X1  g541(.A1(new_n742), .A2(new_n727), .B1(new_n725), .B2(new_n724), .ZN(new_n743));
  OAI211_X1 g542(.A(new_n738), .B(new_n739), .C1(new_n743), .C2(new_n729), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(G1337gat));
  OAI21_X1  g544(.A(G99gat), .B1(new_n713), .B2(new_n629), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n405), .A2(new_n524), .A3(new_n610), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n746), .B1(new_n721), .B2(new_n747), .ZN(G1338gat));
  NAND4_X1  g547(.A1(new_n654), .A2(new_n708), .A3(new_n655), .A4(new_n712), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n749), .A2(G106gat), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT117), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n378), .A2(G106gat), .A3(new_n611), .ZN(new_n753));
  AOI21_X1  g552(.A(new_n752), .B1(new_n720), .B2(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n753), .ZN(new_n755));
  NOR3_X1   g554(.A1(new_n721), .A2(KEYINPUT117), .A3(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n751), .B1(new_n754), .B2(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n740), .A2(new_n741), .A3(new_n755), .ZN(new_n758));
  OAI21_X1  g557(.A(KEYINPUT53), .B1(new_n750), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n757), .A2(new_n759), .ZN(G1339gat));
  INV_X1    g559(.A(G113gat), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n607), .B1(new_n603), .B2(new_n583), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n596), .B1(new_n762), .B2(new_n597), .ZN(new_n763));
  INV_X1    g562(.A(KEYINPUT54), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n593), .A2(KEYINPUT106), .A3(new_n594), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n763), .A2(new_n764), .A3(new_n765), .ZN(new_n766));
  AOI21_X1  g565(.A(new_n764), .B1(new_n593), .B2(new_n594), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n590), .A2(new_n597), .A3(new_n592), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n581), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n766), .A2(new_n769), .A3(KEYINPUT55), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(new_n609), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT55), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n595), .A2(new_n598), .A3(KEYINPUT54), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n608), .A2(KEYINPUT54), .A3(new_n768), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n582), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n772), .B1(new_n773), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n511), .A2(new_n771), .A3(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n488), .B1(new_n497), .B2(new_n486), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n487), .A2(new_n489), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n506), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n780), .A2(KEYINPUT118), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(KEYINPUT118), .ZN(new_n782));
  AND3_X1   g581(.A1(new_n781), .A2(new_n510), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n610), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n554), .B1(new_n777), .B2(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n554), .A2(new_n783), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n771), .A2(new_n776), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  OAI21_X1  g587(.A(new_n577), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n615), .A2(new_n647), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n708), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n692), .A2(new_n440), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n792), .A2(new_n631), .ZN(new_n793));
  AND2_X1   g592(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n761), .B1(new_n794), .B2(new_n511), .ZN(new_n795));
  XOR2_X1   g594(.A(new_n795), .B(KEYINPUT119), .Z(new_n796));
  AOI21_X1  g595(.A(new_n618), .B1(new_n789), .B2(new_n790), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n408), .A2(new_n409), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n800), .A2(new_n761), .A3(new_n511), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n796), .A2(new_n801), .ZN(G1340gat));
  AOI21_X1  g601(.A(G120gat), .B1(new_n800), .B2(new_n610), .ZN(new_n803));
  AND2_X1   g602(.A1(new_n610), .A2(G120gat), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n803), .B1(new_n794), .B2(new_n804), .ZN(G1341gat));
  INV_X1    g604(.A(new_n794), .ZN(new_n806));
  OAI21_X1  g605(.A(G127gat), .B1(new_n806), .B2(new_n577), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n800), .A2(new_n212), .A3(new_n711), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(G1342gat));
  NOR3_X1   g608(.A1(new_n799), .A2(G134gat), .A3(new_n661), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n811), .A2(KEYINPUT56), .ZN(new_n812));
  OAI21_X1  g611(.A(G134gat), .B1(new_n806), .B2(new_n661), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n811), .A2(KEYINPUT56), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n812), .A2(new_n813), .A3(new_n814), .ZN(G1343gat));
  NOR3_X1   g614(.A1(new_n628), .A2(new_n378), .A3(new_n409), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n797), .A2(new_n816), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n817), .A2(G141gat), .A3(new_n647), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n628), .A2(new_n792), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n789), .A2(new_n790), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n820), .A2(new_n708), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n821), .B2(KEYINPUT57), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n766), .A2(new_n769), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n823), .B1(new_n824), .B2(new_n772), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT120), .B(KEYINPUT55), .C1(new_n766), .C2(new_n769), .ZN(new_n826));
  OAI211_X1 g625(.A(new_n771), .B(KEYINPUT121), .C1(new_n825), .C2(new_n826), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(new_n511), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n776), .A2(KEYINPUT120), .ZN(new_n829));
  NAND3_X1  g628(.A1(new_n824), .A2(new_n823), .A3(new_n772), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI21_X1  g630(.A(KEYINPUT121), .B1(new_n831), .B2(new_n771), .ZN(new_n832));
  OAI21_X1  g631(.A(new_n784), .B1(new_n828), .B2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(KEYINPUT122), .ZN(new_n834));
  INV_X1    g633(.A(KEYINPUT122), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n835), .B(new_n784), .C1(new_n828), .C2(new_n832), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n834), .A2(new_n661), .A3(new_n836), .ZN(new_n837));
  INV_X1    g636(.A(new_n788), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n711), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  INV_X1    g638(.A(new_n790), .ZN(new_n840));
  OAI21_X1  g639(.A(new_n708), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  AOI21_X1  g640(.A(new_n822), .B1(new_n841), .B2(KEYINPUT57), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n511), .ZN(new_n843));
  AOI21_X1  g642(.A(new_n818), .B1(new_n843), .B2(G141gat), .ZN(new_n844));
  XOR2_X1   g643(.A(KEYINPUT123), .B(KEYINPUT58), .Z(new_n845));
  XNOR2_X1  g644(.A(new_n844), .B(new_n845), .ZN(G1344gat));
  INV_X1    g645(.A(new_n817), .ZN(new_n847));
  INV_X1    g646(.A(G148gat), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n847), .A2(new_n848), .A3(new_n610), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT59), .ZN(new_n850));
  NOR2_X1   g649(.A1(new_n378), .A2(KEYINPUT57), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n616), .A2(new_n647), .A3(new_n614), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n839), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n821), .A2(KEYINPUT57), .ZN(new_n854));
  AND2_X1   g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n855), .A2(new_n610), .A3(new_n819), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n850), .B1(new_n856), .B2(G148gat), .ZN(new_n857));
  AOI211_X1 g656(.A(KEYINPUT59), .B(new_n848), .C1(new_n842), .C2(new_n610), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n849), .B1(new_n857), .B2(new_n858), .ZN(G1345gat));
  NAND3_X1  g658(.A1(new_n847), .A2(new_n219), .A3(new_n711), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n842), .A2(new_n711), .ZN(new_n861));
  OAI21_X1  g660(.A(new_n860), .B1(new_n861), .B2(new_n219), .ZN(G1346gat));
  AOI21_X1  g661(.A(G162gat), .B1(new_n847), .B2(new_n554), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n661), .A2(new_n220), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n863), .B1(new_n842), .B2(new_n864), .ZN(G1347gat));
  AOI21_X1  g664(.A(new_n692), .B1(new_n789), .B2(new_n790), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n408), .A2(new_n440), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(G169gat), .B1(new_n869), .B2(new_n511), .ZN(new_n870));
  AND4_X1   g669(.A1(new_n618), .A2(new_n791), .A3(new_n409), .A4(new_n405), .ZN(new_n871));
  AND2_X1   g670(.A1(new_n511), .A2(G169gat), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n870), .B1(new_n871), .B2(new_n872), .ZN(G1348gat));
  NAND3_X1  g672(.A1(new_n871), .A2(G176gat), .A3(new_n610), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n875));
  NOR2_X1   g674(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n876));
  AOI21_X1  g675(.A(G176gat), .B1(new_n869), .B2(new_n610), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(G1349gat));
  NOR3_X1   g677(.A1(new_n868), .A2(new_n275), .A3(new_n577), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n871), .A2(new_n711), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(new_n880), .B2(new_n283), .ZN(new_n881));
  XOR2_X1   g680(.A(new_n881), .B(KEYINPUT60), .Z(G1350gat));
  AOI21_X1  g681(.A(new_n278), .B1(new_n871), .B2(new_n554), .ZN(new_n883));
  XOR2_X1   g682(.A(new_n883), .B(KEYINPUT61), .Z(new_n884));
  NAND3_X1  g683(.A1(new_n869), .A2(new_n278), .A3(new_n554), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(G1351gat));
  NOR3_X1   g685(.A1(new_n628), .A2(new_n692), .A3(new_n440), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n855), .A2(new_n887), .ZN(new_n888));
  INV_X1    g687(.A(G197gat), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n888), .A2(new_n889), .A3(new_n647), .ZN(new_n890));
  NOR3_X1   g689(.A1(new_n628), .A2(new_n378), .A3(new_n440), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n866), .A2(new_n891), .ZN(new_n892));
  INV_X1    g691(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g692(.A(G197gat), .B1(new_n893), .B2(new_n511), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n890), .A2(new_n894), .ZN(G1352gat));
  NAND4_X1  g694(.A1(new_n853), .A2(new_n610), .A3(new_n854), .A4(new_n887), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n896), .A2(G204gat), .ZN(new_n897));
  NOR2_X1   g696(.A1(new_n611), .A2(G204gat), .ZN(new_n898));
  INV_X1    g697(.A(new_n898), .ZN(new_n899));
  OAI21_X1  g698(.A(KEYINPUT125), .B1(new_n892), .B2(new_n899), .ZN(new_n900));
  INV_X1    g699(.A(KEYINPUT125), .ZN(new_n901));
  NAND4_X1  g700(.A1(new_n866), .A2(new_n901), .A3(new_n891), .A4(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT62), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n900), .A2(KEYINPUT62), .A3(new_n902), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n897), .A2(new_n905), .A3(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT126), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n907), .B(new_n908), .ZN(G1353gat));
  NAND3_X1  g708(.A1(new_n893), .A2(new_n267), .A3(new_n711), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n853), .A2(new_n711), .A3(new_n854), .A4(new_n887), .ZN(new_n911));
  AND3_X1   g710(.A1(new_n911), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n912));
  AOI21_X1  g711(.A(KEYINPUT63), .B1(new_n911), .B2(G211gat), .ZN(new_n913));
  OAI21_X1  g712(.A(new_n910), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n914), .A2(KEYINPUT127), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT127), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n916), .B(new_n910), .C1(new_n912), .C2(new_n913), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n915), .A2(new_n917), .ZN(G1354gat));
  OAI21_X1  g717(.A(G218gat), .B1(new_n888), .B2(new_n661), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n893), .A2(new_n268), .A3(new_n554), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(G1355gat));
endmodule


