

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594;

  XNOR2_X1 U321 ( .A(n457), .B(n456), .ZN(n473) );
  NOR2_X1 U322 ( .A1(n557), .A2(n401), .ZN(n544) );
  XNOR2_X1 U323 ( .A(n415), .B(KEYINPUT37), .ZN(n416) );
  XNOR2_X1 U324 ( .A(n332), .B(n331), .ZN(n572) );
  INV_X1 U325 ( .A(n558), .ZN(n559) );
  XNOR2_X1 U326 ( .A(n399), .B(n398), .ZN(n532) );
  XNOR2_X1 U327 ( .A(n442), .B(G204GAT), .ZN(n443) );
  INV_X1 U328 ( .A(KEYINPUT65), .ZN(n312) );
  INV_X1 U329 ( .A(KEYINPUT100), .ZN(n389) );
  XNOR2_X1 U330 ( .A(n444), .B(n443), .ZN(n448) );
  XNOR2_X1 U331 ( .A(n313), .B(n312), .ZN(n314) );
  XNOR2_X1 U332 ( .A(n390), .B(n389), .ZN(n391) );
  NOR2_X1 U333 ( .A1(n579), .A2(n482), .ZN(n484) );
  XNOR2_X1 U334 ( .A(n315), .B(n314), .ZN(n316) );
  INV_X1 U335 ( .A(KEYINPUT112), .ZN(n415) );
  XNOR2_X1 U336 ( .A(n392), .B(n391), .ZN(n395) );
  XNOR2_X1 U337 ( .A(n330), .B(n457), .ZN(n331) );
  XNOR2_X1 U338 ( .A(n417), .B(n416), .ZN(n528) );
  XOR2_X1 U339 ( .A(n473), .B(KEYINPUT41), .Z(n563) );
  INV_X1 U340 ( .A(G50GAT), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U342 ( .A(n459), .B(KEYINPUT114), .ZN(n460) );
  XNOR2_X1 U343 ( .A(n493), .B(n492), .ZN(G1349GAT) );
  XNOR2_X1 U344 ( .A(n461), .B(n460), .ZN(G1331GAT) );
  XOR2_X1 U345 ( .A(KEYINPUT93), .B(KEYINPUT24), .Z(n290) );
  XNOR2_X1 U346 ( .A(KEYINPUT92), .B(KEYINPUT23), .ZN(n289) );
  XNOR2_X1 U347 ( .A(n290), .B(n289), .ZN(n291) );
  XOR2_X1 U348 ( .A(KEYINPUT87), .B(n291), .Z(n293) );
  NAND2_X1 U349 ( .A1(G228GAT), .A2(G233GAT), .ZN(n292) );
  XNOR2_X1 U350 ( .A(n293), .B(n292), .ZN(n294) );
  XOR2_X1 U351 ( .A(n294), .B(KEYINPUT91), .Z(n299) );
  XOR2_X1 U352 ( .A(KEYINPUT90), .B(KEYINPUT2), .Z(n296) );
  XNOR2_X1 U353 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n295) );
  XNOR2_X1 U354 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U355 ( .A(G141GAT), .B(n297), .Z(n377) );
  XNOR2_X1 U356 ( .A(n377), .B(KEYINPUT22), .ZN(n298) );
  XNOR2_X1 U357 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U358 ( .A(G106GAT), .B(G218GAT), .Z(n301) );
  XOR2_X1 U359 ( .A(G148GAT), .B(G78GAT), .Z(n450) );
  XOR2_X1 U360 ( .A(G22GAT), .B(G155GAT), .Z(n347) );
  XNOR2_X1 U361 ( .A(n450), .B(n347), .ZN(n300) );
  XNOR2_X1 U362 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U363 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U364 ( .A(KEYINPUT88), .B(G211GAT), .Z(n305) );
  XNOR2_X1 U365 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n304) );
  XNOR2_X1 U366 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U367 ( .A(G197GAT), .B(n306), .Z(n397) );
  XOR2_X1 U368 ( .A(G50GAT), .B(G162GAT), .Z(n323) );
  XNOR2_X1 U369 ( .A(n397), .B(n323), .ZN(n307) );
  XNOR2_X1 U370 ( .A(n308), .B(n307), .ZN(n482) );
  XOR2_X1 U371 ( .A(n482), .B(KEYINPUT28), .Z(n538) );
  XNOR2_X1 U372 ( .A(KEYINPUT36), .B(KEYINPUT111), .ZN(n333) );
  XOR2_X1 U373 ( .A(KEYINPUT8), .B(KEYINPUT7), .Z(n310) );
  XNOR2_X1 U374 ( .A(G43GAT), .B(G29GAT), .ZN(n309) );
  XNOR2_X1 U375 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U376 ( .A(KEYINPUT69), .B(n311), .Z(n435) );
  INV_X1 U377 ( .A(n435), .ZN(n315) );
  XOR2_X1 U378 ( .A(KEYINPUT9), .B(KEYINPUT11), .Z(n313) );
  XOR2_X1 U379 ( .A(n316), .B(KEYINPUT80), .Z(n332) );
  XOR2_X1 U380 ( .A(KEYINPUT79), .B(G92GAT), .Z(n318) );
  XNOR2_X1 U381 ( .A(G190GAT), .B(G218GAT), .ZN(n317) );
  XNOR2_X1 U382 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U383 ( .A(G36GAT), .B(n319), .ZN(n398) );
  XOR2_X1 U384 ( .A(KEYINPUT78), .B(KEYINPUT10), .Z(n321) );
  XNOR2_X1 U385 ( .A(G134GAT), .B(KEYINPUT77), .ZN(n320) );
  XNOR2_X1 U386 ( .A(n321), .B(n320), .ZN(n322) );
  XOR2_X1 U387 ( .A(n323), .B(n322), .Z(n325) );
  NAND2_X1 U388 ( .A1(G232GAT), .A2(G233GAT), .ZN(n324) );
  XNOR2_X1 U389 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U390 ( .A(n398), .B(n326), .Z(n330) );
  XOR2_X1 U391 ( .A(KEYINPUT74), .B(KEYINPUT75), .Z(n328) );
  XNOR2_X1 U392 ( .A(G106GAT), .B(G85GAT), .ZN(n327) );
  XNOR2_X1 U393 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U394 ( .A(G99GAT), .B(n329), .ZN(n457) );
  XNOR2_X1 U395 ( .A(KEYINPUT81), .B(n572), .ZN(n553) );
  XNOR2_X1 U396 ( .A(n333), .B(n553), .ZN(n471) );
  XOR2_X1 U397 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n335) );
  XNOR2_X1 U398 ( .A(G64GAT), .B(KEYINPUT83), .ZN(n334) );
  XNOR2_X1 U399 ( .A(n335), .B(n334), .ZN(n351) );
  XOR2_X1 U400 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n337) );
  NAND2_X1 U401 ( .A1(G231GAT), .A2(G233GAT), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U403 ( .A(n338), .B(KEYINPUT12), .Z(n342) );
  XNOR2_X1 U404 ( .A(G57GAT), .B(KEYINPUT71), .ZN(n339) );
  XNOR2_X1 U405 ( .A(n339), .B(KEYINPUT13), .ZN(n439) );
  XNOR2_X1 U406 ( .A(G8GAT), .B(G183GAT), .ZN(n340) );
  XNOR2_X1 U407 ( .A(n340), .B(KEYINPUT82), .ZN(n388) );
  XNOR2_X1 U408 ( .A(n439), .B(n388), .ZN(n341) );
  XNOR2_X1 U409 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U410 ( .A(G78GAT), .B(G211GAT), .Z(n344) );
  XNOR2_X1 U411 ( .A(G71GAT), .B(G127GAT), .ZN(n343) );
  XNOR2_X1 U412 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U413 ( .A(n346), .B(n345), .Z(n349) );
  XOR2_X1 U414 ( .A(G15GAT), .B(G1GAT), .Z(n429) );
  XNOR2_X1 U415 ( .A(n429), .B(n347), .ZN(n348) );
  XNOR2_X1 U416 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U417 ( .A(n351), .B(n350), .ZN(n569) );
  XOR2_X1 U418 ( .A(KEYINPUT20), .B(G176GAT), .Z(n353) );
  XNOR2_X1 U419 ( .A(G15GAT), .B(G190GAT), .ZN(n352) );
  XNOR2_X1 U420 ( .A(n353), .B(n352), .ZN(n362) );
  XOR2_X1 U421 ( .A(G127GAT), .B(KEYINPUT0), .Z(n355) );
  XNOR2_X1 U422 ( .A(G113GAT), .B(G134GAT), .ZN(n354) );
  XNOR2_X1 U423 ( .A(n355), .B(n354), .ZN(n373) );
  XOR2_X1 U424 ( .A(n373), .B(G183GAT), .Z(n357) );
  NAND2_X1 U425 ( .A1(G227GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U426 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U427 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U428 ( .A(n358), .B(n437), .Z(n360) );
  XNOR2_X1 U429 ( .A(G43GAT), .B(G99GAT), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U431 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U432 ( .A(KEYINPUT18), .B(KEYINPUT17), .Z(n364) );
  XNOR2_X1 U433 ( .A(G169GAT), .B(KEYINPUT19), .ZN(n363) );
  XOR2_X1 U434 ( .A(n364), .B(n363), .Z(n393) );
  INV_X1 U435 ( .A(n393), .ZN(n365) );
  XOR2_X1 U436 ( .A(n366), .B(n365), .Z(n543) );
  INV_X1 U437 ( .A(n543), .ZN(n535) );
  XOR2_X1 U438 ( .A(G57GAT), .B(KEYINPUT94), .Z(n368) );
  XNOR2_X1 U439 ( .A(KEYINPUT98), .B(KEYINPUT1), .ZN(n367) );
  XNOR2_X1 U440 ( .A(n368), .B(n367), .ZN(n372) );
  XOR2_X1 U441 ( .A(KEYINPUT5), .B(KEYINPUT96), .Z(n370) );
  XNOR2_X1 U442 ( .A(KEYINPUT97), .B(KEYINPUT95), .ZN(n369) );
  XNOR2_X1 U443 ( .A(n370), .B(n369), .ZN(n371) );
  XOR2_X1 U444 ( .A(n372), .B(n371), .Z(n379) );
  XOR2_X1 U445 ( .A(n373), .B(KEYINPUT4), .Z(n375) );
  NAND2_X1 U446 ( .A1(G225GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U448 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U449 ( .A(n379), .B(n378), .ZN(n387) );
  XOR2_X1 U450 ( .A(KEYINPUT6), .B(G155GAT), .Z(n381) );
  XNOR2_X1 U451 ( .A(G1GAT), .B(G148GAT), .ZN(n380) );
  XNOR2_X1 U452 ( .A(n381), .B(n380), .ZN(n385) );
  XOR2_X1 U453 ( .A(G85GAT), .B(G162GAT), .Z(n383) );
  XNOR2_X1 U454 ( .A(G29GAT), .B(G120GAT), .ZN(n382) );
  XNOR2_X1 U455 ( .A(n383), .B(n382), .ZN(n384) );
  XOR2_X1 U456 ( .A(n385), .B(n384), .Z(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n530) );
  XOR2_X1 U458 ( .A(G176GAT), .B(G64GAT), .Z(n449) );
  XOR2_X1 U459 ( .A(n388), .B(n449), .Z(n392) );
  NAND2_X1 U460 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XOR2_X1 U461 ( .A(n393), .B(KEYINPUT99), .Z(n394) );
  XNOR2_X1 U462 ( .A(n395), .B(n394), .ZN(n396) );
  XNOR2_X1 U463 ( .A(n397), .B(n396), .ZN(n399) );
  XNOR2_X1 U464 ( .A(KEYINPUT27), .B(n532), .ZN(n405) );
  NOR2_X1 U465 ( .A1(n530), .A2(n405), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n400), .B(KEYINPUT101), .ZN(n557) );
  INV_X1 U467 ( .A(n538), .ZN(n401) );
  XNOR2_X1 U468 ( .A(n544), .B(KEYINPUT102), .ZN(n402) );
  NAND2_X1 U469 ( .A1(n535), .A2(n402), .ZN(n413) );
  XOR2_X1 U470 ( .A(KEYINPUT103), .B(KEYINPUT26), .Z(n404) );
  NAND2_X1 U471 ( .A1(n482), .A2(n535), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n580) );
  NOR2_X1 U473 ( .A1(n580), .A2(n405), .ZN(n406) );
  XOR2_X1 U474 ( .A(KEYINPUT104), .B(n406), .Z(n410) );
  NOR2_X1 U475 ( .A1(n535), .A2(n532), .ZN(n407) );
  NOR2_X1 U476 ( .A1(n482), .A2(n407), .ZN(n408) );
  XNOR2_X1 U477 ( .A(KEYINPUT25), .B(n408), .ZN(n409) );
  NAND2_X1 U478 ( .A1(n410), .A2(n409), .ZN(n411) );
  NAND2_X1 U479 ( .A1(n411), .A2(n530), .ZN(n412) );
  NAND2_X1 U480 ( .A1(n413), .A2(n412), .ZN(n496) );
  NAND2_X1 U481 ( .A1(n569), .A2(n496), .ZN(n414) );
  NOR2_X1 U482 ( .A1(n471), .A2(n414), .ZN(n417) );
  XOR2_X1 U483 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n419) );
  XNOR2_X1 U484 ( .A(KEYINPUT68), .B(KEYINPUT66), .ZN(n418) );
  XNOR2_X1 U485 ( .A(n419), .B(n418), .ZN(n433) );
  XOR2_X1 U486 ( .A(G113GAT), .B(G36GAT), .Z(n421) );
  XNOR2_X1 U487 ( .A(G169GAT), .B(G50GAT), .ZN(n420) );
  XNOR2_X1 U488 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U489 ( .A(G8GAT), .B(G141GAT), .Z(n423) );
  XNOR2_X1 U490 ( .A(G22GAT), .B(G197GAT), .ZN(n422) );
  XNOR2_X1 U491 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U492 ( .A(n425), .B(n424), .Z(n431) );
  XOR2_X1 U493 ( .A(KEYINPUT30), .B(KEYINPUT70), .Z(n427) );
  NAND2_X1 U494 ( .A1(G229GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U495 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U496 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U497 ( .A(n431), .B(n430), .ZN(n432) );
  XNOR2_X1 U498 ( .A(n433), .B(n432), .ZN(n434) );
  XOR2_X1 U499 ( .A(n435), .B(n434), .Z(n581) );
  INV_X1 U500 ( .A(n581), .ZN(n561) );
  INV_X1 U501 ( .A(n439), .ZN(n436) );
  NAND2_X1 U502 ( .A1(n436), .A2(n437), .ZN(n441) );
  INV_X1 U503 ( .A(n437), .ZN(n438) );
  NAND2_X1 U504 ( .A1(n439), .A2(n438), .ZN(n440) );
  NAND2_X1 U505 ( .A1(n441), .A2(n440), .ZN(n444) );
  NAND2_X1 U506 ( .A1(G230GAT), .A2(G233GAT), .ZN(n442) );
  XOR2_X1 U507 ( .A(KEYINPUT73), .B(KEYINPUT72), .Z(n446) );
  XNOR2_X1 U508 ( .A(KEYINPUT33), .B(KEYINPUT31), .ZN(n445) );
  XNOR2_X1 U509 ( .A(n446), .B(n445), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n448), .B(n447), .ZN(n455) );
  XOR2_X1 U511 ( .A(KEYINPUT76), .B(KEYINPUT32), .Z(n452) );
  XNOR2_X1 U512 ( .A(n450), .B(n449), .ZN(n451) );
  XNOR2_X1 U513 ( .A(n452), .B(n451), .ZN(n453) );
  XOR2_X1 U514 ( .A(n453), .B(G92GAT), .Z(n454) );
  XNOR2_X1 U515 ( .A(n455), .B(n454), .ZN(n456) );
  INV_X1 U516 ( .A(n473), .ZN(n585) );
  NOR2_X1 U517 ( .A1(n561), .A2(n585), .ZN(n498) );
  NAND2_X1 U518 ( .A1(n528), .A2(n498), .ZN(n458) );
  XNOR2_X1 U519 ( .A(n458), .B(KEYINPUT38), .ZN(n516) );
  NOR2_X1 U520 ( .A1(n538), .A2(n516), .ZN(n461) );
  INV_X1 U521 ( .A(n569), .ZN(n588) );
  NOR2_X1 U522 ( .A1(n561), .A2(n563), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n462), .B(KEYINPUT46), .ZN(n463) );
  NOR2_X2 U524 ( .A1(n588), .A2(n463), .ZN(n464) );
  NAND2_X1 U525 ( .A1(n464), .A2(KEYINPUT118), .ZN(n468) );
  INV_X1 U526 ( .A(KEYINPUT118), .ZN(n466) );
  INV_X1 U527 ( .A(n464), .ZN(n465) );
  NAND2_X1 U528 ( .A1(n466), .A2(n465), .ZN(n467) );
  NAND2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  NAND2_X1 U530 ( .A1(n469), .A2(n572), .ZN(n470) );
  XNOR2_X1 U531 ( .A(n470), .B(KEYINPUT47), .ZN(n477) );
  NOR2_X1 U532 ( .A1(n471), .A2(n569), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(KEYINPUT45), .ZN(n474) );
  NAND2_X1 U534 ( .A1(n474), .A2(n473), .ZN(n475) );
  NOR2_X1 U535 ( .A1(n581), .A2(n475), .ZN(n476) );
  NOR2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n478) );
  XNOR2_X1 U537 ( .A(n478), .B(KEYINPUT64), .ZN(n479) );
  XNOR2_X1 U538 ( .A(n479), .B(KEYINPUT48), .ZN(n542) );
  NOR2_X1 U539 ( .A1(n542), .A2(n532), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n480), .B(KEYINPUT54), .ZN(n481) );
  NAND2_X1 U541 ( .A1(n481), .A2(n530), .ZN(n579) );
  XNOR2_X1 U542 ( .A(KEYINPUT55), .B(KEYINPUT123), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(n485) );
  NAND2_X1 U544 ( .A1(n543), .A2(n485), .ZN(n486) );
  XOR2_X2 U545 ( .A(KEYINPUT124), .B(n486), .Z(n576) );
  NAND2_X1 U546 ( .A1(n576), .A2(n553), .ZN(n490) );
  XOR2_X1 U547 ( .A(KEYINPUT58), .B(KEYINPUT126), .Z(n488) );
  INV_X1 U548 ( .A(G190GAT), .ZN(n487) );
  XNOR2_X1 U549 ( .A(n490), .B(n489), .ZN(G1351GAT) );
  INV_X1 U550 ( .A(n563), .ZN(n547) );
  NAND2_X1 U551 ( .A1(n547), .A2(n576), .ZN(n493) );
  XOR2_X1 U552 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G176GAT), .ZN(n492) );
  NOR2_X1 U554 ( .A1(n553), .A2(n569), .ZN(n495) );
  XNOR2_X1 U555 ( .A(KEYINPUT86), .B(KEYINPUT16), .ZN(n494) );
  XNOR2_X1 U556 ( .A(n495), .B(n494), .ZN(n497) );
  AND2_X1 U557 ( .A1(n497), .A2(n496), .ZN(n519) );
  NAND2_X1 U558 ( .A1(n498), .A2(n519), .ZN(n508) );
  NOR2_X1 U559 ( .A1(n530), .A2(n508), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT107), .B(KEYINPUT34), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n501) );
  XOR2_X1 U562 ( .A(n501), .B(KEYINPUT106), .Z(n503) );
  XNOR2_X1 U563 ( .A(G1GAT), .B(KEYINPUT105), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n503), .B(n502), .ZN(G1324GAT) );
  NOR2_X1 U565 ( .A1(n532), .A2(n508), .ZN(n504) );
  XOR2_X1 U566 ( .A(KEYINPUT108), .B(n504), .Z(n505) );
  XNOR2_X1 U567 ( .A(G8GAT), .B(n505), .ZN(G1325GAT) );
  NOR2_X1 U568 ( .A1(n535), .A2(n508), .ZN(n507) );
  XNOR2_X1 U569 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n506) );
  XNOR2_X1 U570 ( .A(n507), .B(n506), .ZN(G1326GAT) );
  NOR2_X1 U571 ( .A1(n538), .A2(n508), .ZN(n510) );
  XNOR2_X1 U572 ( .A(KEYINPUT109), .B(KEYINPUT110), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U574 ( .A(G22GAT), .B(n511), .ZN(G1327GAT) );
  NOR2_X1 U575 ( .A1(n516), .A2(n530), .ZN(n513) );
  XNOR2_X1 U576 ( .A(KEYINPUT113), .B(KEYINPUT39), .ZN(n512) );
  XNOR2_X1 U577 ( .A(n513), .B(n512), .ZN(n514) );
  XOR2_X1 U578 ( .A(G29GAT), .B(n514), .Z(G1328GAT) );
  NOR2_X1 U579 ( .A1(n516), .A2(n532), .ZN(n515) );
  XOR2_X1 U580 ( .A(G36GAT), .B(n515), .Z(G1329GAT) );
  NOR2_X1 U581 ( .A1(n535), .A2(n516), .ZN(n517) );
  XOR2_X1 U582 ( .A(KEYINPUT40), .B(n517), .Z(n518) );
  XNOR2_X1 U583 ( .A(G43GAT), .B(n518), .ZN(G1330GAT) );
  NOR2_X1 U584 ( .A1(n581), .A2(n563), .ZN(n529) );
  NAND2_X1 U585 ( .A1(n529), .A2(n519), .ZN(n524) );
  NOR2_X1 U586 ( .A1(n530), .A2(n524), .ZN(n520) );
  XOR2_X1 U587 ( .A(G57GAT), .B(n520), .Z(n521) );
  XNOR2_X1 U588 ( .A(KEYINPUT42), .B(n521), .ZN(G1332GAT) );
  NOR2_X1 U589 ( .A1(n532), .A2(n524), .ZN(n522) );
  XOR2_X1 U590 ( .A(G64GAT), .B(n522), .Z(G1333GAT) );
  NOR2_X1 U591 ( .A1(n535), .A2(n524), .ZN(n523) );
  XOR2_X1 U592 ( .A(G71GAT), .B(n523), .Z(G1334GAT) );
  NOR2_X1 U593 ( .A1(n538), .A2(n524), .ZN(n526) );
  XNOR2_X1 U594 ( .A(KEYINPUT115), .B(KEYINPUT43), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U596 ( .A(G78GAT), .B(n527), .Z(G1335GAT) );
  NAND2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n537) );
  NOR2_X1 U598 ( .A1(n530), .A2(n537), .ZN(n531) );
  XOR2_X1 U599 ( .A(G85GAT), .B(n531), .Z(G1336GAT) );
  NOR2_X1 U600 ( .A1(n532), .A2(n537), .ZN(n533) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(n533), .Z(n534) );
  XNOR2_X1 U602 ( .A(G92GAT), .B(n534), .ZN(G1337GAT) );
  NOR2_X1 U603 ( .A1(n535), .A2(n537), .ZN(n536) );
  XOR2_X1 U604 ( .A(G99GAT), .B(n536), .Z(G1338GAT) );
  NOR2_X1 U605 ( .A1(n538), .A2(n537), .ZN(n540) );
  XNOR2_X1 U606 ( .A(KEYINPUT117), .B(KEYINPUT44), .ZN(n539) );
  XNOR2_X1 U607 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U608 ( .A(G106GAT), .B(n541), .ZN(G1339GAT) );
  BUF_X1 U609 ( .A(n542), .Z(n558) );
  NAND2_X1 U610 ( .A1(n544), .A2(n543), .ZN(n545) );
  NOR2_X1 U611 ( .A1(n558), .A2(n545), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n581), .A2(n554), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n546), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U614 ( .A(G120GAT), .B(KEYINPUT49), .Z(n549) );
  NAND2_X1 U615 ( .A1(n554), .A2(n547), .ZN(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(G1341GAT) );
  XOR2_X1 U617 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n551) );
  NAND2_X1 U618 ( .A1(n554), .A2(n588), .ZN(n550) );
  XNOR2_X1 U619 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U620 ( .A(G127GAT), .B(n552), .ZN(G1342GAT) );
  XOR2_X1 U621 ( .A(G134GAT), .B(KEYINPUT51), .Z(n556) );
  NAND2_X1 U622 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1343GAT) );
  NOR2_X1 U624 ( .A1(n580), .A2(n557), .ZN(n560) );
  NAND2_X1 U625 ( .A1(n560), .A2(n559), .ZN(n571) );
  NOR2_X1 U626 ( .A1(n561), .A2(n571), .ZN(n562) );
  XOR2_X1 U627 ( .A(G141GAT), .B(n562), .Z(G1344GAT) );
  NOR2_X1 U628 ( .A1(n563), .A2(n571), .ZN(n568) );
  XOR2_X1 U629 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n565) );
  XNOR2_X1 U630 ( .A(G148GAT), .B(KEYINPUT52), .ZN(n564) );
  XNOR2_X1 U631 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U632 ( .A(KEYINPUT53), .B(n566), .ZN(n567) );
  XNOR2_X1 U633 ( .A(n568), .B(n567), .ZN(G1345GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n571), .ZN(n570) );
  XOR2_X1 U635 ( .A(G155GAT), .B(n570), .Z(G1346GAT) );
  NOR2_X1 U636 ( .A1(n572), .A2(n571), .ZN(n573) );
  XOR2_X1 U637 ( .A(KEYINPUT122), .B(n573), .Z(n574) );
  XNOR2_X1 U638 ( .A(G162GAT), .B(n574), .ZN(G1347GAT) );
  NAND2_X1 U639 ( .A1(n576), .A2(n581), .ZN(n575) );
  XNOR2_X1 U640 ( .A(n575), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U641 ( .A(G183GAT), .B(KEYINPUT125), .Z(n578) );
  NAND2_X1 U642 ( .A1(n588), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(G1350GAT) );
  XOR2_X1 U644 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n583) );
  NOR2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n591) );
  NAND2_X1 U646 ( .A1(n591), .A2(n581), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(G204GAT), .B(KEYINPUT61), .Z(n587) );
  NAND2_X1 U650 ( .A1(n591), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n587), .B(n586), .ZN(G1353GAT) );
  XOR2_X1 U652 ( .A(G211GAT), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U653 ( .A1(n591), .A2(n588), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(G1354GAT) );
  INV_X1 U655 ( .A(n591), .ZN(n592) );
  NOR2_X1 U656 ( .A1(n471), .A2(n592), .ZN(n593) );
  XOR2_X1 U657 ( .A(KEYINPUT62), .B(n593), .Z(n594) );
  XNOR2_X1 U658 ( .A(G218GAT), .B(n594), .ZN(G1355GAT) );
endmodule

