

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  XOR2_X1 U548 ( .A(KEYINPUT1), .B(n520), .Z(n792) );
  XNOR2_X1 U549 ( .A(KEYINPUT66), .B(G543), .ZN(n516) );
  XOR2_X1 U550 ( .A(KEYINPUT92), .B(n738), .Z(n514) );
  INV_X1 U551 ( .A(n1008), .ZN(n618) );
  INV_X1 U552 ( .A(n666), .ZN(n643) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n641) );
  XNOR2_X1 U554 ( .A(n642), .B(n641), .ZN(n647) );
  AND2_X1 U555 ( .A1(n673), .A2(n672), .ZN(n674) );
  INV_X1 U556 ( .A(G2104), .ZN(n579) );
  NOR2_X2 U557 ( .A1(G2105), .A2(n579), .ZN(n886) );
  INV_X1 U558 ( .A(KEYINPUT109), .ZN(n742) );
  INV_X1 U559 ( .A(KEYINPUT0), .ZN(n515) );
  NOR2_X1 U560 ( .A1(G651), .A2(n551), .ZN(n791) );
  INV_X1 U561 ( .A(KEYINPUT91), .ZN(n589) );
  XNOR2_X1 U562 ( .A(n516), .B(n515), .ZN(n551) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n797) );
  NAND2_X1 U564 ( .A1(n797), .A2(G91), .ZN(n518) );
  XNOR2_X1 U565 ( .A(KEYINPUT67), .B(G651), .ZN(n519) );
  NOR2_X1 U566 ( .A1(n551), .A2(n519), .ZN(n795) );
  NAND2_X1 U567 ( .A1(G78), .A2(n795), .ZN(n517) );
  NAND2_X1 U568 ( .A1(n518), .A2(n517), .ZN(n524) );
  NAND2_X1 U569 ( .A1(n791), .A2(G53), .ZN(n522) );
  NOR2_X1 U570 ( .A1(G543), .A2(n519), .ZN(n520) );
  NAND2_X1 U571 ( .A1(G65), .A2(n792), .ZN(n521) );
  NAND2_X1 U572 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U573 ( .A1(n524), .A2(n523), .ZN(n525) );
  XOR2_X1 U574 ( .A(KEYINPUT70), .B(n525), .Z(G299) );
  NAND2_X1 U575 ( .A1(n792), .A2(G64), .ZN(n526) );
  XNOR2_X1 U576 ( .A(n526), .B(KEYINPUT68), .ZN(n529) );
  NAND2_X1 U577 ( .A1(G52), .A2(n791), .ZN(n527) );
  XOR2_X1 U578 ( .A(KEYINPUT69), .B(n527), .Z(n528) );
  NAND2_X1 U579 ( .A1(n529), .A2(n528), .ZN(n534) );
  NAND2_X1 U580 ( .A1(n797), .A2(G90), .ZN(n531) );
  NAND2_X1 U581 ( .A1(G77), .A2(n795), .ZN(n530) );
  NAND2_X1 U582 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U583 ( .A(KEYINPUT9), .B(n532), .Z(n533) );
  NOR2_X1 U584 ( .A1(n534), .A2(n533), .ZN(G171) );
  NAND2_X1 U585 ( .A1(n791), .A2(G51), .ZN(n536) );
  NAND2_X1 U586 ( .A1(G63), .A2(n792), .ZN(n535) );
  NAND2_X1 U587 ( .A1(n536), .A2(n535), .ZN(n537) );
  XNOR2_X1 U588 ( .A(KEYINPUT6), .B(n537), .ZN(n544) );
  NAND2_X1 U589 ( .A1(n797), .A2(G89), .ZN(n538) );
  XNOR2_X1 U590 ( .A(n538), .B(KEYINPUT4), .ZN(n540) );
  NAND2_X1 U591 ( .A1(G76), .A2(n795), .ZN(n539) );
  NAND2_X1 U592 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U593 ( .A(KEYINPUT5), .B(n541), .Z(n542) );
  XNOR2_X1 U594 ( .A(KEYINPUT74), .B(n542), .ZN(n543) );
  NOR2_X1 U595 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U596 ( .A(KEYINPUT7), .B(n545), .Z(G168) );
  NAND2_X1 U597 ( .A1(n791), .A2(G49), .ZN(n546) );
  XNOR2_X1 U598 ( .A(n546), .B(KEYINPUT80), .ZN(n548) );
  NAND2_X1 U599 ( .A1(G74), .A2(G651), .ZN(n547) );
  NAND2_X1 U600 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U601 ( .A(KEYINPUT81), .B(n549), .Z(n550) );
  NOR2_X1 U602 ( .A1(n792), .A2(n550), .ZN(n553) );
  NAND2_X1 U603 ( .A1(G87), .A2(n551), .ZN(n552) );
  NAND2_X1 U604 ( .A1(n553), .A2(n552), .ZN(G288) );
  XOR2_X1 U605 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U606 ( .A1(n797), .A2(G88), .ZN(n555) );
  NAND2_X1 U607 ( .A1(G75), .A2(n795), .ZN(n554) );
  NAND2_X1 U608 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U609 ( .A1(n791), .A2(G50), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G62), .A2(n792), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U612 ( .A(KEYINPUT83), .B(n558), .Z(n559) );
  NOR2_X1 U613 ( .A1(n560), .A2(n559), .ZN(G166) );
  INV_X1 U614 ( .A(G166), .ZN(G303) );
  NAND2_X1 U615 ( .A1(n795), .A2(G73), .ZN(n561) );
  XNOR2_X1 U616 ( .A(n561), .B(KEYINPUT2), .ZN(n568) );
  NAND2_X1 U617 ( .A1(n797), .A2(G86), .ZN(n563) );
  NAND2_X1 U618 ( .A1(G61), .A2(n792), .ZN(n562) );
  NAND2_X1 U619 ( .A1(n563), .A2(n562), .ZN(n566) );
  NAND2_X1 U620 ( .A1(n791), .A2(G48), .ZN(n564) );
  XOR2_X1 U621 ( .A(KEYINPUT82), .B(n564), .Z(n565) );
  NOR2_X1 U622 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U623 ( .A1(n568), .A2(n567), .ZN(G305) );
  NAND2_X1 U624 ( .A1(n797), .A2(G85), .ZN(n570) );
  NAND2_X1 U625 ( .A1(G72), .A2(n795), .ZN(n569) );
  NAND2_X1 U626 ( .A1(n570), .A2(n569), .ZN(n574) );
  NAND2_X1 U627 ( .A1(n791), .A2(G47), .ZN(n572) );
  NAND2_X1 U628 ( .A1(G60), .A2(n792), .ZN(n571) );
  NAND2_X1 U629 ( .A1(n572), .A2(n571), .ZN(n573) );
  OR2_X1 U630 ( .A1(n574), .A2(n573), .ZN(G290) );
  NOR2_X1 U631 ( .A1(G2105), .A2(G2104), .ZN(n575) );
  XOR2_X1 U632 ( .A(KEYINPUT17), .B(n575), .Z(n707) );
  NAND2_X1 U633 ( .A1(n707), .A2(G137), .ZN(n578) );
  NAND2_X1 U634 ( .A1(G101), .A2(n886), .ZN(n576) );
  XOR2_X1 U635 ( .A(KEYINPUT23), .B(n576), .Z(n577) );
  NAND2_X1 U636 ( .A1(n578), .A2(n577), .ZN(n584) );
  AND2_X1 U637 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U638 ( .A1(G113), .A2(n882), .ZN(n582) );
  NAND2_X1 U639 ( .A1(n579), .A2(G2105), .ZN(n580) );
  XNOR2_X2 U640 ( .A(n580), .B(KEYINPUT65), .ZN(n883) );
  NAND2_X1 U641 ( .A1(G125), .A2(n883), .ZN(n581) );
  NAND2_X1 U642 ( .A1(n582), .A2(n581), .ZN(n583) );
  NOR2_X1 U643 ( .A1(n584), .A2(n583), .ZN(n760) );
  NAND2_X1 U644 ( .A1(n760), .A2(G40), .ZN(n705) );
  INV_X1 U645 ( .A(n705), .ZN(n593) );
  NAND2_X1 U646 ( .A1(G114), .A2(n882), .ZN(n586) );
  NAND2_X1 U647 ( .A1(G126), .A2(n883), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n592) );
  NAND2_X1 U649 ( .A1(G102), .A2(n886), .ZN(n588) );
  NAND2_X1 U650 ( .A1(G138), .A2(n707), .ZN(n587) );
  NAND2_X1 U651 ( .A1(n588), .A2(n587), .ZN(n590) );
  XNOR2_X1 U652 ( .A(n590), .B(n589), .ZN(n591) );
  NOR2_X1 U653 ( .A1(n592), .A2(n591), .ZN(n761) );
  NOR2_X2 U654 ( .A1(n761), .A2(G1384), .ZN(n706) );
  NAND2_X2 U655 ( .A1(n593), .A2(n706), .ZN(n666) );
  NOR2_X1 U656 ( .A1(G2084), .A2(n666), .ZN(n648) );
  NAND2_X1 U657 ( .A1(G8), .A2(n648), .ZN(n663) );
  NAND2_X1 U658 ( .A1(G8), .A2(n666), .ZN(n701) );
  NOR2_X1 U659 ( .A1(G1966), .A2(n701), .ZN(n649) );
  INV_X1 U660 ( .A(n649), .ZN(n661) );
  NAND2_X1 U661 ( .A1(n791), .A2(G54), .ZN(n595) );
  NAND2_X1 U662 ( .A1(G66), .A2(n792), .ZN(n594) );
  NAND2_X1 U663 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U664 ( .A1(n797), .A2(G92), .ZN(n597) );
  NAND2_X1 U665 ( .A1(G79), .A2(n795), .ZN(n596) );
  NAND2_X1 U666 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U667 ( .A1(n599), .A2(n598), .ZN(n600) );
  XNOR2_X1 U668 ( .A(n600), .B(KEYINPUT15), .ZN(n768) );
  NAND2_X1 U669 ( .A1(G1996), .A2(n643), .ZN(n601) );
  XNOR2_X1 U670 ( .A(n601), .B(KEYINPUT26), .ZN(n603) );
  NAND2_X1 U671 ( .A1(G1341), .A2(n666), .ZN(n602) );
  NAND2_X1 U672 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT104), .ZN(n605) );
  INV_X1 U674 ( .A(n605), .ZN(n619) );
  NAND2_X1 U675 ( .A1(G81), .A2(n797), .ZN(n606) );
  XNOR2_X1 U676 ( .A(n606), .B(KEYINPUT12), .ZN(n607) );
  XNOR2_X1 U677 ( .A(n607), .B(KEYINPUT72), .ZN(n609) );
  NAND2_X1 U678 ( .A1(n795), .A2(G68), .ZN(n608) );
  NAND2_X1 U679 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U680 ( .A(KEYINPUT13), .B(n610), .ZN(n614) );
  XOR2_X1 U681 ( .A(KEYINPUT71), .B(KEYINPUT14), .Z(n612) );
  NAND2_X1 U682 ( .A1(G56), .A2(n792), .ZN(n611) );
  XNOR2_X1 U683 ( .A(n612), .B(n611), .ZN(n613) );
  NAND2_X1 U684 ( .A1(n614), .A2(n613), .ZN(n615) );
  XNOR2_X1 U685 ( .A(n615), .B(KEYINPUT73), .ZN(n617) );
  NAND2_X1 U686 ( .A1(n791), .A2(G43), .ZN(n616) );
  NAND2_X1 U687 ( .A1(n617), .A2(n616), .ZN(n1008) );
  NAND2_X1 U688 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U689 ( .A(n620), .B(KEYINPUT64), .ZN(n625) );
  OR2_X1 U690 ( .A1(n768), .A2(n625), .ZN(n624) );
  NOR2_X1 U691 ( .A1(n643), .A2(G1348), .ZN(n622) );
  NOR2_X1 U692 ( .A1(G2067), .A2(n666), .ZN(n621) );
  NOR2_X1 U693 ( .A1(n622), .A2(n621), .ZN(n623) );
  NAND2_X1 U694 ( .A1(n624), .A2(n623), .ZN(n627) );
  NAND2_X1 U695 ( .A1(n625), .A2(n768), .ZN(n626) );
  NAND2_X1 U696 ( .A1(n627), .A2(n626), .ZN(n634) );
  NAND2_X1 U697 ( .A1(G2072), .A2(n643), .ZN(n628) );
  XOR2_X1 U698 ( .A(KEYINPUT101), .B(n628), .Z(n629) );
  XNOR2_X1 U699 ( .A(KEYINPUT27), .B(n629), .ZN(n632) );
  NAND2_X1 U700 ( .A1(G1956), .A2(n666), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT102), .B(n630), .Z(n631) );
  NOR2_X1 U702 ( .A1(n632), .A2(n631), .ZN(n636) );
  INV_X1 U703 ( .A(G299), .ZN(n635) );
  NAND2_X1 U704 ( .A1(n636), .A2(n635), .ZN(n633) );
  NAND2_X1 U705 ( .A1(n634), .A2(n633), .ZN(n640) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n638) );
  XNOR2_X1 U707 ( .A(KEYINPUT103), .B(KEYINPUT28), .ZN(n637) );
  XNOR2_X1 U708 ( .A(n638), .B(n637), .ZN(n639) );
  NAND2_X1 U709 ( .A1(n640), .A2(n639), .ZN(n642) );
  INV_X1 U710 ( .A(G1961), .ZN(n968) );
  NAND2_X1 U711 ( .A1(n666), .A2(n968), .ZN(n645) );
  XNOR2_X1 U712 ( .A(G2078), .B(KEYINPUT25), .ZN(n929) );
  NAND2_X1 U713 ( .A1(n643), .A2(n929), .ZN(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n655) );
  NAND2_X1 U715 ( .A1(n655), .A2(G171), .ZN(n646) );
  NAND2_X1 U716 ( .A1(n647), .A2(n646), .ZN(n660) );
  NOR2_X1 U717 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U718 ( .A1(G8), .A2(n650), .ZN(n651) );
  XNOR2_X1 U719 ( .A(KEYINPUT106), .B(n651), .ZN(n653) );
  XOR2_X1 U720 ( .A(KEYINPUT30), .B(KEYINPUT105), .Z(n652) );
  XNOR2_X1 U721 ( .A(n653), .B(n652), .ZN(n654) );
  NOR2_X1 U722 ( .A1(G168), .A2(n654), .ZN(n657) );
  NOR2_X1 U723 ( .A1(G171), .A2(n655), .ZN(n656) );
  NOR2_X1 U724 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U725 ( .A(KEYINPUT31), .B(n658), .Z(n659) );
  NAND2_X1 U726 ( .A1(n660), .A2(n659), .ZN(n665) );
  AND2_X1 U727 ( .A1(n661), .A2(n665), .ZN(n662) );
  NAND2_X1 U728 ( .A1(n663), .A2(n662), .ZN(n691) );
  INV_X1 U729 ( .A(n701), .ZN(n664) );
  NAND2_X1 U730 ( .A1(G1976), .A2(G288), .ZN(n993) );
  AND2_X1 U731 ( .A1(n664), .A2(n993), .ZN(n676) );
  AND2_X1 U732 ( .A1(n691), .A2(n676), .ZN(n675) );
  NAND2_X1 U733 ( .A1(n665), .A2(G286), .ZN(n673) );
  INV_X1 U734 ( .A(G8), .ZN(n671) );
  NOR2_X1 U735 ( .A1(G1971), .A2(n701), .ZN(n668) );
  NOR2_X1 U736 ( .A1(G2090), .A2(n666), .ZN(n667) );
  NOR2_X1 U737 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n669), .A2(G303), .ZN(n670) );
  OR2_X1 U739 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U740 ( .A(n674), .B(KEYINPUT32), .ZN(n690) );
  AND2_X1 U741 ( .A1(n675), .A2(n690), .ZN(n682) );
  INV_X1 U742 ( .A(n676), .ZN(n678) );
  NOR2_X1 U743 ( .A1(G1976), .A2(G288), .ZN(n683) );
  NOR2_X1 U744 ( .A1(G1971), .A2(G303), .ZN(n677) );
  NOR2_X1 U745 ( .A1(n683), .A2(n677), .ZN(n994) );
  OR2_X1 U746 ( .A1(n678), .A2(n994), .ZN(n680) );
  INV_X1 U747 ( .A(KEYINPUT33), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U749 ( .A1(n682), .A2(n681), .ZN(n686) );
  NAND2_X1 U750 ( .A1(n683), .A2(KEYINPUT33), .ZN(n684) );
  NOR2_X1 U751 ( .A1(n701), .A2(n684), .ZN(n685) );
  NOR2_X1 U752 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U753 ( .A(G1981), .B(G305), .Z(n1005) );
  NAND2_X1 U754 ( .A1(n687), .A2(n1005), .ZN(n696) );
  NOR2_X1 U755 ( .A1(G2090), .A2(G303), .ZN(n688) );
  XOR2_X1 U756 ( .A(KEYINPUT107), .B(n688), .Z(n689) );
  NAND2_X1 U757 ( .A1(G8), .A2(n689), .ZN(n693) );
  NAND2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  NAND2_X1 U759 ( .A1(n693), .A2(n692), .ZN(n694) );
  NAND2_X1 U760 ( .A1(n694), .A2(n701), .ZN(n695) );
  NAND2_X1 U761 ( .A1(n696), .A2(n695), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n697), .B(KEYINPUT108), .ZN(n703) );
  NOR2_X1 U763 ( .A1(G1981), .A2(G305), .ZN(n698) );
  XOR2_X1 U764 ( .A(n698), .B(KEYINPUT100), .Z(n699) );
  XNOR2_X1 U765 ( .A(KEYINPUT24), .B(n699), .ZN(n700) );
  NOR2_X1 U766 ( .A1(n701), .A2(n700), .ZN(n702) );
  NOR2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n704) );
  INV_X1 U768 ( .A(n704), .ZN(n741) );
  NOR2_X1 U769 ( .A1(n706), .A2(n705), .ZN(n755) );
  BUF_X1 U770 ( .A(n707), .Z(n887) );
  NAND2_X1 U771 ( .A1(G141), .A2(n887), .ZN(n709) );
  NAND2_X1 U772 ( .A1(G129), .A2(n883), .ZN(n708) );
  NAND2_X1 U773 ( .A1(n709), .A2(n708), .ZN(n712) );
  NAND2_X1 U774 ( .A1(n886), .A2(G105), .ZN(n710) );
  XOR2_X1 U775 ( .A(KEYINPUT38), .B(n710), .Z(n711) );
  NOR2_X1 U776 ( .A1(n712), .A2(n711), .ZN(n714) );
  NAND2_X1 U777 ( .A1(n882), .A2(G117), .ZN(n713) );
  NAND2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n899) );
  NAND2_X1 U779 ( .A1(G1996), .A2(n899), .ZN(n715) );
  XNOR2_X1 U780 ( .A(n715), .B(KEYINPUT98), .ZN(n725) );
  NAND2_X1 U781 ( .A1(G95), .A2(n886), .ZN(n717) );
  NAND2_X1 U782 ( .A1(G131), .A2(n887), .ZN(n716) );
  NAND2_X1 U783 ( .A1(n717), .A2(n716), .ZN(n722) );
  NAND2_X1 U784 ( .A1(G107), .A2(n882), .ZN(n719) );
  NAND2_X1 U785 ( .A1(G119), .A2(n883), .ZN(n718) );
  NAND2_X1 U786 ( .A1(n719), .A2(n718), .ZN(n720) );
  XOR2_X1 U787 ( .A(KEYINPUT95), .B(n720), .Z(n721) );
  NOR2_X1 U788 ( .A1(n722), .A2(n721), .ZN(n723) );
  XOR2_X1 U789 ( .A(KEYINPUT96), .B(n723), .Z(n896) );
  XOR2_X1 U790 ( .A(KEYINPUT97), .B(G1991), .Z(n924) );
  NAND2_X1 U791 ( .A1(n896), .A2(n924), .ZN(n724) );
  NAND2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n951) );
  NAND2_X1 U793 ( .A1(n755), .A2(n951), .ZN(n744) );
  NAND2_X1 U794 ( .A1(G104), .A2(n886), .ZN(n727) );
  NAND2_X1 U795 ( .A1(G140), .A2(n887), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n728) );
  XNOR2_X1 U797 ( .A(KEYINPUT34), .B(n728), .ZN(n734) );
  NAND2_X1 U798 ( .A1(G116), .A2(n882), .ZN(n730) );
  NAND2_X1 U799 ( .A1(G128), .A2(n883), .ZN(n729) );
  NAND2_X1 U800 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U801 ( .A(KEYINPUT93), .B(n731), .ZN(n732) );
  XNOR2_X1 U802 ( .A(KEYINPUT35), .B(n732), .ZN(n733) );
  NOR2_X1 U803 ( .A1(n734), .A2(n733), .ZN(n735) );
  XNOR2_X1 U804 ( .A(n735), .B(KEYINPUT36), .ZN(n736) );
  XNOR2_X1 U805 ( .A(n736), .B(KEYINPUT94), .ZN(n879) );
  XNOR2_X1 U806 ( .A(KEYINPUT37), .B(G2067), .ZN(n753) );
  NOR2_X1 U807 ( .A1(n879), .A2(n753), .ZN(n956) );
  NAND2_X1 U808 ( .A1(n755), .A2(n956), .ZN(n751) );
  NAND2_X1 U809 ( .A1(n744), .A2(n751), .ZN(n737) );
  XOR2_X1 U810 ( .A(KEYINPUT99), .B(n737), .Z(n739) );
  XNOR2_X1 U811 ( .A(G1986), .B(G290), .ZN(n1001) );
  NAND2_X1 U812 ( .A1(n755), .A2(n1001), .ZN(n738) );
  NOR2_X1 U813 ( .A1(n739), .A2(n514), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n741), .A2(n740), .ZN(n743) );
  XNOR2_X1 U815 ( .A(n743), .B(n742), .ZN(n758) );
  NOR2_X1 U816 ( .A1(G1996), .A2(n899), .ZN(n945) );
  INV_X1 U817 ( .A(n744), .ZN(n747) );
  NOR2_X1 U818 ( .A1(G1986), .A2(G290), .ZN(n745) );
  NOR2_X1 U819 ( .A1(n924), .A2(n896), .ZN(n952) );
  NOR2_X1 U820 ( .A1(n745), .A2(n952), .ZN(n746) );
  NOR2_X1 U821 ( .A1(n747), .A2(n746), .ZN(n748) );
  NOR2_X1 U822 ( .A1(n945), .A2(n748), .ZN(n749) );
  XNOR2_X1 U823 ( .A(KEYINPUT110), .B(n749), .ZN(n750) );
  XNOR2_X1 U824 ( .A(n750), .B(KEYINPUT39), .ZN(n752) );
  NAND2_X1 U825 ( .A1(n752), .A2(n751), .ZN(n754) );
  NAND2_X1 U826 ( .A1(n879), .A2(n753), .ZN(n959) );
  NAND2_X1 U827 ( .A1(n754), .A2(n959), .ZN(n756) );
  NAND2_X1 U828 ( .A1(n756), .A2(n755), .ZN(n757) );
  NAND2_X1 U829 ( .A1(n758), .A2(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n759), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U831 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U832 ( .A(G132), .ZN(G219) );
  INV_X1 U833 ( .A(G82), .ZN(G220) );
  INV_X1 U834 ( .A(G120), .ZN(G236) );
  INV_X1 U835 ( .A(G69), .ZN(G235) );
  INV_X1 U836 ( .A(G108), .ZN(G238) );
  BUF_X1 U837 ( .A(n760), .Z(G160) );
  BUF_X1 U838 ( .A(n761), .Z(G164) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U840 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U841 ( .A(G223), .ZN(n835) );
  NAND2_X1 U842 ( .A1(n835), .A2(G567), .ZN(n763) );
  XOR2_X1 U843 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  INV_X1 U844 ( .A(G860), .ZN(n842) );
  OR2_X1 U845 ( .A1(n1008), .A2(n842), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  NAND2_X1 U847 ( .A1(G868), .A2(G301), .ZN(n765) );
  INV_X1 U848 ( .A(G868), .ZN(n806) );
  NAND2_X1 U849 ( .A1(n768), .A2(n806), .ZN(n764) );
  NAND2_X1 U850 ( .A1(n765), .A2(n764), .ZN(G284) );
  NOR2_X1 U851 ( .A1(G286), .A2(n806), .ZN(n767) );
  NOR2_X1 U852 ( .A1(G299), .A2(G868), .ZN(n766) );
  NOR2_X1 U853 ( .A1(n767), .A2(n766), .ZN(G297) );
  NAND2_X1 U854 ( .A1(n842), .A2(G559), .ZN(n769) );
  INV_X1 U855 ( .A(n768), .ZN(n997) );
  NAND2_X1 U856 ( .A1(n769), .A2(n997), .ZN(n770) );
  XNOR2_X1 U857 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n1008), .ZN(n773) );
  NAND2_X1 U859 ( .A1(G868), .A2(n997), .ZN(n771) );
  NOR2_X1 U860 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U861 ( .A1(n773), .A2(n772), .ZN(G282) );
  XOR2_X1 U862 ( .A(G2100), .B(KEYINPUT76), .Z(n783) );
  NAND2_X1 U863 ( .A1(n883), .A2(G123), .ZN(n774) );
  XNOR2_X1 U864 ( .A(n774), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U865 ( .A1(G135), .A2(n887), .ZN(n775) );
  NAND2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n781) );
  NAND2_X1 U867 ( .A1(G99), .A2(n886), .ZN(n778) );
  NAND2_X1 U868 ( .A1(G111), .A2(n882), .ZN(n777) );
  NAND2_X1 U869 ( .A1(n778), .A2(n777), .ZN(n779) );
  XOR2_X1 U870 ( .A(KEYINPUT75), .B(n779), .Z(n780) );
  NOR2_X1 U871 ( .A1(n781), .A2(n780), .ZN(n950) );
  XNOR2_X1 U872 ( .A(G2096), .B(n950), .ZN(n782) );
  NAND2_X1 U873 ( .A1(n783), .A2(n782), .ZN(G156) );
  NAND2_X1 U874 ( .A1(G559), .A2(n997), .ZN(n784) );
  XOR2_X1 U875 ( .A(n1008), .B(n784), .Z(n841) );
  XNOR2_X1 U876 ( .A(KEYINPUT84), .B(KEYINPUT19), .ZN(n786) );
  XNOR2_X1 U877 ( .A(G290), .B(KEYINPUT85), .ZN(n785) );
  XNOR2_X1 U878 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U879 ( .A(G299), .B(n787), .ZN(n789) );
  XNOR2_X1 U880 ( .A(G305), .B(G166), .ZN(n788) );
  XNOR2_X1 U881 ( .A(n789), .B(n788), .ZN(n790) );
  XNOR2_X1 U882 ( .A(n790), .B(G288), .ZN(n804) );
  NAND2_X1 U883 ( .A1(n791), .A2(G55), .ZN(n794) );
  NAND2_X1 U884 ( .A1(G67), .A2(n792), .ZN(n793) );
  NAND2_X1 U885 ( .A1(n794), .A2(n793), .ZN(n802) );
  NAND2_X1 U886 ( .A1(G80), .A2(n795), .ZN(n796) );
  XOR2_X1 U887 ( .A(KEYINPUT77), .B(n796), .Z(n799) );
  NAND2_X1 U888 ( .A1(n797), .A2(G93), .ZN(n798) );
  NAND2_X1 U889 ( .A1(n799), .A2(n798), .ZN(n800) );
  XNOR2_X1 U890 ( .A(KEYINPUT78), .B(n800), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n803) );
  XNOR2_X1 U892 ( .A(n803), .B(KEYINPUT79), .ZN(n843) );
  XNOR2_X1 U893 ( .A(n804), .B(n843), .ZN(n908) );
  XNOR2_X1 U894 ( .A(n841), .B(n908), .ZN(n805) );
  NAND2_X1 U895 ( .A1(n805), .A2(G868), .ZN(n808) );
  NAND2_X1 U896 ( .A1(n806), .A2(n843), .ZN(n807) );
  NAND2_X1 U897 ( .A1(n808), .A2(n807), .ZN(G295) );
  NAND2_X1 U898 ( .A1(G2078), .A2(G2084), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n809) );
  XNOR2_X1 U900 ( .A(n810), .B(n809), .ZN(n811) );
  NAND2_X1 U901 ( .A1(G2090), .A2(n811), .ZN(n812) );
  XNOR2_X1 U902 ( .A(KEYINPUT21), .B(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n813), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U904 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U905 ( .A1(G235), .A2(G236), .ZN(n814) );
  XOR2_X1 U906 ( .A(KEYINPUT88), .B(n814), .Z(n815) );
  NOR2_X1 U907 ( .A1(G238), .A2(n815), .ZN(n816) );
  NAND2_X1 U908 ( .A1(G57), .A2(n816), .ZN(n839) );
  NAND2_X1 U909 ( .A1(G567), .A2(n839), .ZN(n822) );
  NOR2_X1 U910 ( .A1(G220), .A2(G219), .ZN(n817) );
  XNOR2_X1 U911 ( .A(KEYINPUT22), .B(n817), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n818), .A2(G96), .ZN(n819) );
  NOR2_X1 U913 ( .A1(n819), .A2(G218), .ZN(n820) );
  XNOR2_X1 U914 ( .A(n820), .B(KEYINPUT87), .ZN(n840) );
  NAND2_X1 U915 ( .A1(G2106), .A2(n840), .ZN(n821) );
  NAND2_X1 U916 ( .A1(n822), .A2(n821), .ZN(n845) );
  NAND2_X1 U917 ( .A1(G661), .A2(G483), .ZN(n823) );
  XOR2_X1 U918 ( .A(KEYINPUT89), .B(n823), .Z(n824) );
  NOR2_X1 U919 ( .A1(n845), .A2(n824), .ZN(n825) );
  XNOR2_X1 U920 ( .A(KEYINPUT90), .B(n825), .ZN(n838) );
  NAND2_X1 U921 ( .A1(G36), .A2(n838), .ZN(G176) );
  XNOR2_X1 U922 ( .A(G1341), .B(G2454), .ZN(n826) );
  XNOR2_X1 U923 ( .A(n826), .B(G2430), .ZN(n827) );
  XNOR2_X1 U924 ( .A(n827), .B(G1348), .ZN(n833) );
  XOR2_X1 U925 ( .A(G2443), .B(G2427), .Z(n829) );
  XNOR2_X1 U926 ( .A(G2438), .B(G2446), .ZN(n828) );
  XNOR2_X1 U927 ( .A(n829), .B(n828), .ZN(n831) );
  XOR2_X1 U928 ( .A(G2451), .B(G2435), .Z(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(n832) );
  XNOR2_X1 U930 ( .A(n833), .B(n832), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n834), .A2(G14), .ZN(n912) );
  XNOR2_X1 U932 ( .A(KEYINPUT111), .B(n912), .ZN(G401) );
  NAND2_X1 U933 ( .A1(G2106), .A2(n835), .ZN(G217) );
  AND2_X1 U934 ( .A1(G15), .A2(G2), .ZN(n836) );
  NAND2_X1 U935 ( .A1(G661), .A2(n836), .ZN(G259) );
  NAND2_X1 U936 ( .A1(G3), .A2(G1), .ZN(n837) );
  NAND2_X1 U937 ( .A1(n838), .A2(n837), .ZN(G188) );
  INV_X1 U939 ( .A(G96), .ZN(G221) );
  NOR2_X1 U940 ( .A1(n840), .A2(n839), .ZN(G325) );
  INV_X1 U941 ( .A(G325), .ZN(G261) );
  NAND2_X1 U942 ( .A1(n842), .A2(n841), .ZN(n844) );
  XNOR2_X1 U943 ( .A(n844), .B(n843), .ZN(G145) );
  XOR2_X1 U944 ( .A(KEYINPUT112), .B(n845), .Z(G319) );
  XOR2_X1 U945 ( .A(G2096), .B(G2100), .Z(n847) );
  XNOR2_X1 U946 ( .A(KEYINPUT42), .B(G2678), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n847), .B(n846), .ZN(n851) );
  XOR2_X1 U948 ( .A(KEYINPUT43), .B(G2072), .Z(n849) );
  XNOR2_X1 U949 ( .A(G2067), .B(G2090), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(n850) );
  XOR2_X1 U951 ( .A(n851), .B(n850), .Z(n853) );
  XNOR2_X1 U952 ( .A(G2078), .B(G2084), .ZN(n852) );
  XNOR2_X1 U953 ( .A(n853), .B(n852), .ZN(G227) );
  XOR2_X1 U954 ( .A(G1976), .B(G1971), .Z(n855) );
  XNOR2_X1 U955 ( .A(G1986), .B(G1956), .ZN(n854) );
  XNOR2_X1 U956 ( .A(n855), .B(n854), .ZN(n856) );
  XOR2_X1 U957 ( .A(n856), .B(G2474), .Z(n858) );
  XNOR2_X1 U958 ( .A(G1966), .B(G1961), .ZN(n857) );
  XNOR2_X1 U959 ( .A(n858), .B(n857), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT41), .B(G1981), .Z(n860) );
  XNOR2_X1 U961 ( .A(G1996), .B(G1991), .ZN(n859) );
  XNOR2_X1 U962 ( .A(n860), .B(n859), .ZN(n861) );
  XNOR2_X1 U963 ( .A(n862), .B(n861), .ZN(G229) );
  NAND2_X1 U964 ( .A1(G136), .A2(n887), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G112), .A2(n882), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n870) );
  NAND2_X1 U967 ( .A1(G124), .A2(n883), .ZN(n865) );
  XNOR2_X1 U968 ( .A(n865), .B(KEYINPUT44), .ZN(n868) );
  NAND2_X1 U969 ( .A1(G100), .A2(n886), .ZN(n866) );
  XOR2_X1 U970 ( .A(KEYINPUT113), .B(n866), .Z(n867) );
  NAND2_X1 U971 ( .A1(n868), .A2(n867), .ZN(n869) );
  NOR2_X1 U972 ( .A1(n870), .A2(n869), .ZN(G162) );
  NAND2_X1 U973 ( .A1(G103), .A2(n886), .ZN(n872) );
  NAND2_X1 U974 ( .A1(G139), .A2(n887), .ZN(n871) );
  NAND2_X1 U975 ( .A1(n872), .A2(n871), .ZN(n878) );
  NAND2_X1 U976 ( .A1(n882), .A2(G115), .ZN(n873) );
  XNOR2_X1 U977 ( .A(n873), .B(KEYINPUT116), .ZN(n875) );
  NAND2_X1 U978 ( .A1(G127), .A2(n883), .ZN(n874) );
  NAND2_X1 U979 ( .A1(n875), .A2(n874), .ZN(n876) );
  XOR2_X1 U980 ( .A(KEYINPUT47), .B(n876), .Z(n877) );
  NOR2_X1 U981 ( .A1(n878), .A2(n877), .ZN(n940) );
  XOR2_X1 U982 ( .A(n940), .B(n950), .Z(n881) );
  XNOR2_X1 U983 ( .A(G160), .B(n879), .ZN(n880) );
  XNOR2_X1 U984 ( .A(n881), .B(n880), .ZN(n895) );
  NAND2_X1 U985 ( .A1(G118), .A2(n882), .ZN(n885) );
  NAND2_X1 U986 ( .A1(G130), .A2(n883), .ZN(n884) );
  NAND2_X1 U987 ( .A1(n885), .A2(n884), .ZN(n893) );
  NAND2_X1 U988 ( .A1(G106), .A2(n886), .ZN(n889) );
  NAND2_X1 U989 ( .A1(G142), .A2(n887), .ZN(n888) );
  NAND2_X1 U990 ( .A1(n889), .A2(n888), .ZN(n890) );
  XOR2_X1 U991 ( .A(KEYINPUT114), .B(n890), .Z(n891) );
  XNOR2_X1 U992 ( .A(KEYINPUT45), .B(n891), .ZN(n892) );
  NOR2_X1 U993 ( .A1(n893), .A2(n892), .ZN(n894) );
  XOR2_X1 U994 ( .A(n895), .B(n894), .Z(n898) );
  XNOR2_X1 U995 ( .A(n896), .B(G162), .ZN(n897) );
  XNOR2_X1 U996 ( .A(n898), .B(n897), .ZN(n904) );
  XNOR2_X1 U997 ( .A(KEYINPUT46), .B(KEYINPUT115), .ZN(n901) );
  XNOR2_X1 U998 ( .A(n899), .B(KEYINPUT48), .ZN(n900) );
  XNOR2_X1 U999 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1000 ( .A(G164), .B(n902), .Z(n903) );
  XNOR2_X1 U1001 ( .A(n904), .B(n903), .ZN(n905) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n905), .ZN(G395) );
  XOR2_X1 U1003 ( .A(KEYINPUT117), .B(G286), .Z(n907) );
  XNOR2_X1 U1004 ( .A(G171), .B(n997), .ZN(n906) );
  XNOR2_X1 U1005 ( .A(n907), .B(n906), .ZN(n910) );
  XNOR2_X1 U1006 ( .A(n1008), .B(n908), .ZN(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  NOR2_X1 U1008 ( .A1(G37), .A2(n911), .ZN(G397) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n912), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G57), .ZN(G237) );
  XOR2_X1 U1017 ( .A(G2090), .B(G35), .Z(n920) );
  XOR2_X1 U1018 ( .A(KEYINPUT54), .B(G34), .Z(n918) );
  XNOR2_X1 U1019 ( .A(G2084), .B(n918), .ZN(n919) );
  NAND2_X1 U1020 ( .A1(n920), .A2(n919), .ZN(n934) );
  XNOR2_X1 U1021 ( .A(G2067), .B(G26), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(G1996), .B(G32), .ZN(n921) );
  NOR2_X1 U1023 ( .A1(n922), .A2(n921), .ZN(n928) );
  XOR2_X1 U1024 ( .A(G2072), .B(G33), .Z(n923) );
  NAND2_X1 U1025 ( .A1(n923), .A2(G28), .ZN(n926) );
  XNOR2_X1 U1026 ( .A(G25), .B(n924), .ZN(n925) );
  NOR2_X1 U1027 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n931) );
  XOR2_X1 U1029 ( .A(G27), .B(n929), .Z(n930) );
  NOR2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT53), .ZN(n933) );
  NOR2_X1 U1032 ( .A1(n934), .A2(n933), .ZN(n935) );
  XNOR2_X1 U1033 ( .A(KEYINPUT55), .B(n935), .ZN(n937) );
  INV_X1 U1034 ( .A(G29), .ZN(n936) );
  NAND2_X1 U1035 ( .A1(n937), .A2(n936), .ZN(n938) );
  NAND2_X1 U1036 ( .A1(n938), .A2(G11), .ZN(n939) );
  XNOR2_X1 U1037 ( .A(n939), .B(KEYINPUT119), .ZN(n967) );
  XOR2_X1 U1038 ( .A(G2072), .B(n940), .Z(n942) );
  XOR2_X1 U1039 ( .A(G164), .B(G2078), .Z(n941) );
  NOR2_X1 U1040 ( .A1(n942), .A2(n941), .ZN(n943) );
  XNOR2_X1 U1041 ( .A(KEYINPUT50), .B(n943), .ZN(n948) );
  XOR2_X1 U1042 ( .A(G2090), .B(G162), .Z(n944) );
  NOR2_X1 U1043 ( .A1(n945), .A2(n944), .ZN(n946) );
  XOR2_X1 U1044 ( .A(KEYINPUT51), .B(n946), .Z(n947) );
  NAND2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n961) );
  XOR2_X1 U1046 ( .A(G160), .B(G2084), .Z(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n954) );
  NOR2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  NOR2_X1 U1050 ( .A1(n956), .A2(n955), .ZN(n957) );
  XNOR2_X1 U1051 ( .A(n957), .B(KEYINPUT118), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  NOR2_X1 U1053 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(KEYINPUT52), .B(n962), .ZN(n964) );
  INV_X1 U1055 ( .A(KEYINPUT55), .ZN(n963) );
  NAND2_X1 U1056 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1057 ( .A1(n965), .A2(G29), .ZN(n966) );
  NAND2_X1 U1058 ( .A1(n967), .A2(n966), .ZN(n1022) );
  XNOR2_X1 U1059 ( .A(n968), .B(G5), .ZN(n989) );
  XOR2_X1 U1060 ( .A(G1966), .B(G21), .Z(n977) );
  XOR2_X1 U1061 ( .A(G1986), .B(G24), .Z(n971) );
  XOR2_X1 U1062 ( .A(G22), .B(KEYINPUT122), .Z(n969) );
  XNOR2_X1 U1063 ( .A(n969), .B(G1971), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n974) );
  XOR2_X1 U1065 ( .A(KEYINPUT123), .B(G1976), .Z(n972) );
  XNOR2_X1 U1066 ( .A(G23), .B(n972), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n975) );
  XNOR2_X1 U1068 ( .A(KEYINPUT58), .B(n975), .ZN(n976) );
  NAND2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n987) );
  XOR2_X1 U1070 ( .A(G1348), .B(KEYINPUT59), .Z(n978) );
  XNOR2_X1 U1071 ( .A(G4), .B(n978), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(G20), .B(G1956), .ZN(n979) );
  NOR2_X1 U1073 ( .A1(n980), .A2(n979), .ZN(n984) );
  XNOR2_X1 U1074 ( .A(G1981), .B(G6), .ZN(n982) );
  XNOR2_X1 U1075 ( .A(G1341), .B(G19), .ZN(n981) );
  NOR2_X1 U1076 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1077 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1078 ( .A(KEYINPUT60), .B(n985), .ZN(n986) );
  NOR2_X1 U1079 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1080 ( .A1(n989), .A2(n988), .ZN(n990) );
  XNOR2_X1 U1081 ( .A(n990), .B(KEYINPUT61), .ZN(n991) );
  XNOR2_X1 U1082 ( .A(n991), .B(KEYINPUT124), .ZN(n992) );
  NOR2_X1 U1083 ( .A1(G16), .A2(n992), .ZN(n1019) );
  XOR2_X1 U1084 ( .A(G16), .B(KEYINPUT56), .Z(n1017) );
  NAND2_X1 U1085 ( .A1(n994), .A2(n993), .ZN(n996) );
  XNOR2_X1 U1086 ( .A(G1956), .B(G299), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n1014) );
  XNOR2_X1 U1088 ( .A(G1348), .B(n997), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(G1961), .B(G171), .ZN(n999) );
  NAND2_X1 U1090 ( .A1(G1971), .A2(G303), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NOR2_X1 U1092 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G1966), .B(G168), .ZN(n1004) );
  XNOR2_X1 U1095 ( .A(n1004), .B(KEYINPUT120), .ZN(n1006) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(n1007), .B(KEYINPUT57), .ZN(n1010) );
  XOR2_X1 U1098 ( .A(G1341), .B(n1008), .Z(n1009) );
  NAND2_X1 U1099 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NOR2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(n1015), .B(KEYINPUT121), .ZN(n1016) );
  NOR2_X1 U1103 ( .A1(n1017), .A2(n1016), .ZN(n1018) );
  NOR2_X1 U1104 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  XNOR2_X1 U1105 ( .A(n1020), .B(KEYINPUT125), .ZN(n1021) );
  NOR2_X1 U1106 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  XNOR2_X1 U1107 ( .A(n1023), .B(KEYINPUT62), .ZN(n1024) );
  XNOR2_X1 U1108 ( .A(n1024), .B(KEYINPUT126), .ZN(G311) );
  XNOR2_X1 U1109 ( .A(KEYINPUT127), .B(G311), .ZN(G150) );
endmodule

