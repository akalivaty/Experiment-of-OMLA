

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587;

  AND2_X1 U324 ( .A1(n388), .A2(n387), .ZN(n389) );
  XOR2_X1 U325 ( .A(n553), .B(KEYINPUT36), .Z(n584) );
  AND2_X1 U326 ( .A1(n576), .A2(n391), .ZN(n292) );
  XOR2_X1 U327 ( .A(n375), .B(n374), .Z(n293) );
  NOR2_X1 U328 ( .A1(n533), .A2(n453), .ZN(n562) );
  XNOR2_X1 U329 ( .A(KEYINPUT46), .B(KEYINPUT107), .ZN(n349) );
  XNOR2_X1 U330 ( .A(n350), .B(n349), .ZN(n369) );
  XNOR2_X1 U331 ( .A(n315), .B(n314), .ZN(n316) );
  INV_X1 U332 ( .A(n553), .ZN(n387) );
  AND2_X1 U333 ( .A1(n392), .A2(n292), .ZN(n393) );
  XNOR2_X1 U334 ( .A(KEYINPUT48), .B(KEYINPUT110), .ZN(n396) );
  XNOR2_X1 U335 ( .A(n398), .B(n363), .ZN(n328) );
  XNOR2_X1 U336 ( .A(n293), .B(n376), .ZN(n377) );
  XNOR2_X1 U337 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U338 ( .A(n378), .B(n377), .ZN(n382) );
  INV_X1 U339 ( .A(n330), .ZN(n576) );
  XOR2_X1 U340 ( .A(n386), .B(n385), .Z(n553) );
  XNOR2_X1 U341 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n456) );
  XNOR2_X1 U342 ( .A(n457), .B(n456), .ZN(G1351GAT) );
  XNOR2_X1 U343 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n294), .B(KEYINPUT17), .ZN(n295) );
  XOR2_X1 U345 ( .A(n295), .B(KEYINPUT83), .Z(n297) );
  XNOR2_X1 U346 ( .A(G169GAT), .B(G183GAT), .ZN(n296) );
  XNOR2_X1 U347 ( .A(n297), .B(n296), .ZN(n409) );
  XOR2_X1 U348 ( .A(KEYINPUT82), .B(KEYINPUT20), .Z(n299) );
  XNOR2_X1 U349 ( .A(G43GAT), .B(G99GAT), .ZN(n298) );
  XNOR2_X1 U350 ( .A(n299), .B(n298), .ZN(n300) );
  XNOR2_X1 U351 ( .A(n300), .B(G176GAT), .ZN(n304) );
  XOR2_X1 U352 ( .A(G113GAT), .B(KEYINPUT0), .Z(n419) );
  XOR2_X1 U353 ( .A(G120GAT), .B(G71GAT), .Z(n309) );
  XOR2_X1 U354 ( .A(n419), .B(n309), .Z(n302) );
  NAND2_X1 U355 ( .A1(G227GAT), .A2(G233GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X1 U358 ( .A(G15GAT), .B(G127GAT), .Z(n356) );
  XOR2_X1 U359 ( .A(n305), .B(n356), .Z(n307) );
  XNOR2_X1 U360 ( .A(G134GAT), .B(G190GAT), .ZN(n306) );
  XNOR2_X1 U361 ( .A(n307), .B(n306), .ZN(n308) );
  XNOR2_X1 U362 ( .A(n409), .B(n308), .ZN(n533) );
  XOR2_X2 U363 ( .A(G99GAT), .B(G85GAT), .Z(n371) );
  XOR2_X1 U364 ( .A(KEYINPUT71), .B(n371), .Z(n311) );
  XNOR2_X1 U365 ( .A(n309), .B(G204GAT), .ZN(n310) );
  XNOR2_X1 U366 ( .A(n311), .B(n310), .ZN(n317) );
  XOR2_X1 U367 ( .A(KEYINPUT70), .B(KEYINPUT33), .Z(n313) );
  XNOR2_X1 U368 ( .A(KEYINPUT31), .B(KEYINPUT32), .ZN(n312) );
  XOR2_X1 U369 ( .A(n313), .B(n312), .Z(n315) );
  NAND2_X1 U370 ( .A1(G230GAT), .A2(G233GAT), .ZN(n314) );
  XNOR2_X1 U371 ( .A(n317), .B(n316), .ZN(n320) );
  INV_X1 U372 ( .A(n320), .ZN(n318) );
  NAND2_X1 U373 ( .A1(n318), .A2(KEYINPUT72), .ZN(n322) );
  INV_X1 U374 ( .A(KEYINPUT72), .ZN(n319) );
  NAND2_X1 U375 ( .A1(n320), .A2(n319), .ZN(n321) );
  NAND2_X1 U376 ( .A1(n322), .A2(n321), .ZN(n325) );
  XNOR2_X1 U377 ( .A(G106GAT), .B(G78GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n323), .B(G148GAT), .ZN(n439) );
  XNOR2_X1 U379 ( .A(n439), .B(KEYINPUT69), .ZN(n324) );
  XNOR2_X1 U380 ( .A(n325), .B(n324), .ZN(n329) );
  XOR2_X1 U381 ( .A(G176GAT), .B(G92GAT), .Z(n326) );
  XOR2_X1 U382 ( .A(G64GAT), .B(n326), .Z(n398) );
  XNOR2_X1 U383 ( .A(G57GAT), .B(KEYINPUT68), .ZN(n327) );
  XNOR2_X1 U384 ( .A(n327), .B(KEYINPUT13), .ZN(n363) );
  XNOR2_X1 U385 ( .A(KEYINPUT41), .B(n576), .ZN(n563) );
  XOR2_X1 U386 ( .A(KEYINPUT66), .B(G141GAT), .Z(n332) );
  XNOR2_X1 U387 ( .A(G15GAT), .B(G197GAT), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n332), .B(n331), .ZN(n336) );
  XOR2_X1 U389 ( .A(KEYINPUT67), .B(KEYINPUT65), .Z(n334) );
  XNOR2_X1 U390 ( .A(KEYINPUT64), .B(KEYINPUT30), .ZN(n333) );
  XNOR2_X1 U391 ( .A(n334), .B(n333), .ZN(n335) );
  XNOR2_X1 U392 ( .A(n336), .B(n335), .ZN(n348) );
  XNOR2_X1 U393 ( .A(G113GAT), .B(G36GAT), .ZN(n337) );
  XNOR2_X1 U394 ( .A(n337), .B(G50GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(G22GAT), .B(G1GAT), .ZN(n338) );
  XNOR2_X1 U396 ( .A(n338), .B(G8GAT), .ZN(n364) );
  XOR2_X1 U397 ( .A(n339), .B(n364), .Z(n346) );
  XOR2_X1 U398 ( .A(G29GAT), .B(G43GAT), .Z(n341) );
  XNOR2_X1 U399 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n340) );
  XNOR2_X1 U400 ( .A(n341), .B(n340), .ZN(n384) );
  XOR2_X1 U401 ( .A(n384), .B(KEYINPUT29), .Z(n343) );
  NAND2_X1 U402 ( .A1(G229GAT), .A2(G233GAT), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XNOR2_X1 U404 ( .A(G169GAT), .B(n344), .ZN(n345) );
  XNOR2_X1 U405 ( .A(n346), .B(n345), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n573) );
  NAND2_X1 U407 ( .A1(n563), .A2(n573), .ZN(n350) );
  XOR2_X1 U408 ( .A(G64GAT), .B(KEYINPUT12), .Z(n352) );
  XNOR2_X1 U409 ( .A(G155GAT), .B(KEYINPUT14), .ZN(n351) );
  XNOR2_X1 U410 ( .A(n352), .B(n351), .ZN(n368) );
  XOR2_X1 U411 ( .A(G78GAT), .B(G211GAT), .Z(n354) );
  XNOR2_X1 U412 ( .A(G183GAT), .B(G71GAT), .ZN(n353) );
  XNOR2_X1 U413 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U414 ( .A(n356), .B(n355), .Z(n358) );
  NAND2_X1 U415 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n362) );
  XOR2_X1 U417 ( .A(KEYINPUT15), .B(KEYINPUT81), .Z(n360) );
  XNOR2_X1 U418 ( .A(KEYINPUT80), .B(KEYINPUT79), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U420 ( .A(n362), .B(n361), .Z(n366) );
  XNOR2_X1 U421 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U422 ( .A(n366), .B(n365), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n368), .B(n367), .ZN(n487) );
  INV_X1 U424 ( .A(n487), .ZN(n579) );
  NOR2_X1 U425 ( .A1(n369), .A2(n579), .ZN(n370) );
  XNOR2_X1 U426 ( .A(n370), .B(KEYINPUT108), .ZN(n388) );
  XOR2_X1 U427 ( .A(KEYINPUT11), .B(n371), .Z(n373) );
  XOR2_X1 U428 ( .A(G36GAT), .B(G190GAT), .Z(n399) );
  XNOR2_X1 U429 ( .A(G218GAT), .B(n399), .ZN(n372) );
  XNOR2_X1 U430 ( .A(n373), .B(n372), .ZN(n378) );
  XOR2_X1 U431 ( .A(KEYINPUT76), .B(G92GAT), .Z(n375) );
  NAND2_X1 U432 ( .A1(G232GAT), .A2(G233GAT), .ZN(n374) );
  XOR2_X1 U433 ( .A(G134GAT), .B(KEYINPUT77), .Z(n418) );
  XNOR2_X1 U434 ( .A(G106GAT), .B(n418), .ZN(n376) );
  XOR2_X1 U435 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n380) );
  XNOR2_X1 U436 ( .A(KEYINPUT9), .B(KEYINPUT10), .ZN(n379) );
  XNOR2_X1 U437 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U438 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U439 ( .A(G50GAT), .B(KEYINPUT74), .ZN(n383) );
  XNOR2_X1 U440 ( .A(n383), .B(G162GAT), .ZN(n442) );
  XNOR2_X1 U441 ( .A(n384), .B(n442), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n389), .B(KEYINPUT47), .ZN(n395) );
  NOR2_X1 U443 ( .A1(n487), .A2(n584), .ZN(n390) );
  XNOR2_X1 U444 ( .A(n390), .B(KEYINPUT45), .ZN(n392) );
  INV_X1 U445 ( .A(n573), .ZN(n391) );
  XNOR2_X1 U446 ( .A(KEYINPUT109), .B(n393), .ZN(n394) );
  AND2_X1 U447 ( .A1(n395), .A2(n394), .ZN(n397) );
  XNOR2_X1 U448 ( .A(n397), .B(n396), .ZN(n529) );
  XOR2_X1 U449 ( .A(KEYINPUT89), .B(n398), .Z(n401) );
  XNOR2_X1 U450 ( .A(G8GAT), .B(n399), .ZN(n400) );
  XNOR2_X1 U451 ( .A(n401), .B(n400), .ZN(n413) );
  XOR2_X1 U452 ( .A(KEYINPUT92), .B(KEYINPUT90), .Z(n403) );
  NAND2_X1 U453 ( .A1(G226GAT), .A2(G233GAT), .ZN(n402) );
  XNOR2_X1 U454 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U455 ( .A(n404), .B(KEYINPUT91), .Z(n411) );
  XNOR2_X1 U456 ( .A(G211GAT), .B(G218GAT), .ZN(n405) );
  XNOR2_X1 U457 ( .A(n405), .B(KEYINPUT21), .ZN(n406) );
  XOR2_X1 U458 ( .A(n406), .B(KEYINPUT85), .Z(n408) );
  XNOR2_X1 U459 ( .A(G197GAT), .B(G204GAT), .ZN(n407) );
  XNOR2_X1 U460 ( .A(n408), .B(n407), .ZN(n451) );
  XNOR2_X1 U461 ( .A(n409), .B(n451), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n412) );
  XOR2_X1 U463 ( .A(n413), .B(n412), .Z(n463) );
  NOR2_X1 U464 ( .A1(n529), .A2(n463), .ZN(n415) );
  INV_X1 U465 ( .A(KEYINPUT54), .ZN(n414) );
  XNOR2_X1 U466 ( .A(n415), .B(n414), .ZN(n438) );
  XOR2_X1 U467 ( .A(KEYINPUT5), .B(KEYINPUT1), .Z(n417) );
  XNOR2_X1 U468 ( .A(KEYINPUT87), .B(KEYINPUT6), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n417), .B(n416), .ZN(n423) );
  XOR2_X1 U470 ( .A(G85GAT), .B(n418), .Z(n421) );
  XNOR2_X1 U471 ( .A(n419), .B(G162GAT), .ZN(n420) );
  XNOR2_X1 U472 ( .A(n421), .B(n420), .ZN(n422) );
  XOR2_X1 U473 ( .A(n423), .B(n422), .Z(n425) );
  NAND2_X1 U474 ( .A1(G225GAT), .A2(G233GAT), .ZN(n424) );
  XNOR2_X1 U475 ( .A(n425), .B(n424), .ZN(n429) );
  XOR2_X1 U476 ( .A(G148GAT), .B(G120GAT), .Z(n427) );
  XNOR2_X1 U477 ( .A(G29GAT), .B(G127GAT), .ZN(n426) );
  XNOR2_X1 U478 ( .A(n427), .B(n426), .ZN(n428) );
  XOR2_X1 U479 ( .A(n429), .B(n428), .Z(n437) );
  XOR2_X1 U480 ( .A(KEYINPUT2), .B(KEYINPUT86), .Z(n431) );
  XNOR2_X1 U481 ( .A(KEYINPUT3), .B(G155GAT), .ZN(n430) );
  XNOR2_X1 U482 ( .A(n431), .B(n430), .ZN(n432) );
  XOR2_X1 U483 ( .A(G141GAT), .B(n432), .Z(n447) );
  XOR2_X1 U484 ( .A(KEYINPUT4), .B(G57GAT), .Z(n434) );
  XNOR2_X1 U485 ( .A(G1GAT), .B(KEYINPUT88), .ZN(n433) );
  XNOR2_X1 U486 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U487 ( .A(n447), .B(n435), .ZN(n436) );
  XNOR2_X1 U488 ( .A(n437), .B(n436), .ZN(n516) );
  NOR2_X1 U489 ( .A1(n438), .A2(n516), .ZN(n571) );
  XOR2_X1 U490 ( .A(KEYINPUT84), .B(KEYINPUT24), .Z(n441) );
  XNOR2_X1 U491 ( .A(KEYINPUT23), .B(n439), .ZN(n440) );
  XNOR2_X1 U492 ( .A(n441), .B(n440), .ZN(n446) );
  XOR2_X1 U493 ( .A(n442), .B(KEYINPUT22), .Z(n444) );
  NAND2_X1 U494 ( .A1(G228GAT), .A2(G233GAT), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n445) );
  XOR2_X1 U496 ( .A(n446), .B(n445), .Z(n449) );
  XNOR2_X1 U497 ( .A(G22GAT), .B(n447), .ZN(n448) );
  XNOR2_X1 U498 ( .A(n449), .B(n448), .ZN(n450) );
  XNOR2_X1 U499 ( .A(n451), .B(n450), .ZN(n470) );
  AND2_X1 U500 ( .A1(n571), .A2(n470), .ZN(n452) );
  XNOR2_X1 U501 ( .A(n452), .B(KEYINPUT55), .ZN(n453) );
  NAND2_X1 U502 ( .A1(n562), .A2(n573), .ZN(n455) );
  XNOR2_X1 U503 ( .A(G169GAT), .B(KEYINPUT118), .ZN(n454) );
  XNOR2_X1 U504 ( .A(n455), .B(n454), .ZN(G1348GAT) );
  NAND2_X1 U505 ( .A1(n553), .A2(n562), .ZN(n457) );
  XNOR2_X1 U506 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n478) );
  NAND2_X1 U507 ( .A1(n576), .A2(n573), .ZN(n458) );
  XOR2_X1 U508 ( .A(KEYINPUT73), .B(n458), .Z(n491) );
  NOR2_X1 U509 ( .A1(n553), .A2(n487), .ZN(n459) );
  XNOR2_X1 U510 ( .A(n459), .B(KEYINPUT16), .ZN(n476) );
  INV_X1 U511 ( .A(n533), .ZN(n520) );
  NOR2_X1 U512 ( .A1(n520), .A2(n470), .ZN(n461) );
  XNOR2_X1 U513 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n460) );
  XOR2_X1 U514 ( .A(n461), .B(n460), .Z(n572) );
  XNOR2_X1 U515 ( .A(n463), .B(KEYINPUT93), .ZN(n462) );
  XNOR2_X1 U516 ( .A(n462), .B(KEYINPUT27), .ZN(n471) );
  NAND2_X1 U517 ( .A1(n572), .A2(n471), .ZN(n467) );
  INV_X1 U518 ( .A(n463), .ZN(n518) );
  NAND2_X1 U519 ( .A1(n520), .A2(n518), .ZN(n464) );
  NAND2_X1 U520 ( .A1(n470), .A2(n464), .ZN(n465) );
  XOR2_X1 U521 ( .A(KEYINPUT25), .B(n465), .Z(n466) );
  NAND2_X1 U522 ( .A1(n467), .A2(n466), .ZN(n469) );
  INV_X1 U523 ( .A(n516), .ZN(n468) );
  NAND2_X1 U524 ( .A1(n469), .A2(n468), .ZN(n475) );
  XNOR2_X1 U525 ( .A(KEYINPUT28), .B(n470), .ZN(n531) );
  NAND2_X1 U526 ( .A1(n471), .A2(n516), .ZN(n472) );
  XNOR2_X1 U527 ( .A(n472), .B(KEYINPUT94), .ZN(n528) );
  NOR2_X1 U528 ( .A1(n528), .A2(n520), .ZN(n473) );
  NAND2_X1 U529 ( .A1(n531), .A2(n473), .ZN(n474) );
  NAND2_X1 U530 ( .A1(n475), .A2(n474), .ZN(n486) );
  NAND2_X1 U531 ( .A1(n476), .A2(n486), .ZN(n501) );
  NOR2_X1 U532 ( .A1(n491), .A2(n501), .ZN(n483) );
  NAND2_X1 U533 ( .A1(n516), .A2(n483), .ZN(n477) );
  XNOR2_X1 U534 ( .A(n478), .B(n477), .ZN(G1324GAT) );
  NAND2_X1 U535 ( .A1(n518), .A2(n483), .ZN(n479) );
  XNOR2_X1 U536 ( .A(n479), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT96), .B(KEYINPUT35), .Z(n481) );
  NAND2_X1 U538 ( .A1(n483), .A2(n520), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G15GAT), .B(n482), .ZN(G1326GAT) );
  XOR2_X1 U541 ( .A(G22GAT), .B(KEYINPUT97), .Z(n485) );
  INV_X1 U542 ( .A(n531), .ZN(n522) );
  NAND2_X1 U543 ( .A1(n483), .A2(n522), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(G1327GAT) );
  XOR2_X1 U545 ( .A(G29GAT), .B(KEYINPUT39), .Z(n494) );
  NAND2_X1 U546 ( .A1(n487), .A2(n486), .ZN(n488) );
  XNOR2_X1 U547 ( .A(KEYINPUT98), .B(n488), .ZN(n489) );
  NOR2_X1 U548 ( .A1(n584), .A2(n489), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT37), .B(n490), .ZN(n514) );
  NOR2_X1 U550 ( .A1(n491), .A2(n514), .ZN(n492) );
  XNOR2_X1 U551 ( .A(n492), .B(KEYINPUT38), .ZN(n498) );
  NAND2_X1 U552 ( .A1(n516), .A2(n498), .ZN(n493) );
  XNOR2_X1 U553 ( .A(n494), .B(n493), .ZN(G1328GAT) );
  NAND2_X1 U554 ( .A1(n498), .A2(n518), .ZN(n495) );
  XNOR2_X1 U555 ( .A(n495), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U556 ( .A1(n498), .A2(n520), .ZN(n496) );
  XNOR2_X1 U557 ( .A(n496), .B(KEYINPUT40), .ZN(n497) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NAND2_X1 U559 ( .A1(n522), .A2(n498), .ZN(n499) );
  XNOR2_X1 U560 ( .A(G50GAT), .B(n499), .ZN(G1331GAT) );
  NAND2_X1 U561 ( .A1(n391), .A2(n563), .ZN(n500) );
  XNOR2_X1 U562 ( .A(n500), .B(KEYINPUT100), .ZN(n515) );
  NOR2_X1 U563 ( .A1(n515), .A2(n501), .ZN(n502) );
  XOR2_X1 U564 ( .A(KEYINPUT101), .B(n502), .Z(n509) );
  NAND2_X1 U565 ( .A1(n509), .A2(n516), .ZN(n506) );
  XOR2_X1 U566 ( .A(KEYINPUT102), .B(KEYINPUT42), .Z(n504) );
  XNOR2_X1 U567 ( .A(G57GAT), .B(KEYINPUT99), .ZN(n503) );
  XNOR2_X1 U568 ( .A(n504), .B(n503), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(G1332GAT) );
  NAND2_X1 U570 ( .A1(n518), .A2(n509), .ZN(n507) );
  XNOR2_X1 U571 ( .A(n507), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U572 ( .A1(n509), .A2(n520), .ZN(n508) );
  XNOR2_X1 U573 ( .A(n508), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT104), .B(KEYINPUT43), .Z(n511) );
  NAND2_X1 U575 ( .A1(n509), .A2(n522), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(n513) );
  XOR2_X1 U577 ( .A(G78GAT), .B(KEYINPUT103), .Z(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NOR2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n523) );
  NAND2_X1 U580 ( .A1(n523), .A2(n516), .ZN(n517) );
  XNOR2_X1 U581 ( .A(n517), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U582 ( .A1(n518), .A2(n523), .ZN(n519) );
  XNOR2_X1 U583 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U584 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U586 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n527) );
  XOR2_X1 U587 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n525) );
  NAND2_X1 U588 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U589 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U590 ( .A(n527), .B(n526), .ZN(G1339GAT) );
  NOR2_X1 U591 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U592 ( .A(KEYINPUT111), .B(n530), .Z(n547) );
  NAND2_X1 U593 ( .A1(n547), .A2(n531), .ZN(n532) );
  NOR2_X1 U594 ( .A1(n533), .A2(n532), .ZN(n544) );
  NAND2_X1 U595 ( .A1(n544), .A2(n573), .ZN(n534) );
  XNOR2_X1 U596 ( .A(n534), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT49), .B(KEYINPUT113), .Z(n536) );
  NAND2_X1 U598 ( .A1(n544), .A2(n563), .ZN(n535) );
  XNOR2_X1 U599 ( .A(n536), .B(n535), .ZN(n538) );
  XOR2_X1 U600 ( .A(G120GAT), .B(KEYINPUT112), .Z(n537) );
  XNOR2_X1 U601 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  NAND2_X1 U602 ( .A1(n544), .A2(n579), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n539), .B(KEYINPUT50), .ZN(n540) );
  XNOR2_X1 U604 ( .A(G127GAT), .B(n540), .ZN(G1342GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n542) );
  XNOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U608 ( .A(KEYINPUT114), .B(n543), .Z(n546) );
  NAND2_X1 U609 ( .A1(n544), .A2(n553), .ZN(n545) );
  XNOR2_X1 U610 ( .A(n546), .B(n545), .ZN(G1343GAT) );
  AND2_X1 U611 ( .A1(n572), .A2(n547), .ZN(n554) );
  NAND2_X1 U612 ( .A1(n573), .A2(n554), .ZN(n548) );
  XNOR2_X1 U613 ( .A(G141GAT), .B(n548), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n550) );
  NAND2_X1 U615 ( .A1(n554), .A2(n563), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U618 ( .A1(n554), .A2(n579), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(G155GAT), .ZN(G1346GAT) );
  XOR2_X1 U620 ( .A(G162GAT), .B(KEYINPUT117), .Z(n556) );
  NAND2_X1 U621 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U622 ( .A(n556), .B(n555), .ZN(G1347GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT119), .B(KEYINPUT120), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XOR2_X1 U626 ( .A(n559), .B(KEYINPUT122), .Z(n561) );
  XNOR2_X1 U627 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n565) );
  NAND2_X1 U629 ( .A1(n562), .A2(n563), .ZN(n564) );
  XOR2_X1 U630 ( .A(n565), .B(n564), .Z(G1349GAT) );
  XOR2_X1 U631 ( .A(G183GAT), .B(KEYINPUT123), .Z(n567) );
  NAND2_X1 U632 ( .A1(n562), .A2(n579), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT125), .B(KEYINPUT60), .Z(n569) );
  XNOR2_X1 U635 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n570) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(n570), .Z(n575) );
  NAND2_X1 U638 ( .A1(n572), .A2(n571), .ZN(n583) );
  INV_X1 U639 ( .A(n583), .ZN(n580) );
  NAND2_X1 U640 ( .A1(n580), .A2(n573), .ZN(n574) );
  XNOR2_X1 U641 ( .A(n575), .B(n574), .ZN(G1352GAT) );
  XOR2_X1 U642 ( .A(G204GAT), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U643 ( .A1(n580), .A2(n330), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(G1353GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n581), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U647 ( .A(G211GAT), .B(n582), .ZN(G1354GAT) );
  NOR2_X1 U648 ( .A1(n584), .A2(n583), .ZN(n586) );
  XNOR2_X1 U649 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(n587) );
  XNOR2_X1 U651 ( .A(G218GAT), .B(n587), .ZN(G1355GAT) );
endmodule

