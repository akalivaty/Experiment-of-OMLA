//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 1 1 1 0 1 0 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:54 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n753, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n856, new_n857,
    new_n858, new_n859, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n899, new_n900, new_n902, new_n903,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943;
  XNOR2_X1  g000(.A(G78gat), .B(G106gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G22gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n206), .A2(KEYINPUT86), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n205), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(G228gat), .A2(G233gat), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT3), .ZN(new_n211));
  XNOR2_X1  g010(.A(G211gat), .B(G218gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT71), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(G197gat), .B(G204gat), .ZN(new_n215));
  INV_X1    g014(.A(G211gat), .ZN(new_n216));
  INV_X1    g015(.A(G218gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  OAI21_X1  g017(.A(new_n215), .B1(KEYINPUT22), .B2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n214), .B(new_n219), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n211), .B1(new_n220), .B2(KEYINPUT29), .ZN(new_n221));
  NAND2_X1  g020(.A1(G155gat), .A2(G162gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT76), .ZN(new_n223));
  NOR3_X1   g022(.A1(new_n223), .A2(G155gat), .A3(G162gat), .ZN(new_n224));
  INV_X1    g023(.A(G155gat), .ZN(new_n225));
  INV_X1    g024(.A(G162gat), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT76), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(new_n222), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT77), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G148gat), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n231), .A2(G141gat), .ZN(new_n232));
  INV_X1    g031(.A(G141gat), .ZN(new_n233));
  NOR2_X1   g032(.A1(new_n233), .A2(G148gat), .ZN(new_n234));
  INV_X1    g033(.A(new_n222), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT2), .ZN(new_n236));
  OAI22_X1  g035(.A1(new_n232), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n225), .A2(new_n226), .A3(KEYINPUT76), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n223), .B1(G155gat), .B2(G162gat), .ZN(new_n239));
  AOI21_X1  g038(.A(new_n235), .B1(new_n238), .B2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(KEYINPUT77), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n230), .A2(new_n237), .A3(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(KEYINPUT79), .B(G162gat), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n236), .B1(new_n243), .B2(G155gat), .ZN(new_n244));
  INV_X1    g043(.A(new_n244), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT78), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(new_n233), .B2(G148gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n231), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n232), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  NOR2_X1   g049(.A1(G155gat), .A2(G162gat), .ZN(new_n251));
  NOR2_X1   g050(.A1(new_n235), .A2(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n245), .A2(new_n250), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n242), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n221), .A2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(KEYINPUT84), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n210), .B1(new_n256), .B2(new_n257), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT80), .B(KEYINPUT3), .Z(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  NAND3_X1  g059(.A1(new_n242), .A2(new_n254), .A3(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT29), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n263), .A2(new_n220), .ZN(new_n264));
  NAND3_X1  g063(.A1(new_n221), .A2(KEYINPUT84), .A3(new_n255), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n258), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(KEYINPUT85), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT85), .ZN(new_n268));
  NAND4_X1  g067(.A1(new_n258), .A2(new_n268), .A3(new_n264), .A4(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g069(.A1(new_n219), .A2(new_n212), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n262), .B1(new_n219), .B2(new_n212), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n260), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n255), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n264), .A2(new_n274), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(new_n210), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n209), .B1(new_n270), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n276), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n278), .B(new_n208), .C1(new_n267), .C2(new_n269), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n277), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT30), .ZN(new_n281));
  INV_X1    g080(.A(G183gat), .ZN(new_n282));
  INV_X1    g081(.A(G190gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT24), .ZN(new_n285));
  AOI21_X1  g084(.A(new_n285), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G183gat), .A2(G190gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n284), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(G169gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  NOR2_X1   g091(.A1(KEYINPUT64), .A2(G176gat), .ZN(new_n293));
  OAI211_X1 g092(.A(KEYINPUT23), .B(new_n290), .C1(new_n292), .C2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(new_n294), .A3(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n303), .A3(new_n285), .ZN(new_n304));
  OAI211_X1 g103(.A(G183gat), .B(G190gat), .C1(KEYINPUT65), .C2(KEYINPUT24), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n304), .A2(new_n284), .A3(new_n305), .ZN(new_n306));
  AOI21_X1  g105(.A(new_n301), .B1(new_n295), .B2(KEYINPUT23), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n306), .A2(new_n299), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT66), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n306), .A2(KEYINPUT66), .A3(new_n299), .A4(new_n307), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n302), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT28), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n315));
  OR2_X1    g114(.A1(new_n314), .A2(KEYINPUT67), .ZN(new_n316));
  XNOR2_X1  g115(.A(KEYINPUT27), .B(G183gat), .ZN(new_n317));
  INV_X1    g116(.A(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n315), .B(new_n316), .C1(new_n318), .C2(G190gat), .ZN(new_n319));
  NAND4_X1  g118(.A1(new_n317), .A2(KEYINPUT67), .A3(new_n314), .A4(new_n283), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n296), .A2(KEYINPUT26), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT26), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n295), .A2(new_n322), .ZN(new_n323));
  NAND3_X1  g122(.A1(new_n321), .A2(new_n297), .A3(new_n323), .ZN(new_n324));
  NAND4_X1  g123(.A1(new_n319), .A2(new_n287), .A3(new_n320), .A4(new_n324), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n312), .A2(new_n313), .A3(new_n325), .ZN(new_n326));
  AOI22_X1  g125(.A1(new_n312), .A2(new_n325), .B1(new_n262), .B2(new_n313), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n220), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n310), .A2(new_n311), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT64), .ZN(new_n330));
  INV_X1    g129(.A(G176gat), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AOI21_X1  g131(.A(G169gat), .B1(new_n332), .B2(new_n291), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n287), .A2(KEYINPUT24), .ZN(new_n334));
  NAND3_X1  g133(.A1(new_n285), .A2(G183gat), .A3(G190gat), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  AOI22_X1  g135(.A1(KEYINPUT23), .A2(new_n333), .B1(new_n336), .B2(new_n284), .ZN(new_n337));
  AOI21_X1  g136(.A(KEYINPUT25), .B1(new_n337), .B2(new_n299), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n325), .B1(new_n329), .B2(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n313), .A2(new_n262), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n312), .A2(new_n313), .A3(new_n325), .ZN(new_n342));
  INV_X1    g141(.A(new_n220), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  NAND3_X1  g143(.A1(new_n328), .A2(KEYINPUT72), .A3(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(KEYINPUT72), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n220), .C1(new_n326), .C2(new_n327), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  XNOR2_X1  g147(.A(G8gat), .B(G36gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n349), .B(KEYINPUT73), .ZN(new_n350));
  XNOR2_X1  g149(.A(G64gat), .B(G92gat), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n350), .B(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT75), .B1(new_n348), .B2(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT75), .ZN(new_n354));
  INV_X1    g153(.A(new_n352), .ZN(new_n355));
  AOI211_X1 g154(.A(new_n354), .B(new_n355), .C1(new_n345), .C2(new_n347), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n281), .B1(new_n353), .B2(new_n356), .ZN(new_n357));
  XNOR2_X1  g156(.A(new_n352), .B(KEYINPUT74), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n348), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(new_n355), .B1(new_n345), .B2(new_n347), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n359), .B1(KEYINPUT30), .B2(new_n360), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n357), .A2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT40), .ZN(new_n363));
  NAND2_X1  g162(.A1(G225gat), .A2(G233gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(KEYINPUT68), .A2(G134gat), .ZN(new_n365));
  INV_X1    g164(.A(G120gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G113gat), .ZN(new_n367));
  INV_X1    g166(.A(G113gat), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n368), .A2(G120gat), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n367), .A2(new_n369), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT1), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n365), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  AOI211_X1 g171(.A(KEYINPUT1), .B(G134gat), .C1(new_n367), .C2(new_n369), .ZN(new_n373));
  OAI21_X1  g172(.A(G127gat), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  INV_X1    g173(.A(new_n365), .ZN(new_n375));
  XNOR2_X1  g174(.A(G113gat), .B(G120gat), .ZN(new_n376));
  OAI21_X1  g175(.A(new_n375), .B1(new_n376), .B2(KEYINPUT1), .ZN(new_n377));
  INV_X1    g176(.A(G134gat), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n370), .A2(new_n371), .A3(new_n378), .ZN(new_n379));
  INV_X1    g178(.A(G127gat), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n377), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n374), .A2(new_n381), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n382), .B1(new_n255), .B2(KEYINPUT3), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT4), .ZN(new_n384));
  INV_X1    g183(.A(new_n381), .ZN(new_n385));
  AOI21_X1  g184(.A(new_n380), .B1(new_n377), .B2(new_n379), .ZN(new_n386));
  OAI211_X1 g185(.A(new_n242), .B(new_n254), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AOI22_X1  g186(.A1(new_n383), .A2(new_n261), .B1(new_n384), .B2(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT82), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g189(.A1(new_n382), .A2(KEYINPUT82), .A3(new_n254), .A4(new_n242), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n364), .B1(new_n388), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n390), .A2(new_n391), .ZN(new_n394));
  INV_X1    g193(.A(new_n382), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n255), .ZN(new_n396));
  AND3_X1   g195(.A1(new_n394), .A2(new_n364), .A3(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT39), .ZN(new_n398));
  NOR3_X1   g197(.A1(new_n393), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  INV_X1    g198(.A(new_n364), .ZN(new_n400));
  AND3_X1   g199(.A1(new_n390), .A2(KEYINPUT4), .A3(new_n391), .ZN(new_n401));
  NOR3_X1   g200(.A1(new_n244), .A2(new_n252), .A3(new_n249), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n240), .A2(KEYINPUT77), .ZN(new_n403));
  AOI211_X1 g202(.A(new_n229), .B(new_n235), .C1(new_n238), .C2(new_n239), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n403), .A2(new_n404), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n402), .B1(new_n405), .B2(new_n237), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n395), .B(new_n261), .C1(new_n406), .C2(new_n211), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n387), .A2(new_n384), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n398), .B(new_n400), .C1(new_n401), .C2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G1gat), .B(G29gat), .ZN(new_n411));
  INV_X1    g210(.A(G85gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n413), .B(new_n414), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT87), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n410), .A2(new_n416), .ZN(new_n417));
  OAI21_X1  g216(.A(new_n363), .B1(new_n399), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n400), .B1(new_n401), .B2(new_n409), .ZN(new_n419));
  INV_X1    g218(.A(new_n391), .ZN(new_n420));
  AOI21_X1  g219(.A(KEYINPUT82), .B1(new_n406), .B2(new_n382), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n396), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI211_X1 g221(.A(new_n419), .B(KEYINPUT39), .C1(new_n400), .C2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n416), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n424), .B1(new_n393), .B2(new_n398), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n423), .A2(new_n425), .A3(KEYINPUT40), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n400), .A2(KEYINPUT5), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n388), .A2(new_n392), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n407), .A2(new_n364), .ZN(new_n429));
  AND3_X1   g228(.A1(new_n387), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n430));
  AOI21_X1  g229(.A(KEYINPUT81), .B1(new_n387), .B2(KEYINPUT4), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n390), .A2(new_n384), .A3(new_n391), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n429), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n390), .A2(new_n391), .B1(new_n255), .B2(new_n395), .ZN(new_n435));
  OAI21_X1  g234(.A(KEYINPUT5), .B1(new_n435), .B2(new_n364), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n428), .B1(new_n434), .B2(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n437), .A2(new_n424), .ZN(new_n438));
  AND3_X1   g237(.A1(new_n418), .A2(new_n426), .A3(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n280), .B1(new_n362), .B2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT89), .ZN(new_n441));
  AOI21_X1  g240(.A(KEYINPUT37), .B1(new_n345), .B2(new_n347), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n345), .A2(KEYINPUT37), .A3(new_n347), .ZN(new_n444));
  NAND4_X1  g243(.A1(new_n443), .A2(KEYINPUT38), .A3(new_n355), .A4(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT37), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n343), .B1(new_n341), .B2(new_n342), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n447), .B1(KEYINPUT88), .B2(new_n344), .ZN(new_n448));
  OR2_X1    g247(.A1(new_n344), .A2(KEYINPUT88), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n446), .B1(new_n448), .B2(new_n449), .ZN(new_n450));
  NOR3_X1   g249(.A1(new_n450), .A2(new_n442), .A3(new_n358), .ZN(new_n451));
  OAI21_X1  g250(.A(new_n445), .B1(new_n451), .B2(KEYINPUT38), .ZN(new_n452));
  AND3_X1   g251(.A1(new_n388), .A2(new_n392), .A3(new_n427), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n387), .A2(KEYINPUT4), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT81), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n387), .A2(KEYINPUT81), .A3(KEYINPUT4), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n433), .A2(new_n456), .A3(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n429), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT5), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n422), .B2(new_n400), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n453), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(KEYINPUT6), .B1(new_n463), .B2(new_n415), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n460), .A2(new_n462), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n415), .B1(new_n465), .B2(new_n428), .ZN(new_n466));
  AOI22_X1  g265(.A1(new_n464), .A2(new_n438), .B1(new_n466), .B2(KEYINPUT6), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n360), .B(KEYINPUT75), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n452), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n440), .A2(new_n441), .A3(new_n469), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n441), .B1(new_n440), .B2(new_n469), .ZN(new_n471));
  XNOR2_X1  g270(.A(new_n339), .B(new_n382), .ZN(new_n472));
  AND2_X1   g271(.A1(G227gat), .A2(G233gat), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  XNOR2_X1  g274(.A(G15gat), .B(G43gat), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT69), .B(KEYINPUT70), .ZN(new_n477));
  XNOR2_X1  g276(.A(new_n476), .B(new_n477), .ZN(new_n478));
  XOR2_X1   g277(.A(G71gat), .B(G99gat), .Z(new_n479));
  XNOR2_X1  g278(.A(new_n478), .B(new_n479), .ZN(new_n480));
  INV_X1    g279(.A(new_n480), .ZN(new_n481));
  NOR2_X1   g280(.A1(new_n472), .A2(new_n474), .ZN(new_n482));
  OAI211_X1 g281(.A(new_n475), .B(new_n481), .C1(new_n482), .C2(KEYINPUT33), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT33), .ZN(new_n484));
  OAI211_X1 g283(.A(new_n472), .B(new_n474), .C1(new_n484), .C2(new_n480), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n483), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT32), .ZN(new_n487));
  OAI21_X1  g286(.A(KEYINPUT34), .B1(new_n482), .B2(new_n487), .ZN(new_n488));
  INV_X1    g287(.A(KEYINPUT34), .ZN(new_n489));
  OAI211_X1 g288(.A(KEYINPUT32), .B(new_n489), .C1(new_n472), .C2(new_n474), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n486), .A2(new_n491), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n483), .A2(new_n488), .A3(new_n490), .A4(new_n485), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  XNOR2_X1  g293(.A(new_n494), .B(KEYINPUT36), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n470), .A2(new_n471), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT83), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n348), .A2(new_n352), .ZN(new_n498));
  OAI22_X1  g297(.A1(new_n498), .A2(new_n281), .B1(new_n348), .B2(new_n358), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n499), .B1(new_n468), .B2(new_n281), .ZN(new_n500));
  INV_X1    g299(.A(new_n415), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n437), .A2(KEYINPUT6), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g301(.A(new_n415), .B(new_n428), .C1(new_n434), .C2(new_n436), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT6), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n502), .B1(new_n505), .B2(new_n466), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n497), .B1(new_n500), .B2(new_n506), .ZN(new_n507));
  AND4_X1   g306(.A1(new_n497), .A2(new_n506), .A3(new_n357), .A4(new_n361), .ZN(new_n508));
  OAI21_X1  g307(.A(new_n280), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n496), .A2(new_n509), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n463), .A2(new_n504), .A3(new_n415), .ZN(new_n511));
  INV_X1    g310(.A(new_n466), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n511), .B1(new_n512), .B2(new_n464), .ZN(new_n513));
  OAI21_X1  g312(.A(KEYINPUT83), .B1(new_n513), .B2(new_n362), .ZN(new_n514));
  NAND4_X1  g313(.A1(new_n506), .A2(new_n497), .A3(new_n357), .A4(new_n361), .ZN(new_n515));
  NOR2_X1   g314(.A1(new_n280), .A2(new_n494), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n514), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n463), .A2(new_n416), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n502), .B1(new_n518), .B2(new_n505), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n519), .A2(KEYINPUT90), .A3(new_n357), .A4(new_n361), .ZN(new_n520));
  AND2_X1   g319(.A1(new_n520), .A2(new_n516), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n519), .A2(new_n357), .A3(new_n361), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT90), .ZN(new_n523));
  AOI21_X1  g322(.A(KEYINPUT35), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AOI22_X1  g323(.A1(KEYINPUT35), .A2(new_n517), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n526), .ZN(new_n527));
  NAND3_X1  g326(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n528));
  XNOR2_X1  g327(.A(KEYINPUT98), .B(KEYINPUT7), .ZN(new_n529));
  AND2_X1   g328(.A1(G85gat), .A2(G92gat), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n529), .B(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G99gat), .ZN(new_n532));
  INV_X1    g331(.A(G106gat), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT99), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT99), .B1(new_n532), .B2(new_n533), .ZN(new_n535));
  NAND3_X1  g334(.A1(new_n534), .A2(KEYINPUT8), .A3(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n531), .B(new_n536), .C1(G85gat), .C2(G92gat), .ZN(new_n537));
  XOR2_X1   g336(.A(G99gat), .B(G106gat), .Z(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G43gat), .B(G50gat), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT14), .ZN(new_n542));
  INV_X1    g341(.A(G29gat), .ZN(new_n543));
  INV_X1    g342(.A(G36gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(new_n543), .A3(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT92), .ZN(new_n548));
  NAND2_X1  g347(.A1(G29gat), .A2(G36gat), .ZN(new_n549));
  XNOR2_X1  g348(.A(new_n549), .B(KEYINPUT93), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n540), .A2(KEYINPUT15), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n541), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g352(.A1(new_n547), .A2(KEYINPUT15), .A3(new_n540), .A4(new_n549), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n528), .B1(new_n539), .B2(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT100), .ZN(new_n557));
  OR2_X1    g356(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(KEYINPUT17), .ZN(new_n559));
  NAND3_X1  g358(.A1(new_n558), .A2(new_n539), .A3(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n557), .A2(new_n560), .ZN(new_n561));
  XOR2_X1   g360(.A(G190gat), .B(G218gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G134gat), .B(G162gat), .Z(new_n564));
  AOI21_X1  g363(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n565));
  XNOR2_X1  g364(.A(new_n564), .B(new_n565), .ZN(new_n566));
  AND2_X1   g365(.A1(new_n563), .A2(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n563), .A2(new_n566), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g368(.A(G15gat), .B(G22gat), .ZN(new_n570));
  INV_X1    g369(.A(G1gat), .ZN(new_n571));
  NAND3_X1  g370(.A1(new_n570), .A2(KEYINPUT16), .A3(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(G8gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n573), .A2(KEYINPUT94), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n572), .B(new_n574), .C1(new_n571), .C2(new_n570), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n573), .A2(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT21), .ZN(new_n578));
  OAI21_X1  g377(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n579));
  XNOR2_X1  g378(.A(G57gat), .B(G64gat), .ZN(new_n580));
  AOI21_X1  g379(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  XOR2_X1   g381(.A(G71gat), .B(G78gat), .Z(new_n583));
  XNOR2_X1  g382(.A(new_n582), .B(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n577), .B1(new_n578), .B2(new_n585), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n586), .B(KEYINPUT97), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  NOR2_X1   g388(.A1(new_n584), .A2(KEYINPUT21), .ZN(new_n590));
  XOR2_X1   g389(.A(G183gat), .B(G211gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n592), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n589), .B(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G231gat), .A2(G233gat), .ZN(new_n596));
  XOR2_X1   g395(.A(new_n595), .B(new_n596), .Z(new_n597));
  INV_X1    g396(.A(new_n597), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n594), .B(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G120gat), .B(G148gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(G176gat), .B(G204gat), .ZN(new_n601));
  XNOR2_X1  g400(.A(new_n600), .B(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G230gat), .A2(G233gat), .ZN(new_n603));
  INV_X1    g402(.A(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(new_n539), .B(new_n584), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT10), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  OR3_X1    g406(.A1(new_n539), .A2(new_n606), .A3(new_n585), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n604), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n605), .A2(new_n603), .ZN(new_n610));
  OAI21_X1  g409(.A(new_n602), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT102), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n609), .B1(KEYINPUT101), .B2(new_n610), .ZN(new_n614));
  NOR2_X1   g413(.A1(new_n610), .A2(KEYINPUT101), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n615), .A2(new_n602), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  AND2_X1   g416(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND3_X1  g417(.A1(new_n569), .A2(new_n599), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g418(.A(KEYINPUT91), .B(KEYINPUT11), .Z(new_n620));
  XNOR2_X1  g419(.A(G113gat), .B(G141gat), .ZN(new_n621));
  XNOR2_X1  g420(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XOR2_X1   g421(.A(G169gat), .B(G197gat), .Z(new_n623));
  XNOR2_X1  g422(.A(new_n622), .B(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT12), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n555), .A2(new_n577), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n559), .A2(new_n577), .ZN(new_n627));
  AOI21_X1  g426(.A(new_n626), .B1(new_n627), .B2(new_n558), .ZN(new_n628));
  NAND2_X1  g427(.A1(G229gat), .A2(G233gat), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT18), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n625), .B1(new_n632), .B2(KEYINPUT95), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n555), .B(new_n577), .ZN(new_n634));
  XOR2_X1   g433(.A(new_n629), .B(KEYINPUT13), .Z(new_n635));
  NAND2_X1  g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n628), .A2(KEYINPUT18), .A3(new_n629), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n632), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OR2_X1    g437(.A1(new_n633), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(new_n633), .A2(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n619), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n527), .A2(new_n643), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n644), .A2(new_n506), .ZN(new_n645));
  XNOR2_X1  g444(.A(new_n645), .B(new_n571), .ZN(G1324gat));
  NOR2_X1   g445(.A1(new_n644), .A2(new_n500), .ZN(new_n647));
  OAI21_X1  g446(.A(new_n573), .B1(new_n647), .B2(KEYINPUT42), .ZN(new_n648));
  INV_X1    g447(.A(KEYINPUT42), .ZN(new_n649));
  NAND2_X1  g448(.A1(new_n649), .A2(KEYINPUT103), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n647), .A2(new_n651), .ZN(new_n652));
  MUX2_X1   g451(.A(new_n573), .B(new_n648), .S(new_n652), .Z(G1325gat));
  INV_X1    g452(.A(new_n644), .ZN(new_n654));
  AND3_X1   g453(.A1(new_n654), .A2(G15gat), .A3(new_n495), .ZN(new_n655));
  INV_X1    g454(.A(new_n494), .ZN(new_n656));
  AOI21_X1  g455(.A(G15gat), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n657), .ZN(G1326gat));
  INV_X1    g457(.A(new_n280), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n644), .A2(new_n659), .ZN(new_n660));
  XOR2_X1   g459(.A(KEYINPUT104), .B(KEYINPUT105), .Z(new_n661));
  XNOR2_X1  g460(.A(new_n660), .B(new_n661), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT43), .B(G22gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1327gat));
  NOR2_X1   g463(.A1(new_n567), .A2(new_n568), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT44), .ZN(new_n666));
  NAND2_X1  g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n509), .A2(KEYINPUT106), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n514), .A2(new_n515), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT106), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n280), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n471), .ZN(new_n673));
  INV_X1    g472(.A(new_n495), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n440), .A2(new_n441), .A3(new_n469), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n673), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n526), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(KEYINPUT107), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR2_X1   g478(.A1(new_n470), .A2(new_n471), .ZN(new_n680));
  NAND4_X1  g479(.A1(new_n680), .A2(new_n668), .A3(new_n674), .A4(new_n671), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n681), .A2(KEYINPUT107), .A3(new_n526), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n667), .B1(new_n679), .B2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n569), .B1(new_n510), .B2(new_n526), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n684), .A2(new_n666), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n683), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  XNOR2_X1  g486(.A(new_n594), .B(new_n597), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n618), .A2(new_n688), .A3(new_n641), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(KEYINPUT108), .B1(new_n691), .B2(new_n506), .ZN(new_n692));
  NOR2_X1   g491(.A1(new_n686), .A2(new_n689), .ZN(new_n693));
  INV_X1    g492(.A(KEYINPUT108), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n693), .A2(new_n694), .A3(new_n513), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n692), .A2(G29gat), .A3(new_n695), .ZN(new_n696));
  AND2_X1   g495(.A1(new_n684), .A2(new_n690), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n697), .A2(new_n543), .A3(new_n513), .ZN(new_n698));
  XNOR2_X1  g497(.A(new_n698), .B(KEYINPUT45), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n696), .A2(new_n699), .ZN(G1328gat));
  OAI21_X1  g499(.A(G36gat), .B1(new_n691), .B2(new_n500), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n697), .A2(new_n544), .A3(new_n362), .ZN(new_n702));
  AND2_X1   g501(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n703));
  NOR2_X1   g502(.A1(KEYINPUT109), .A2(KEYINPUT46), .ZN(new_n704));
  OAI21_X1  g503(.A(new_n702), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  OAI211_X1 g504(.A(new_n701), .B(new_n705), .C1(new_n703), .C2(new_n702), .ZN(G1329gat));
  NAND3_X1  g505(.A1(new_n693), .A2(G43gat), .A3(new_n495), .ZN(new_n707));
  AND2_X1   g506(.A1(new_n697), .A2(new_n656), .ZN(new_n708));
  OR2_X1    g507(.A1(new_n708), .A2(G43gat), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT47), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT47), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n707), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1330gat));
  OAI21_X1  g513(.A(G50gat), .B1(new_n691), .B2(new_n659), .ZN(new_n715));
  INV_X1    g514(.A(G50gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n280), .A2(new_n716), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(KEYINPUT110), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n697), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n715), .A2(KEYINPUT48), .A3(new_n719), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT48), .ZN(new_n721));
  AOI21_X1  g520(.A(new_n716), .B1(new_n693), .B2(new_n280), .ZN(new_n722));
  INV_X1    g521(.A(new_n719), .ZN(new_n723));
  OAI21_X1  g522(.A(new_n721), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n720), .A2(new_n724), .ZN(G1331gat));
  NOR3_X1   g524(.A1(new_n618), .A2(new_n665), .A3(new_n688), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n670), .B1(new_n669), .B2(new_n280), .ZN(new_n727));
  AOI211_X1 g526(.A(KEYINPUT106), .B(new_n659), .C1(new_n514), .C2(new_n515), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n678), .B(new_n525), .C1(new_n729), .C2(new_n496), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT107), .B1(new_n681), .B2(new_n526), .ZN(new_n731));
  OAI211_X1 g530(.A(new_n642), .B(new_n726), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n506), .ZN(new_n733));
  XOR2_X1   g532(.A(new_n733), .B(G57gat), .Z(G1332gat));
  INV_X1    g533(.A(KEYINPUT111), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n679), .A2(new_n682), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(KEYINPUT111), .A3(new_n642), .A4(new_n726), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n500), .B1(new_n736), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g538(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n740));
  AND2_X1   g539(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n742), .B1(new_n739), .B2(new_n740), .ZN(G1333gat));
  OR3_X1    g542(.A1(new_n732), .A2(G71gat), .A3(new_n494), .ZN(new_n744));
  AOI21_X1  g543(.A(new_n674), .B1(new_n736), .B2(new_n738), .ZN(new_n745));
  INV_X1    g544(.A(G71gat), .ZN(new_n746));
  OAI21_X1  g545(.A(new_n744), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  XOR2_X1   g546(.A(KEYINPUT112), .B(KEYINPUT50), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n748), .ZN(new_n750));
  OAI211_X1 g549(.A(new_n744), .B(new_n750), .C1(new_n745), .C2(new_n746), .ZN(new_n751));
  AND2_X1   g550(.A1(new_n749), .A2(new_n751), .ZN(G1334gat));
  AOI21_X1  g551(.A(new_n659), .B1(new_n736), .B2(new_n738), .ZN(new_n753));
  XOR2_X1   g552(.A(new_n753), .B(G78gat), .Z(G1335gat));
  NOR3_X1   g553(.A1(new_n599), .A2(new_n641), .A3(KEYINPUT113), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  OAI21_X1  g555(.A(KEYINPUT113), .B1(new_n599), .B2(new_n641), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n618), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n687), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n506), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n525), .B1(new_n729), .B2(new_n496), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n762));
  INV_X1    g561(.A(new_n757), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n665), .B1(new_n763), .B2(new_n755), .ZN(new_n764));
  NOR3_X1   g563(.A1(new_n761), .A2(new_n762), .A3(new_n764), .ZN(new_n765));
  AOI21_X1  g564(.A(new_n569), .B1(new_n756), .B2(new_n757), .ZN(new_n766));
  AOI21_X1  g565(.A(KEYINPUT51), .B1(new_n677), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n765), .A2(new_n767), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n768), .A2(new_n618), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n769), .A2(new_n412), .A3(new_n513), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n760), .A2(new_n770), .ZN(G1336gat));
  NAND2_X1  g570(.A1(new_n613), .A2(new_n617), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n500), .A2(G92gat), .ZN(new_n773));
  AND2_X1   g572(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n762), .B1(new_n761), .B2(new_n764), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n677), .A2(KEYINPUT51), .A3(new_n766), .ZN(new_n776));
  AOI21_X1  g575(.A(KEYINPUT114), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n767), .A2(new_n778), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n774), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n362), .B(new_n758), .C1(new_n683), .C2(new_n685), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G92gat), .ZN(new_n784));
  OAI211_X1 g583(.A(KEYINPUT115), .B(new_n774), .C1(new_n777), .C2(new_n779), .ZN(new_n785));
  NAND3_X1  g584(.A1(new_n782), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT52), .ZN(new_n787));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(new_n769), .B2(new_n773), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(new_n784), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1337gat));
  OAI21_X1  g589(.A(G99gat), .B1(new_n759), .B2(new_n674), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n772), .A2(new_n656), .A3(new_n532), .ZN(new_n792));
  XNOR2_X1  g591(.A(new_n792), .B(KEYINPUT116), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n791), .B1(new_n768), .B2(new_n793), .ZN(G1338gat));
  INV_X1    g593(.A(KEYINPUT118), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT53), .ZN(new_n796));
  OAI211_X1 g595(.A(new_n280), .B(new_n758), .C1(new_n683), .C2(new_n685), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(G106gat), .ZN(new_n798));
  NOR3_X1   g597(.A1(new_n618), .A2(G106gat), .A3(new_n659), .ZN(new_n799));
  INV_X1    g598(.A(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT117), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(new_n801), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n802), .B(new_n804), .C1(new_n777), .C2(new_n779), .ZN(new_n805));
  AOI21_X1  g604(.A(new_n796), .B1(new_n798), .B2(new_n805), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n796), .B1(new_n768), .B2(new_n800), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n807), .B1(G106gat), .B2(new_n797), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n795), .B1(new_n806), .B2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n807), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n798), .A2(new_n810), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n778), .B1(new_n765), .B2(new_n767), .ZN(new_n812));
  NAND2_X1  g611(.A1(new_n775), .A2(KEYINPUT114), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n803), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  AOI22_X1  g613(.A1(new_n814), .A2(new_n802), .B1(new_n797), .B2(G106gat), .ZN(new_n815));
  OAI211_X1 g614(.A(KEYINPUT118), .B(new_n811), .C1(new_n815), .C2(new_n796), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n809), .A2(new_n816), .ZN(G1339gat));
  NOR2_X1   g616(.A1(new_n619), .A2(new_n641), .ZN(new_n818));
  NAND4_X1  g617(.A1(new_n632), .A2(new_n625), .A3(new_n636), .A4(new_n637), .ZN(new_n819));
  NOR2_X1   g618(.A1(new_n628), .A2(new_n629), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n634), .A2(new_n635), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n624), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AND2_X1   g621(.A1(new_n819), .A2(new_n822), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n665), .B1(new_n772), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT54), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n609), .A2(new_n825), .ZN(new_n826));
  NAND3_X1  g625(.A1(new_n607), .A2(new_n604), .A3(new_n608), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT54), .ZN(new_n828));
  OAI211_X1 g627(.A(new_n826), .B(new_n602), .C1(new_n828), .C2(new_n609), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT55), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n617), .B1(new_n829), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n833), .A2(new_n641), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n599), .B1(new_n824), .B2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n833), .A2(new_n823), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(new_n665), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n818), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NOR3_X1   g637(.A1(new_n838), .A2(new_n280), .A3(new_n494), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n362), .A2(new_n506), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  INV_X1    g640(.A(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n641), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n368), .A2(KEYINPUT119), .ZN(new_n844));
  AND2_X1   g643(.A1(new_n368), .A2(KEYINPUT119), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n846), .B1(new_n843), .B2(new_n844), .ZN(G1340gat));
  NOR2_X1   g646(.A1(new_n841), .A2(new_n618), .ZN(new_n848));
  XNOR2_X1  g647(.A(new_n848), .B(new_n366), .ZN(G1341gat));
  OR3_X1    g648(.A1(new_n841), .A2(KEYINPUT120), .A3(new_n688), .ZN(new_n850));
  OAI21_X1  g649(.A(KEYINPUT120), .B1(new_n841), .B2(new_n688), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g651(.A(KEYINPUT68), .B(G127gat), .ZN(new_n853));
  INV_X1    g652(.A(new_n853), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n852), .B(new_n854), .ZN(G1342gat));
  NAND2_X1  g654(.A1(new_n842), .A2(new_n665), .ZN(new_n856));
  OR3_X1    g655(.A1(new_n856), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(G134gat), .ZN(new_n858));
  OAI21_X1  g657(.A(KEYINPUT56), .B1(new_n856), .B2(G134gat), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n857), .A2(new_n858), .A3(new_n859), .ZN(G1343gat));
  NAND2_X1  g659(.A1(new_n674), .A2(new_n840), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n772), .A2(new_n823), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n834), .A2(new_n569), .A3(new_n862), .ZN(new_n863));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n863), .A2(new_n837), .A3(new_n864), .A4(new_n688), .ZN(new_n865));
  INV_X1    g664(.A(new_n818), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n864), .B1(new_n835), .B2(new_n837), .ZN(new_n868));
  OAI211_X1 g667(.A(KEYINPUT57), .B(new_n280), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  XOR2_X1   g668(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n871), .B1(new_n838), .B2(new_n659), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n861), .B1(new_n869), .B2(new_n872), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n873), .A2(G141gat), .A3(new_n641), .ZN(new_n874));
  NOR2_X1   g673(.A1(new_n838), .A2(new_n659), .ZN(new_n875));
  NAND4_X1  g674(.A1(new_n875), .A2(new_n674), .A3(new_n641), .A4(new_n840), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n233), .ZN(new_n877));
  AOI21_X1  g676(.A(KEYINPUT123), .B1(new_n874), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT124), .B(KEYINPUT58), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n879), .ZN(new_n881));
  AOI211_X1 g680(.A(KEYINPUT123), .B(new_n881), .C1(new_n874), .C2(new_n877), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n882), .ZN(G1344gat));
  AND2_X1   g682(.A1(new_n835), .A2(new_n837), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n280), .B1(new_n884), .B2(new_n818), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n885), .A2(new_n861), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n886), .A2(new_n231), .A3(new_n772), .ZN(new_n887));
  XOR2_X1   g686(.A(new_n887), .B(KEYINPUT125), .Z(new_n888));
  INV_X1    g687(.A(KEYINPUT59), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n885), .A2(KEYINPUT57), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n875), .A2(new_n871), .ZN(new_n891));
  AND2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n861), .A2(KEYINPUT126), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n861), .A2(KEYINPUT126), .ZN(new_n894));
  NAND4_X1  g693(.A1(new_n892), .A2(new_n772), .A3(new_n893), .A4(new_n894), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n889), .B1(new_n895), .B2(G148gat), .ZN(new_n896));
  AOI211_X1 g695(.A(KEYINPUT59), .B(new_n231), .C1(new_n873), .C2(new_n772), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(G1345gat));
  AOI21_X1  g697(.A(G155gat), .B1(new_n886), .B2(new_n599), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n688), .A2(new_n225), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n899), .B1(new_n873), .B2(new_n900), .ZN(G1346gat));
  AOI21_X1  g700(.A(new_n243), .B1(new_n886), .B2(new_n665), .ZN(new_n902));
  AND2_X1   g701(.A1(new_n665), .A2(new_n243), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n902), .B1(new_n873), .B2(new_n903), .ZN(G1347gat));
  NOR2_X1   g703(.A1(new_n500), .A2(new_n513), .ZN(new_n905));
  AND2_X1   g704(.A1(new_n839), .A2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n641), .ZN(new_n907));
  XNOR2_X1  g706(.A(new_n907), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g707(.A1(new_n906), .A2(new_n772), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n909), .A2(G176gat), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n292), .A2(new_n293), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n911), .B2(new_n909), .ZN(G1349gat));
  AND3_X1   g711(.A1(new_n906), .A2(new_n317), .A3(new_n599), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n282), .B1(new_n906), .B2(new_n599), .ZN(new_n914));
  OR3_X1    g713(.A1(new_n913), .A2(new_n914), .A3(KEYINPUT60), .ZN(new_n915));
  OAI21_X1  g714(.A(KEYINPUT60), .B1(new_n913), .B2(new_n914), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n915), .A2(new_n916), .ZN(G1350gat));
  NAND2_X1  g716(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n918));
  XNOR2_X1  g717(.A(KEYINPUT61), .B(G190gat), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n906), .A2(new_n665), .ZN(new_n920));
  MUX2_X1   g719(.A(new_n918), .B(new_n919), .S(new_n920), .Z(G1351gat));
  NAND2_X1  g720(.A1(new_n674), .A2(new_n905), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n885), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT127), .ZN(new_n924));
  INV_X1    g723(.A(G197gat), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n924), .A2(new_n925), .A3(new_n641), .ZN(new_n926));
  INV_X1    g725(.A(new_n922), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n892), .A2(new_n927), .ZN(new_n928));
  OAI21_X1  g727(.A(G197gat), .B1(new_n928), .B2(new_n642), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n926), .A2(new_n929), .ZN(G1352gat));
  OAI21_X1  g729(.A(G204gat), .B1(new_n928), .B2(new_n618), .ZN(new_n931));
  NOR4_X1   g730(.A1(new_n885), .A2(G204gat), .A3(new_n618), .A4(new_n922), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT62), .ZN(new_n933));
  OR2_X1    g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n933), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n931), .A2(new_n934), .A3(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n216), .A3(new_n599), .ZN(new_n937));
  NAND4_X1  g736(.A1(new_n890), .A2(new_n891), .A3(new_n599), .A4(new_n927), .ZN(new_n938));
  AOI21_X1  g737(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  AOI21_X1  g740(.A(G218gat), .B1(new_n924), .B2(new_n665), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n928), .A2(new_n217), .A3(new_n569), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n942), .A2(new_n943), .ZN(G1355gat));
endmodule


