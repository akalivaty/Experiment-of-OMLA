

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, n775,
         n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786,
         n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U554 ( .A1(G651), .A2(n622), .ZN(n652) );
  INV_X1 U555 ( .A(n714), .ZN(n701) );
  XOR2_X1 U556 ( .A(KEYINPUT1), .B(n542), .Z(n644) );
  XNOR2_X1 U557 ( .A(n718), .B(n717), .ZN(n719) );
  XNOR2_X1 U558 ( .A(n761), .B(KEYINPUT101), .ZN(n765) );
  AND2_X1 U559 ( .A1(n697), .A2(n973), .ZN(n519) );
  OR2_X1 U560 ( .A1(n764), .A2(n763), .ZN(n520) );
  XNOR2_X1 U561 ( .A(KEYINPUT30), .B(KEYINPUT98), .ZN(n717) );
  INV_X1 U562 ( .A(KEYINPUT31), .ZN(n723) );
  AND2_X1 U563 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U564 ( .A1(n765), .A2(n520), .ZN(n803) );
  NOR2_X2 U565 ( .A1(G2105), .A2(n521), .ZN(n888) );
  INV_X1 U566 ( .A(G2104), .ZN(n521) );
  NAND2_X1 U567 ( .A1(G101), .A2(n888), .ZN(n522) );
  XNOR2_X1 U568 ( .A(KEYINPUT23), .B(n522), .ZN(n529) );
  AND2_X1 U569 ( .A1(G2104), .A2(G2105), .ZN(n884) );
  NAND2_X1 U570 ( .A1(G113), .A2(n884), .ZN(n527) );
  INV_X1 U571 ( .A(G137), .ZN(n525) );
  XNOR2_X1 U572 ( .A(KEYINPUT17), .B(KEYINPUT67), .ZN(n524) );
  NOR2_X1 U573 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XNOR2_X1 U574 ( .A(n524), .B(n523), .ZN(n534) );
  INV_X1 U575 ( .A(n534), .ZN(n602) );
  OR2_X1 U576 ( .A1(n525), .A2(n602), .ZN(n526) );
  NAND2_X1 U577 ( .A1(n527), .A2(n526), .ZN(n528) );
  NOR2_X1 U578 ( .A1(n529), .A2(n528), .ZN(n533) );
  NAND2_X1 U579 ( .A1(n521), .A2(G2105), .ZN(n530) );
  XNOR2_X2 U580 ( .A(n530), .B(KEYINPUT65), .ZN(n885) );
  NAND2_X1 U581 ( .A1(G125), .A2(n885), .ZN(n531) );
  XNOR2_X1 U582 ( .A(n531), .B(KEYINPUT66), .ZN(n532) );
  AND2_X1 U583 ( .A1(n533), .A2(n532), .ZN(G160) );
  NAND2_X1 U584 ( .A1(G138), .A2(n534), .ZN(n535) );
  XNOR2_X1 U585 ( .A(n535), .B(KEYINPUT86), .ZN(n541) );
  NAND2_X1 U586 ( .A1(G114), .A2(n884), .ZN(n537) );
  NAND2_X1 U587 ( .A1(G102), .A2(n888), .ZN(n536) );
  NAND2_X1 U588 ( .A1(n537), .A2(n536), .ZN(n539) );
  AND2_X1 U589 ( .A1(n885), .A2(G126), .ZN(n538) );
  NOR2_X1 U590 ( .A1(n539), .A2(n538), .ZN(n540) );
  AND2_X1 U591 ( .A1(n541), .A2(n540), .ZN(G164) );
  INV_X1 U592 ( .A(G651), .ZN(n544) );
  NOR2_X1 U593 ( .A1(G543), .A2(n544), .ZN(n542) );
  NAND2_X1 U594 ( .A1(G64), .A2(n644), .ZN(n543) );
  XNOR2_X1 U595 ( .A(n543), .B(KEYINPUT69), .ZN(n551) );
  NOR2_X1 U596 ( .A1(G543), .A2(G651), .ZN(n643) );
  NAND2_X1 U597 ( .A1(G90), .A2(n643), .ZN(n546) );
  XOR2_X1 U598 ( .A(G543), .B(KEYINPUT0), .Z(n622) );
  NOR2_X1 U599 ( .A1(n622), .A2(n544), .ZN(n647) );
  NAND2_X1 U600 ( .A1(G77), .A2(n647), .ZN(n545) );
  NAND2_X1 U601 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U602 ( .A(n547), .B(KEYINPUT9), .ZN(n549) );
  NAND2_X1 U603 ( .A1(G52), .A2(n652), .ZN(n548) );
  NAND2_X1 U604 ( .A1(n549), .A2(n548), .ZN(n550) );
  NOR2_X1 U605 ( .A1(n551), .A2(n550), .ZN(G171) );
  AND2_X1 U606 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U607 ( .A(G57), .ZN(G237) );
  INV_X1 U608 ( .A(G120), .ZN(G236) );
  NAND2_X1 U609 ( .A1(n643), .A2(G89), .ZN(n552) );
  XNOR2_X1 U610 ( .A(n552), .B(KEYINPUT4), .ZN(n554) );
  NAND2_X1 U611 ( .A1(G76), .A2(n647), .ZN(n553) );
  NAND2_X1 U612 ( .A1(n554), .A2(n553), .ZN(n555) );
  XNOR2_X1 U613 ( .A(n555), .B(KEYINPUT5), .ZN(n560) );
  NAND2_X1 U614 ( .A1(G51), .A2(n652), .ZN(n557) );
  NAND2_X1 U615 ( .A1(G63), .A2(n644), .ZN(n556) );
  NAND2_X1 U616 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U617 ( .A(KEYINPUT6), .B(n558), .Z(n559) );
  NAND2_X1 U618 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U619 ( .A(n561), .B(KEYINPUT7), .ZN(G168) );
  XOR2_X1 U620 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U621 ( .A1(G7), .A2(G661), .ZN(n562) );
  XNOR2_X1 U622 ( .A(n562), .B(KEYINPUT10), .ZN(n563) );
  XNOR2_X1 U623 ( .A(KEYINPUT74), .B(n563), .ZN(G223) );
  INV_X1 U624 ( .A(G223), .ZN(n832) );
  NAND2_X1 U625 ( .A1(n832), .A2(G567), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(n564), .Z(G234) );
  NAND2_X1 U627 ( .A1(n643), .A2(G81), .ZN(n565) );
  XNOR2_X1 U628 ( .A(n565), .B(KEYINPUT12), .ZN(n567) );
  NAND2_X1 U629 ( .A1(G68), .A2(n647), .ZN(n566) );
  NAND2_X1 U630 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U631 ( .A(n568), .B(KEYINPUT13), .ZN(n570) );
  NAND2_X1 U632 ( .A1(G43), .A2(n652), .ZN(n569) );
  NAND2_X1 U633 ( .A1(n570), .A2(n569), .ZN(n573) );
  NAND2_X1 U634 ( .A1(n644), .A2(G56), .ZN(n571) );
  XOR2_X1 U635 ( .A(KEYINPUT14), .B(n571), .Z(n572) );
  NOR2_X2 U636 ( .A1(n573), .A2(n572), .ZN(n985) );
  NAND2_X1 U637 ( .A1(n985), .A2(G860), .ZN(G153) );
  INV_X1 U638 ( .A(G171), .ZN(G301) );
  NAND2_X1 U639 ( .A1(G868), .A2(G301), .ZN(n582) );
  NAND2_X1 U640 ( .A1(G54), .A2(n652), .ZN(n575) );
  NAND2_X1 U641 ( .A1(G66), .A2(n644), .ZN(n574) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n579) );
  NAND2_X1 U643 ( .A1(G92), .A2(n643), .ZN(n577) );
  NAND2_X1 U644 ( .A1(G79), .A2(n647), .ZN(n576) );
  NAND2_X1 U645 ( .A1(n577), .A2(n576), .ZN(n578) );
  NOR2_X1 U646 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U647 ( .A(n580), .B(KEYINPUT15), .ZN(n973) );
  INV_X1 U648 ( .A(G868), .ZN(n665) );
  NAND2_X1 U649 ( .A1(n973), .A2(n665), .ZN(n581) );
  NAND2_X1 U650 ( .A1(n582), .A2(n581), .ZN(G284) );
  NAND2_X1 U651 ( .A1(n644), .A2(G65), .ZN(n583) );
  XNOR2_X1 U652 ( .A(n583), .B(KEYINPUT72), .ZN(n585) );
  NAND2_X1 U653 ( .A1(G53), .A2(n652), .ZN(n584) );
  NAND2_X1 U654 ( .A1(n585), .A2(n584), .ZN(n586) );
  XNOR2_X1 U655 ( .A(KEYINPUT73), .B(n586), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n647), .A2(G78), .ZN(n587) );
  XNOR2_X1 U657 ( .A(n587), .B(KEYINPUT70), .ZN(n589) );
  NAND2_X1 U658 ( .A1(G91), .A2(n643), .ZN(n588) );
  NAND2_X1 U659 ( .A1(n589), .A2(n588), .ZN(n590) );
  XNOR2_X1 U660 ( .A(KEYINPUT71), .B(n590), .ZN(n591) );
  NAND2_X1 U661 ( .A1(n592), .A2(n591), .ZN(G299) );
  NOR2_X1 U662 ( .A1(G286), .A2(n665), .ZN(n594) );
  NOR2_X1 U663 ( .A1(G868), .A2(G299), .ZN(n593) );
  NOR2_X1 U664 ( .A1(n594), .A2(n593), .ZN(G297) );
  INV_X1 U665 ( .A(G860), .ZN(n595) );
  NAND2_X1 U666 ( .A1(n595), .A2(G559), .ZN(n596) );
  INV_X1 U667 ( .A(n973), .ZN(n619) );
  NAND2_X1 U668 ( .A1(n596), .A2(n619), .ZN(n597) );
  XNOR2_X1 U669 ( .A(n597), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U670 ( .A1(n619), .A2(G868), .ZN(n598) );
  NOR2_X1 U671 ( .A1(G559), .A2(n598), .ZN(n600) );
  AND2_X1 U672 ( .A1(n665), .A2(n985), .ZN(n599) );
  NOR2_X1 U673 ( .A1(n600), .A2(n599), .ZN(G282) );
  NAND2_X1 U674 ( .A1(n885), .A2(G123), .ZN(n601) );
  XNOR2_X1 U675 ( .A(n601), .B(KEYINPUT18), .ZN(n604) );
  INV_X1 U676 ( .A(n602), .ZN(n889) );
  NAND2_X1 U677 ( .A1(G135), .A2(n889), .ZN(n603) );
  NAND2_X1 U678 ( .A1(n604), .A2(n603), .ZN(n609) );
  NAND2_X1 U679 ( .A1(G111), .A2(n884), .ZN(n606) );
  NAND2_X1 U680 ( .A1(G99), .A2(n888), .ZN(n605) );
  NAND2_X1 U681 ( .A1(n606), .A2(n605), .ZN(n607) );
  XOR2_X1 U682 ( .A(KEYINPUT75), .B(n607), .Z(n608) );
  NOR2_X1 U683 ( .A1(n609), .A2(n608), .ZN(n610) );
  XNOR2_X1 U684 ( .A(KEYINPUT76), .B(n610), .ZN(n923) );
  XNOR2_X1 U685 ( .A(n923), .B(G2096), .ZN(n612) );
  INV_X1 U686 ( .A(G2100), .ZN(n611) );
  NAND2_X1 U687 ( .A1(n612), .A2(n611), .ZN(G156) );
  NAND2_X1 U688 ( .A1(G93), .A2(n643), .ZN(n614) );
  NAND2_X1 U689 ( .A1(G80), .A2(n647), .ZN(n613) );
  NAND2_X1 U690 ( .A1(n614), .A2(n613), .ZN(n618) );
  NAND2_X1 U691 ( .A1(G55), .A2(n652), .ZN(n616) );
  NAND2_X1 U692 ( .A1(G67), .A2(n644), .ZN(n615) );
  NAND2_X1 U693 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U694 ( .A1(n618), .A2(n617), .ZN(n664) );
  NAND2_X1 U695 ( .A1(n619), .A2(G559), .ZN(n662) );
  XOR2_X1 U696 ( .A(n985), .B(n662), .Z(n620) );
  NOR2_X1 U697 ( .A1(G860), .A2(n620), .ZN(n621) );
  XOR2_X1 U698 ( .A(n664), .B(n621), .Z(G145) );
  NAND2_X1 U699 ( .A1(G49), .A2(n652), .ZN(n624) );
  NAND2_X1 U700 ( .A1(G87), .A2(n622), .ZN(n623) );
  NAND2_X1 U701 ( .A1(n624), .A2(n623), .ZN(n625) );
  NOR2_X1 U702 ( .A1(n644), .A2(n625), .ZN(n628) );
  NAND2_X1 U703 ( .A1(G74), .A2(G651), .ZN(n626) );
  XOR2_X1 U704 ( .A(KEYINPUT77), .B(n626), .Z(n627) );
  NAND2_X1 U705 ( .A1(n628), .A2(n627), .ZN(G288) );
  NAND2_X1 U706 ( .A1(G85), .A2(n643), .ZN(n630) );
  NAND2_X1 U707 ( .A1(G72), .A2(n647), .ZN(n629) );
  NAND2_X1 U708 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U709 ( .A(KEYINPUT68), .B(n631), .Z(n635) );
  NAND2_X1 U710 ( .A1(G47), .A2(n652), .ZN(n633) );
  NAND2_X1 U711 ( .A1(G60), .A2(n644), .ZN(n632) );
  AND2_X1 U712 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U713 ( .A1(n635), .A2(n634), .ZN(G290) );
  NAND2_X1 U714 ( .A1(G50), .A2(n652), .ZN(n637) );
  NAND2_X1 U715 ( .A1(G62), .A2(n644), .ZN(n636) );
  NAND2_X1 U716 ( .A1(n637), .A2(n636), .ZN(n642) );
  NAND2_X1 U717 ( .A1(G88), .A2(n643), .ZN(n639) );
  NAND2_X1 U718 ( .A1(G75), .A2(n647), .ZN(n638) );
  NAND2_X1 U719 ( .A1(n639), .A2(n638), .ZN(n640) );
  XOR2_X1 U720 ( .A(KEYINPUT79), .B(n640), .Z(n641) );
  NOR2_X1 U721 ( .A1(n642), .A2(n641), .ZN(G166) );
  NAND2_X1 U722 ( .A1(G86), .A2(n643), .ZN(n646) );
  NAND2_X1 U723 ( .A1(G61), .A2(n644), .ZN(n645) );
  NAND2_X1 U724 ( .A1(n646), .A2(n645), .ZN(n650) );
  NAND2_X1 U725 ( .A1(n647), .A2(G73), .ZN(n648) );
  XOR2_X1 U726 ( .A(KEYINPUT2), .B(n648), .Z(n649) );
  NOR2_X1 U727 ( .A1(n650), .A2(n649), .ZN(n651) );
  XNOR2_X1 U728 ( .A(n651), .B(KEYINPUT78), .ZN(n654) );
  NAND2_X1 U729 ( .A1(G48), .A2(n652), .ZN(n653) );
  NAND2_X1 U730 ( .A1(n654), .A2(n653), .ZN(G305) );
  XNOR2_X1 U731 ( .A(KEYINPUT19), .B(KEYINPUT80), .ZN(n656) );
  XNOR2_X1 U732 ( .A(G288), .B(n985), .ZN(n655) );
  XNOR2_X1 U733 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U734 ( .A(n664), .B(n657), .Z(n659) );
  XNOR2_X1 U735 ( .A(G290), .B(G166), .ZN(n658) );
  XNOR2_X1 U736 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U737 ( .A(n660), .B(G305), .ZN(n661) );
  XNOR2_X1 U738 ( .A(n661), .B(G299), .ZN(n904) );
  XNOR2_X1 U739 ( .A(n662), .B(n904), .ZN(n663) );
  NAND2_X1 U740 ( .A1(n663), .A2(G868), .ZN(n667) );
  NAND2_X1 U741 ( .A1(n665), .A2(n664), .ZN(n666) );
  NAND2_X1 U742 ( .A1(n667), .A2(n666), .ZN(G295) );
  NAND2_X1 U743 ( .A1(G2078), .A2(G2084), .ZN(n668) );
  XOR2_X1 U744 ( .A(KEYINPUT20), .B(n668), .Z(n669) );
  NAND2_X1 U745 ( .A1(G2090), .A2(n669), .ZN(n670) );
  XNOR2_X1 U746 ( .A(KEYINPUT21), .B(n670), .ZN(n671) );
  NAND2_X1 U747 ( .A1(n671), .A2(G2072), .ZN(G158) );
  XOR2_X1 U748 ( .A(KEYINPUT81), .B(G44), .Z(n672) );
  XNOR2_X1 U749 ( .A(KEYINPUT3), .B(n672), .ZN(G218) );
  NAND2_X1 U750 ( .A1(G132), .A2(G82), .ZN(n673) );
  XNOR2_X1 U751 ( .A(n673), .B(KEYINPUT22), .ZN(n674) );
  XNOR2_X1 U752 ( .A(n674), .B(KEYINPUT82), .ZN(n675) );
  NOR2_X1 U753 ( .A1(G218), .A2(n675), .ZN(n676) );
  NAND2_X1 U754 ( .A1(G96), .A2(n676), .ZN(n836) );
  NAND2_X1 U755 ( .A1(n836), .A2(G2106), .ZN(n682) );
  NOR2_X1 U756 ( .A1(G236), .A2(G237), .ZN(n677) );
  NAND2_X1 U757 ( .A1(G69), .A2(n677), .ZN(n678) );
  XNOR2_X1 U758 ( .A(KEYINPUT83), .B(n678), .ZN(n679) );
  NAND2_X1 U759 ( .A1(n679), .A2(G108), .ZN(n680) );
  XNOR2_X1 U760 ( .A(KEYINPUT84), .B(n680), .ZN(n837) );
  NAND2_X1 U761 ( .A1(n837), .A2(G567), .ZN(n681) );
  NAND2_X1 U762 ( .A1(n682), .A2(n681), .ZN(n838) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n683) );
  XOR2_X1 U764 ( .A(KEYINPUT85), .B(n683), .Z(n684) );
  NOR2_X1 U765 ( .A1(n838), .A2(n684), .ZN(n835) );
  NAND2_X1 U766 ( .A1(n835), .A2(G36), .ZN(G176) );
  XNOR2_X1 U767 ( .A(KEYINPUT87), .B(G166), .ZN(G303) );
  NOR2_X1 U768 ( .A1(G164), .A2(G1384), .ZN(n766) );
  AND2_X1 U769 ( .A1(G160), .A2(G40), .ZN(n685) );
  NAND2_X1 U770 ( .A1(n766), .A2(n685), .ZN(n714) );
  XNOR2_X1 U771 ( .A(G2078), .B(KEYINPUT25), .ZN(n953) );
  NOR2_X1 U772 ( .A1(n714), .A2(n953), .ZN(n687) );
  INV_X1 U773 ( .A(G1961), .ZN(n1008) );
  NOR2_X1 U774 ( .A1(n701), .A2(n1008), .ZN(n686) );
  NOR2_X1 U775 ( .A1(n687), .A2(n686), .ZN(n720) );
  NAND2_X1 U776 ( .A1(G171), .A2(n720), .ZN(n713) );
  NAND2_X1 U777 ( .A1(n701), .A2(G1996), .ZN(n688) );
  XNOR2_X1 U778 ( .A(n688), .B(KEYINPUT26), .ZN(n689) );
  XNOR2_X1 U779 ( .A(n689), .B(KEYINPUT64), .ZN(n696) );
  NAND2_X1 U780 ( .A1(G1348), .A2(n714), .ZN(n691) );
  NAND2_X1 U781 ( .A1(G2067), .A2(n701), .ZN(n690) );
  NAND2_X1 U782 ( .A1(n691), .A2(n690), .ZN(n697) );
  NAND2_X1 U783 ( .A1(n714), .A2(G1341), .ZN(n692) );
  XOR2_X1 U784 ( .A(KEYINPUT97), .B(n692), .Z(n693) );
  NAND2_X1 U785 ( .A1(n985), .A2(n693), .ZN(n694) );
  NOR2_X1 U786 ( .A1(n519), .A2(n694), .ZN(n695) );
  AND2_X1 U787 ( .A1(n696), .A2(n695), .ZN(n699) );
  NOR2_X1 U788 ( .A1(n697), .A2(n973), .ZN(n698) );
  NOR2_X1 U789 ( .A1(n699), .A2(n698), .ZN(n705) );
  INV_X1 U790 ( .A(G299), .ZN(n969) );
  NAND2_X1 U791 ( .A1(n701), .A2(G2072), .ZN(n700) );
  XNOR2_X1 U792 ( .A(n700), .B(KEYINPUT27), .ZN(n703) );
  INV_X1 U793 ( .A(G1956), .ZN(n999) );
  NOR2_X1 U794 ( .A1(n999), .A2(n701), .ZN(n702) );
  NOR2_X1 U795 ( .A1(n703), .A2(n702), .ZN(n706) );
  NAND2_X1 U796 ( .A1(n969), .A2(n706), .ZN(n704) );
  NAND2_X1 U797 ( .A1(n705), .A2(n704), .ZN(n710) );
  NOR2_X1 U798 ( .A1(n969), .A2(n706), .ZN(n708) );
  XOR2_X1 U799 ( .A(KEYINPUT96), .B(KEYINPUT28), .Z(n707) );
  XNOR2_X1 U800 ( .A(n708), .B(n707), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  XOR2_X1 U802 ( .A(KEYINPUT29), .B(n711), .Z(n712) );
  NAND2_X1 U803 ( .A1(n713), .A2(n712), .ZN(n726) );
  NAND2_X1 U804 ( .A1(G8), .A2(n714), .ZN(n764) );
  NOR2_X1 U805 ( .A1(G1966), .A2(n764), .ZN(n738) );
  NOR2_X1 U806 ( .A1(G2084), .A2(n714), .ZN(n735) );
  INV_X1 U807 ( .A(n735), .ZN(n715) );
  NAND2_X1 U808 ( .A1(G8), .A2(n715), .ZN(n716) );
  OR2_X1 U809 ( .A1(n738), .A2(n716), .ZN(n718) );
  NOR2_X1 U810 ( .A1(G168), .A2(n719), .ZN(n722) );
  NOR2_X1 U811 ( .A1(G171), .A2(n720), .ZN(n721) );
  NOR2_X1 U812 ( .A1(n722), .A2(n721), .ZN(n724) );
  XNOR2_X1 U813 ( .A(n724), .B(n723), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n726), .A2(n725), .ZN(n736) );
  NAND2_X1 U815 ( .A1(n736), .A2(G286), .ZN(n733) );
  INV_X1 U816 ( .A(G8), .ZN(n731) );
  NOR2_X1 U817 ( .A1(G1971), .A2(n764), .ZN(n728) );
  NOR2_X1 U818 ( .A1(G2090), .A2(n714), .ZN(n727) );
  NOR2_X1 U819 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U820 ( .A1(n729), .A2(G303), .ZN(n730) );
  OR2_X1 U821 ( .A1(n731), .A2(n730), .ZN(n732) );
  XNOR2_X1 U822 ( .A(n734), .B(KEYINPUT32), .ZN(n742) );
  NAND2_X1 U823 ( .A1(G8), .A2(n735), .ZN(n740) );
  INV_X1 U824 ( .A(n736), .ZN(n737) );
  NOR2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n739) );
  NAND2_X1 U826 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U827 ( .A1(n742), .A2(n741), .ZN(n757) );
  NOR2_X1 U828 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NOR2_X1 U829 ( .A1(G1971), .A2(G303), .ZN(n743) );
  NOR2_X1 U830 ( .A1(n748), .A2(n743), .ZN(n981) );
  NAND2_X1 U831 ( .A1(n757), .A2(n981), .ZN(n744) );
  NAND2_X1 U832 ( .A1(G1976), .A2(G288), .ZN(n972) );
  NAND2_X1 U833 ( .A1(n744), .A2(n972), .ZN(n745) );
  NOR2_X1 U834 ( .A1(KEYINPUT33), .A2(n745), .ZN(n746) );
  INV_X1 U835 ( .A(n764), .ZN(n747) );
  NAND2_X1 U836 ( .A1(n746), .A2(n747), .ZN(n751) );
  NAND2_X1 U837 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U838 ( .A1(n749), .A2(KEYINPUT33), .ZN(n750) );
  NAND2_X1 U839 ( .A1(n751), .A2(n750), .ZN(n752) );
  XOR2_X1 U840 ( .A(KEYINPUT99), .B(n752), .Z(n754) );
  XOR2_X1 U841 ( .A(G1981), .B(KEYINPUT100), .Z(n753) );
  XNOR2_X1 U842 ( .A(G305), .B(n753), .ZN(n966) );
  NAND2_X1 U843 ( .A1(n754), .A2(n966), .ZN(n760) );
  NOR2_X1 U844 ( .A1(G2090), .A2(G303), .ZN(n755) );
  NAND2_X1 U845 ( .A1(G8), .A2(n755), .ZN(n756) );
  NAND2_X1 U846 ( .A1(n757), .A2(n756), .ZN(n758) );
  NAND2_X1 U847 ( .A1(n758), .A2(n764), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n762) );
  XOR2_X1 U850 ( .A(n762), .B(KEYINPUT24), .Z(n763) );
  NAND2_X1 U851 ( .A1(G160), .A2(G40), .ZN(n767) );
  NOR2_X1 U852 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U853 ( .A(n768), .B(KEYINPUT88), .Z(n799) );
  INV_X1 U854 ( .A(n799), .ZN(n816) );
  XOR2_X1 U855 ( .A(G2067), .B(KEYINPUT37), .Z(n814) );
  NAND2_X1 U856 ( .A1(n889), .A2(G140), .ZN(n769) );
  XOR2_X1 U857 ( .A(KEYINPUT89), .B(n769), .Z(n771) );
  NAND2_X1 U858 ( .A1(n888), .A2(G104), .ZN(n770) );
  NAND2_X1 U859 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n772), .ZN(n777) );
  NAND2_X1 U861 ( .A1(G116), .A2(n884), .ZN(n774) );
  NAND2_X1 U862 ( .A1(G128), .A2(n885), .ZN(n773) );
  NAND2_X1 U863 ( .A1(n774), .A2(n773), .ZN(n775) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n775), .Z(n776) );
  NOR2_X1 U865 ( .A1(n777), .A2(n776), .ZN(n778) );
  XOR2_X1 U866 ( .A(KEYINPUT36), .B(n778), .Z(n900) );
  NAND2_X1 U867 ( .A1(n814), .A2(n900), .ZN(n779) );
  XOR2_X1 U868 ( .A(KEYINPUT90), .B(n779), .Z(n937) );
  NAND2_X1 U869 ( .A1(n816), .A2(n937), .ZN(n812) );
  NAND2_X1 U870 ( .A1(G105), .A2(n888), .ZN(n780) );
  XOR2_X1 U871 ( .A(KEYINPUT38), .B(n780), .Z(n785) );
  NAND2_X1 U872 ( .A1(G117), .A2(n884), .ZN(n782) );
  NAND2_X1 U873 ( .A1(G129), .A2(n885), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  XOR2_X1 U875 ( .A(KEYINPUT93), .B(n783), .Z(n784) );
  NOR2_X1 U876 ( .A1(n785), .A2(n784), .ZN(n787) );
  NAND2_X1 U877 ( .A1(n889), .A2(G141), .ZN(n786) );
  NAND2_X1 U878 ( .A1(n787), .A2(n786), .ZN(n878) );
  NAND2_X1 U879 ( .A1(G1996), .A2(n878), .ZN(n788) );
  XOR2_X1 U880 ( .A(KEYINPUT94), .B(n788), .Z(n798) );
  NAND2_X1 U881 ( .A1(G119), .A2(n885), .ZN(n795) );
  NAND2_X1 U882 ( .A1(G107), .A2(n884), .ZN(n790) );
  NAND2_X1 U883 ( .A1(G95), .A2(n888), .ZN(n789) );
  NAND2_X1 U884 ( .A1(n790), .A2(n789), .ZN(n793) );
  NAND2_X1 U885 ( .A1(G131), .A2(n889), .ZN(n791) );
  XNOR2_X1 U886 ( .A(KEYINPUT91), .B(n791), .ZN(n792) );
  NOR2_X1 U887 ( .A1(n793), .A2(n792), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(n796), .B(KEYINPUT92), .ZN(n880) );
  AND2_X1 U890 ( .A1(G1991), .A2(n880), .ZN(n797) );
  NOR2_X1 U891 ( .A1(n798), .A2(n797), .ZN(n935) );
  NOR2_X1 U892 ( .A1(n799), .A2(n935), .ZN(n809) );
  INV_X1 U893 ( .A(n809), .ZN(n800) );
  NAND2_X1 U894 ( .A1(n812), .A2(n800), .ZN(n801) );
  XOR2_X1 U895 ( .A(KEYINPUT95), .B(n801), .Z(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n805) );
  XNOR2_X1 U897 ( .A(G1986), .B(G290), .ZN(n979) );
  NAND2_X1 U898 ( .A1(n979), .A2(n816), .ZN(n804) );
  NAND2_X1 U899 ( .A1(n805), .A2(n804), .ZN(n819) );
  NOR2_X1 U900 ( .A1(G1996), .A2(n878), .ZN(n806) );
  XNOR2_X1 U901 ( .A(KEYINPUT102), .B(n806), .ZN(n929) );
  NOR2_X1 U902 ( .A1(G1986), .A2(G290), .ZN(n807) );
  NOR2_X1 U903 ( .A1(G1991), .A2(n880), .ZN(n924) );
  NOR2_X1 U904 ( .A1(n807), .A2(n924), .ZN(n808) );
  NOR2_X1 U905 ( .A1(n809), .A2(n808), .ZN(n810) );
  NOR2_X1 U906 ( .A1(n929), .A2(n810), .ZN(n811) );
  XNOR2_X1 U907 ( .A(KEYINPUT39), .B(n811), .ZN(n813) );
  NAND2_X1 U908 ( .A1(n813), .A2(n812), .ZN(n815) );
  OR2_X1 U909 ( .A1(n814), .A2(n900), .ZN(n921) );
  NAND2_X1 U910 ( .A1(n815), .A2(n921), .ZN(n817) );
  NAND2_X1 U911 ( .A1(n817), .A2(n816), .ZN(n818) );
  NAND2_X1 U912 ( .A1(n819), .A2(n818), .ZN(n820) );
  XNOR2_X1 U913 ( .A(n820), .B(KEYINPUT40), .ZN(G329) );
  XNOR2_X1 U914 ( .A(G2443), .B(G2454), .ZN(n830) );
  XOR2_X1 U915 ( .A(G2430), .B(KEYINPUT104), .Z(n822) );
  XNOR2_X1 U916 ( .A(G2446), .B(KEYINPUT103), .ZN(n821) );
  XNOR2_X1 U917 ( .A(n822), .B(n821), .ZN(n826) );
  XOR2_X1 U918 ( .A(G2451), .B(G2427), .Z(n824) );
  XNOR2_X1 U919 ( .A(G1348), .B(G1341), .ZN(n823) );
  XNOR2_X1 U920 ( .A(n824), .B(n823), .ZN(n825) );
  XOR2_X1 U921 ( .A(n826), .B(n825), .Z(n828) );
  XNOR2_X1 U922 ( .A(G2438), .B(G2435), .ZN(n827) );
  XNOR2_X1 U923 ( .A(n828), .B(n827), .ZN(n829) );
  XNOR2_X1 U924 ( .A(n830), .B(n829), .ZN(n831) );
  NAND2_X1 U925 ( .A1(n831), .A2(G14), .ZN(n910) );
  XNOR2_X1 U926 ( .A(KEYINPUT105), .B(n910), .ZN(G401) );
  NAND2_X1 U927 ( .A1(G2106), .A2(n832), .ZN(G217) );
  AND2_X1 U928 ( .A1(G15), .A2(G2), .ZN(n833) );
  NAND2_X1 U929 ( .A1(G661), .A2(n833), .ZN(G259) );
  NAND2_X1 U930 ( .A1(G3), .A2(G1), .ZN(n834) );
  NAND2_X1 U931 ( .A1(n835), .A2(n834), .ZN(G188) );
  INV_X1 U933 ( .A(G132), .ZN(G219) );
  INV_X1 U934 ( .A(G108), .ZN(G238) );
  INV_X1 U935 ( .A(G82), .ZN(G220) );
  NOR2_X1 U936 ( .A1(n837), .A2(n836), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  INV_X1 U938 ( .A(n838), .ZN(G319) );
  XOR2_X1 U939 ( .A(KEYINPUT109), .B(G1961), .Z(n840) );
  XNOR2_X1 U940 ( .A(G1996), .B(G1991), .ZN(n839) );
  XNOR2_X1 U941 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U942 ( .A(n841), .B(KEYINPUT41), .Z(n843) );
  XNOR2_X1 U943 ( .A(G1981), .B(G1966), .ZN(n842) );
  XNOR2_X1 U944 ( .A(n843), .B(n842), .ZN(n847) );
  XOR2_X1 U945 ( .A(G1956), .B(G1971), .Z(n845) );
  XNOR2_X1 U946 ( .A(G1986), .B(G1976), .ZN(n844) );
  XNOR2_X1 U947 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U948 ( .A(n847), .B(n846), .Z(n849) );
  XNOR2_X1 U949 ( .A(KEYINPUT108), .B(G2474), .ZN(n848) );
  XNOR2_X1 U950 ( .A(n849), .B(n848), .ZN(G229) );
  XOR2_X1 U951 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n851) );
  XNOR2_X1 U952 ( .A(G2678), .B(KEYINPUT43), .ZN(n850) );
  XNOR2_X1 U953 ( .A(n851), .B(n850), .ZN(n855) );
  XOR2_X1 U954 ( .A(KEYINPUT42), .B(G2090), .Z(n853) );
  XNOR2_X1 U955 ( .A(G2067), .B(G2072), .ZN(n852) );
  XNOR2_X1 U956 ( .A(n853), .B(n852), .ZN(n854) );
  XOR2_X1 U957 ( .A(n855), .B(n854), .Z(n857) );
  XNOR2_X1 U958 ( .A(G2096), .B(G2100), .ZN(n856) );
  XNOR2_X1 U959 ( .A(n857), .B(n856), .ZN(n859) );
  XOR2_X1 U960 ( .A(G2078), .B(G2084), .Z(n858) );
  XNOR2_X1 U961 ( .A(n859), .B(n858), .ZN(G227) );
  NAND2_X1 U962 ( .A1(G112), .A2(n884), .ZN(n861) );
  NAND2_X1 U963 ( .A1(G100), .A2(n888), .ZN(n860) );
  NAND2_X1 U964 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U965 ( .A(KEYINPUT110), .B(n862), .ZN(n867) );
  NAND2_X1 U966 ( .A1(n885), .A2(G124), .ZN(n863) );
  XNOR2_X1 U967 ( .A(n863), .B(KEYINPUT44), .ZN(n865) );
  NAND2_X1 U968 ( .A1(G136), .A2(n889), .ZN(n864) );
  NAND2_X1 U969 ( .A1(n865), .A2(n864), .ZN(n866) );
  NOR2_X1 U970 ( .A1(n867), .A2(n866), .ZN(G162) );
  NAND2_X1 U971 ( .A1(G103), .A2(n888), .ZN(n876) );
  NAND2_X1 U972 ( .A1(n889), .A2(G139), .ZN(n868) );
  XNOR2_X1 U973 ( .A(KEYINPUT111), .B(n868), .ZN(n874) );
  NAND2_X1 U974 ( .A1(G115), .A2(n884), .ZN(n870) );
  NAND2_X1 U975 ( .A1(G127), .A2(n885), .ZN(n869) );
  NAND2_X1 U976 ( .A1(n870), .A2(n869), .ZN(n871) );
  XOR2_X1 U977 ( .A(KEYINPUT47), .B(n871), .Z(n872) );
  XNOR2_X1 U978 ( .A(KEYINPUT112), .B(n872), .ZN(n873) );
  NOR2_X1 U979 ( .A1(n874), .A2(n873), .ZN(n875) );
  NAND2_X1 U980 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(n877), .B(KEYINPUT113), .ZN(n916) );
  XNOR2_X1 U982 ( .A(n916), .B(n878), .ZN(n879) );
  XNOR2_X1 U983 ( .A(n879), .B(n923), .ZN(n881) );
  XOR2_X1 U984 ( .A(n881), .B(n880), .Z(n883) );
  XNOR2_X1 U985 ( .A(G164), .B(G160), .ZN(n882) );
  XNOR2_X1 U986 ( .A(n883), .B(n882), .ZN(n902) );
  NAND2_X1 U987 ( .A1(G118), .A2(n884), .ZN(n887) );
  NAND2_X1 U988 ( .A1(G130), .A2(n885), .ZN(n886) );
  NAND2_X1 U989 ( .A1(n887), .A2(n886), .ZN(n894) );
  NAND2_X1 U990 ( .A1(G106), .A2(n888), .ZN(n891) );
  NAND2_X1 U991 ( .A1(G142), .A2(n889), .ZN(n890) );
  NAND2_X1 U992 ( .A1(n891), .A2(n890), .ZN(n892) );
  XOR2_X1 U993 ( .A(n892), .B(KEYINPUT45), .Z(n893) );
  NOR2_X1 U994 ( .A1(n894), .A2(n893), .ZN(n895) );
  XOR2_X1 U995 ( .A(KEYINPUT114), .B(n895), .Z(n896) );
  XOR2_X1 U996 ( .A(n896), .B(KEYINPUT46), .Z(n898) );
  XNOR2_X1 U997 ( .A(G162), .B(KEYINPUT48), .ZN(n897) );
  XNOR2_X1 U998 ( .A(n898), .B(n897), .ZN(n899) );
  XNOR2_X1 U999 ( .A(n900), .B(n899), .ZN(n901) );
  XNOR2_X1 U1000 ( .A(n902), .B(n901), .ZN(n903) );
  NOR2_X1 U1001 ( .A1(G37), .A2(n903), .ZN(G395) );
  XNOR2_X1 U1002 ( .A(KEYINPUT116), .B(KEYINPUT115), .ZN(n906) );
  XNOR2_X1 U1003 ( .A(n973), .B(n904), .ZN(n905) );
  XNOR2_X1 U1004 ( .A(n906), .B(n905), .ZN(n908) );
  XOR2_X1 U1005 ( .A(G286), .B(G171), .Z(n907) );
  XNOR2_X1 U1006 ( .A(n908), .B(n907), .ZN(n909) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n909), .ZN(G397) );
  NAND2_X1 U1008 ( .A1(G319), .A2(n910), .ZN(n913) );
  NOR2_X1 U1009 ( .A1(G229), .A2(G227), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(KEYINPUT49), .B(n911), .ZN(n912) );
  NOR2_X1 U1011 ( .A1(n913), .A2(n912), .ZN(n915) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n914) );
  NAND2_X1 U1013 ( .A1(n915), .A2(n914), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G69), .ZN(G235) );
  INV_X1 U1016 ( .A(G96), .ZN(G221) );
  XOR2_X1 U1017 ( .A(G2072), .B(n916), .Z(n918) );
  XOR2_X1 U1018 ( .A(G164), .B(G2078), .Z(n917) );
  NOR2_X1 U1019 ( .A1(n918), .A2(n917), .ZN(n919) );
  XNOR2_X1 U1020 ( .A(KEYINPUT120), .B(n919), .ZN(n920) );
  XNOR2_X1 U1021 ( .A(n920), .B(KEYINPUT50), .ZN(n922) );
  NAND2_X1 U1022 ( .A1(n922), .A2(n921), .ZN(n940) );
  NOR2_X1 U1023 ( .A1(n924), .A2(n923), .ZN(n927) );
  XOR2_X1 U1024 ( .A(G160), .B(G2084), .Z(n925) );
  XNOR2_X1 U1025 ( .A(KEYINPUT117), .B(n925), .ZN(n926) );
  NAND2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n933) );
  XOR2_X1 U1027 ( .A(G2090), .B(G162), .Z(n928) );
  NOR2_X1 U1028 ( .A1(n929), .A2(n928), .ZN(n930) );
  XOR2_X1 U1029 ( .A(KEYINPUT118), .B(n930), .Z(n931) );
  XOR2_X1 U1030 ( .A(KEYINPUT51), .B(n931), .Z(n932) );
  NOR2_X1 U1031 ( .A1(n933), .A2(n932), .ZN(n934) );
  NAND2_X1 U1032 ( .A1(n935), .A2(n934), .ZN(n936) );
  NOR2_X1 U1033 ( .A1(n937), .A2(n936), .ZN(n938) );
  XNOR2_X1 U1034 ( .A(n938), .B(KEYINPUT119), .ZN(n939) );
  NOR2_X1 U1035 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1036 ( .A(KEYINPUT52), .B(n941), .Z(n942) );
  NOR2_X1 U1037 ( .A1(KEYINPUT55), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT121), .B(n943), .ZN(n944) );
  NAND2_X1 U1039 ( .A1(n944), .A2(G29), .ZN(n1024) );
  XNOR2_X1 U1040 ( .A(G1991), .B(G25), .ZN(n946) );
  XNOR2_X1 U1041 ( .A(G33), .B(G2072), .ZN(n945) );
  NOR2_X1 U1042 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1043 ( .A(G1996), .B(G32), .Z(n947) );
  NAND2_X1 U1044 ( .A1(n947), .A2(G28), .ZN(n950) );
  XNOR2_X1 U1045 ( .A(KEYINPUT122), .B(G2067), .ZN(n948) );
  XNOR2_X1 U1046 ( .A(G26), .B(n948), .ZN(n949) );
  NOR2_X1 U1047 ( .A1(n950), .A2(n949), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XOR2_X1 U1049 ( .A(G27), .B(n953), .Z(n954) );
  NOR2_X1 U1050 ( .A1(n955), .A2(n954), .ZN(n956) );
  XOR2_X1 U1051 ( .A(KEYINPUT53), .B(n956), .Z(n959) );
  XOR2_X1 U1052 ( .A(KEYINPUT54), .B(G34), .Z(n957) );
  XNOR2_X1 U1053 ( .A(G2084), .B(n957), .ZN(n958) );
  NAND2_X1 U1054 ( .A1(n959), .A2(n958), .ZN(n961) );
  XNOR2_X1 U1055 ( .A(G35), .B(G2090), .ZN(n960) );
  NOR2_X1 U1056 ( .A1(n961), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1057 ( .A(KEYINPUT55), .B(n962), .ZN(n964) );
  INV_X1 U1058 ( .A(G29), .ZN(n963) );
  NAND2_X1 U1059 ( .A1(n964), .A2(n963), .ZN(n965) );
  NAND2_X1 U1060 ( .A1(n965), .A2(G11), .ZN(n1022) );
  XNOR2_X1 U1061 ( .A(G16), .B(KEYINPUT56), .ZN(n992) );
  XNOR2_X1 U1062 ( .A(G168), .B(G1966), .ZN(n967) );
  NAND2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  XNOR2_X1 U1064 ( .A(KEYINPUT57), .B(n968), .ZN(n990) );
  XNOR2_X1 U1065 ( .A(n999), .B(n969), .ZN(n970) );
  XNOR2_X1 U1066 ( .A(n970), .B(KEYINPUT123), .ZN(n977) );
  NAND2_X1 U1067 ( .A1(G1971), .A2(G303), .ZN(n971) );
  NAND2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n975) );
  XNOR2_X1 U1069 ( .A(G1348), .B(n973), .ZN(n974) );
  NOR2_X1 U1070 ( .A1(n975), .A2(n974), .ZN(n976) );
  NAND2_X1 U1071 ( .A1(n977), .A2(n976), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(G1961), .B(G301), .ZN(n978) );
  NOR2_X1 U1073 ( .A1(n979), .A2(n978), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(KEYINPUT124), .B(n984), .ZN(n987) );
  XNOR2_X1 U1077 ( .A(n985), .B(G1341), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XNOR2_X1 U1079 ( .A(KEYINPUT125), .B(n988), .ZN(n989) );
  NAND2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n1020) );
  INV_X1 U1082 ( .A(G16), .ZN(n1018) );
  XOR2_X1 U1083 ( .A(G1971), .B(G22), .Z(n995) );
  XNOR2_X1 U1084 ( .A(G1986), .B(KEYINPUT127), .ZN(n993) );
  XNOR2_X1 U1085 ( .A(n993), .B(G24), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n995), .A2(n994), .ZN(n997) );
  XNOR2_X1 U1087 ( .A(G23), .B(G1976), .ZN(n996) );
  NOR2_X1 U1088 ( .A1(n997), .A2(n996), .ZN(n998) );
  XOR2_X1 U1089 ( .A(KEYINPUT58), .B(n998), .Z(n1015) );
  XNOR2_X1 U1090 ( .A(G20), .B(n999), .ZN(n1003) );
  XNOR2_X1 U1091 ( .A(G1981), .B(G6), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(G19), .B(G1341), .ZN(n1000) );
  NOR2_X1 U1093 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NAND2_X1 U1094 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1095 ( .A(KEYINPUT59), .B(G1348), .Z(n1004) );
  XNOR2_X1 U1096 ( .A(G4), .B(n1004), .ZN(n1005) );
  NOR2_X1 U1097 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1098 ( .A(KEYINPUT60), .B(n1007), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(n1008), .B(G5), .ZN(n1009) );
  NAND2_X1 U1100 ( .A1(n1010), .A2(n1009), .ZN(n1012) );
  XNOR2_X1 U1101 ( .A(G21), .B(G1966), .ZN(n1011) );
  NOR2_X1 U1102 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  XOR2_X1 U1103 ( .A(KEYINPUT126), .B(n1013), .Z(n1014) );
  NOR2_X1 U1104 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(KEYINPUT61), .B(n1016), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NAND2_X1 U1107 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  NOR2_X1 U1108 ( .A1(n1022), .A2(n1021), .ZN(n1023) );
  NAND2_X1 U1109 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  XOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1025), .Z(G311) );
  INV_X1 U1111 ( .A(G311), .ZN(G150) );
endmodule

