

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597;

  NOR2_X1 U324 ( .A1(n404), .A2(n403), .ZN(n406) );
  INV_X1 U325 ( .A(n591), .ZN(n466) );
  XNOR2_X1 U326 ( .A(n586), .B(n483), .ZN(n545) );
  XOR2_X1 U327 ( .A(KEYINPUT102), .B(n481), .Z(n292) );
  INV_X1 U328 ( .A(KEYINPUT91), .ZN(n405) );
  XNOR2_X1 U329 ( .A(n406), .B(n405), .ZN(n407) );
  XNOR2_X1 U330 ( .A(n373), .B(n372), .ZN(n375) );
  XNOR2_X1 U331 ( .A(n303), .B(G120GAT), .ZN(n373) );
  INV_X1 U332 ( .A(KEYINPUT75), .ZN(n328) );
  OR2_X1 U333 ( .A1(n595), .A2(n466), .ZN(n467) );
  XNOR2_X1 U334 ( .A(n329), .B(n328), .ZN(n330) );
  INV_X1 U335 ( .A(KEYINPUT65), .ZN(n482) );
  XNOR2_X1 U336 ( .A(n331), .B(n330), .ZN(n336) );
  XNOR2_X1 U337 ( .A(n482), .B(KEYINPUT41), .ZN(n483) );
  AND2_X1 U338 ( .A1(n563), .A2(n562), .ZN(n576) );
  XNOR2_X1 U339 ( .A(n471), .B(KEYINPUT38), .ZN(n480) );
  XOR2_X1 U340 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n294) );
  XNOR2_X1 U341 ( .A(G1GAT), .B(KEYINPUT94), .ZN(n293) );
  XNOR2_X1 U342 ( .A(n294), .B(n293), .ZN(n456) );
  XOR2_X1 U343 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n296) );
  XNOR2_X1 U344 ( .A(KEYINPUT5), .B(KEYINPUT86), .ZN(n295) );
  XNOR2_X1 U345 ( .A(n296), .B(n295), .ZN(n314) );
  XOR2_X1 U346 ( .A(G155GAT), .B(G148GAT), .Z(n298) );
  XNOR2_X1 U347 ( .A(G29GAT), .B(G127GAT), .ZN(n297) );
  XNOR2_X1 U348 ( .A(n298), .B(n297), .ZN(n302) );
  XOR2_X1 U349 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n300) );
  XNOR2_X1 U350 ( .A(G57GAT), .B(G1GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n300), .B(n299), .ZN(n301) );
  XOR2_X1 U352 ( .A(n302), .B(n301), .Z(n312) );
  XNOR2_X1 U353 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n303) );
  XOR2_X1 U354 ( .A(n373), .B(KEYINPUT4), .Z(n305) );
  NAND2_X1 U355 ( .A1(G225GAT), .A2(G233GAT), .ZN(n304) );
  XNOR2_X1 U356 ( .A(n305), .B(n304), .ZN(n310) );
  XNOR2_X1 U357 ( .A(G141GAT), .B(KEYINPUT3), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n306), .B(KEYINPUT2), .ZN(n386) );
  XOR2_X1 U359 ( .A(n386), .B(G162GAT), .Z(n308) );
  XOR2_X1 U360 ( .A(KEYINPUT77), .B(G134GAT), .Z(n418) );
  XNOR2_X1 U361 ( .A(G85GAT), .B(n418), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n309) );
  XNOR2_X1 U363 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n314), .B(n313), .ZN(n558) );
  XOR2_X1 U366 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n316) );
  NAND2_X1 U367 ( .A1(G230GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U368 ( .A(n316), .B(n315), .ZN(n318) );
  INV_X1 U369 ( .A(KEYINPUT33), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n327) );
  INV_X1 U371 ( .A(G176GAT), .ZN(n319) );
  NAND2_X1 U372 ( .A1(G204GAT), .A2(n319), .ZN(n322) );
  INV_X1 U373 ( .A(G204GAT), .ZN(n320) );
  NAND2_X1 U374 ( .A1(n320), .A2(G176GAT), .ZN(n321) );
  NAND2_X1 U375 ( .A1(n322), .A2(n321), .ZN(n324) );
  XNOR2_X1 U376 ( .A(G92GAT), .B(G64GAT), .ZN(n323) );
  XNOR2_X1 U377 ( .A(n324), .B(n323), .ZN(n359) );
  XNOR2_X1 U378 ( .A(G85GAT), .B(KEYINPUT74), .ZN(n325) );
  XNOR2_X1 U379 ( .A(n325), .B(G99GAT), .ZN(n430) );
  XNOR2_X1 U380 ( .A(n359), .B(n430), .ZN(n326) );
  XNOR2_X1 U381 ( .A(n327), .B(n326), .ZN(n331) );
  XOR2_X1 U382 ( .A(G148GAT), .B(G106GAT), .Z(n383) );
  XNOR2_X1 U383 ( .A(G120GAT), .B(n383), .ZN(n329) );
  XOR2_X1 U384 ( .A(G78GAT), .B(G71GAT), .Z(n333) );
  XNOR2_X1 U385 ( .A(KEYINPUT13), .B(KEYINPUT73), .ZN(n332) );
  XNOR2_X1 U386 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U387 ( .A(G57GAT), .B(n334), .Z(n447) );
  INV_X1 U388 ( .A(n447), .ZN(n335) );
  XNOR2_X1 U389 ( .A(n336), .B(n335), .ZN(n586) );
  XOR2_X1 U390 ( .A(KEYINPUT29), .B(G197GAT), .Z(n338) );
  XNOR2_X1 U391 ( .A(G8GAT), .B(G22GAT), .ZN(n337) );
  XNOR2_X1 U392 ( .A(n338), .B(n337), .ZN(n354) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G15GAT), .Z(n340) );
  XNOR2_X1 U394 ( .A(G36GAT), .B(G50GAT), .ZN(n339) );
  XNOR2_X1 U395 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U396 ( .A(G1GAT), .B(KEYINPUT71), .Z(n437) );
  XOR2_X1 U397 ( .A(n341), .B(n437), .Z(n343) );
  XNOR2_X1 U398 ( .A(G113GAT), .B(G141GAT), .ZN(n342) );
  XNOR2_X1 U399 ( .A(n343), .B(n342), .ZN(n347) );
  XOR2_X1 U400 ( .A(KEYINPUT69), .B(KEYINPUT72), .Z(n345) );
  NAND2_X1 U401 ( .A1(G229GAT), .A2(G233GAT), .ZN(n344) );
  XNOR2_X1 U402 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U403 ( .A(n347), .B(n346), .Z(n352) );
  XOR2_X1 U404 ( .A(KEYINPUT70), .B(KEYINPUT8), .Z(n349) );
  XNOR2_X1 U405 ( .A(KEYINPUT7), .B(G43GAT), .ZN(n348) );
  XNOR2_X1 U406 ( .A(n349), .B(n348), .ZN(n350) );
  XOR2_X1 U407 ( .A(G29GAT), .B(n350), .Z(n422) );
  XNOR2_X1 U408 ( .A(n422), .B(KEYINPUT30), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n353) );
  XNOR2_X1 U410 ( .A(n354), .B(n353), .ZN(n581) );
  NOR2_X1 U411 ( .A1(n586), .A2(n581), .ZN(n470) );
  INV_X1 U412 ( .A(n558), .ZN(n501) );
  XOR2_X1 U413 ( .A(KEYINPUT21), .B(G197GAT), .Z(n382) );
  XOR2_X1 U414 ( .A(KEYINPUT89), .B(n382), .Z(n356) );
  NAND2_X1 U415 ( .A1(G226GAT), .A2(G233GAT), .ZN(n355) );
  XNOR2_X1 U416 ( .A(n356), .B(n355), .ZN(n365) );
  XOR2_X1 U417 ( .A(G169GAT), .B(KEYINPUT19), .Z(n358) );
  XNOR2_X1 U418 ( .A(KEYINPUT18), .B(KEYINPUT17), .ZN(n357) );
  XNOR2_X1 U419 ( .A(n358), .B(n357), .ZN(n376) );
  XOR2_X1 U420 ( .A(n359), .B(n376), .Z(n363) );
  XNOR2_X1 U421 ( .A(G218GAT), .B(G36GAT), .ZN(n360) );
  XNOR2_X1 U422 ( .A(n360), .B(G190GAT), .ZN(n417) );
  XNOR2_X1 U423 ( .A(G183GAT), .B(G211GAT), .ZN(n361) );
  XNOR2_X1 U424 ( .A(n361), .B(G8GAT), .ZN(n443) );
  XNOR2_X1 U425 ( .A(n417), .B(n443), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U427 ( .A(n365), .B(n364), .Z(n474) );
  XNOR2_X1 U428 ( .A(n474), .B(KEYINPUT27), .ZN(n409) );
  XOR2_X1 U429 ( .A(G190GAT), .B(G99GAT), .Z(n367) );
  XNOR2_X1 U430 ( .A(G134GAT), .B(G43GAT), .ZN(n366) );
  XNOR2_X1 U431 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U432 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n369) );
  XNOR2_X1 U433 ( .A(G183GAT), .B(KEYINPUT66), .ZN(n368) );
  XNOR2_X1 U434 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n381) );
  XOR2_X1 U436 ( .A(G127GAT), .B(G15GAT), .Z(n441) );
  INV_X1 U437 ( .A(n441), .ZN(n372) );
  NAND2_X1 U438 ( .A1(G227GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U439 ( .A(n375), .B(n374), .ZN(n377) );
  XOR2_X1 U440 ( .A(n377), .B(n376), .Z(n379) );
  XNOR2_X1 U441 ( .A(G71GAT), .B(G176GAT), .ZN(n378) );
  XNOR2_X1 U442 ( .A(n379), .B(n378), .ZN(n380) );
  XNOR2_X1 U443 ( .A(n381), .B(n380), .ZN(n563) );
  XOR2_X1 U444 ( .A(n383), .B(n382), .Z(n385) );
  XOR2_X1 U445 ( .A(G162GAT), .B(G50GAT), .Z(n426) );
  XOR2_X1 U446 ( .A(G155GAT), .B(G22GAT), .Z(n438) );
  XNOR2_X1 U447 ( .A(n426), .B(n438), .ZN(n384) );
  XNOR2_X1 U448 ( .A(n385), .B(n384), .ZN(n390) );
  XOR2_X1 U449 ( .A(G78GAT), .B(n386), .Z(n388) );
  NAND2_X1 U450 ( .A1(G228GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U452 ( .A(n390), .B(n389), .Z(n398) );
  XOR2_X1 U453 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n392) );
  XNOR2_X1 U454 ( .A(G218GAT), .B(KEYINPUT23), .ZN(n391) );
  XNOR2_X1 U455 ( .A(n392), .B(n391), .ZN(n396) );
  XOR2_X1 U456 ( .A(KEYINPUT85), .B(KEYINPUT84), .Z(n394) );
  XNOR2_X1 U457 ( .A(G211GAT), .B(G204GAT), .ZN(n393) );
  XNOR2_X1 U458 ( .A(n394), .B(n393), .ZN(n395) );
  XNOR2_X1 U459 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U460 ( .A(n398), .B(n397), .ZN(n410) );
  INV_X1 U461 ( .A(n410), .ZN(n399) );
  OR2_X1 U462 ( .A1(n563), .A2(n399), .ZN(n400) );
  XNOR2_X1 U463 ( .A(n400), .B(KEYINPUT26), .ZN(n541) );
  NOR2_X1 U464 ( .A1(n409), .A2(n541), .ZN(n404) );
  INV_X1 U465 ( .A(n474), .ZN(n553) );
  NAND2_X1 U466 ( .A1(n563), .A2(n553), .ZN(n401) );
  NAND2_X1 U467 ( .A1(n399), .A2(n401), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n402), .B(KEYINPUT25), .ZN(n403) );
  NOR2_X1 U469 ( .A1(n501), .A2(n407), .ZN(n408) );
  XNOR2_X1 U470 ( .A(n408), .B(KEYINPUT92), .ZN(n415) );
  NOR2_X1 U471 ( .A1(n558), .A2(n409), .ZN(n524) );
  XOR2_X1 U472 ( .A(n410), .B(KEYINPUT68), .Z(n411) );
  XNOR2_X1 U473 ( .A(KEYINPUT28), .B(n411), .ZN(n526) );
  NAND2_X1 U474 ( .A1(n524), .A2(n526), .ZN(n412) );
  NOR2_X1 U475 ( .A1(n563), .A2(n412), .ZN(n413) );
  XNOR2_X1 U476 ( .A(KEYINPUT90), .B(n413), .ZN(n414) );
  NOR2_X1 U477 ( .A1(n415), .A2(n414), .ZN(n416) );
  XOR2_X1 U478 ( .A(KEYINPUT93), .B(n416), .Z(n468) );
  XOR2_X1 U479 ( .A(n418), .B(n417), .Z(n420) );
  NAND2_X1 U480 ( .A1(G232GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U481 ( .A(n420), .B(n419), .ZN(n421) );
  XNOR2_X1 U482 ( .A(n422), .B(n421), .ZN(n434) );
  XOR2_X1 U483 ( .A(KEYINPUT76), .B(KEYINPUT9), .Z(n424) );
  XNOR2_X1 U484 ( .A(G106GAT), .B(G92GAT), .ZN(n423) );
  XNOR2_X1 U485 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U486 ( .A(n425), .B(KEYINPUT11), .Z(n428) );
  XNOR2_X1 U487 ( .A(n426), .B(KEYINPUT78), .ZN(n427) );
  XNOR2_X1 U488 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U489 ( .A(n429), .B(KEYINPUT67), .Z(n432) );
  XNOR2_X1 U490 ( .A(n430), .B(KEYINPUT10), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n575) );
  XOR2_X1 U493 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n436) );
  XNOR2_X1 U494 ( .A(KEYINPUT81), .B(KEYINPUT15), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n451) );
  XOR2_X1 U496 ( .A(KEYINPUT79), .B(G64GAT), .Z(n440) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U498 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U499 ( .A(n442), .B(n441), .Z(n449) );
  XOR2_X1 U500 ( .A(KEYINPUT14), .B(n443), .Z(n445) );
  NAND2_X1 U501 ( .A1(G231GAT), .A2(G233GAT), .ZN(n444) );
  XNOR2_X1 U502 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U503 ( .A(n447), .B(n446), .ZN(n448) );
  XNOR2_X1 U504 ( .A(n449), .B(n448), .ZN(n450) );
  XOR2_X1 U505 ( .A(n451), .B(n450), .Z(n591) );
  NOR2_X1 U506 ( .A1(n575), .A2(n591), .ZN(n452) );
  XOR2_X1 U507 ( .A(KEYINPUT82), .B(n452), .Z(n453) );
  XNOR2_X1 U508 ( .A(KEYINPUT16), .B(n453), .ZN(n454) );
  NOR2_X1 U509 ( .A1(n468), .A2(n454), .ZN(n484) );
  NAND2_X1 U510 ( .A1(n470), .A2(n484), .ZN(n461) );
  NOR2_X1 U511 ( .A1(n558), .A2(n461), .ZN(n455) );
  XOR2_X1 U512 ( .A(n456), .B(n455), .Z(G1324GAT) );
  NOR2_X1 U513 ( .A1(n474), .A2(n461), .ZN(n457) );
  XOR2_X1 U514 ( .A(G8GAT), .B(n457), .Z(G1325GAT) );
  INV_X1 U515 ( .A(n563), .ZN(n528) );
  NOR2_X1 U516 ( .A1(n528), .A2(n461), .ZN(n459) );
  XNOR2_X1 U517 ( .A(KEYINPUT35), .B(KEYINPUT96), .ZN(n458) );
  XNOR2_X1 U518 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U519 ( .A(G15GAT), .B(n460), .ZN(G1326GAT) );
  NOR2_X1 U520 ( .A1(n526), .A2(n461), .ZN(n463) );
  XNOR2_X1 U521 ( .A(KEYINPUT97), .B(KEYINPUT98), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U523 ( .A(G22GAT), .B(n464), .ZN(G1327GAT) );
  XNOR2_X1 U524 ( .A(n575), .B(KEYINPUT99), .ZN(n465) );
  XNOR2_X1 U525 ( .A(n465), .B(KEYINPUT36), .ZN(n595) );
  OR2_X1 U526 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U527 ( .A(KEYINPUT37), .B(n469), .ZN(n499) );
  NAND2_X1 U528 ( .A1(n470), .A2(n499), .ZN(n471) );
  NOR2_X1 U529 ( .A1(n480), .A2(n558), .ZN(n472) );
  XNOR2_X1 U530 ( .A(G29GAT), .B(n472), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT39), .ZN(G1328GAT) );
  NOR2_X1 U532 ( .A1(n474), .A2(n480), .ZN(n475) );
  XOR2_X1 U533 ( .A(G36GAT), .B(n475), .Z(G1329GAT) );
  XOR2_X1 U534 ( .A(KEYINPUT40), .B(KEYINPUT101), .Z(n477) );
  XNOR2_X1 U535 ( .A(G43GAT), .B(KEYINPUT100), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n477), .B(n476), .ZN(n479) );
  NOR2_X1 U537 ( .A1(n480), .A2(n528), .ZN(n478) );
  XOR2_X1 U538 ( .A(n479), .B(n478), .Z(G1330GAT) );
  NOR2_X1 U539 ( .A1(n480), .A2(n526), .ZN(n481) );
  XNOR2_X1 U540 ( .A(G50GAT), .B(n292), .ZN(G1331GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT42), .B(KEYINPUT104), .Z(n487) );
  INV_X1 U542 ( .A(n581), .ZN(n564) );
  NOR2_X1 U543 ( .A1(n564), .A2(n545), .ZN(n498) );
  NAND2_X1 U544 ( .A1(n498), .A2(n484), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT103), .B(n485), .ZN(n493) );
  NAND2_X1 U546 ( .A1(n493), .A2(n501), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n488) );
  XOR2_X1 U548 ( .A(G57GAT), .B(n488), .Z(G1332GAT) );
  XOR2_X1 U549 ( .A(G64GAT), .B(KEYINPUT105), .Z(n490) );
  NAND2_X1 U550 ( .A1(n493), .A2(n553), .ZN(n489) );
  XNOR2_X1 U551 ( .A(n490), .B(n489), .ZN(G1333GAT) );
  NAND2_X1 U552 ( .A1(n493), .A2(n563), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(KEYINPUT106), .ZN(n492) );
  XNOR2_X1 U554 ( .A(G71GAT), .B(n492), .ZN(G1334GAT) );
  XOR2_X1 U555 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n495) );
  INV_X1 U556 ( .A(n526), .ZN(n508) );
  NAND2_X1 U557 ( .A1(n493), .A2(n508), .ZN(n494) );
  XNOR2_X1 U558 ( .A(n495), .B(n494), .ZN(n497) );
  XOR2_X1 U559 ( .A(G78GAT), .B(KEYINPUT107), .Z(n496) );
  XNOR2_X1 U560 ( .A(n497), .B(n496), .ZN(G1335GAT) );
  NAND2_X1 U561 ( .A1(n499), .A2(n498), .ZN(n500) );
  XNOR2_X1 U562 ( .A(KEYINPUT109), .B(n500), .ZN(n509) );
  NAND2_X1 U563 ( .A1(n509), .A2(n501), .ZN(n502) );
  XNOR2_X1 U564 ( .A(n502), .B(KEYINPUT110), .ZN(n503) );
  XNOR2_X1 U565 ( .A(G85GAT), .B(n503), .ZN(G1336GAT) );
  NAND2_X1 U566 ( .A1(n553), .A2(n509), .ZN(n504) );
  XNOR2_X1 U567 ( .A(n504), .B(G92GAT), .ZN(G1337GAT) );
  XOR2_X1 U568 ( .A(KEYINPUT111), .B(KEYINPUT112), .Z(n506) );
  NAND2_X1 U569 ( .A1(n509), .A2(n563), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G99GAT), .B(n507), .ZN(G1338GAT) );
  XOR2_X1 U572 ( .A(KEYINPUT44), .B(KEYINPUT113), .Z(n511) );
  NAND2_X1 U573 ( .A1(n509), .A2(n508), .ZN(n510) );
  XNOR2_X1 U574 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U575 ( .A(G106GAT), .B(n512), .ZN(G1339GAT) );
  NOR2_X1 U576 ( .A1(n581), .A2(n545), .ZN(n513) );
  XNOR2_X1 U577 ( .A(n513), .B(KEYINPUT46), .ZN(n514) );
  NOR2_X1 U578 ( .A1(n575), .A2(n514), .ZN(n515) );
  XNOR2_X1 U579 ( .A(n591), .B(KEYINPUT114), .ZN(n573) );
  NAND2_X1 U580 ( .A1(n515), .A2(n573), .ZN(n516) );
  XNOR2_X1 U581 ( .A(n516), .B(KEYINPUT47), .ZN(n521) );
  NOR2_X1 U582 ( .A1(n595), .A2(n591), .ZN(n517) );
  XNOR2_X1 U583 ( .A(n517), .B(KEYINPUT45), .ZN(n518) );
  NAND2_X1 U584 ( .A1(n518), .A2(n581), .ZN(n519) );
  NOR2_X1 U585 ( .A1(n519), .A2(n586), .ZN(n520) );
  NOR2_X1 U586 ( .A1(n521), .A2(n520), .ZN(n523) );
  XNOR2_X1 U587 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n523), .B(n522), .ZN(n555) );
  INV_X1 U589 ( .A(n524), .ZN(n525) );
  NOR2_X1 U590 ( .A1(n555), .A2(n525), .ZN(n542) );
  NAND2_X1 U591 ( .A1(n542), .A2(n526), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n528), .A2(n527), .ZN(n538) );
  NAND2_X1 U593 ( .A1(n564), .A2(n538), .ZN(n529) );
  XNOR2_X1 U594 ( .A(G113GAT), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT49), .B(KEYINPUT116), .Z(n531) );
  INV_X1 U596 ( .A(n545), .ZN(n567) );
  NAND2_X1 U597 ( .A1(n538), .A2(n567), .ZN(n530) );
  XNOR2_X1 U598 ( .A(n531), .B(n530), .ZN(n533) );
  XOR2_X1 U599 ( .A(G120GAT), .B(KEYINPUT115), .Z(n532) );
  XNOR2_X1 U600 ( .A(n533), .B(n532), .ZN(G1341GAT) );
  INV_X1 U601 ( .A(n538), .ZN(n534) );
  NOR2_X1 U602 ( .A1(n573), .A2(n534), .ZN(n536) );
  XNOR2_X1 U603 ( .A(KEYINPUT50), .B(KEYINPUT117), .ZN(n535) );
  XNOR2_X1 U604 ( .A(n536), .B(n535), .ZN(n537) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n537), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(G134GAT), .B(KEYINPUT51), .Z(n540) );
  NAND2_X1 U607 ( .A1(n538), .A2(n575), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(G1343GAT) );
  INV_X1 U609 ( .A(n541), .ZN(n579) );
  NAND2_X1 U610 ( .A1(n542), .A2(n579), .ZN(n550) );
  NOR2_X1 U611 ( .A1(n581), .A2(n550), .ZN(n543) );
  XOR2_X1 U612 ( .A(G141GAT), .B(n543), .Z(n544) );
  XNOR2_X1 U613 ( .A(KEYINPUT118), .B(n544), .ZN(G1344GAT) );
  NOR2_X1 U614 ( .A1(n545), .A2(n550), .ZN(n547) );
  XNOR2_X1 U615 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n546) );
  XNOR2_X1 U616 ( .A(n547), .B(n546), .ZN(n548) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(n548), .ZN(G1345GAT) );
  NOR2_X1 U618 ( .A1(n591), .A2(n550), .ZN(n549) );
  XOR2_X1 U619 ( .A(G155GAT), .B(n549), .Z(G1346GAT) );
  INV_X1 U620 ( .A(n575), .ZN(n551) );
  NOR2_X1 U621 ( .A1(n551), .A2(n550), .ZN(n552) );
  XOR2_X1 U622 ( .A(G162GAT), .B(n552), .Z(G1347GAT) );
  XOR2_X1 U623 ( .A(KEYINPUT120), .B(KEYINPUT121), .Z(n560) );
  XNOR2_X1 U624 ( .A(KEYINPUT119), .B(n553), .ZN(n554) );
  NOR2_X1 U625 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U626 ( .A(n556), .B(KEYINPUT54), .ZN(n557) );
  AND2_X1 U627 ( .A1(n558), .A2(n557), .ZN(n580) );
  NAND2_X1 U628 ( .A1(n580), .A2(n399), .ZN(n559) );
  XNOR2_X1 U629 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U630 ( .A(KEYINPUT55), .B(n561), .ZN(n562) );
  NAND2_X1 U631 ( .A1(n576), .A2(n564), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(KEYINPUT122), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G169GAT), .B(n566), .ZN(G1348GAT) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT57), .Z(n569) );
  NAND2_X1 U635 ( .A1(n576), .A2(n567), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n571) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT123), .Z(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(G1349GAT) );
  INV_X1 U639 ( .A(n576), .ZN(n572) );
  NOR2_X1 U640 ( .A1(n573), .A2(n572), .ZN(n574) );
  XOR2_X1 U641 ( .A(G183GAT), .B(n574), .Z(G1350GAT) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n577), .B(KEYINPUT58), .ZN(n578) );
  XNOR2_X1 U644 ( .A(G190GAT), .B(n578), .ZN(G1351GAT) );
  NAND2_X1 U645 ( .A1(n580), .A2(n579), .ZN(n594) );
  NOR2_X1 U646 ( .A1(n581), .A2(n594), .ZN(n585) );
  XNOR2_X1 U647 ( .A(G197GAT), .B(KEYINPUT59), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n582), .B(KEYINPUT60), .ZN(n583) );
  XNOR2_X1 U649 ( .A(KEYINPUT124), .B(n583), .ZN(n584) );
  XNOR2_X1 U650 ( .A(n585), .B(n584), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n589) );
  INV_X1 U652 ( .A(n594), .ZN(n587) );
  NAND2_X1 U653 ( .A1(n587), .A2(n586), .ZN(n588) );
  XNOR2_X1 U654 ( .A(n589), .B(n588), .ZN(n590) );
  XOR2_X1 U655 ( .A(G204GAT), .B(n590), .Z(G1353GAT) );
  NOR2_X1 U656 ( .A1(n591), .A2(n594), .ZN(n592) );
  XOR2_X1 U657 ( .A(KEYINPUT126), .B(n592), .Z(n593) );
  XNOR2_X1 U658 ( .A(G211GAT), .B(n593), .ZN(G1354GAT) );
  NOR2_X1 U659 ( .A1(n595), .A2(n594), .ZN(n596) );
  XOR2_X1 U660 ( .A(KEYINPUT62), .B(n596), .Z(n597) );
  XNOR2_X1 U661 ( .A(G218GAT), .B(n597), .ZN(G1355GAT) );
endmodule

