

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788;

  OR2_X1 U378 ( .A1(n588), .A2(n572), .ZN(n691) );
  OR2_X1 U379 ( .A1(n613), .A2(n527), .ZN(n530) );
  AND2_X2 U380 ( .A1(n576), .A2(n577), .ZN(n565) );
  NOR2_X1 U381 ( .A1(G902), .A2(n742), .ZN(n466) );
  BUF_X1 U382 ( .A(G953), .Z(n783) );
  NAND2_X2 U383 ( .A1(n388), .A2(n387), .ZN(n666) );
  AND2_X2 U384 ( .A1(n389), .A2(n425), .ZN(n388) );
  XNOR2_X2 U385 ( .A(n456), .B(KEYINPUT67), .ZN(n382) );
  OR2_X1 U386 ( .A1(n365), .A2(n366), .ZN(n683) );
  NAND2_X2 U387 ( .A1(n430), .A2(n426), .ZN(n621) );
  AND2_X1 U388 ( .A1(n381), .A2(n401), .ZN(n399) );
  NAND2_X1 U389 ( .A1(n585), .A2(n363), .ZN(n589) );
  XNOR2_X1 U390 ( .A(n630), .B(n629), .ZN(n692) );
  XNOR2_X1 U391 ( .A(n550), .B(n506), .ZN(n613) );
  OR2_X1 U392 ( .A1(n532), .A2(n644), .ZN(n535) );
  XNOR2_X1 U393 ( .A(n707), .B(n708), .ZN(n709) );
  XOR2_X1 U394 ( .A(n747), .B(KEYINPUT59), .Z(n748) );
  XNOR2_X1 U395 ( .A(n477), .B(n478), .ZN(n714) );
  XNOR2_X1 U396 ( .A(G137), .B(KEYINPUT68), .ZN(n457) );
  INV_X1 U397 ( .A(n550), .ZN(n355) );
  XNOR2_X1 U398 ( .A(n505), .B(n362), .ZN(n361) );
  NOR2_X2 U399 ( .A1(n695), .A2(n672), .ZN(n674) );
  INV_X4 U400 ( .A(G953), .ZN(n779) );
  INV_X1 U401 ( .A(KEYINPUT99), .ZN(n418) );
  XNOR2_X1 U402 ( .A(G119), .B(G116), .ZN(n473) );
  NAND2_X1 U403 ( .A1(n621), .A2(n660), .ZN(n609) );
  INV_X1 U404 ( .A(G472), .ZN(n429) );
  NAND2_X1 U405 ( .A1(G902), .A2(G472), .ZN(n431) );
  XNOR2_X1 U406 ( .A(G119), .B(G128), .ZN(n444) );
  XNOR2_X1 U407 ( .A(n394), .B(n393), .ZN(n392) );
  XNOR2_X1 U408 ( .A(KEYINPUT23), .B(KEYINPUT96), .ZN(n393) );
  XNOR2_X1 U409 ( .A(n457), .B(KEYINPUT24), .ZN(n394) );
  XOR2_X1 U410 ( .A(G131), .B(G140), .Z(n520) );
  XNOR2_X1 U411 ( .A(n519), .B(n414), .ZN(n522) );
  XNOR2_X1 U412 ( .A(n518), .B(n415), .ZN(n414) );
  XNOR2_X1 U413 ( .A(G143), .B(G122), .ZN(n516) );
  XNOR2_X1 U414 ( .A(n494), .B(KEYINPUT10), .ZN(n774) );
  XNOR2_X1 U415 ( .A(n411), .B(n410), .ZN(n577) );
  XNOR2_X1 U416 ( .A(n525), .B(G475), .ZN(n410) );
  OR2_X1 U417 ( .A1(n747), .A2(G902), .ZN(n411) );
  XOR2_X1 U418 ( .A(KEYINPUT98), .B(G131), .Z(n468) );
  XOR2_X1 U419 ( .A(KEYINPUT5), .B(G137), .Z(n470) );
  NAND2_X1 U420 ( .A1(n779), .A2(n412), .ZN(n415) );
  NOR2_X1 U421 ( .A1(n413), .A2(G237), .ZN(n412) );
  INV_X1 U422 ( .A(G214), .ZN(n413) );
  XOR2_X1 U423 ( .A(KEYINPUT12), .B(KEYINPUT11), .Z(n518) );
  XOR2_X1 U424 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n517) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n442) );
  INV_X1 U426 ( .A(G237), .ZN(n502) );
  XNOR2_X1 U427 ( .A(G902), .B(KEYINPUT15), .ZN(n699) );
  INV_X1 U428 ( .A(n536), .ZN(n576) );
  XNOR2_X1 U429 ( .A(G110), .B(KEYINPUT78), .ZN(n459) );
  XNOR2_X1 U430 ( .A(KEYINPUT16), .B(G122), .ZN(n499) );
  XNOR2_X1 U431 ( .A(G122), .B(KEYINPUT104), .ZN(n507) );
  XOR2_X1 U432 ( .A(KEYINPUT103), .B(KEYINPUT9), .Z(n508) );
  NAND2_X1 U433 ( .A1(n526), .A2(G214), .ZN(n660) );
  NAND2_X1 U434 ( .A1(n613), .A2(KEYINPUT39), .ZN(n425) );
  INV_X1 U435 ( .A(KEYINPUT31), .ZN(n439) );
  AND2_X1 U436 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U437 ( .A1(n429), .A2(n428), .ZN(n427) );
  XNOR2_X1 U438 ( .A(n714), .B(KEYINPUT62), .ZN(n715) );
  XNOR2_X1 U439 ( .A(n391), .B(n390), .ZN(n757) );
  XNOR2_X1 U440 ( .A(n446), .B(n774), .ZN(n390) );
  XNOR2_X1 U441 ( .A(n441), .B(n392), .ZN(n391) );
  XNOR2_X1 U442 ( .A(n524), .B(n523), .ZN(n747) );
  XNOR2_X1 U443 ( .A(n522), .B(n521), .ZN(n524) );
  AND2_X1 U444 ( .A1(n711), .A2(n783), .ZN(n761) );
  AND2_X1 U445 ( .A1(n635), .A2(n634), .ZN(n724) );
  INV_X1 U446 ( .A(n361), .ZN(n550) );
  AND2_X1 U447 ( .A1(n691), .A2(KEYINPUT107), .ZN(n356) );
  AND2_X1 U448 ( .A1(n620), .A2(n619), .ZN(n357) );
  NAND2_X1 U449 ( .A1(n643), .A2(n642), .ZN(n358) );
  INV_X1 U450 ( .A(G902), .ZN(n428) );
  INV_X1 U451 ( .A(KEYINPUT107), .ZN(n436) );
  INV_X1 U452 ( .A(KEYINPUT73), .ZN(n591) );
  XOR2_X1 U453 ( .A(n359), .B(n360), .Z(n364) );
  XNOR2_X1 U454 ( .A(n509), .B(KEYINPUT7), .ZN(n359) );
  XOR2_X1 U455 ( .A(G116), .B(G107), .Z(n360) );
  XOR2_X1 U456 ( .A(n504), .B(n503), .Z(n362) );
  XNOR2_X1 U457 ( .A(n440), .B(n439), .ZN(n563) );
  NAND2_X1 U458 ( .A1(n384), .A2(n383), .ZN(n405) );
  NOR2_X1 U459 ( .A1(n587), .A2(n380), .ZN(n363) );
  XNOR2_X1 U460 ( .A(n405), .B(n631), .ZN(n404) );
  XNOR2_X1 U461 ( .A(n364), .B(n510), .ZN(n513) );
  XNOR2_X1 U462 ( .A(n515), .B(n514), .ZN(n536) );
  NAND2_X1 U463 ( .A1(n563), .A2(n562), .ZN(n419) );
  XNOR2_X1 U464 ( .A(n520), .B(n457), .ZN(n775) );
  INV_X1 U465 ( .A(n403), .ZN(n398) );
  NOR2_X2 U466 ( .A1(n617), .A2(n610), .ZN(n611) );
  NAND2_X1 U467 ( .A1(n680), .A2(n679), .ZN(n365) );
  OR2_X1 U468 ( .A1(n783), .A2(n681), .ZN(n366) );
  NAND2_X1 U469 ( .A1(n496), .A2(n495), .ZN(n369) );
  NAND2_X1 U470 ( .A1(n367), .A2(n368), .ZN(n370) );
  NAND2_X1 U471 ( .A1(n370), .A2(n369), .ZN(n498) );
  INV_X1 U472 ( .A(n496), .ZN(n367) );
  INV_X1 U473 ( .A(n495), .ZN(n368) );
  NAND2_X1 U474 ( .A1(n417), .A2(n636), .ZN(n371) );
  XNOR2_X2 U475 ( .A(n419), .B(n418), .ZN(n417) );
  NAND2_X1 U476 ( .A1(n564), .A2(n560), .ZN(n440) );
  BUF_X1 U477 ( .A(n564), .Z(n573) );
  XNOR2_X1 U478 ( .A(n416), .B(KEYINPUT106), .ZN(n372) );
  XNOR2_X1 U479 ( .A(n371), .B(KEYINPUT106), .ZN(n438) );
  BUF_X1 U480 ( .A(n746), .Z(n756) );
  BUF_X1 U481 ( .A(n695), .Z(n778) );
  NAND2_X1 U482 ( .A1(n668), .A2(n667), .ZN(n695) );
  XNOR2_X1 U483 ( .A(n420), .B(KEYINPUT89), .ZN(n668) );
  INV_X1 U484 ( .A(n692), .ZN(n383) );
  AND2_X1 U485 ( .A1(n581), .A2(n435), .ZN(n373) );
  XNOR2_X1 U486 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n374) );
  XNOR2_X1 U487 ( .A(n580), .B(n579), .ZN(n375) );
  XNOR2_X1 U488 ( .A(n580), .B(n579), .ZN(n788) );
  BUF_X1 U489 ( .A(n563), .Z(n376) );
  NAND2_X1 U490 ( .A1(n703), .A2(n702), .ZN(n705) );
  AND2_X2 U491 ( .A1(n705), .A2(n704), .ZN(n746) );
  XNOR2_X2 U492 ( .A(n377), .B(n378), .ZN(n564) );
  NOR2_X2 U493 ( .A1(n632), .A2(n558), .ZN(n377) );
  XOR2_X1 U494 ( .A(n559), .B(KEYINPUT0), .Z(n378) );
  NAND2_X1 U495 ( .A1(n734), .A2(n409), .ZN(n408) );
  XNOR2_X2 U496 ( .A(n776), .B(G146), .ZN(n478) );
  XNOR2_X1 U497 ( .A(n379), .B(KEYINPUT108), .ZN(n645) );
  NAND2_X1 U498 ( .A1(n380), .A2(n357), .ZN(n379) );
  INV_X1 U499 ( .A(n644), .ZN(n380) );
  XNOR2_X1 U500 ( .A(n551), .B(KEYINPUT91), .ZN(n647) );
  NAND2_X1 U501 ( .A1(n398), .A2(n396), .ZN(n395) );
  NAND2_X1 U502 ( .A1(n581), .A2(n435), .ZN(n434) );
  INV_X1 U503 ( .A(n691), .ZN(n437) );
  NAND2_X1 U504 ( .A1(n400), .A2(n582), .ZN(n381) );
  NAND2_X1 U505 ( .A1(n417), .A2(n636), .ZN(n416) );
  NAND2_X1 U506 ( .A1(n382), .A2(n624), .ZN(n605) );
  NAND2_X1 U507 ( .A1(n663), .A2(n382), .ZN(n532) );
  NOR2_X1 U508 ( .A1(n663), .A2(n382), .ZN(n481) );
  INV_X1 U509 ( .A(n385), .ZN(n384) );
  XNOR2_X1 U510 ( .A(n385), .B(G131), .ZN(n787) );
  XNOR2_X2 U511 ( .A(n616), .B(n615), .ZN(n385) );
  NAND2_X1 U512 ( .A1(n612), .A2(n611), .ZN(n657) );
  NAND2_X1 U513 ( .A1(n612), .A2(n386), .ZN(n389) );
  AND2_X1 U514 ( .A1(n424), .A2(n611), .ZN(n386) );
  NAND2_X1 U515 ( .A1(n657), .A2(KEYINPUT39), .ZN(n387) );
  NAND2_X1 U516 ( .A1(n399), .A2(n395), .ZN(n602) );
  AND2_X1 U517 ( .A1(n402), .A2(n397), .ZN(n396) );
  NOR2_X1 U518 ( .A1(n434), .A2(n582), .ZN(n397) );
  NAND2_X1 U519 ( .A1(n373), .A2(n402), .ZN(n400) );
  NAND2_X1 U520 ( .A1(n403), .A2(n582), .ZN(n401) );
  NAND2_X1 U521 ( .A1(n438), .A2(n356), .ZN(n402) );
  NOR2_X2 U522 ( .A1(n372), .A2(KEYINPUT107), .ZN(n403) );
  NAND2_X1 U523 ( .A1(n406), .A2(n404), .ZN(n422) );
  AND2_X1 U524 ( .A1(n407), .A2(n358), .ZN(n406) );
  NOR2_X1 U525 ( .A1(n658), .A2(n408), .ZN(n407) );
  INV_X1 U526 ( .A(n729), .ZN(n409) );
  NOR2_X1 U527 ( .A1(n783), .A2(G237), .ZN(n423) );
  NAND2_X1 U528 ( .A1(n421), .A2(n737), .ZN(n420) );
  XNOR2_X1 U529 ( .A(n422), .B(n659), .ZN(n421) );
  NAND2_X1 U530 ( .A1(n423), .A2(G210), .ZN(n469) );
  NAND2_X1 U531 ( .A1(n666), .A2(n731), .ZN(n616) );
  NOR2_X1 U532 ( .A1(n613), .A2(KEYINPUT39), .ZN(n424) );
  NAND2_X1 U533 ( .A1(n714), .A2(G472), .ZN(n432) );
  OR2_X1 U534 ( .A1(n714), .A2(n427), .ZN(n426) );
  XNOR2_X1 U535 ( .A(n488), .B(n433), .ZN(n492) );
  XNOR2_X2 U536 ( .A(KEYINPUT18), .B(KEYINPUT81), .ZN(n433) );
  XNOR2_X2 U537 ( .A(KEYINPUT64), .B(KEYINPUT4), .ZN(n488) );
  NAND2_X1 U538 ( .A1(n437), .A2(n436), .ZN(n435) );
  INV_X1 U539 ( .A(n376), .ZN(n685) );
  XNOR2_X1 U540 ( .A(n647), .B(KEYINPUT19), .ZN(n632) );
  AND2_X1 U541 ( .A1(n564), .A2(n561), .ZN(n720) );
  AND2_X1 U542 ( .A1(n511), .A2(G221), .ZN(n441) );
  INV_X1 U543 ( .A(n720), .ZN(n562) );
  INV_X1 U544 ( .A(KEYINPUT46), .ZN(n631) );
  XNOR2_X1 U545 ( .A(n592), .B(n591), .ZN(n594) );
  XNOR2_X1 U546 ( .A(n533), .B(KEYINPUT93), .ZN(n534) );
  XNOR2_X1 U547 ( .A(n442), .B(KEYINPUT14), .ZN(n443) );
  XNOR2_X1 U548 ( .A(KEYINPUT76), .B(n443), .ZN(n552) );
  NAND2_X1 U549 ( .A1(G952), .A2(n552), .ZN(n555) );
  XOR2_X1 U550 ( .A(G110), .B(G140), .Z(n445) );
  XNOR2_X1 U551 ( .A(n445), .B(n444), .ZN(n446) );
  XNOR2_X1 U552 ( .A(G146), .B(G125), .ZN(n494) );
  NAND2_X1 U553 ( .A1(G234), .A2(n779), .ZN(n447) );
  XOR2_X1 U554 ( .A(KEYINPUT8), .B(n447), .Z(n511) );
  NOR2_X1 U555 ( .A1(n757), .A2(G902), .ZN(n453) );
  XOR2_X1 U556 ( .A(KEYINPUT25), .B(KEYINPUT80), .Z(n451) );
  XOR2_X1 U557 ( .A(KEYINPUT97), .B(KEYINPUT20), .Z(n449) );
  NAND2_X1 U558 ( .A1(G234), .A2(n699), .ZN(n448) );
  XNOR2_X1 U559 ( .A(n449), .B(n448), .ZN(n454) );
  AND2_X1 U560 ( .A1(n454), .A2(G217), .ZN(n450) );
  XNOR2_X1 U561 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X2 U562 ( .A(n453), .B(n452), .ZN(n618) );
  AND2_X1 U563 ( .A1(n454), .A2(G221), .ZN(n455) );
  XNOR2_X1 U564 ( .A(n455), .B(KEYINPUT21), .ZN(n619) );
  NAND2_X1 U565 ( .A1(n618), .A2(n619), .ZN(n456) );
  NAND2_X1 U566 ( .A1(G227), .A2(n779), .ZN(n458) );
  XNOR2_X1 U567 ( .A(n775), .B(n458), .ZN(n463) );
  INV_X1 U568 ( .A(n459), .ZN(n461) );
  XNOR2_X1 U569 ( .A(G107), .B(G104), .ZN(n460) );
  XNOR2_X1 U570 ( .A(n461), .B(n460), .ZN(n767) );
  XNOR2_X1 U571 ( .A(KEYINPUT66), .B(G101), .ZN(n467) );
  XNOR2_X1 U572 ( .A(n467), .B(KEYINPUT71), .ZN(n462) );
  XNOR2_X1 U573 ( .A(n767), .B(n462), .ZN(n497) );
  XNOR2_X1 U574 ( .A(n463), .B(n497), .ZN(n464) );
  XNOR2_X2 U575 ( .A(G143), .B(G128), .ZN(n493) );
  XNOR2_X1 U576 ( .A(n493), .B(G134), .ZN(n510) );
  XNOR2_X1 U577 ( .A(n374), .B(n510), .ZN(n776) );
  XNOR2_X1 U578 ( .A(n464), .B(n478), .ZN(n742) );
  XNOR2_X1 U579 ( .A(KEYINPUT69), .B(G469), .ZN(n465) );
  XNOR2_X2 U580 ( .A(n466), .B(n465), .ZN(n624) );
  XNOR2_X2 U581 ( .A(n624), .B(KEYINPUT1), .ZN(n663) );
  XNOR2_X1 U582 ( .A(n468), .B(n467), .ZN(n472) );
  XNOR2_X1 U583 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U584 ( .A(n472), .B(n471), .ZN(n476) );
  XNOR2_X1 U585 ( .A(n473), .B(KEYINPUT3), .ZN(n475) );
  XNOR2_X1 U586 ( .A(G113), .B(KEYINPUT70), .ZN(n474) );
  XNOR2_X1 U587 ( .A(n475), .B(n474), .ZN(n500) );
  XNOR2_X1 U588 ( .A(n476), .B(n500), .ZN(n477) );
  INV_X1 U589 ( .A(n621), .ZN(n479) );
  NOR2_X1 U590 ( .A1(n532), .A2(n479), .ZN(n560) );
  NOR2_X1 U591 ( .A1(n618), .A2(n619), .ZN(n480) );
  XNOR2_X1 U592 ( .A(KEYINPUT49), .B(n480), .ZN(n484) );
  XOR2_X1 U593 ( .A(KEYINPUT50), .B(n481), .Z(n482) );
  XNOR2_X1 U594 ( .A(KEYINPUT122), .B(n482), .ZN(n483) );
  NAND2_X1 U595 ( .A1(n484), .A2(n483), .ZN(n485) );
  NOR2_X1 U596 ( .A1(n621), .A2(n485), .ZN(n486) );
  NOR2_X1 U597 ( .A1(n560), .A2(n486), .ZN(n487) );
  XNOR2_X1 U598 ( .A(KEYINPUT51), .B(n487), .ZN(n531) );
  NAND2_X1 U599 ( .A1(n779), .A2(G224), .ZN(n490) );
  XNOR2_X2 U600 ( .A(KEYINPUT94), .B(KEYINPUT17), .ZN(n489) );
  XNOR2_X1 U601 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U602 ( .A(n491), .B(n492), .ZN(n496) );
  XNOR2_X1 U603 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U604 ( .A(n498), .B(n497), .ZN(n501) );
  XNOR2_X1 U605 ( .A(n500), .B(n499), .ZN(n769) );
  XNOR2_X1 U606 ( .A(n501), .B(n769), .ZN(n706) );
  NAND2_X1 U607 ( .A1(n706), .A2(n699), .ZN(n505) );
  NAND2_X1 U608 ( .A1(n428), .A2(n502), .ZN(n526) );
  NAND2_X1 U609 ( .A1(n526), .A2(G210), .ZN(n504) );
  INV_X1 U610 ( .A(KEYINPUT83), .ZN(n503) );
  XNOR2_X1 U611 ( .A(KEYINPUT77), .B(KEYINPUT38), .ZN(n506) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n509) );
  NAND2_X1 U613 ( .A1(G217), .A2(n511), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n513), .B(n512), .ZN(n752) );
  NOR2_X1 U615 ( .A1(G902), .A2(n752), .ZN(n515) );
  INV_X1 U616 ( .A(G478), .ZN(n514) );
  XNOR2_X1 U617 ( .A(KEYINPUT102), .B(KEYINPUT13), .ZN(n525) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n519) );
  XOR2_X1 U619 ( .A(n520), .B(G104), .Z(n521) );
  XNOR2_X1 U620 ( .A(n774), .B(G113), .ZN(n523) );
  NAND2_X1 U621 ( .A1(n565), .A2(n660), .ZN(n527) );
  INV_X1 U622 ( .A(KEYINPUT113), .ZN(n528) );
  XNOR2_X1 U623 ( .A(n528), .B(KEYINPUT41), .ZN(n529) );
  XNOR2_X2 U624 ( .A(n530), .B(n529), .ZN(n677) );
  NAND2_X1 U625 ( .A1(n531), .A2(n677), .ZN(n547) );
  XNOR2_X1 U626 ( .A(n621), .B(KEYINPUT6), .ZN(n644) );
  XOR2_X1 U627 ( .A(KEYINPUT33), .B(KEYINPUT72), .Z(n533) );
  XNOR2_X2 U628 ( .A(n535), .B(n534), .ZN(n678) );
  AND2_X1 U629 ( .A1(n577), .A2(n536), .ZN(n725) );
  INV_X1 U630 ( .A(n725), .ZN(n537) );
  OR2_X1 U631 ( .A1(n577), .A2(n536), .ZN(n646) );
  NAND2_X1 U632 ( .A1(n537), .A2(n646), .ZN(n538) );
  XNOR2_X1 U633 ( .A(n538), .B(KEYINPUT105), .ZN(n650) );
  INV_X1 U634 ( .A(n660), .ZN(n541) );
  NOR2_X1 U635 ( .A1(n650), .A2(n541), .ZN(n540) );
  INV_X1 U636 ( .A(n613), .ZN(n539) );
  NAND2_X1 U637 ( .A1(n540), .A2(n539), .ZN(n544) );
  NAND2_X1 U638 ( .A1(n613), .A2(n541), .ZN(n542) );
  NAND2_X1 U639 ( .A1(n542), .A2(n565), .ZN(n543) );
  NAND2_X1 U640 ( .A1(n544), .A2(n543), .ZN(n545) );
  NAND2_X1 U641 ( .A1(n678), .A2(n545), .ZN(n546) );
  NAND2_X1 U642 ( .A1(n547), .A2(n546), .ZN(n548) );
  XOR2_X1 U643 ( .A(KEYINPUT52), .B(n548), .Z(n549) );
  NOR2_X1 U644 ( .A1(n555), .A2(n549), .ZN(n681) );
  NAND2_X1 U645 ( .A1(n361), .A2(n660), .ZN(n551) );
  AND2_X1 U646 ( .A1(n552), .A2(n783), .ZN(n553) );
  NAND2_X1 U647 ( .A1(G902), .A2(n553), .ZN(n606) );
  NOR2_X1 U648 ( .A1(G898), .A2(n606), .ZN(n554) );
  XNOR2_X1 U649 ( .A(n554), .B(KEYINPUT95), .ZN(n557) );
  NOR2_X1 U650 ( .A1(n555), .A2(n783), .ZN(n608) );
  INV_X1 U651 ( .A(n608), .ZN(n556) );
  AND2_X1 U652 ( .A1(n557), .A2(n556), .ZN(n558) );
  INV_X1 U653 ( .A(KEYINPUT92), .ZN(n559) );
  NOR2_X1 U654 ( .A1(n605), .A2(n621), .ZN(n561) );
  INV_X1 U655 ( .A(n565), .ZN(n567) );
  INV_X1 U656 ( .A(n619), .ZN(n566) );
  NOR2_X1 U657 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U658 ( .A1(n573), .A2(n568), .ZN(n570) );
  XNOR2_X1 U659 ( .A(KEYINPUT74), .B(KEYINPUT22), .ZN(n569) );
  XNOR2_X1 U660 ( .A(n570), .B(n569), .ZN(n588) );
  INV_X1 U661 ( .A(n618), .ZN(n586) );
  NOR2_X1 U662 ( .A1(n586), .A2(n663), .ZN(n571) );
  NAND2_X1 U663 ( .A1(n571), .A2(n644), .ZN(n572) );
  NAND2_X1 U664 ( .A1(n678), .A2(n573), .ZN(n575) );
  XOR2_X1 U665 ( .A(KEYINPUT34), .B(KEYINPUT82), .Z(n574) );
  XNOR2_X1 U666 ( .A(n575), .B(n574), .ZN(n578) );
  NOR2_X1 U667 ( .A1(n577), .A2(n576), .ZN(n655) );
  NAND2_X1 U668 ( .A1(n578), .A2(n655), .ZN(n580) );
  XNOR2_X1 U669 ( .A(KEYINPUT88), .B(KEYINPUT35), .ZN(n579) );
  NAND2_X1 U670 ( .A1(n788), .A2(KEYINPUT44), .ZN(n581) );
  INV_X1 U671 ( .A(KEYINPUT90), .ZN(n582) );
  INV_X1 U672 ( .A(n588), .ZN(n585) );
  OR2_X1 U673 ( .A1(n618), .A2(n621), .ZN(n583) );
  NOR2_X1 U674 ( .A1(n663), .A2(n583), .ZN(n584) );
  AND2_X1 U675 ( .A1(n585), .A2(n584), .ZN(n690) );
  NOR2_X1 U676 ( .A1(n375), .A2(n690), .ZN(n590) );
  NAND2_X1 U677 ( .A1(n586), .A2(n663), .ZN(n587) );
  XNOR2_X2 U678 ( .A(n589), .B(KEYINPUT32), .ZN(n693) );
  NAND2_X1 U679 ( .A1(n590), .A2(n693), .ZN(n592) );
  INV_X1 U680 ( .A(KEYINPUT44), .ZN(n593) );
  NAND2_X1 U681 ( .A1(n594), .A2(n593), .ZN(n600) );
  INV_X1 U682 ( .A(n693), .ZN(n598) );
  INV_X1 U683 ( .A(n690), .ZN(n596) );
  AND2_X1 U684 ( .A1(n591), .A2(KEYINPUT44), .ZN(n595) );
  NAND2_X1 U685 ( .A1(n596), .A2(n595), .ZN(n597) );
  OR2_X1 U686 ( .A1(n598), .A2(n597), .ZN(n599) );
  NAND2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n601) );
  NAND2_X1 U688 ( .A1(n602), .A2(n601), .ZN(n604) );
  INV_X1 U689 ( .A(KEYINPUT45), .ZN(n603) );
  XNOR2_X2 U690 ( .A(n604), .B(n603), .ZN(n694) );
  INV_X1 U691 ( .A(n694), .ZN(n762) );
  XNOR2_X1 U692 ( .A(KEYINPUT109), .B(n605), .ZN(n612) );
  NOR2_X1 U693 ( .A1(G900), .A2(n606), .ZN(n607) );
  NOR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n617) );
  XNOR2_X1 U695 ( .A(KEYINPUT30), .B(n609), .ZN(n610) );
  INV_X1 U696 ( .A(n646), .ZN(n731) );
  INV_X1 U697 ( .A(KEYINPUT112), .ZN(n614) );
  XNOR2_X1 U698 ( .A(n614), .B(KEYINPUT40), .ZN(n615) );
  XOR2_X1 U699 ( .A(KEYINPUT110), .B(KEYINPUT28), .Z(n623) );
  NOR2_X1 U700 ( .A1(n618), .A2(n617), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n357), .A2(n621), .ZN(n622) );
  XNOR2_X1 U702 ( .A(n623), .B(n622), .ZN(n625) );
  AND2_X1 U703 ( .A1(n625), .A2(n624), .ZN(n627) );
  INV_X1 U704 ( .A(KEYINPUT111), .ZN(n626) );
  XNOR2_X1 U705 ( .A(n627), .B(n626), .ZN(n635) );
  NAND2_X1 U706 ( .A1(n635), .A2(n677), .ZN(n630) );
  INV_X1 U707 ( .A(KEYINPUT114), .ZN(n628) );
  XNOR2_X1 U708 ( .A(n628), .B(KEYINPUT42), .ZN(n629) );
  BUF_X1 U709 ( .A(n632), .Z(n633) );
  INV_X1 U710 ( .A(n633), .ZN(n634) );
  INV_X1 U711 ( .A(n650), .ZN(n636) );
  AND2_X1 U712 ( .A1(n724), .A2(n636), .ZN(n639) );
  INV_X1 U713 ( .A(KEYINPUT75), .ZN(n640) );
  INV_X1 U714 ( .A(KEYINPUT47), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n640), .A2(n637), .ZN(n638) );
  NAND2_X1 U716 ( .A1(n639), .A2(n638), .ZN(n643) );
  INV_X1 U717 ( .A(n639), .ZN(n641) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n646), .A2(n645), .ZN(n661) );
  AND2_X1 U720 ( .A1(n647), .A2(n661), .ZN(n648) );
  XNOR2_X1 U721 ( .A(n648), .B(KEYINPUT36), .ZN(n649) );
  NAND2_X1 U722 ( .A1(n649), .A2(n663), .ZN(n734) );
  NAND2_X1 U723 ( .A1(n650), .A2(KEYINPUT47), .ZN(n651) );
  XOR2_X1 U724 ( .A(n651), .B(KEYINPUT85), .Z(n654) );
  NAND2_X1 U725 ( .A1(n724), .A2(n640), .ZN(n652) );
  NAND2_X1 U726 ( .A1(n652), .A2(KEYINPUT47), .ZN(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n655), .A2(n355), .ZN(n656) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n729) );
  INV_X1 U730 ( .A(KEYINPUT48), .ZN(n659) );
  NAND2_X1 U731 ( .A1(n661), .A2(n660), .ZN(n662) );
  OR2_X1 U732 ( .A1(n663), .A2(n662), .ZN(n664) );
  XNOR2_X1 U733 ( .A(n664), .B(KEYINPUT43), .ZN(n665) );
  NAND2_X1 U734 ( .A1(n665), .A2(n550), .ZN(n737) );
  AND2_X1 U735 ( .A1(n666), .A2(n725), .ZN(n736) );
  INV_X1 U736 ( .A(n736), .ZN(n667) );
  INV_X1 U737 ( .A(n778), .ZN(n669) );
  NAND2_X1 U738 ( .A1(n762), .A2(n669), .ZN(n670) );
  INV_X1 U739 ( .A(KEYINPUT2), .ZN(n672) );
  NAND2_X1 U740 ( .A1(n670), .A2(n672), .ZN(n671) );
  XNOR2_X1 U741 ( .A(n671), .B(KEYINPUT84), .ZN(n676) );
  INV_X1 U742 ( .A(KEYINPUT87), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n674), .B(n673), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(n762), .ZN(n704) );
  NAND2_X1 U745 ( .A1(n676), .A2(n704), .ZN(n680) );
  NAND2_X1 U746 ( .A1(n678), .A2(n677), .ZN(n679) );
  INV_X1 U747 ( .A(KEYINPUT53), .ZN(n682) );
  XNOR2_X1 U748 ( .A(n683), .B(n682), .ZN(G75) );
  NAND2_X1 U749 ( .A1(n720), .A2(n731), .ZN(n684) );
  XNOR2_X1 U750 ( .A(n684), .B(G104), .ZN(G6) );
  NAND2_X1 U751 ( .A1(n685), .A2(n731), .ZN(n686) );
  XNOR2_X1 U752 ( .A(n686), .B(G113), .ZN(G15) );
  NAND2_X1 U753 ( .A1(n685), .A2(n725), .ZN(n688) );
  XOR2_X1 U754 ( .A(G116), .B(KEYINPUT119), .Z(n687) );
  XNOR2_X1 U755 ( .A(n688), .B(n687), .ZN(G18) );
  XOR2_X1 U756 ( .A(G110), .B(KEYINPUT116), .Z(n689) );
  XNOR2_X1 U757 ( .A(n690), .B(n689), .ZN(G12) );
  XNOR2_X1 U758 ( .A(n691), .B(G101), .ZN(G3) );
  XOR2_X1 U759 ( .A(G137), .B(n692), .Z(G39) );
  XNOR2_X1 U760 ( .A(n693), .B(G119), .ZN(G21) );
  NOR2_X2 U761 ( .A1(n694), .A2(n699), .ZN(n697) );
  XNOR2_X1 U762 ( .A(n695), .B(KEYINPUT79), .ZN(n696) );
  NAND2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n703) );
  INV_X1 U764 ( .A(KEYINPUT86), .ZN(n698) );
  XNOR2_X1 U765 ( .A(n699), .B(n698), .ZN(n700) );
  AND2_X1 U766 ( .A1(n700), .A2(KEYINPUT2), .ZN(n701) );
  XNOR2_X1 U767 ( .A(n701), .B(KEYINPUT65), .ZN(n702) );
  NAND2_X1 U768 ( .A1(n746), .A2(G210), .ZN(n710) );
  BUF_X1 U769 ( .A(n706), .Z(n707) );
  XNOR2_X1 U770 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n708) );
  XNOR2_X1 U771 ( .A(n710), .B(n709), .ZN(n712) );
  INV_X1 U772 ( .A(G952), .ZN(n711) );
  NOR2_X2 U773 ( .A1(n712), .A2(n761), .ZN(n713) );
  XNOR2_X1 U774 ( .A(n713), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U775 ( .A1(n746), .A2(G472), .ZN(n716) );
  XNOR2_X1 U776 ( .A(n716), .B(n715), .ZN(n717) );
  NOR2_X2 U777 ( .A1(n717), .A2(n761), .ZN(n719) );
  XNOR2_X1 U778 ( .A(KEYINPUT115), .B(KEYINPUT63), .ZN(n718) );
  XNOR2_X1 U779 ( .A(n719), .B(n718), .ZN(G57) );
  NAND2_X1 U780 ( .A1(n720), .A2(n725), .ZN(n722) );
  XOR2_X1 U781 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n721) );
  XNOR2_X1 U782 ( .A(n722), .B(n721), .ZN(n723) );
  XNOR2_X1 U783 ( .A(G107), .B(n723), .ZN(G9) );
  XOR2_X1 U784 ( .A(KEYINPUT117), .B(KEYINPUT29), .Z(n727) );
  NAND2_X1 U785 ( .A1(n724), .A2(n725), .ZN(n726) );
  XNOR2_X1 U786 ( .A(n727), .B(n726), .ZN(n728) );
  XOR2_X1 U787 ( .A(G128), .B(n728), .Z(G30) );
  XOR2_X1 U788 ( .A(G143), .B(n729), .Z(n730) );
  XNOR2_X1 U789 ( .A(KEYINPUT118), .B(n730), .ZN(G45) );
  NAND2_X1 U790 ( .A1(n724), .A2(n731), .ZN(n732) );
  XNOR2_X1 U791 ( .A(n732), .B(G146), .ZN(G48) );
  XOR2_X1 U792 ( .A(KEYINPUT120), .B(KEYINPUT37), .Z(n733) );
  XNOR2_X1 U793 ( .A(n734), .B(n733), .ZN(n735) );
  XNOR2_X1 U794 ( .A(G125), .B(n735), .ZN(G27) );
  XOR2_X1 U795 ( .A(G134), .B(n736), .Z(G36) );
  XOR2_X1 U796 ( .A(G140), .B(n737), .Z(n738) );
  XNOR2_X1 U797 ( .A(n738), .B(KEYINPUT121), .ZN(G42) );
  NAND2_X1 U798 ( .A1(n756), .A2(G469), .ZN(n744) );
  XOR2_X1 U799 ( .A(KEYINPUT58), .B(KEYINPUT57), .Z(n740) );
  XNOR2_X1 U800 ( .A(KEYINPUT124), .B(KEYINPUT123), .ZN(n739) );
  XNOR2_X1 U801 ( .A(n740), .B(n739), .ZN(n741) );
  XOR2_X1 U802 ( .A(n742), .B(n741), .Z(n743) );
  XNOR2_X1 U803 ( .A(n744), .B(n743), .ZN(n745) );
  NOR2_X1 U804 ( .A1(n761), .A2(n745), .ZN(G54) );
  NAND2_X1 U805 ( .A1(n746), .A2(G475), .ZN(n749) );
  XNOR2_X1 U806 ( .A(n749), .B(n748), .ZN(n750) );
  NOR2_X2 U807 ( .A1(n750), .A2(n761), .ZN(n751) );
  XNOR2_X1 U808 ( .A(n751), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U809 ( .A1(n756), .A2(G478), .ZN(n754) );
  XOR2_X1 U810 ( .A(n752), .B(KEYINPUT125), .Z(n753) );
  XNOR2_X1 U811 ( .A(n754), .B(n753), .ZN(n755) );
  NOR2_X1 U812 ( .A1(n761), .A2(n755), .ZN(G63) );
  NAND2_X1 U813 ( .A1(n756), .A2(G217), .ZN(n759) );
  XNOR2_X1 U814 ( .A(n757), .B(KEYINPUT126), .ZN(n758) );
  XNOR2_X1 U815 ( .A(n759), .B(n758), .ZN(n760) );
  NOR2_X1 U816 ( .A1(n761), .A2(n760), .ZN(G66) );
  NAND2_X1 U817 ( .A1(n762), .A2(n779), .ZN(n766) );
  NAND2_X1 U818 ( .A1(n783), .A2(G224), .ZN(n763) );
  XNOR2_X1 U819 ( .A(KEYINPUT61), .B(n763), .ZN(n764) );
  NAND2_X1 U820 ( .A1(n764), .A2(G898), .ZN(n765) );
  NAND2_X1 U821 ( .A1(n766), .A2(n765), .ZN(n773) );
  XOR2_X1 U822 ( .A(G101), .B(n767), .Z(n768) );
  XNOR2_X1 U823 ( .A(n769), .B(n768), .ZN(n771) );
  NOR2_X1 U824 ( .A1(G898), .A2(n779), .ZN(n770) );
  NOR2_X1 U825 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U826 ( .A(n773), .B(n772), .ZN(G69) );
  XNOR2_X1 U827 ( .A(n775), .B(n774), .ZN(n777) );
  XNOR2_X1 U828 ( .A(n777), .B(n776), .ZN(n781) );
  XNOR2_X1 U829 ( .A(n778), .B(n781), .ZN(n780) );
  NAND2_X1 U830 ( .A1(n780), .A2(n779), .ZN(n786) );
  XNOR2_X1 U831 ( .A(G227), .B(n781), .ZN(n782) );
  NAND2_X1 U832 ( .A1(n782), .A2(G900), .ZN(n784) );
  NAND2_X1 U833 ( .A1(n784), .A2(n783), .ZN(n785) );
  NAND2_X1 U834 ( .A1(n786), .A2(n785), .ZN(G72) );
  XNOR2_X1 U835 ( .A(n787), .B(KEYINPUT127), .ZN(G33) );
  XOR2_X1 U836 ( .A(G122), .B(n375), .Z(G24) );
endmodule

