

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582;

  XNOR2_X1 U321 ( .A(n304), .B(n303), .ZN(n305) );
  XNOR2_X2 U322 ( .A(n306), .B(n305), .ZN(n555) );
  XNOR2_X1 U323 ( .A(n302), .B(n290), .ZN(n303) );
  XNOR2_X1 U324 ( .A(KEYINPUT64), .B(KEYINPUT41), .ZN(n394) );
  XOR2_X1 U325 ( .A(n343), .B(n296), .Z(n289) );
  XOR2_X1 U326 ( .A(n301), .B(n300), .Z(n290) );
  XNOR2_X1 U327 ( .A(KEYINPUT48), .B(KEYINPUT117), .ZN(n423) );
  XNOR2_X1 U328 ( .A(n388), .B(n387), .ZN(n389) );
  XNOR2_X1 U329 ( .A(n390), .B(n389), .ZN(n393) );
  NOR2_X1 U330 ( .A1(n464), .A2(n566), .ZN(n447) );
  XNOR2_X1 U331 ( .A(n572), .B(n394), .ZN(n534) );
  XOR2_X1 U332 ( .A(KEYINPUT94), .B(n462), .Z(n547) );
  XNOR2_X1 U333 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n449) );
  XNOR2_X1 U334 ( .A(n450), .B(n449), .ZN(G1351GAT) );
  XNOR2_X1 U335 ( .A(G43GAT), .B(KEYINPUT8), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n291), .B(KEYINPUT7), .ZN(n370) );
  XOR2_X1 U337 ( .A(G92GAT), .B(KEYINPUT75), .Z(n293) );
  XNOR2_X1 U338 ( .A(G99GAT), .B(G106GAT), .ZN(n292) );
  XNOR2_X1 U339 ( .A(n293), .B(n292), .ZN(n384) );
  XNOR2_X1 U340 ( .A(n370), .B(n384), .ZN(n306) );
  XOR2_X1 U341 ( .A(G50GAT), .B(G162GAT), .Z(n343) );
  XOR2_X1 U342 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n295) );
  XNOR2_X1 U343 ( .A(KEYINPUT11), .B(KEYINPUT9), .ZN(n294) );
  XNOR2_X1 U344 ( .A(n295), .B(n294), .ZN(n296) );
  NAND2_X1 U345 ( .A1(G232GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n289), .B(n297), .ZN(n304) );
  XNOR2_X1 U347 ( .A(G36GAT), .B(G190GAT), .ZN(n298) );
  XNOR2_X1 U348 ( .A(n298), .B(G218GAT), .ZN(n347) );
  XNOR2_X1 U349 ( .A(G29GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U350 ( .A(n299), .B(G85GAT), .ZN(n435) );
  XNOR2_X1 U351 ( .A(n347), .B(n435), .ZN(n302) );
  XOR2_X1 U352 ( .A(KEYINPUT76), .B(KEYINPUT66), .Z(n301) );
  XNOR2_X1 U353 ( .A(KEYINPUT65), .B(KEYINPUT77), .ZN(n300) );
  XNOR2_X1 U354 ( .A(KEYINPUT78), .B(n555), .ZN(n540) );
  XOR2_X1 U355 ( .A(G176GAT), .B(KEYINPUT20), .Z(n308) );
  XNOR2_X1 U356 ( .A(G43GAT), .B(G99GAT), .ZN(n307) );
  XNOR2_X1 U357 ( .A(n308), .B(n307), .ZN(n318) );
  XOR2_X1 U358 ( .A(G120GAT), .B(KEYINPUT82), .Z(n310) );
  XNOR2_X1 U359 ( .A(G15GAT), .B(G71GAT), .ZN(n309) );
  XNOR2_X1 U360 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U361 ( .A(G134GAT), .B(G190GAT), .Z(n312) );
  XOR2_X1 U362 ( .A(KEYINPUT0), .B(G127GAT), .Z(n436) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(n436), .ZN(n311) );
  XNOR2_X1 U364 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U365 ( .A(n314), .B(n313), .Z(n316) );
  NAND2_X1 U366 ( .A1(G227GAT), .A2(G233GAT), .ZN(n315) );
  XNOR2_X1 U367 ( .A(n316), .B(n315), .ZN(n317) );
  XNOR2_X1 U368 ( .A(n318), .B(n317), .ZN(n323) );
  XOR2_X1 U369 ( .A(KEYINPUT81), .B(G183GAT), .Z(n320) );
  XNOR2_X1 U370 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n319) );
  XNOR2_X1 U371 ( .A(n320), .B(n319), .ZN(n322) );
  XOR2_X1 U372 ( .A(KEYINPUT19), .B(KEYINPUT17), .Z(n321) );
  XOR2_X1 U373 ( .A(n322), .B(n321), .Z(n351) );
  XNOR2_X1 U374 ( .A(n323), .B(n351), .ZN(n467) );
  INV_X1 U375 ( .A(n467), .ZN(n529) );
  XOR2_X1 U376 ( .A(KEYINPUT86), .B(G211GAT), .Z(n325) );
  XNOR2_X1 U377 ( .A(KEYINPUT21), .B(G204GAT), .ZN(n324) );
  XNOR2_X1 U378 ( .A(n325), .B(n324), .ZN(n326) );
  XOR2_X1 U379 ( .A(G197GAT), .B(n326), .Z(n352) );
  XOR2_X1 U380 ( .A(KEYINPUT84), .B(KEYINPUT89), .Z(n328) );
  XNOR2_X1 U381 ( .A(KEYINPUT22), .B(KEYINPUT23), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n329) );
  XOR2_X1 U383 ( .A(G22GAT), .B(n329), .Z(n331) );
  NAND2_X1 U384 ( .A1(G228GAT), .A2(G233GAT), .ZN(n330) );
  XNOR2_X1 U385 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U386 ( .A(n332), .B(KEYINPUT85), .Z(n338) );
  XNOR2_X1 U387 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n333) );
  XNOR2_X1 U388 ( .A(n333), .B(KEYINPUT87), .ZN(n334) );
  XOR2_X1 U389 ( .A(n334), .B(KEYINPUT3), .Z(n336) );
  XNOR2_X1 U390 ( .A(G141GAT), .B(G148GAT), .ZN(n335) );
  XNOR2_X1 U391 ( .A(n336), .B(n335), .ZN(n443) );
  XNOR2_X1 U392 ( .A(n443), .B(KEYINPUT24), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT88), .B(KEYINPUT83), .Z(n340) );
  XNOR2_X1 U395 ( .A(G218GAT), .B(G106GAT), .ZN(n339) );
  XNOR2_X1 U396 ( .A(n340), .B(n339), .ZN(n341) );
  XOR2_X1 U397 ( .A(n342), .B(n341), .Z(n345) );
  XOR2_X1 U398 ( .A(KEYINPUT74), .B(G78GAT), .Z(n376) );
  XNOR2_X1 U399 ( .A(n343), .B(n376), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U401 ( .A(n352), .B(n346), .ZN(n464) );
  XOR2_X1 U402 ( .A(n347), .B(KEYINPUT95), .Z(n349) );
  NAND2_X1 U403 ( .A1(G226GAT), .A2(G233GAT), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U405 ( .A(n351), .B(n350), .ZN(n356) );
  XOR2_X1 U406 ( .A(G176GAT), .B(G64GAT), .Z(n391) );
  XOR2_X1 U407 ( .A(n391), .B(G92GAT), .Z(n354) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(n352), .ZN(n353) );
  XNOR2_X1 U409 ( .A(n354), .B(n353), .ZN(n355) );
  XNOR2_X1 U410 ( .A(n356), .B(n355), .ZN(n474) );
  XOR2_X1 U411 ( .A(KEYINPUT71), .B(KEYINPUT70), .Z(n358) );
  XNOR2_X1 U412 ( .A(KEYINPUT69), .B(KEYINPUT72), .ZN(n357) );
  XNOR2_X1 U413 ( .A(n358), .B(n357), .ZN(n365) );
  XOR2_X1 U414 ( .A(G141GAT), .B(G197GAT), .Z(n360) );
  XNOR2_X1 U415 ( .A(G50GAT), .B(G36GAT), .ZN(n359) );
  XNOR2_X1 U416 ( .A(n360), .B(n359), .ZN(n361) );
  XOR2_X1 U417 ( .A(n361), .B(G29GAT), .Z(n363) );
  XOR2_X1 U418 ( .A(G113GAT), .B(G1GAT), .Z(n430) );
  XNOR2_X1 U419 ( .A(G169GAT), .B(n430), .ZN(n362) );
  XNOR2_X1 U420 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U421 ( .A(n365), .B(n364), .ZN(n374) );
  XOR2_X1 U422 ( .A(KEYINPUT68), .B(KEYINPUT30), .Z(n367) );
  NAND2_X1 U423 ( .A1(G229GAT), .A2(G233GAT), .ZN(n366) );
  XNOR2_X1 U424 ( .A(n367), .B(n366), .ZN(n368) );
  XOR2_X1 U425 ( .A(n368), .B(KEYINPUT29), .Z(n372) );
  XNOR2_X1 U426 ( .A(G15GAT), .B(G22GAT), .ZN(n369) );
  XNOR2_X1 U427 ( .A(n369), .B(G8GAT), .ZN(n405) );
  XNOR2_X1 U428 ( .A(n370), .B(n405), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U430 ( .A(n374), .B(n373), .ZN(n502) );
  XNOR2_X1 U431 ( .A(G71GAT), .B(KEYINPUT73), .ZN(n375) );
  XNOR2_X1 U432 ( .A(n375), .B(KEYINPUT13), .ZN(n402) );
  XNOR2_X1 U433 ( .A(n402), .B(n376), .ZN(n380) );
  INV_X1 U434 ( .A(n380), .ZN(n378) );
  AND2_X1 U435 ( .A1(G230GAT), .A2(G233GAT), .ZN(n379) );
  INV_X1 U436 ( .A(n379), .ZN(n377) );
  NAND2_X1 U437 ( .A1(n378), .A2(n377), .ZN(n382) );
  NAND2_X1 U438 ( .A1(n380), .A2(n379), .ZN(n381) );
  NAND2_X1 U439 ( .A1(n382), .A2(n381), .ZN(n383) );
  XOR2_X1 U440 ( .A(n383), .B(KEYINPUT31), .Z(n390) );
  XNOR2_X1 U441 ( .A(n384), .B(KEYINPUT33), .ZN(n388) );
  XOR2_X1 U442 ( .A(KEYINPUT32), .B(G85GAT), .Z(n386) );
  XNOR2_X1 U443 ( .A(G204GAT), .B(G148GAT), .ZN(n385) );
  XNOR2_X1 U444 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U445 ( .A(G120GAT), .B(G57GAT), .Z(n433) );
  XOR2_X1 U446 ( .A(n391), .B(n433), .Z(n392) );
  XNOR2_X1 U447 ( .A(n393), .B(n392), .ZN(n572) );
  NOR2_X1 U448 ( .A1(n502), .A2(n534), .ZN(n395) );
  XNOR2_X1 U449 ( .A(n395), .B(KEYINPUT46), .ZN(n413) );
  XOR2_X1 U450 ( .A(G64GAT), .B(KEYINPUT14), .Z(n397) );
  XNOR2_X1 U451 ( .A(G1GAT), .B(G155GAT), .ZN(n396) );
  XNOR2_X1 U452 ( .A(n397), .B(n396), .ZN(n401) );
  XOR2_X1 U453 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n399) );
  XNOR2_X1 U454 ( .A(KEYINPUT12), .B(KEYINPUT15), .ZN(n398) );
  XNOR2_X1 U455 ( .A(n399), .B(n398), .ZN(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n412) );
  XOR2_X1 U457 ( .A(n402), .B(G78GAT), .Z(n404) );
  XNOR2_X1 U458 ( .A(G183GAT), .B(G127GAT), .ZN(n403) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n410) );
  XOR2_X1 U460 ( .A(n405), .B(G57GAT), .Z(n407) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U462 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U463 ( .A(G211GAT), .B(n408), .Z(n409) );
  XNOR2_X1 U464 ( .A(n410), .B(n409), .ZN(n411) );
  XNOR2_X1 U465 ( .A(n412), .B(n411), .ZN(n576) );
  NOR2_X1 U466 ( .A1(n413), .A2(n576), .ZN(n414) );
  XNOR2_X1 U467 ( .A(n414), .B(KEYINPUT115), .ZN(n415) );
  NOR2_X1 U468 ( .A1(n415), .A2(n555), .ZN(n416) );
  XNOR2_X1 U469 ( .A(n416), .B(KEYINPUT47), .ZN(n422) );
  INV_X1 U470 ( .A(n576), .ZN(n484) );
  XOR2_X1 U471 ( .A(KEYINPUT36), .B(n540), .Z(n579) );
  NOR2_X1 U472 ( .A1(n484), .A2(n579), .ZN(n417) );
  XNOR2_X1 U473 ( .A(n417), .B(KEYINPUT45), .ZN(n418) );
  NAND2_X1 U474 ( .A1(n418), .A2(n502), .ZN(n419) );
  NOR2_X1 U475 ( .A1(n572), .A2(n419), .ZN(n420) );
  XOR2_X1 U476 ( .A(KEYINPUT116), .B(n420), .Z(n421) );
  AND2_X1 U477 ( .A1(n422), .A2(n421), .ZN(n424) );
  XNOR2_X1 U478 ( .A(n424), .B(n423), .ZN(n530) );
  NAND2_X1 U479 ( .A1(n474), .A2(n530), .ZN(n425) );
  XNOR2_X1 U480 ( .A(n425), .B(KEYINPUT54), .ZN(n426) );
  XNOR2_X1 U481 ( .A(n426), .B(KEYINPUT123), .ZN(n446) );
  XOR2_X1 U482 ( .A(KEYINPUT1), .B(KEYINPUT93), .Z(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT90), .B(KEYINPUT4), .ZN(n427) );
  XNOR2_X1 U484 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U485 ( .A(n429), .B(KEYINPUT6), .Z(n432) );
  XNOR2_X1 U486 ( .A(n430), .B(G162GAT), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n434) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U490 ( .A(n438), .B(n437), .ZN(n442) );
  XOR2_X1 U491 ( .A(KEYINPUT91), .B(KEYINPUT5), .Z(n440) );
  NAND2_X1 U492 ( .A1(G225GAT), .A2(G233GAT), .ZN(n439) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XOR2_X1 U494 ( .A(n442), .B(n441), .Z(n445) );
  XNOR2_X1 U495 ( .A(n443), .B(KEYINPUT92), .ZN(n444) );
  XNOR2_X1 U496 ( .A(n445), .B(n444), .ZN(n462) );
  NAND2_X1 U497 ( .A1(n446), .A2(n547), .ZN(n566) );
  XNOR2_X1 U498 ( .A(n447), .B(KEYINPUT55), .ZN(n448) );
  NOR2_X2 U499 ( .A1(n529), .A2(n448), .ZN(n560) );
  NAND2_X1 U500 ( .A1(n540), .A2(n560), .ZN(n450) );
  NAND2_X1 U501 ( .A1(n576), .A2(n560), .ZN(n452) );
  XNOR2_X1 U502 ( .A(KEYINPUT124), .B(G183GAT), .ZN(n451) );
  XNOR2_X1 U503 ( .A(n452), .B(n451), .ZN(G1350GAT) );
  NOR2_X1 U504 ( .A1(n502), .A2(n572), .ZN(n489) );
  XOR2_X1 U505 ( .A(KEYINPUT26), .B(KEYINPUT97), .Z(n454) );
  NAND2_X1 U506 ( .A1(n464), .A2(n529), .ZN(n453) );
  XNOR2_X1 U507 ( .A(n454), .B(n453), .ZN(n567) );
  XOR2_X1 U508 ( .A(n474), .B(KEYINPUT96), .Z(n455) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n455), .ZN(n463) );
  NOR2_X1 U510 ( .A1(n567), .A2(n463), .ZN(n545) );
  NAND2_X1 U511 ( .A1(n467), .A2(n474), .ZN(n456) );
  XOR2_X1 U512 ( .A(KEYINPUT98), .B(n456), .Z(n457) );
  NOR2_X1 U513 ( .A1(n464), .A2(n457), .ZN(n458) );
  XOR2_X1 U514 ( .A(KEYINPUT25), .B(n458), .Z(n459) );
  NOR2_X1 U515 ( .A1(n545), .A2(n459), .ZN(n460) );
  XOR2_X1 U516 ( .A(KEYINPUT99), .B(n460), .Z(n461) );
  NOR2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n469) );
  INV_X1 U518 ( .A(n463), .ZN(n466) );
  XNOR2_X1 U519 ( .A(KEYINPUT28), .B(n464), .ZN(n479) );
  NOR2_X1 U520 ( .A1(n547), .A2(n479), .ZN(n465) );
  NAND2_X1 U521 ( .A1(n466), .A2(n465), .ZN(n528) );
  NOR2_X1 U522 ( .A1(n467), .A2(n528), .ZN(n468) );
  NOR2_X1 U523 ( .A1(n469), .A2(n468), .ZN(n483) );
  NOR2_X1 U524 ( .A1(n484), .A2(n540), .ZN(n470) );
  XOR2_X1 U525 ( .A(KEYINPUT16), .B(n470), .Z(n471) );
  NOR2_X1 U526 ( .A1(n483), .A2(n471), .ZN(n503) );
  NAND2_X1 U527 ( .A1(n489), .A2(n503), .ZN(n480) );
  NOR2_X1 U528 ( .A1(n547), .A2(n480), .ZN(n472) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(n472), .Z(n473) );
  XNOR2_X1 U530 ( .A(G1GAT), .B(n473), .ZN(G1324GAT) );
  INV_X1 U531 ( .A(n474), .ZN(n518) );
  NOR2_X1 U532 ( .A1(n518), .A2(n480), .ZN(n475) );
  XOR2_X1 U533 ( .A(KEYINPUT100), .B(n475), .Z(n476) );
  XNOR2_X1 U534 ( .A(G8GAT), .B(n476), .ZN(G1325GAT) );
  NOR2_X1 U535 ( .A1(n529), .A2(n480), .ZN(n478) );
  XNOR2_X1 U536 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n477) );
  XNOR2_X1 U537 ( .A(n478), .B(n477), .ZN(G1326GAT) );
  INV_X1 U538 ( .A(n479), .ZN(n524) );
  NOR2_X1 U539 ( .A1(n524), .A2(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G22GAT), .B(KEYINPUT101), .ZN(n481) );
  XNOR2_X1 U541 ( .A(n482), .B(n481), .ZN(G1327GAT) );
  XNOR2_X1 U542 ( .A(KEYINPUT102), .B(KEYINPUT39), .ZN(n493) );
  XOR2_X1 U543 ( .A(KEYINPUT105), .B(KEYINPUT38), .Z(n491) );
  NOR2_X1 U544 ( .A1(n483), .A2(n579), .ZN(n485) );
  NAND2_X1 U545 ( .A1(n485), .A2(n484), .ZN(n488) );
  XOR2_X1 U546 ( .A(KEYINPUT104), .B(KEYINPUT37), .Z(n486) );
  XNOR2_X1 U547 ( .A(KEYINPUT103), .B(n486), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(n514) );
  NAND2_X1 U549 ( .A1(n489), .A2(n514), .ZN(n490) );
  XNOR2_X1 U550 ( .A(n491), .B(n490), .ZN(n498) );
  NOR2_X1 U551 ( .A1(n547), .A2(n498), .ZN(n492) );
  XNOR2_X1 U552 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U553 ( .A(G29GAT), .B(n494), .ZN(G1328GAT) );
  NOR2_X1 U554 ( .A1(n498), .A2(n518), .ZN(n495) );
  XOR2_X1 U555 ( .A(G36GAT), .B(n495), .Z(G1329GAT) );
  NOR2_X1 U556 ( .A1(n498), .A2(n529), .ZN(n496) );
  XOR2_X1 U557 ( .A(KEYINPUT40), .B(n496), .Z(n497) );
  XNOR2_X1 U558 ( .A(G43GAT), .B(n497), .ZN(G1330GAT) );
  NOR2_X1 U559 ( .A1(n498), .A2(n524), .ZN(n499) );
  XOR2_X1 U560 ( .A(G50GAT), .B(n499), .Z(G1331GAT) );
  XOR2_X1 U561 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n501) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT107), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n501), .B(n500), .ZN(n505) );
  INV_X1 U564 ( .A(n502), .ZN(n569) );
  NOR2_X1 U565 ( .A1(n534), .A2(n569), .ZN(n515) );
  NAND2_X1 U566 ( .A1(n515), .A2(n503), .ZN(n508) );
  NOR2_X1 U567 ( .A1(n547), .A2(n508), .ZN(n504) );
  XOR2_X1 U568 ( .A(n505), .B(n504), .Z(G1332GAT) );
  NOR2_X1 U569 ( .A1(n518), .A2(n508), .ZN(n506) );
  XOR2_X1 U570 ( .A(G64GAT), .B(n506), .Z(G1333GAT) );
  NOR2_X1 U571 ( .A1(n529), .A2(n508), .ZN(n507) );
  XOR2_X1 U572 ( .A(G71GAT), .B(n507), .Z(G1334GAT) );
  NOR2_X1 U573 ( .A1(n524), .A2(n508), .ZN(n513) );
  XOR2_X1 U574 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n510) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n509) );
  XNOR2_X1 U576 ( .A(n510), .B(n509), .ZN(n511) );
  XNOR2_X1 U577 ( .A(KEYINPUT108), .B(n511), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1335GAT) );
  NAND2_X1 U579 ( .A1(n515), .A2(n514), .ZN(n523) );
  NOR2_X1 U580 ( .A1(n547), .A2(n523), .ZN(n517) );
  XNOR2_X1 U581 ( .A(G85GAT), .B(KEYINPUT111), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(G1336GAT) );
  NOR2_X1 U583 ( .A1(n518), .A2(n523), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT112), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G92GAT), .B(n520), .ZN(G1337GAT) );
  NOR2_X1 U586 ( .A1(n529), .A2(n523), .ZN(n522) );
  XNOR2_X1 U587 ( .A(G99GAT), .B(KEYINPUT113), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n522), .B(n521), .ZN(G1338GAT) );
  NOR2_X1 U589 ( .A1(n524), .A2(n523), .ZN(n526) );
  XNOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT114), .ZN(n525) );
  XNOR2_X1 U591 ( .A(n526), .B(n525), .ZN(n527) );
  XOR2_X1 U592 ( .A(G106GAT), .B(n527), .Z(G1339GAT) );
  NOR2_X1 U593 ( .A1(n529), .A2(n528), .ZN(n531) );
  NAND2_X1 U594 ( .A1(n531), .A2(n530), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT118), .B(n532), .Z(n541) );
  NAND2_X1 U596 ( .A1(n541), .A2(n569), .ZN(n533) );
  XNOR2_X1 U597 ( .A(n533), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U598 ( .A(G120GAT), .B(KEYINPUT49), .Z(n536) );
  INV_X1 U599 ( .A(n534), .ZN(n559) );
  NAND2_X1 U600 ( .A1(n541), .A2(n559), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n536), .B(n535), .ZN(G1341GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT50), .B(KEYINPUT119), .Z(n538) );
  NAND2_X1 U603 ( .A1(n541), .A2(n576), .ZN(n537) );
  XNOR2_X1 U604 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(G127GAT), .B(n539), .ZN(G1342GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT120), .B(KEYINPUT51), .Z(n543) );
  NAND2_X1 U607 ( .A1(n541), .A2(n540), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G134GAT), .B(n544), .ZN(G1343GAT) );
  NAND2_X1 U610 ( .A1(n530), .A2(n545), .ZN(n546) );
  NOR2_X1 U611 ( .A1(n547), .A2(n546), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n569), .A2(n556), .ZN(n548) );
  XNOR2_X1 U613 ( .A(n548), .B(G141GAT), .ZN(G1344GAT) );
  XOR2_X1 U614 ( .A(KEYINPUT52), .B(KEYINPUT121), .Z(n550) );
  NAND2_X1 U615 ( .A1(n556), .A2(n559), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n550), .B(n549), .ZN(n552) );
  XOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT53), .Z(n551) );
  XNOR2_X1 U618 ( .A(n552), .B(n551), .ZN(G1345GAT) );
  NAND2_X1 U619 ( .A1(n576), .A2(n556), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n553), .B(KEYINPUT122), .ZN(n554) );
  XNOR2_X1 U621 ( .A(G155GAT), .B(n554), .ZN(G1346GAT) );
  NAND2_X1 U622 ( .A1(n556), .A2(n555), .ZN(n557) );
  XNOR2_X1 U623 ( .A(n557), .B(G162GAT), .ZN(G1347GAT) );
  NAND2_X1 U624 ( .A1(n569), .A2(n560), .ZN(n558) );
  XNOR2_X1 U625 ( .A(n558), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U626 ( .A1(n560), .A2(n559), .ZN(n562) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n561) );
  XNOR2_X1 U628 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U629 ( .A(G176GAT), .B(n563), .ZN(G1349GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n565) );
  XNOR2_X1 U631 ( .A(G197GAT), .B(KEYINPUT125), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n571) );
  NOR2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n568) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n570) );
  XOR2_X1 U635 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U636 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n574) );
  NAND2_X1 U637 ( .A1(n568), .A2(n572), .ZN(n573) );
  XNOR2_X1 U638 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U639 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  NAND2_X1 U640 ( .A1(n576), .A2(n568), .ZN(n577) );
  XNOR2_X1 U641 ( .A(n577), .B(G211GAT), .ZN(G1354GAT) );
  INV_X1 U642 ( .A(n568), .ZN(n578) );
  NOR2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n581) );
  XNOR2_X1 U644 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n581), .B(n580), .ZN(n582) );
  XNOR2_X1 U646 ( .A(G218GAT), .B(n582), .ZN(G1355GAT) );
endmodule

