//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 0 0 1 0 0 0 0 1 0 1 1 1 1 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:31 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n444, new_n448, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n530, new_n531, new_n532, new_n533, new_n535,
    new_n536, new_n537, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n545, new_n546, new_n548, new_n549, new_n550, new_n551, new_n552,
    new_n553, new_n554, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n567, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n590, new_n593, new_n594, new_n596, new_n597, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT66), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT67), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n442));
  XOR2_X1   g017(.A(new_n442), .B(KEYINPUT68), .Z(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(new_n444));
  XNOR2_X1  g019(.A(new_n444), .B(KEYINPUT69), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(G261));
  INV_X1    g030(.A(G261), .ZN(G325));
  INV_X1    g031(.A(G2106), .ZN(new_n457));
  INV_X1    g032(.A(G567), .ZN(new_n458));
  OAI22_X1  g033(.A1(new_n453), .A2(new_n457), .B1(new_n458), .B2(new_n454), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G125), .ZN(new_n463));
  NAND2_X1  g038(.A1(G113), .A2(G2104), .ZN(new_n464));
  INV_X1    g039(.A(KEYINPUT70), .ZN(new_n465));
  XNOR2_X1  g040(.A(new_n464), .B(new_n465), .ZN(new_n466));
  AOI21_X1  g041(.A(new_n461), .B1(new_n463), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n461), .A2(G2104), .ZN(new_n468));
  INV_X1    g043(.A(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(G101), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n462), .A2(new_n461), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n470), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(new_n473), .ZN(G160));
  OAI21_X1  g049(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n475));
  INV_X1    g050(.A(G112), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n475), .B1(new_n476), .B2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n471), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G136), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g057(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n483));
  AOI21_X1  g058(.A(new_n461), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  XOR2_X1   g059(.A(new_n484), .B(KEYINPUT71), .Z(new_n485));
  AOI211_X1 g060(.A(new_n477), .B(new_n480), .C1(new_n485), .C2(G124), .ZN(G162));
  AND2_X1   g061(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n487));
  OAI211_X1 g062(.A(G126), .B(G2105), .C1(new_n487), .C2(new_n481), .ZN(new_n488));
  INV_X1    g063(.A(G114), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n490), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n494), .B(new_n496), .C1(new_n481), .C2(new_n487), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n494), .B1(new_n487), .B2(new_n481), .ZN(new_n498));
  INV_X1    g073(.A(new_n496), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(new_n492), .B1(new_n497), .B2(new_n500), .ZN(G164));
  INV_X1    g076(.A(G543), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  OAI21_X1  g078(.A(new_n502), .B1(new_n503), .B2(KEYINPUT73), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT73), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .A3(G543), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  AOI22_X1  g082(.A1(new_n507), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n508));
  INV_X1    g083(.A(G651), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g085(.A(KEYINPUT6), .B(G651), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(new_n511), .ZN(new_n512));
  INV_X1    g087(.A(G88), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n511), .A2(G543), .ZN(new_n514));
  INV_X1    g089(.A(G50), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  OR2_X1    g091(.A1(new_n510), .A2(new_n516), .ZN(G303));
  INV_X1    g092(.A(G303), .ZN(G166));
  INV_X1    g093(.A(G51), .ZN(new_n519));
  INV_X1    g094(.A(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n514), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g096(.A1(new_n511), .A2(KEYINPUT74), .A3(G543), .ZN(new_n522));
  AOI21_X1  g097(.A(new_n519), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g098(.A1(new_n507), .A2(G63), .A3(G651), .ZN(new_n524));
  NAND3_X1  g099(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n525));
  XNOR2_X1  g100(.A(new_n525), .B(KEYINPUT7), .ZN(new_n526));
  INV_X1    g101(.A(G89), .ZN(new_n527));
  OAI211_X1 g102(.A(new_n524), .B(new_n526), .C1(new_n512), .C2(new_n527), .ZN(new_n528));
  NOR2_X1   g103(.A1(new_n523), .A2(new_n528), .ZN(G168));
  AOI22_X1  g104(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n530));
  INV_X1    g105(.A(G90), .ZN(new_n531));
  OAI22_X1  g106(.A1(new_n530), .A2(new_n509), .B1(new_n531), .B2(new_n512), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n521), .A2(new_n522), .ZN(new_n533));
  AOI21_X1  g108(.A(new_n532), .B1(G52), .B2(new_n533), .ZN(G171));
  NAND2_X1  g109(.A1(new_n533), .A2(G43), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n509), .ZN(new_n537));
  INV_X1    g112(.A(new_n512), .ZN(new_n538));
  XOR2_X1   g113(.A(KEYINPUT75), .B(G81), .Z(new_n539));
  NAND2_X1  g114(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  NAND3_X1  g115(.A1(new_n535), .A2(new_n537), .A3(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  NAND4_X1  g118(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g119(.A1(G1), .A2(G3), .ZN(new_n545));
  XNOR2_X1  g120(.A(new_n545), .B(KEYINPUT8), .ZN(new_n546));
  NAND4_X1  g121(.A1(G319), .A2(G483), .A3(G661), .A4(new_n546), .ZN(G188));
  NAND2_X1  g122(.A1(G78), .A2(G543), .ZN(new_n548));
  INV_X1    g123(.A(new_n507), .ZN(new_n549));
  INV_X1    g124(.A(G65), .ZN(new_n550));
  OAI21_X1  g125(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  AOI22_X1  g126(.A1(new_n551), .A2(G651), .B1(new_n538), .B2(G91), .ZN(new_n552));
  NAND3_X1  g127(.A1(new_n511), .A2(G53), .A3(G543), .ZN(new_n553));
  XNOR2_X1  g128(.A(new_n553), .B(KEYINPUT9), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n552), .A2(new_n554), .ZN(G299));
  INV_X1    g130(.A(G171), .ZN(G301));
  INV_X1    g131(.A(G168), .ZN(G286));
  OAI21_X1  g132(.A(G651), .B1(new_n507), .B2(G74), .ZN(new_n558));
  NAND3_X1  g133(.A1(new_n507), .A2(G87), .A3(new_n511), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n511), .A2(G49), .A3(G543), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n558), .A2(new_n559), .A3(new_n560), .ZN(G288));
  INV_X1    g136(.A(new_n514), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n538), .A2(G86), .B1(new_n562), .B2(G48), .ZN(new_n563));
  AND2_X1   g138(.A1(new_n507), .A2(G61), .ZN(new_n564));
  NAND2_X1  g139(.A1(G73), .A2(G543), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT76), .Z(new_n566));
  OAI21_X1  g141(.A(G651), .B1(new_n564), .B2(new_n566), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G305));
  AOI22_X1  g143(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n569));
  XOR2_X1   g144(.A(KEYINPUT78), .B(G85), .Z(new_n570));
  OAI22_X1  g145(.A1(new_n569), .A2(new_n509), .B1(new_n512), .B2(new_n570), .ZN(new_n571));
  XOR2_X1   g146(.A(KEYINPUT77), .B(G47), .Z(new_n572));
  AOI21_X1  g147(.A(new_n572), .B1(new_n521), .B2(new_n522), .ZN(new_n573));
  NOR2_X1   g148(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(new_n574), .ZN(G290));
  NAND2_X1  g150(.A1(G79), .A2(G543), .ZN(new_n576));
  INV_X1    g151(.A(G66), .ZN(new_n577));
  OAI21_X1  g152(.A(new_n576), .B1(new_n549), .B2(new_n577), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n533), .A2(G54), .B1(new_n578), .B2(G651), .ZN(new_n579));
  NAND3_X1  g154(.A1(new_n538), .A2(KEYINPUT10), .A3(G92), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT10), .ZN(new_n581));
  INV_X1    g156(.A(G92), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n581), .B1(new_n512), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n579), .A2(new_n584), .ZN(new_n585));
  INV_X1    g160(.A(G868), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g162(.A(new_n587), .B1(new_n586), .B2(G171), .ZN(G284));
  OAI21_X1  g163(.A(new_n587), .B1(new_n586), .B2(G171), .ZN(G321));
  NAND2_X1  g164(.A1(G299), .A2(new_n586), .ZN(new_n590));
  OAI21_X1  g165(.A(new_n590), .B1(new_n586), .B2(G168), .ZN(G297));
  XNOR2_X1  g166(.A(G297), .B(KEYINPUT79), .ZN(G280));
  INV_X1    g167(.A(new_n585), .ZN(new_n593));
  INV_X1    g168(.A(G559), .ZN(new_n594));
  OAI21_X1  g169(.A(new_n593), .B1(new_n594), .B2(G860), .ZN(G148));
  NAND2_X1  g170(.A1(new_n541), .A2(new_n586), .ZN(new_n596));
  NOR2_X1   g171(.A1(new_n585), .A2(G559), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n596), .B1(new_n597), .B2(new_n586), .ZN(G323));
  XNOR2_X1  g173(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g174(.A1(new_n462), .A2(new_n469), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT12), .ZN(new_n601));
  XNOR2_X1  g176(.A(new_n601), .B(KEYINPUT13), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n478), .A2(G135), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n461), .A2(G111), .ZN(new_n605));
  OAI21_X1  g180(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n606));
  XNOR2_X1  g181(.A(new_n484), .B(KEYINPUT71), .ZN(new_n607));
  INV_X1    g182(.A(G123), .ZN(new_n608));
  OAI221_X1 g183(.A(new_n604), .B1(new_n605), .B2(new_n606), .C1(new_n607), .C2(new_n608), .ZN(new_n609));
  AOI22_X1  g184(.A1(new_n603), .A2(G2100), .B1(G2096), .B2(new_n609), .ZN(new_n610));
  OR2_X1    g185(.A1(new_n609), .A2(G2096), .ZN(new_n611));
  OAI211_X1 g186(.A(new_n610), .B(new_n611), .C1(G2100), .C2(new_n603), .ZN(G156));
  XOR2_X1   g187(.A(G2451), .B(G2454), .Z(new_n613));
  XNOR2_X1  g188(.A(new_n613), .B(KEYINPUT16), .ZN(new_n614));
  XNOR2_X1  g189(.A(G1341), .B(G1348), .ZN(new_n615));
  XNOR2_X1  g190(.A(new_n614), .B(new_n615), .ZN(new_n616));
  INV_X1    g191(.A(KEYINPUT14), .ZN(new_n617));
  XNOR2_X1  g192(.A(G2427), .B(G2438), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(G2430), .ZN(new_n619));
  XNOR2_X1  g194(.A(KEYINPUT15), .B(G2435), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n621), .B1(new_n620), .B2(new_n619), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n616), .B(new_n622), .ZN(new_n623));
  XNOR2_X1  g198(.A(G2443), .B(G2446), .ZN(new_n624));
  INV_X1    g199(.A(new_n624), .ZN(new_n625));
  OR2_X1    g200(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n623), .A2(new_n625), .ZN(new_n627));
  NAND3_X1  g202(.A1(new_n626), .A2(G14), .A3(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(new_n628), .ZN(G401));
  XOR2_X1   g204(.A(G2084), .B(G2090), .Z(new_n630));
  XNOR2_X1  g205(.A(G2067), .B(G2678), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2072), .B(G2078), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  XOR2_X1   g208(.A(new_n633), .B(KEYINPUT18), .Z(new_n634));
  INV_X1    g209(.A(new_n631), .ZN(new_n635));
  INV_X1    g210(.A(new_n632), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n630), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(KEYINPUT80), .B(KEYINPUT17), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n638), .B(new_n632), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n637), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  NAND3_X1  g215(.A1(new_n639), .A2(new_n635), .A3(new_n630), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n634), .A2(new_n640), .A3(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(KEYINPUT81), .ZN(new_n643));
  XOR2_X1   g218(.A(G2096), .B(G2100), .Z(new_n644));
  XNOR2_X1  g219(.A(new_n643), .B(new_n644), .ZN(G227));
  XOR2_X1   g220(.A(G1971), .B(G1976), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT19), .ZN(new_n647));
  XOR2_X1   g222(.A(G1956), .B(G2474), .Z(new_n648));
  XOR2_X1   g223(.A(G1961), .B(G1966), .Z(new_n649));
  NOR2_X1   g224(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(new_n649), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n647), .A2(new_n652), .A3(new_n650), .ZN(new_n653));
  NAND2_X1  g228(.A1(new_n647), .A2(new_n652), .ZN(new_n654));
  XOR2_X1   g229(.A(KEYINPUT82), .B(KEYINPUT20), .Z(new_n655));
  AOI211_X1 g230(.A(new_n651), .B(new_n653), .C1(new_n654), .C2(new_n655), .ZN(new_n656));
  OAI21_X1  g231(.A(new_n656), .B1(new_n654), .B2(new_n655), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT83), .ZN(new_n658));
  XOR2_X1   g233(.A(G1981), .B(G1986), .Z(new_n659));
  XNOR2_X1  g234(.A(G1991), .B(G1996), .ZN(new_n660));
  XNOR2_X1  g235(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XOR2_X1   g236(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n662));
  XNOR2_X1  g237(.A(new_n661), .B(new_n662), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n658), .B(new_n663), .ZN(new_n664));
  INV_X1    g239(.A(new_n664), .ZN(G229));
  INV_X1    g240(.A(G29), .ZN(new_n666));
  AND2_X1   g241(.A1(new_n666), .A2(G25), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n478), .A2(G131), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n461), .A2(G107), .ZN(new_n669));
  OAI21_X1  g244(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n670));
  INV_X1    g245(.A(G119), .ZN(new_n671));
  OAI221_X1 g246(.A(new_n668), .B1(new_n669), .B2(new_n670), .C1(new_n607), .C2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(KEYINPUT84), .ZN(new_n673));
  AOI21_X1  g248(.A(new_n667), .B1(new_n673), .B2(G29), .ZN(new_n674));
  XOR2_X1   g249(.A(KEYINPUT35), .B(G1991), .Z(new_n675));
  XNOR2_X1  g250(.A(new_n675), .B(KEYINPUT85), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n674), .B(new_n676), .ZN(new_n677));
  INV_X1    g252(.A(G16), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(G24), .ZN(new_n679));
  OAI21_X1  g254(.A(new_n679), .B1(new_n574), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(KEYINPUT86), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n678), .A2(G22), .ZN(new_n683));
  OAI21_X1  g258(.A(new_n683), .B1(G166), .B2(new_n678), .ZN(new_n684));
  INV_X1    g259(.A(G1971), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  NAND2_X1  g261(.A1(G288), .A2(KEYINPUT87), .ZN(new_n687));
  INV_X1    g262(.A(KEYINPUT87), .ZN(new_n688));
  NAND4_X1  g263(.A1(new_n558), .A2(new_n559), .A3(new_n688), .A4(new_n560), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G16), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G16), .B2(G23), .ZN(new_n692));
  XNOR2_X1  g267(.A(KEYINPUT33), .B(G1976), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n692), .A2(new_n693), .ZN(new_n695));
  NOR2_X1   g270(.A1(G6), .A2(G16), .ZN(new_n696));
  INV_X1    g271(.A(G305), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n696), .B1(new_n697), .B2(G16), .ZN(new_n698));
  XOR2_X1   g273(.A(KEYINPUT32), .B(G1981), .Z(new_n699));
  XNOR2_X1  g274(.A(new_n698), .B(new_n699), .ZN(new_n700));
  NAND4_X1  g275(.A1(new_n686), .A2(new_n694), .A3(new_n695), .A4(new_n700), .ZN(new_n701));
  OAI211_X1 g276(.A(new_n677), .B(new_n682), .C1(new_n701), .C2(KEYINPUT34), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n702), .B1(KEYINPUT34), .B2(new_n701), .ZN(new_n703));
  INV_X1    g278(.A(KEYINPUT88), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(KEYINPUT36), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n703), .B(new_n705), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT31), .B(G11), .ZN(new_n707));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n708));
  AND2_X1   g283(.A1(new_n708), .A2(G28), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n666), .B1(new_n708), .B2(G28), .ZN(new_n710));
  OAI221_X1 g285(.A(new_n707), .B1(new_n709), .B2(new_n710), .C1(new_n609), .C2(new_n666), .ZN(new_n711));
  OAI21_X1  g286(.A(G29), .B1(new_n467), .B2(new_n473), .ZN(new_n712));
  INV_X1    g287(.A(KEYINPUT24), .ZN(new_n713));
  INV_X1    g288(.A(G34), .ZN(new_n714));
  AOI21_X1  g289(.A(G29), .B1(new_n713), .B2(new_n714), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  AND2_X1   g291(.A1(new_n712), .A2(new_n716), .ZN(new_n717));
  INV_X1    g292(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n711), .B1(G2084), .B2(new_n718), .ZN(new_n719));
  INV_X1    g294(.A(G2084), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT96), .ZN(new_n722));
  INV_X1    g297(.A(G1966), .ZN(new_n723));
  NOR2_X1   g298(.A1(G168), .A2(new_n678), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(new_n678), .B2(G21), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n719), .B(new_n722), .C1(new_n723), .C2(new_n725), .ZN(new_n726));
  AND2_X1   g301(.A1(new_n666), .A2(G32), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n485), .A2(G129), .ZN(new_n728));
  NAND3_X1  g303(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n729), .B(KEYINPUT26), .ZN(new_n730));
  AND2_X1   g305(.A1(new_n469), .A2(G105), .ZN(new_n731));
  AOI211_X1 g306(.A(new_n730), .B(new_n731), .C1(new_n478), .C2(G141), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n728), .A2(new_n732), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n727), .B1(new_n733), .B2(G29), .ZN(new_n734));
  XNOR2_X1  g309(.A(KEYINPUT27), .B(G1996), .ZN(new_n735));
  AOI22_X1  g310(.A1(new_n725), .A2(new_n723), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  OAI21_X1  g311(.A(new_n736), .B1(new_n734), .B2(new_n735), .ZN(new_n737));
  NOR2_X1   g312(.A1(new_n726), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n678), .A2(G20), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT23), .Z(new_n740));
  AOI21_X1  g315(.A(new_n740), .B1(G299), .B2(G16), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n741), .B(G1956), .ZN(new_n742));
  NOR2_X1   g317(.A1(G29), .A2(G35), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G162), .B2(G29), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT98), .B(KEYINPUT29), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  OAI211_X1 g321(.A(new_n738), .B(new_n742), .C1(G2090), .C2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n746), .A2(G2090), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT99), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n666), .A2(G27), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G164), .B2(new_n666), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n751), .B(KEYINPUT97), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n752), .B(G2078), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n678), .A2(G5), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n754), .B1(G171), .B2(new_n678), .ZN(new_n755));
  INV_X1    g330(.A(G1961), .ZN(new_n756));
  XNOR2_X1  g331(.A(new_n755), .B(new_n756), .ZN(new_n757));
  NAND2_X1  g332(.A1(new_n666), .A2(G33), .ZN(new_n758));
  NAND3_X1  g333(.A1(new_n478), .A2(KEYINPUT93), .A3(G139), .ZN(new_n759));
  NAND3_X1  g334(.A1(new_n461), .A2(G103), .A3(G2104), .ZN(new_n760));
  XOR2_X1   g335(.A(new_n760), .B(KEYINPUT25), .Z(new_n761));
  NAND2_X1  g336(.A1(new_n759), .A2(new_n761), .ZN(new_n762));
  AOI21_X1  g337(.A(KEYINPUT93), .B1(new_n478), .B2(G139), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n762), .A2(KEYINPUT94), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(KEYINPUT94), .B1(new_n762), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n462), .A2(G127), .ZN(new_n767));
  AND2_X1   g342(.A1(G115), .A2(G2104), .ZN(new_n768));
  OAI21_X1  g343(.A(G2105), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n766), .A2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n758), .B1(new_n771), .B2(new_n666), .ZN(new_n772));
  OAI211_X1 g347(.A(new_n753), .B(new_n757), .C1(new_n772), .C2(G2072), .ZN(new_n773));
  NOR3_X1   g348(.A1(new_n747), .A2(new_n749), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n666), .A2(G26), .ZN(new_n775));
  XNOR2_X1  g350(.A(new_n775), .B(KEYINPUT28), .ZN(new_n776));
  OAI21_X1  g351(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n777));
  INV_X1    g352(.A(G116), .ZN(new_n778));
  AOI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(G2105), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n478), .B2(G140), .ZN(new_n780));
  INV_X1    g355(.A(G128), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n780), .B1(new_n607), .B2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(KEYINPUT91), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  OAI21_X1  g359(.A(new_n776), .B1(new_n784), .B2(new_n666), .ZN(new_n785));
  INV_X1    g360(.A(G2067), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NOR2_X1   g362(.A1(G16), .A2(G19), .ZN(new_n788));
  AOI21_X1  g363(.A(new_n788), .B1(new_n542), .B2(G16), .ZN(new_n789));
  XNOR2_X1  g364(.A(KEYINPUT90), .B(G1341), .ZN(new_n790));
  XNOR2_X1  g365(.A(new_n789), .B(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n678), .A2(G4), .ZN(new_n792));
  OAI21_X1  g367(.A(new_n792), .B1(new_n593), .B2(new_n678), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT89), .B(G1348), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NAND3_X1  g370(.A1(new_n787), .A2(new_n791), .A3(new_n795), .ZN(new_n796));
  XOR2_X1   g371(.A(new_n796), .B(KEYINPUT92), .Z(new_n797));
  NAND2_X1  g372(.A1(new_n772), .A2(G2072), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(KEYINPUT95), .ZN(new_n799));
  AND3_X1   g374(.A1(new_n774), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  AND2_X1   g375(.A1(new_n706), .A2(new_n800), .ZN(G311));
  NAND2_X1  g376(.A1(new_n706), .A2(new_n800), .ZN(G150));
  AOI22_X1  g377(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n803));
  INV_X1    g378(.A(G93), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n803), .A2(new_n509), .B1(new_n804), .B2(new_n512), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT100), .B(G55), .Z(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(new_n521), .B2(new_n522), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n805), .A2(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(G860), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT37), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n593), .A2(G559), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n812), .B(KEYINPUT101), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT38), .ZN(new_n814));
  OR2_X1    g389(.A1(new_n805), .A2(new_n807), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n815), .A2(new_n541), .ZN(new_n816));
  NAND4_X1  g391(.A1(new_n808), .A2(new_n535), .A3(new_n537), .A4(new_n540), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n816), .A2(new_n817), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n814), .B(new_n818), .ZN(new_n819));
  AND2_X1   g394(.A1(new_n819), .A2(KEYINPUT39), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n809), .B1(new_n819), .B2(KEYINPUT39), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n811), .B1(new_n820), .B2(new_n821), .ZN(G145));
  XNOR2_X1  g397(.A(new_n609), .B(G160), .ZN(new_n823));
  XOR2_X1   g398(.A(new_n823), .B(G162), .Z(new_n824));
  XNOR2_X1  g399(.A(new_n782), .B(KEYINPUT91), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n825), .A2(new_n733), .ZN(new_n826));
  INV_X1    g401(.A(new_n733), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n784), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g403(.A(new_n770), .B1(new_n826), .B2(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(KEYINPUT102), .ZN(new_n831));
  INV_X1    g406(.A(new_n497), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n496), .B1(new_n462), .B2(new_n494), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n831), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND3_X1  g409(.A1(new_n500), .A2(KEYINPUT102), .A3(new_n497), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n492), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n826), .A2(new_n828), .A3(new_n770), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n830), .A2(new_n836), .A3(new_n837), .ZN(new_n838));
  AND2_X1   g413(.A1(new_n488), .A2(new_n491), .ZN(new_n839));
  AND3_X1   g414(.A1(new_n500), .A2(KEYINPUT102), .A3(new_n497), .ZN(new_n840));
  AOI21_X1  g415(.A(KEYINPUT102), .B1(new_n500), .B2(new_n497), .ZN(new_n841));
  OAI21_X1  g416(.A(new_n839), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(new_n837), .ZN(new_n843));
  OAI21_X1  g418(.A(new_n842), .B1(new_n843), .B2(new_n829), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n838), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n478), .A2(G142), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n461), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G130), .B2(new_n485), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(new_n601), .Z(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(new_n673), .ZN(new_n852));
  AOI21_X1  g427(.A(new_n824), .B1(new_n845), .B2(new_n852), .ZN(new_n853));
  INV_X1    g428(.A(new_n852), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n854), .A2(new_n838), .A3(new_n844), .ZN(new_n855));
  AOI21_X1  g430(.A(G37), .B1(new_n853), .B2(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT103), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n845), .B1(new_n857), .B2(new_n854), .ZN(new_n858));
  NAND4_X1  g433(.A1(new_n838), .A2(new_n844), .A3(KEYINPUT103), .A4(new_n852), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n858), .A2(new_n824), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n856), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(new_n861), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g437(.A1(new_n585), .A2(G299), .ZN(new_n863));
  NAND4_X1  g438(.A1(new_n579), .A2(new_n584), .A3(new_n554), .A4(new_n552), .ZN(new_n864));
  AND3_X1   g439(.A1(new_n863), .A2(KEYINPUT41), .A3(new_n864), .ZN(new_n865));
  AOI21_X1  g440(.A(KEYINPUT41), .B1(new_n863), .B2(new_n864), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n818), .A2(new_n597), .ZN(new_n868));
  OAI211_X1 g443(.A(new_n816), .B(new_n817), .C1(G559), .C2(new_n585), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n867), .A2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(KEYINPUT105), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n871), .B(new_n872), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n690), .B(G303), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n574), .A2(G305), .ZN(new_n875));
  NOR2_X1   g450(.A1(G290), .A2(new_n697), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n874), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(G166), .B(new_n690), .ZN(new_n878));
  NOR2_X1   g453(.A1(new_n876), .A2(new_n875), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT42), .ZN(new_n882));
  NAND4_X1  g457(.A1(new_n868), .A2(new_n863), .A3(new_n864), .A4(new_n869), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT104), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n883), .B(new_n884), .ZN(new_n885));
  AND3_X1   g460(.A1(new_n873), .A2(new_n882), .A3(new_n885), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n882), .B1(new_n873), .B2(new_n885), .ZN(new_n887));
  OAI21_X1  g462(.A(G868), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT106), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n808), .A2(G868), .ZN(new_n890));
  INV_X1    g465(.A(new_n890), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(new_n889), .B1(new_n888), .B2(new_n891), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n893), .ZN(G295));
  NAND2_X1  g469(.A1(new_n888), .A2(new_n891), .ZN(G331));
  INV_X1    g470(.A(KEYINPUT44), .ZN(new_n896));
  AND2_X1   g471(.A1(new_n877), .A2(new_n880), .ZN(new_n897));
  NAND2_X1  g472(.A1(G171), .A2(G168), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n533), .A2(G52), .ZN(new_n899));
  OAI22_X1  g474(.A1(new_n899), .A2(new_n532), .B1(new_n523), .B2(new_n528), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n818), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  NAND4_X1  g478(.A1(new_n816), .A2(new_n898), .A3(new_n817), .A4(new_n900), .ZN(new_n904));
  NAND3_X1  g479(.A1(new_n902), .A2(new_n903), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n818), .A2(new_n901), .A3(KEYINPUT109), .ZN(new_n906));
  AND3_X1   g481(.A1(new_n905), .A2(new_n867), .A3(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n863), .A2(new_n864), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n902), .A2(new_n909), .A3(new_n904), .ZN(new_n910));
  AND2_X1   g485(.A1(new_n898), .A2(new_n900), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n911), .A2(KEYINPUT108), .A3(new_n816), .A4(new_n817), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n908), .B1(new_n910), .B2(new_n912), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n897), .B1(new_n907), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n910), .A2(new_n867), .A3(new_n912), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n905), .A2(new_n906), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n881), .B(new_n915), .C1(new_n916), .C2(new_n908), .ZN(new_n917));
  INV_X1    g492(.A(G37), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n914), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n919), .A2(KEYINPUT43), .ZN(new_n920));
  INV_X1    g495(.A(KEYINPUT111), .ZN(new_n921));
  AND3_X1   g496(.A1(new_n910), .A2(new_n867), .A3(new_n912), .ZN(new_n922));
  AOI21_X1  g497(.A(new_n908), .B1(new_n905), .B2(new_n906), .ZN(new_n923));
  OAI21_X1  g498(.A(new_n897), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AND3_X1   g499(.A1(new_n924), .A2(new_n917), .A3(new_n918), .ZN(new_n925));
  XNOR2_X1  g500(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n926));
  AOI22_X1  g501(.A1(new_n920), .A2(new_n921), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n919), .A2(KEYINPUT111), .A3(KEYINPUT43), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n896), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT110), .ZN(new_n930));
  NAND4_X1  g505(.A1(new_n914), .A2(new_n917), .A3(new_n918), .A4(new_n926), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n930), .B(new_n931), .C1(new_n925), .C2(new_n926), .ZN(new_n932));
  OR2_X1    g507(.A1(new_n931), .A2(new_n930), .ZN(new_n933));
  AOI21_X1  g508(.A(KEYINPUT44), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n929), .A2(new_n934), .ZN(G397));
  XNOR2_X1  g510(.A(new_n673), .B(new_n676), .ZN(new_n936));
  INV_X1    g511(.A(G1996), .ZN(new_n937));
  XNOR2_X1  g512(.A(new_n733), .B(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n825), .A2(G2067), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n784), .A2(new_n786), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n938), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  NOR2_X1   g516(.A1(new_n936), .A2(new_n941), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n574), .B(G1986), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  OAI21_X1  g519(.A(KEYINPUT112), .B1(new_n836), .B2(G1384), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT112), .ZN(new_n946));
  INV_X1    g521(.A(G1384), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n842), .A2(new_n946), .A3(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT45), .ZN(new_n949));
  NAND3_X1  g524(.A1(new_n945), .A2(new_n948), .A3(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G40), .ZN(new_n951));
  NOR3_X1   g526(.A1(new_n467), .A2(new_n473), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(new_n952), .ZN(new_n953));
  NOR2_X1   g528(.A1(new_n950), .A2(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n944), .A2(new_n954), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT126), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT50), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n842), .A2(KEYINPUT114), .A3(new_n957), .A4(new_n947), .ZN(new_n958));
  NOR3_X1   g533(.A1(new_n836), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT114), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n500), .A2(new_n497), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n961), .A2(new_n839), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(new_n947), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n960), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n964));
  OAI211_X1 g539(.A(new_n952), .B(new_n958), .C1(new_n959), .C2(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n952), .B1(new_n963), .B2(new_n949), .ZN(new_n966));
  NAND2_X1  g541(.A1(new_n842), .A2(new_n947), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n966), .B1(new_n949), .B2(new_n967), .ZN(new_n968));
  OAI22_X1  g543(.A1(new_n965), .A2(G2084), .B1(new_n968), .B2(G1966), .ZN(new_n969));
  XNOR2_X1  g544(.A(KEYINPUT115), .B(G8), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(G286), .A3(new_n971), .ZN(new_n972));
  NOR2_X1   g547(.A1(G168), .A2(new_n970), .ZN(new_n973));
  INV_X1    g548(.A(G8), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n842), .A2(new_n957), .A3(new_n947), .ZN(new_n975));
  AOI21_X1  g550(.A(G1384), .B1(new_n961), .B2(new_n839), .ZN(new_n976));
  OAI21_X1  g551(.A(KEYINPUT114), .B1(new_n976), .B2(new_n957), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n953), .B1(new_n975), .B2(new_n977), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n978), .A2(new_n720), .A3(new_n958), .ZN(new_n979));
  NOR2_X1   g554(.A1(new_n836), .A2(G1384), .ZN(new_n980));
  NOR2_X1   g555(.A1(new_n980), .A2(KEYINPUT45), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n723), .B1(new_n981), .B2(new_n966), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n974), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n972), .B(KEYINPUT51), .C1(new_n973), .C2(new_n983), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n970), .B1(new_n979), .B2(new_n982), .ZN(new_n985));
  INV_X1    g560(.A(new_n973), .ZN(new_n986));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n985), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT62), .B1(new_n984), .B2(new_n990), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT49), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n697), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT118), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n567), .A2(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n992), .B1(new_n563), .B2(new_n567), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND4_X1  g572(.A1(new_n993), .A2(G1981), .A3(new_n995), .A4(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n970), .B1(new_n980), .B2(new_n952), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n995), .A2(G1981), .ZN(new_n1000));
  NOR2_X1   g575(.A1(G305), .A2(KEYINPUT49), .ZN(new_n1001));
  OAI21_X1  g576(.A(new_n1000), .B1(new_n1001), .B2(new_n996), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n998), .A2(new_n999), .A3(new_n1002), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n687), .A2(G1976), .A3(new_n689), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT116), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n842), .A2(new_n947), .A3(new_n952), .ZN(new_n1007));
  NAND4_X1  g582(.A1(new_n687), .A2(KEYINPUT116), .A3(G1976), .A4(new_n689), .ZN(new_n1008));
  NAND4_X1  g583(.A1(new_n1006), .A2(new_n971), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n1009), .A2(KEYINPUT52), .ZN(new_n1010));
  XNOR2_X1  g585(.A(KEYINPUT117), .B(G1976), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT52), .B1(G288), .B2(new_n1011), .ZN(new_n1012));
  NAND4_X1  g587(.A1(new_n999), .A2(new_n1006), .A3(new_n1008), .A4(new_n1012), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1003), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1014));
  NAND2_X1  g589(.A1(G303), .A2(G8), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n1015), .B(KEYINPUT55), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(G2090), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n978), .A2(new_n1018), .A3(new_n958), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n976), .B2(KEYINPUT45), .ZN(new_n1021));
  OAI211_X1 g596(.A(KEYINPUT113), .B(new_n949), .C1(G164), .C2(G1384), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n842), .A2(KEYINPUT45), .A3(new_n947), .ZN(new_n1024));
  NAND3_X1  g599(.A1(new_n1023), .A2(new_n952), .A3(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1025), .A2(new_n685), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n974), .B1(new_n1019), .B2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g602(.A(new_n1014), .B1(new_n1017), .B2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G2078), .ZN(new_n1029));
  NAND4_X1  g604(.A1(new_n1023), .A2(new_n1029), .A3(new_n952), .A4(new_n1024), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT53), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n756), .A2(new_n965), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n968), .A2(KEYINPUT53), .A3(new_n1029), .ZN(new_n1033));
  AOI21_X1  g608(.A(G301), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n957), .B1(new_n842), .B2(new_n947), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n952), .B1(new_n963), .B2(KEYINPUT50), .ZN(new_n1036));
  NOR3_X1   g611(.A1(new_n1035), .A2(new_n1036), .A3(G2090), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1037), .B1(new_n685), .B2(new_n1025), .ZN(new_n1038));
  OAI21_X1  g613(.A(new_n1016), .B1(new_n1038), .B2(new_n970), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1028), .A2(new_n1034), .A3(new_n1039), .ZN(new_n1040));
  OAI21_X1  g615(.A(new_n956), .B1(new_n991), .B2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1027), .A2(new_n1017), .ZN(new_n1042));
  AND3_X1   g617(.A1(new_n1003), .A2(new_n1010), .A3(new_n1013), .ZN(new_n1043));
  AND4_X1   g618(.A1(new_n1034), .A2(new_n1042), .A3(new_n1039), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n969), .A2(G8), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n987), .B1(new_n1045), .B2(new_n986), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n989), .B1(new_n1046), .B2(new_n972), .ZN(new_n1047));
  OAI211_X1 g622(.A(KEYINPUT126), .B(new_n1044), .C1(new_n1047), .C2(KEYINPUT62), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1049));
  AND3_X1   g624(.A1(new_n1041), .A2(new_n1048), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(G288), .A2(G1976), .ZN(new_n1051));
  AND2_X1   g626(.A1(new_n1003), .A2(new_n1051), .ZN(new_n1052));
  NOR2_X1   g627(.A1(G305), .A2(G1981), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n999), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(new_n1042), .B2(new_n1014), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n985), .A2(G168), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT63), .ZN(new_n1057));
  NOR2_X1   g632(.A1(new_n1056), .A2(new_n1057), .ZN(new_n1058));
  OAI211_X1 g633(.A(new_n1058), .B(new_n1028), .C1(new_n1017), .C2(new_n1027), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1042), .A2(new_n1039), .A3(new_n1043), .ZN(new_n1060));
  OAI21_X1  g635(.A(new_n1057), .B1(new_n1060), .B2(new_n1056), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1055), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(G1348), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n965), .A2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g639(.A1(new_n1007), .A2(G2067), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(new_n585), .B(KEYINPUT122), .ZN(new_n1067));
  NAND4_X1  g642(.A1(new_n1064), .A2(KEYINPUT60), .A3(new_n1066), .A4(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT60), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1348), .B1(new_n978), .B2(new_n958), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n1069), .B1(new_n1070), .B2(new_n1065), .ZN(new_n1071));
  AOI211_X1 g646(.A(new_n1069), .B(new_n1065), .C1(new_n965), .C2(new_n1063), .ZN(new_n1072));
  OR2_X1    g647(.A1(new_n593), .A2(KEYINPUT122), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(new_n1071), .C1(new_n1072), .C2(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT61), .ZN(new_n1075));
  XNOR2_X1  g650(.A(KEYINPUT56), .B(G2072), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1023), .A2(new_n952), .A3(new_n1024), .A4(new_n1076), .ZN(new_n1077));
  INV_X1    g652(.A(G1956), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1078), .B1(new_n1035), .B2(new_n1036), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1077), .A2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g655(.A(KEYINPUT57), .B1(new_n554), .B2(KEYINPUT119), .ZN(new_n1081));
  NAND2_X1  g656(.A1(G299), .A2(new_n1081), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n552), .B(new_n554), .C1(KEYINPUT119), .C2(KEYINPUT57), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(new_n1084), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1080), .A2(KEYINPUT121), .A3(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1077), .A2(new_n1079), .A3(new_n1084), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(new_n1084), .B1(new_n1077), .B2(new_n1079), .ZN(new_n1090));
  OAI211_X1 g665(.A(new_n1075), .B(new_n1086), .C1(new_n1089), .C2(new_n1090), .ZN(new_n1091));
  XOR2_X1   g666(.A(KEYINPUT58), .B(G1341), .Z(new_n1092));
  NAND2_X1  g667(.A1(new_n1007), .A2(new_n1092), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1093), .B1(new_n1025), .B2(G1996), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1094), .A2(KEYINPUT59), .A3(new_n542), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1094), .A2(new_n542), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1096), .A2(new_n1097), .B1(KEYINPUT61), .B2(new_n1087), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1074), .A2(new_n1091), .A3(new_n1095), .A4(new_n1098), .ZN(new_n1099));
  OR2_X1    g674(.A1(new_n1080), .A2(KEYINPUT120), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n1084), .B1(new_n1080), .B2(KEYINPUT120), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n585), .B1(new_n1064), .B2(new_n1066), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1100), .A2(new_n1101), .B1(new_n1102), .B2(new_n1087), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1099), .A2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT54), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n965), .A2(new_n756), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n463), .A2(new_n466), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n461), .B1(new_n1107), .B2(KEYINPUT123), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(KEYINPUT123), .B2(new_n1107), .ZN(new_n1109));
  NOR4_X1   g684(.A1(new_n473), .A2(new_n1031), .A3(new_n951), .A4(G2078), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n950), .A2(new_n1024), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1112));
  AND4_X1   g687(.A1(G301), .A2(new_n1106), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1105), .B1(new_n1034), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT124), .ZN(new_n1115));
  AOI21_X1  g690(.A(new_n1060), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1104), .A2(new_n1116), .ZN(new_n1117));
  OAI211_X1 g692(.A(KEYINPUT124), .B(new_n1105), .C1(new_n1034), .C2(new_n1113), .ZN(new_n1118));
  INV_X1    g693(.A(KEYINPUT125), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1106), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1120));
  AOI21_X1  g695(.A(new_n1119), .B1(new_n1120), .B2(G171), .ZN(new_n1121));
  NAND3_X1  g696(.A1(new_n1120), .A2(new_n1119), .A3(G171), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1032), .A2(G301), .A3(new_n1033), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1122), .A2(KEYINPUT54), .A3(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1047), .B(new_n1118), .C1(new_n1121), .C2(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1062), .B1(new_n1117), .B2(new_n1125), .ZN(new_n1126));
  OAI21_X1  g701(.A(new_n955), .B1(new_n1050), .B2(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(new_n954), .ZN(new_n1128));
  NOR3_X1   g703(.A1(new_n1128), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT46), .ZN(new_n1130));
  AOI21_X1  g705(.A(new_n1130), .B1(new_n954), .B2(new_n937), .ZN(new_n1131));
  AND3_X1   g706(.A1(new_n939), .A2(new_n940), .A3(new_n827), .ZN(new_n1132));
  OAI22_X1  g707(.A1(new_n1129), .A2(new_n1131), .B1(new_n1128), .B2(new_n1132), .ZN(new_n1133));
  XOR2_X1   g708(.A(new_n1133), .B(KEYINPUT47), .Z(new_n1134));
  OR2_X1    g709(.A1(new_n673), .A2(new_n676), .ZN(new_n1135));
  OAI21_X1  g710(.A(new_n940), .B1(new_n1135), .B2(new_n941), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1136), .A2(new_n954), .ZN(new_n1137));
  OR3_X1    g712(.A1(new_n1128), .A2(G1986), .A3(G290), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT48), .ZN(new_n1139));
  OAI22_X1  g714(.A1(new_n942), .A2(new_n1128), .B1(new_n1138), .B2(new_n1139), .ZN(new_n1140));
  AND2_X1   g715(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1141));
  OAI21_X1  g716(.A(new_n1137), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1134), .A2(new_n1142), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1127), .A2(new_n1143), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g719(.A1(G227), .A2(new_n459), .ZN(new_n1146));
  OR2_X1    g720(.A1(new_n1146), .A2(KEYINPUT127), .ZN(new_n1147));
  NAND2_X1  g721(.A1(new_n1146), .A2(KEYINPUT127), .ZN(new_n1148));
  NAND4_X1  g722(.A1(new_n1147), .A2(new_n664), .A3(new_n628), .A4(new_n1148), .ZN(new_n1149));
  AOI21_X1  g723(.A(new_n1149), .B1(new_n856), .B2(new_n860), .ZN(new_n1150));
  NAND3_X1  g724(.A1(new_n1150), .A2(new_n932), .A3(new_n933), .ZN(G225));
  INV_X1    g725(.A(G225), .ZN(G308));
endmodule


