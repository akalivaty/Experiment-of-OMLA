//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 0 0 0 1 0 0 0 1 0 1 0 0 0 1 0 1 0 1 0 1 0 1 0 0 1 1 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:19 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n779, new_n780, new_n781, new_n782, new_n784, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n791, new_n792, new_n793, new_n794,
    new_n795, new_n796, new_n797, new_n798, new_n799, new_n800, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n877, new_n878, new_n879, new_n881, new_n882, new_n883, new_n885,
    new_n886, new_n887, new_n888, new_n889, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n981, new_n982, new_n984, new_n985, new_n986,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002;
  INV_X1    g000(.A(KEYINPUT5), .ZN(new_n202));
  NAND2_X1  g001(.A1(G155gat), .A2(G162gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT2), .ZN(new_n204));
  INV_X1    g003(.A(G141gat), .ZN(new_n205));
  INV_X1    g004(.A(G148gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g006(.A1(G141gat), .A2(G148gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n204), .A2(new_n207), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT73), .ZN(new_n210));
  XNOR2_X1  g009(.A(G155gat), .B(G162gat), .ZN(new_n211));
  INV_X1    g010(.A(new_n211), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n210), .A2(new_n212), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n209), .A2(KEYINPUT73), .A3(new_n211), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(G127gat), .B(G134gat), .ZN(new_n216));
  INV_X1    g015(.A(new_n216), .ZN(new_n217));
  AND2_X1   g016(.A1(G113gat), .A2(G120gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT1), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n219), .B1(G113gat), .B2(G120gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(G113gat), .ZN(new_n222));
  INV_X1    g021(.A(G120gat), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT1), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT66), .B(G120gat), .ZN(new_n225));
  OAI211_X1 g024(.A(new_n224), .B(new_n216), .C1(new_n225), .C2(new_n222), .ZN(new_n226));
  NAND3_X1  g025(.A1(new_n215), .A2(new_n221), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n216), .A2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n223), .A2(KEYINPUT66), .ZN(new_n229));
  INV_X1    g028(.A(KEYINPUT66), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n230), .A2(G120gat), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n222), .B1(new_n229), .B2(new_n231), .ZN(new_n232));
  NOR2_X1   g031(.A1(new_n220), .A2(new_n218), .ZN(new_n233));
  OAI22_X1  g032(.A1(new_n228), .A2(new_n232), .B1(new_n233), .B2(new_n216), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT74), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n221), .A2(new_n226), .A3(KEYINPUT74), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n227), .B1(new_n238), .B2(new_n215), .ZN(new_n239));
  NAND2_X1  g038(.A1(G225gat), .A2(G233gat), .ZN(new_n240));
  INV_X1    g039(.A(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n202), .B1(new_n239), .B2(new_n241), .ZN(new_n242));
  XOR2_X1   g041(.A(KEYINPUT75), .B(KEYINPUT3), .Z(new_n243));
  AND3_X1   g042(.A1(new_n209), .A2(KEYINPUT73), .A3(new_n211), .ZN(new_n244));
  AOI21_X1  g043(.A(new_n211), .B1(new_n209), .B2(KEYINPUT73), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n213), .A2(KEYINPUT3), .A3(new_n214), .ZN(new_n247));
  NAND4_X1  g046(.A1(new_n246), .A2(new_n247), .A3(new_n236), .A4(new_n237), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n234), .A2(KEYINPUT67), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n221), .A2(new_n226), .A3(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n249), .A2(new_n215), .A3(KEYINPUT4), .A4(new_n251), .ZN(new_n252));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n244), .A2(new_n245), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n253), .B1(new_n254), .B2(new_n234), .ZN(new_n255));
  NAND4_X1  g054(.A1(new_n248), .A2(new_n252), .A3(new_n255), .A4(new_n240), .ZN(new_n256));
  AND3_X1   g055(.A1(new_n248), .A2(new_n202), .A3(new_n240), .ZN(new_n257));
  NAND4_X1  g056(.A1(new_n249), .A2(new_n215), .A3(new_n253), .A4(new_n251), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n254), .A2(new_n234), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n258), .B1(new_n259), .B2(new_n253), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n242), .A2(new_n256), .B1(new_n257), .B2(new_n260), .ZN(new_n261));
  XOR2_X1   g060(.A(G1gat), .B(G29gat), .Z(new_n262));
  XNOR2_X1  g061(.A(new_n262), .B(KEYINPUT0), .ZN(new_n263));
  XNOR2_X1  g062(.A(G57gat), .B(G85gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n263), .B(new_n264), .ZN(new_n265));
  OAI21_X1  g064(.A(KEYINPUT81), .B1(new_n261), .B2(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(KEYINPUT76), .B(KEYINPUT6), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n268), .B1(new_n261), .B2(new_n265), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n239), .A2(new_n241), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n270), .A2(new_n256), .A3(KEYINPUT5), .ZN(new_n271));
  NAND4_X1  g070(.A1(new_n260), .A2(new_n202), .A3(new_n240), .A4(new_n248), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT81), .ZN(new_n274));
  INV_X1    g073(.A(new_n265), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(new_n274), .A3(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(new_n266), .A2(new_n269), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n277), .A2(KEYINPUT82), .ZN(new_n278));
  AOI211_X1 g077(.A(new_n265), .B(new_n267), .C1(new_n271), .C2(new_n272), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT82), .ZN(new_n281));
  NAND4_X1  g080(.A1(new_n266), .A2(new_n269), .A3(new_n276), .A4(new_n281), .ZN(new_n282));
  NAND3_X1  g081(.A1(new_n278), .A2(new_n280), .A3(new_n282), .ZN(new_n283));
  AND2_X1   g082(.A1(G228gat), .A2(G233gat), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT29), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n246), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT70), .ZN(new_n288));
  INV_X1    g087(.A(G197gat), .ZN(new_n289));
  INV_X1    g088(.A(G204gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g090(.A1(G197gat), .A2(G204gat), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT22), .ZN(new_n293));
  NAND2_X1  g092(.A1(G211gat), .A2(G218gat), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n291), .A2(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  XNOR2_X1  g094(.A(G211gat), .B(G218gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n288), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n296), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n295), .B2(KEYINPUT69), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n291), .A2(new_n292), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n294), .A2(new_n293), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n300), .A2(KEYINPUT69), .A3(new_n301), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n297), .B1(new_n299), .B2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT69), .ZN(new_n304));
  XOR2_X1   g103(.A(G197gat), .B(G204gat), .Z(new_n305));
  INV_X1    g104(.A(new_n301), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n300), .A2(KEYINPUT69), .A3(new_n301), .ZN(new_n308));
  NAND4_X1  g107(.A1(new_n307), .A2(new_n288), .A3(new_n298), .A4(new_n308), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n303), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n287), .A2(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n295), .A2(new_n296), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n295), .A2(new_n296), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n286), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n215), .B1(new_n314), .B2(new_n243), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n285), .B1(new_n311), .B2(new_n315), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n285), .B1(new_n287), .B2(new_n310), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n303), .A2(new_n286), .A3(new_n309), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT3), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n215), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  OAI21_X1  g119(.A(new_n317), .B1(new_n320), .B2(KEYINPUT78), .ZN(new_n321));
  INV_X1    g120(.A(KEYINPUT78), .ZN(new_n322));
  AOI211_X1 g121(.A(new_n322), .B(new_n215), .C1(new_n318), .C2(new_n319), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n316), .B1(new_n321), .B2(new_n323), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(G22gat), .ZN(new_n325));
  INV_X1    g124(.A(G22gat), .ZN(new_n326));
  OAI211_X1 g125(.A(new_n316), .B(new_n326), .C1(new_n321), .C2(new_n323), .ZN(new_n327));
  XNOR2_X1  g126(.A(G78gat), .B(G106gat), .ZN(new_n328));
  INV_X1    g127(.A(G50gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(KEYINPUT77), .B(KEYINPUT31), .ZN(new_n331));
  XNOR2_X1  g130(.A(new_n330), .B(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n332), .B1(new_n325), .B2(new_n327), .ZN(new_n334));
  NOR2_X1   g133(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT65), .ZN(new_n336));
  INV_X1    g135(.A(G169gat), .ZN(new_n337));
  INV_X1    g136(.A(G176gat), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(KEYINPUT26), .ZN(new_n340));
  NAND2_X1  g139(.A1(G169gat), .A2(G176gat), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT26), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n336), .A2(new_n342), .A3(new_n337), .A4(new_n338), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  NAND2_X1  g143(.A1(G183gat), .A2(G190gat), .ZN(new_n345));
  INV_X1    g144(.A(G183gat), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n346), .A2(KEYINPUT27), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT27), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n348), .A2(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n347), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n351), .A2(KEYINPUT28), .ZN(new_n352));
  XNOR2_X1  g151(.A(KEYINPUT27), .B(G183gat), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT28), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n350), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n344), .A2(new_n345), .A3(new_n352), .A4(new_n355), .ZN(new_n356));
  OAI21_X1  g155(.A(KEYINPUT64), .B1(G169gat), .B2(G176gat), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT23), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(KEYINPUT64), .B(KEYINPUT23), .C1(G169gat), .C2(G176gat), .ZN(new_n360));
  AND2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT24), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(G183gat), .A3(G190gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n345), .A2(KEYINPUT24), .ZN(new_n364));
  NOR2_X1   g163(.A1(G183gat), .A2(G190gat), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n341), .B(new_n363), .C1(new_n364), .C2(new_n365), .ZN(new_n366));
  INV_X1    g165(.A(KEYINPUT25), .ZN(new_n367));
  NOR3_X1   g166(.A1(new_n361), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n341), .B1(new_n345), .B2(KEYINPUT24), .ZN(new_n369));
  INV_X1    g168(.A(new_n365), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n362), .B1(G183gat), .B2(G190gat), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n369), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n359), .A2(new_n360), .ZN(new_n373));
  AOI21_X1  g172(.A(KEYINPUT25), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n356), .B1(new_n368), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n249), .A2(new_n251), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n375), .A2(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(G227gat), .ZN(new_n378));
  INV_X1    g177(.A(G233gat), .ZN(new_n379));
  NOR2_X1   g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n367), .B1(new_n361), .B2(new_n366), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n372), .A2(KEYINPUT25), .A3(new_n373), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n384), .A2(new_n249), .A3(new_n251), .A4(new_n356), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n377), .A2(new_n381), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT34), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT34), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n377), .A2(new_n388), .A3(new_n385), .A4(new_n381), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  XOR2_X1   g189(.A(KEYINPUT68), .B(G71gat), .Z(new_n391));
  XNOR2_X1  g190(.A(new_n391), .B(G99gat), .ZN(new_n392));
  XOR2_X1   g191(.A(G15gat), .B(G43gat), .Z(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  NOR2_X1   g193(.A1(new_n375), .A2(new_n376), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n384), .A2(new_n356), .B1(new_n249), .B2(new_n251), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n380), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT33), .ZN(new_n398));
  AOI21_X1  g197(.A(new_n394), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n390), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n377), .A2(new_n385), .ZN(new_n401));
  AOI21_X1  g200(.A(KEYINPUT33), .B1(new_n401), .B2(new_n380), .ZN(new_n402));
  OAI211_X1 g201(.A(new_n387), .B(new_n389), .C1(new_n402), .C2(new_n394), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n404));
  INV_X1    g203(.A(new_n404), .ZN(new_n405));
  AND3_X1   g204(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n405), .B1(new_n400), .B2(new_n403), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(new_n310), .ZN(new_n409));
  NAND2_X1  g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  XNOR2_X1  g209(.A(new_n410), .B(KEYINPUT71), .ZN(new_n411));
  AND3_X1   g210(.A1(new_n352), .A2(new_n355), .A3(new_n345), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n344), .A2(new_n412), .B1(new_n382), .B2(new_n383), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n411), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n414));
  INV_X1    g213(.A(new_n410), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n375), .A2(new_n415), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n409), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n375), .B2(new_n286), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n411), .B1(new_n384), .B2(new_n356), .ZN(new_n419));
  NOR3_X1   g218(.A1(new_n418), .A2(new_n310), .A3(new_n419), .ZN(new_n420));
  OAI21_X1  g219(.A(KEYINPUT72), .B1(new_n417), .B2(new_n420), .ZN(new_n421));
  XNOR2_X1  g220(.A(G8gat), .B(G36gat), .ZN(new_n422));
  XNOR2_X1  g221(.A(G64gat), .B(G92gat), .ZN(new_n423));
  XOR2_X1   g222(.A(new_n422), .B(new_n423), .Z(new_n424));
  INV_X1    g223(.A(new_n424), .ZN(new_n425));
  INV_X1    g224(.A(new_n411), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n426), .B1(new_n375), .B2(new_n286), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n413), .A2(new_n410), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n310), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n410), .B1(new_n413), .B2(KEYINPUT29), .ZN(new_n430));
  INV_X1    g229(.A(new_n419), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(new_n409), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT72), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n429), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n421), .A2(new_n425), .A3(new_n434), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n429), .A2(new_n432), .A3(KEYINPUT30), .A4(new_n424), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n429), .A2(new_n432), .A3(new_n424), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n435), .A2(new_n436), .A3(new_n439), .ZN(new_n440));
  NOR2_X1   g239(.A1(new_n440), .A2(KEYINPUT35), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n283), .A2(new_n335), .A3(new_n408), .A4(new_n441), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n273), .A2(new_n275), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n279), .B1(new_n443), .B2(new_n269), .ZN(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n440), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n332), .ZN(new_n448));
  AND2_X1   g247(.A1(new_n318), .A2(new_n319), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n322), .B1(new_n449), .B2(new_n215), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n320), .A2(KEYINPUT78), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n450), .A2(new_n451), .A3(new_n317), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n326), .B1(new_n452), .B2(new_n316), .ZN(new_n453));
  INV_X1    g252(.A(new_n327), .ZN(new_n454));
  OAI21_X1  g253(.A(new_n448), .B1(new_n453), .B2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n400), .A2(new_n403), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n456), .A2(new_n404), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n325), .A2(new_n327), .A3(new_n332), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n400), .A2(new_n403), .A3(new_n405), .ZN(new_n459));
  NAND4_X1  g258(.A1(new_n455), .A2(new_n457), .A3(new_n458), .A4(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT85), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n335), .A2(KEYINPUT85), .A3(new_n408), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n447), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g263(.A(KEYINPUT35), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n442), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  OAI22_X1  g265(.A1(new_n444), .A2(new_n440), .B1(new_n333), .B2(new_n334), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT36), .ZN(new_n468));
  NOR3_X1   g267(.A1(new_n406), .A2(new_n407), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(KEYINPUT36), .B1(new_n457), .B2(new_n459), .ZN(new_n470));
  OAI21_X1  g269(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT79), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n468), .B1(new_n406), .B2(new_n407), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n457), .A2(KEYINPUT36), .A3(new_n459), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT79), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(new_n476), .A3(new_n467), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n240), .B1(new_n260), .B2(new_n248), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n275), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  OR2_X1    g279(.A1(new_n478), .A2(new_n479), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n227), .B(new_n240), .C1(new_n238), .C2(new_n215), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n482), .B(KEYINPUT80), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n480), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n484), .A2(KEYINPUT40), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT40), .ZN(new_n486));
  OAI211_X1 g285(.A(new_n486), .B(new_n480), .C1(new_n481), .C2(new_n483), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(new_n266), .A2(new_n276), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n488), .A2(new_n440), .A3(new_n489), .ZN(new_n490));
  AND3_X1   g289(.A1(new_n421), .A2(KEYINPUT37), .A3(new_n434), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT37), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n429), .A2(new_n432), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n425), .ZN(new_n494));
  OAI21_X1  g293(.A(KEYINPUT38), .B1(new_n491), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(new_n494), .A2(KEYINPUT38), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n409), .B1(new_n430), .B2(new_n431), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT83), .ZN(new_n498));
  AOI21_X1  g297(.A(new_n492), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT84), .ZN(new_n500));
  NAND3_X1  g299(.A1(new_n414), .A2(new_n409), .A3(new_n416), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n310), .B1(new_n418), .B2(new_n419), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT83), .ZN(new_n503));
  AND3_X1   g302(.A1(new_n499), .A2(new_n500), .A3(new_n503), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n500), .B1(new_n499), .B2(new_n503), .ZN(new_n505));
  OAI21_X1  g304(.A(new_n496), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n495), .A2(new_n506), .A3(new_n437), .ZN(new_n507));
  OAI211_X1 g306(.A(new_n335), .B(new_n490), .C1(new_n283), .C2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n472), .A2(new_n477), .A3(new_n508), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n466), .A2(new_n509), .A3(KEYINPUT86), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT86), .B1(new_n466), .B2(new_n509), .ZN(new_n511));
  XNOR2_X1  g310(.A(G15gat), .B(G22gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT92), .ZN(new_n513));
  INV_X1    g312(.A(G1gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(KEYINPUT92), .A3(G1gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT16), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n512), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n519), .A2(G8gat), .ZN(new_n520));
  INV_X1    g319(.A(G8gat), .ZN(new_n521));
  NAND4_X1  g320(.A1(new_n515), .A2(new_n521), .A3(new_n516), .A4(new_n518), .ZN(new_n522));
  AND2_X1   g321(.A1(new_n520), .A2(new_n522), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n329), .A2(G43gat), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n524), .A2(KEYINPUT90), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(KEYINPUT90), .ZN(new_n526));
  INV_X1    g325(.A(G43gat), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n525), .B(new_n526), .C1(new_n527), .C2(G50gat), .ZN(new_n528));
  XOR2_X1   g327(.A(KEYINPUT88), .B(G29gat), .Z(new_n529));
  OAI21_X1  g328(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n530));
  OR3_X1    g329(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n531));
  AOI22_X1  g330(.A1(new_n529), .A2(G36gat), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT15), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n532), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n527), .A2(G50gat), .ZN(new_n536));
  OR3_X1    g335(.A1(new_n524), .A2(new_n536), .A3(new_n533), .ZN(new_n537));
  AND3_X1   g336(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n537), .B1(new_n532), .B2(new_n535), .ZN(new_n539));
  OAI21_X1  g338(.A(new_n534), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n523), .A2(new_n540), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n532), .A2(new_n535), .ZN(new_n542));
  INV_X1    g341(.A(new_n537), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n529), .A2(G36gat), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n531), .A2(new_n530), .ZN(new_n547));
  AND3_X1   g346(.A1(new_n546), .A2(new_n533), .A3(new_n547), .ZN(new_n548));
  AOI22_X1  g347(.A1(new_n544), .A2(new_n545), .B1(new_n528), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n520), .A2(new_n522), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT93), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n541), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n549), .A2(KEYINPUT93), .A3(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(G229gat), .A2(G233gat), .ZN(new_n555));
  XOR2_X1   g354(.A(new_n555), .B(KEYINPUT13), .Z(new_n556));
  AND3_X1   g355(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n558), .B1(new_n540), .B2(KEYINPUT91), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n544), .A2(new_n545), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n561));
  NAND4_X1  g360(.A1(new_n560), .A2(new_n561), .A3(KEYINPUT17), .A4(new_n534), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(new_n523), .ZN(new_n564));
  NAND3_X1  g363(.A1(new_n564), .A2(new_n555), .A3(new_n551), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT18), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n557), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  XNOR2_X1  g366(.A(G113gat), .B(G141gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(G197gat), .ZN(new_n569));
  XOR2_X1   g368(.A(KEYINPUT11), .B(G169gat), .Z(new_n570));
  XNOR2_X1  g369(.A(new_n569), .B(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(KEYINPUT87), .B(KEYINPUT12), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n571), .B(new_n572), .ZN(new_n573));
  NAND4_X1  g372(.A1(new_n564), .A2(KEYINPUT18), .A3(new_n555), .A4(new_n551), .ZN(new_n574));
  AND3_X1   g373(.A1(new_n567), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n573), .B1(new_n567), .B2(new_n574), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NOR3_X1   g376(.A1(new_n510), .A2(new_n511), .A3(new_n577), .ZN(new_n578));
  XOR2_X1   g377(.A(G57gat), .B(G64gat), .Z(new_n579));
  INV_X1    g378(.A(KEYINPUT9), .ZN(new_n580));
  INV_X1    g379(.A(G71gat), .ZN(new_n581));
  INV_X1    g380(.A(G78gat), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n579), .A2(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G71gat), .B(G78gat), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(new_n585), .A3(new_n583), .ZN(new_n588));
  AND3_X1   g387(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(KEYINPUT94), .B1(new_n587), .B2(new_n588), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(KEYINPUT21), .ZN(new_n592));
  NAND2_X1  g391(.A1(G231gat), .A2(G233gat), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g393(.A(new_n593), .B1(new_n591), .B2(new_n592), .ZN(new_n595));
  NOR2_X1   g394(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G127gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g398(.A(new_n523), .B1(new_n591), .B2(new_n592), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT95), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n596), .A2(new_n597), .ZN(new_n603));
  NAND3_X1  g402(.A1(new_n599), .A2(new_n602), .A3(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n603), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n601), .B1(new_n605), .B2(new_n598), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n604), .A2(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n608));
  INV_X1    g407(.A(G155gat), .ZN(new_n609));
  XNOR2_X1  g408(.A(new_n608), .B(new_n609), .ZN(new_n610));
  XNOR2_X1  g409(.A(G183gat), .B(G211gat), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n610), .B(new_n611), .Z(new_n612));
  INV_X1    g411(.A(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n607), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n604), .A2(new_n606), .A3(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n590), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n587), .A2(KEYINPUT94), .A3(new_n588), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G85gat), .A2(G92gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n620), .B(KEYINPUT7), .ZN(new_n621));
  NAND2_X1  g420(.A1(G99gat), .A2(G106gat), .ZN(new_n622));
  INV_X1    g421(.A(G85gat), .ZN(new_n623));
  INV_X1    g422(.A(G92gat), .ZN(new_n624));
  AOI22_X1  g423(.A1(KEYINPUT8), .A2(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  XOR2_X1   g425(.A(G99gat), .B(G106gat), .Z(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n627), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n629), .A2(new_n621), .A3(new_n625), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  INV_X1    g430(.A(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n619), .A2(KEYINPUT10), .A3(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n587), .A2(new_n588), .ZN(new_n634));
  AND3_X1   g433(.A1(new_n634), .A2(new_n630), .A3(new_n628), .ZN(new_n635));
  AOI21_X1  g434(.A(new_n635), .B1(new_n619), .B2(new_n631), .ZN(new_n636));
  XNOR2_X1  g435(.A(KEYINPUT97), .B(KEYINPUT10), .ZN(new_n637));
  OAI211_X1 g436(.A(KEYINPUT98), .B(new_n633), .C1(new_n636), .C2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(KEYINPUT98), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n631), .B1(new_n589), .B2(new_n590), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n632), .A2(new_n634), .ZN(new_n641));
  AOI21_X1  g440(.A(new_n637), .B1(new_n640), .B2(new_n641), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n632), .A2(KEYINPUT10), .ZN(new_n643));
  NOR2_X1   g442(.A1(new_n643), .A2(new_n591), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n639), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(G230gat), .A2(G233gat), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n638), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  XNOR2_X1  g446(.A(G120gat), .B(G148gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(G176gat), .B(G204gat), .ZN(new_n649));
  XOR2_X1   g448(.A(new_n648), .B(new_n649), .Z(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(new_n646), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n651), .B1(new_n636), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n647), .A2(new_n653), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n646), .B1(new_n642), .B2(new_n644), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n652), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  AOI21_X1  g456(.A(KEYINPUT99), .B1(new_n657), .B2(new_n651), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT99), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n659), .B(new_n650), .C1(new_n655), .C2(new_n656), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n654), .B1(new_n658), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n563), .A2(new_n631), .ZN(new_n662));
  XNOR2_X1  g461(.A(G190gat), .B(G218gat), .ZN(new_n663));
  XOR2_X1   g462(.A(new_n663), .B(KEYINPUT96), .Z(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AND2_X1   g464(.A1(G232gat), .A2(G233gat), .ZN(new_n666));
  AOI22_X1  g465(.A1(new_n549), .A2(new_n632), .B1(KEYINPUT41), .B2(new_n666), .ZN(new_n667));
  NAND3_X1  g466(.A1(new_n662), .A2(new_n665), .A3(new_n667), .ZN(new_n668));
  AOI21_X1  g467(.A(new_n632), .B1(new_n559), .B2(new_n562), .ZN(new_n669));
  INV_X1    g468(.A(new_n667), .ZN(new_n670));
  OAI21_X1  g469(.A(new_n664), .B1(new_n669), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g471(.A1(new_n666), .A2(KEYINPUT41), .ZN(new_n673));
  XNOR2_X1  g472(.A(G134gat), .B(G162gat), .ZN(new_n674));
  XNOR2_X1  g473(.A(new_n673), .B(new_n674), .ZN(new_n675));
  INV_X1    g474(.A(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n672), .A2(new_n676), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n668), .A2(new_n675), .A3(new_n671), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n616), .A2(new_n661), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n578), .A2(new_n680), .ZN(new_n681));
  NOR2_X1   g480(.A1(new_n681), .A2(new_n445), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(new_n514), .ZN(G1324gat));
  INV_X1    g482(.A(new_n681), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n521), .B1(new_n684), .B2(new_n440), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT16), .B(G8gat), .ZN(new_n686));
  NOR3_X1   g485(.A1(new_n681), .A2(new_n446), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT42), .B1(new_n685), .B2(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(new_n688), .B1(new_n687), .B2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g488(.A(new_n408), .ZN(new_n690));
  OR3_X1    g489(.A1(new_n681), .A2(G15gat), .A3(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(G15gat), .B1(new_n681), .B2(new_n475), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n691), .A2(new_n692), .ZN(G1326gat));
  INV_X1    g492(.A(new_n335), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n684), .A2(KEYINPUT100), .A3(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT100), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(new_n681), .B2(new_n335), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g497(.A(KEYINPUT43), .B(G22gat), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n698), .B(new_n699), .ZN(G1327gat));
  NAND2_X1  g499(.A1(new_n466), .A2(new_n509), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT86), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n466), .A2(new_n509), .A3(KEYINPUT86), .ZN(new_n704));
  INV_X1    g503(.A(new_n577), .ZN(new_n705));
  INV_X1    g504(.A(new_n616), .ZN(new_n706));
  INV_X1    g505(.A(new_n679), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n706), .A2(new_n661), .A3(new_n707), .ZN(new_n708));
  NAND4_X1  g507(.A1(new_n703), .A2(new_n704), .A3(new_n705), .A4(new_n708), .ZN(new_n709));
  NOR3_X1   g508(.A1(new_n709), .A2(new_n445), .A3(new_n529), .ZN(new_n710));
  XOR2_X1   g509(.A(new_n710), .B(KEYINPUT45), .Z(new_n711));
  NAND4_X1  g510(.A1(new_n703), .A2(KEYINPUT44), .A3(new_n704), .A4(new_n679), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n508), .A2(new_n467), .A3(new_n475), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n707), .B1(new_n466), .B2(new_n713), .ZN(new_n714));
  OR2_X1    g513(.A1(new_n714), .A2(KEYINPUT44), .ZN(new_n715));
  AND2_X1   g514(.A1(new_n712), .A2(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT101), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n616), .A2(new_n717), .ZN(new_n718));
  AOI21_X1  g517(.A(KEYINPUT101), .B1(new_n614), .B2(new_n615), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n577), .A3(new_n661), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n716), .A2(new_n444), .A3(new_n721), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n722), .A2(new_n529), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n711), .A2(new_n723), .ZN(G1328gat));
  INV_X1    g523(.A(KEYINPUT104), .ZN(new_n725));
  NAND4_X1  g524(.A1(new_n712), .A2(new_n715), .A3(new_n440), .A4(new_n721), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G36gat), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n446), .A2(G36gat), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g528(.A1(new_n709), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(KEYINPUT46), .ZN(new_n731));
  AOI21_X1  g530(.A(KEYINPUT103), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT103), .ZN(new_n733));
  NOR4_X1   g532(.A1(new_n709), .A2(new_n733), .A3(KEYINPUT46), .A4(new_n729), .ZN(new_n734));
  OAI21_X1  g533(.A(new_n727), .B1(new_n732), .B2(new_n734), .ZN(new_n735));
  INV_X1    g534(.A(KEYINPUT102), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n510), .A2(new_n511), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n737), .A2(new_n705), .A3(new_n708), .A4(new_n728), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n736), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n739));
  OAI211_X1 g538(.A(new_n736), .B(KEYINPUT46), .C1(new_n709), .C2(new_n729), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g540(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n725), .B1(new_n735), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g542(.A(KEYINPUT102), .B1(new_n730), .B2(new_n731), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n744), .A2(new_n740), .ZN(new_n745));
  OAI21_X1  g544(.A(new_n733), .B1(new_n738), .B2(KEYINPUT46), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n730), .A2(KEYINPUT103), .A3(new_n731), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND4_X1  g547(.A1(new_n745), .A2(new_n748), .A3(KEYINPUT104), .A4(new_n727), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n743), .A2(new_n749), .ZN(G1329gat));
  NOR3_X1   g549(.A1(new_n709), .A2(G43gat), .A3(new_n690), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT47), .ZN(new_n752));
  AOI21_X1  g551(.A(new_n751), .B1(KEYINPUT105), .B2(new_n752), .ZN(new_n753));
  OR2_X1    g552(.A1(new_n752), .A2(KEYINPUT105), .ZN(new_n754));
  INV_X1    g553(.A(new_n475), .ZN(new_n755));
  NAND4_X1  g554(.A1(new_n712), .A2(new_n715), .A3(new_n755), .A4(new_n721), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(G43gat), .ZN(new_n757));
  AND3_X1   g556(.A1(new_n753), .A2(new_n754), .A3(new_n757), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n754), .B1(new_n753), .B2(new_n757), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n758), .A2(new_n759), .ZN(G1330gat));
  NAND4_X1  g559(.A1(new_n712), .A2(new_n715), .A3(new_n694), .A4(new_n721), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(G50gat), .ZN(new_n762));
  AOI21_X1  g561(.A(KEYINPUT48), .B1(new_n762), .B2(KEYINPUT107), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n335), .A2(G50gat), .ZN(new_n764));
  XOR2_X1   g563(.A(new_n764), .B(KEYINPUT106), .Z(new_n765));
  OAI21_X1  g564(.A(new_n762), .B1(new_n709), .B2(new_n765), .ZN(new_n766));
  XNOR2_X1  g565(.A(new_n763), .B(new_n766), .ZN(G1331gat));
  NOR2_X1   g566(.A1(new_n616), .A2(new_n679), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n768), .A2(new_n577), .A3(new_n661), .ZN(new_n769));
  XOR2_X1   g568(.A(new_n769), .B(KEYINPUT108), .Z(new_n770));
  NAND2_X1  g569(.A1(new_n466), .A2(new_n713), .ZN(new_n771));
  AND2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(new_n444), .ZN(new_n773));
  XNOR2_X1  g572(.A(new_n773), .B(G57gat), .ZN(G1332gat));
  AOI21_X1  g573(.A(new_n446), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n772), .A2(new_n775), .ZN(new_n776));
  NOR2_X1   g575(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n777));
  XOR2_X1   g576(.A(new_n776), .B(new_n777), .Z(G1333gat));
  NAND2_X1  g577(.A1(new_n770), .A2(new_n771), .ZN(new_n779));
  OAI21_X1  g578(.A(G71gat), .B1(new_n779), .B2(new_n475), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n408), .A2(new_n581), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n780), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  XOR2_X1   g581(.A(new_n782), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g582(.A1(new_n779), .A2(new_n335), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(new_n582), .ZN(G1335gat));
  INV_X1    g584(.A(new_n661), .ZN(new_n786));
  NOR3_X1   g585(.A1(new_n706), .A2(new_n705), .A3(new_n786), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n716), .A2(new_n444), .A3(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G85gat), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n706), .A2(new_n705), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n714), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT51), .ZN(new_n792));
  AOI21_X1  g591(.A(KEYINPUT110), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT110), .ZN(new_n794));
  AOI211_X1 g593(.A(new_n794), .B(KEYINPUT51), .C1(new_n714), .C2(new_n790), .ZN(new_n795));
  NOR2_X1   g594(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  NAND4_X1  g595(.A1(new_n771), .A2(KEYINPUT51), .A3(new_n679), .A4(new_n790), .ZN(new_n797));
  XNOR2_X1  g596(.A(new_n797), .B(KEYINPUT109), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n661), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n444), .A2(new_n623), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n789), .B1(new_n799), .B2(new_n800), .ZN(G1336gat));
  NAND3_X1  g600(.A1(new_n716), .A2(new_n440), .A3(new_n787), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(G92gat), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT52), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g604(.A1(new_n661), .A2(new_n624), .A3(new_n440), .ZN(new_n806));
  INV_X1    g605(.A(new_n796), .ZN(new_n807));
  INV_X1    g606(.A(new_n798), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n791), .A2(new_n792), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n806), .B1(new_n810), .B2(new_n797), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n811), .B1(new_n802), .B2(G92gat), .ZN(new_n812));
  OAI22_X1  g611(.A1(new_n805), .A2(new_n809), .B1(new_n812), .B2(new_n804), .ZN(G1337gat));
  NOR2_X1   g612(.A1(new_n690), .A2(G99gat), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n661), .B(new_n814), .C1(new_n796), .C2(new_n798), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n712), .A2(new_n715), .A3(new_n755), .A4(new_n787), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(G99gat), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT111), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n815), .A2(KEYINPUT111), .A3(new_n817), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1338gat));
  NAND3_X1  g621(.A1(new_n716), .A2(new_n694), .A3(new_n787), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n823), .A2(G106gat), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT53), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  NOR3_X1   g625(.A1(new_n786), .A2(new_n335), .A3(G106gat), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT112), .Z(new_n828));
  AOI21_X1  g627(.A(new_n828), .B1(new_n807), .B2(new_n808), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n810), .B2(new_n797), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n830), .B1(new_n823), .B2(G106gat), .ZN(new_n831));
  OAI22_X1  g630(.A1(new_n826), .A2(new_n829), .B1(new_n831), .B2(new_n825), .ZN(G1339gat));
  NAND3_X1  g631(.A1(new_n768), .A2(new_n577), .A3(new_n786), .ZN(new_n833));
  AND2_X1   g632(.A1(new_n647), .A2(new_n653), .ZN(new_n834));
  OAI21_X1  g633(.A(new_n651), .B1(new_n655), .B2(KEYINPUT54), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT54), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n642), .A2(new_n644), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n836), .B1(new_n837), .B2(new_n652), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n835), .B1(new_n647), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n834), .B1(new_n839), .B2(KEYINPUT55), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT55), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n647), .A2(new_n838), .ZN(new_n842));
  OAI21_X1  g641(.A(new_n841), .B1(new_n842), .B2(new_n835), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n840), .A2(new_n679), .A3(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n555), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n550), .B1(new_n559), .B2(new_n562), .ZN(new_n846));
  INV_X1    g645(.A(new_n551), .ZN(new_n847));
  OAI21_X1  g646(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n848), .A2(KEYINPUT113), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT113), .ZN(new_n850));
  OAI211_X1 g649(.A(new_n850), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n553), .A2(new_n554), .ZN(new_n852));
  INV_X1    g651(.A(new_n556), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n849), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(new_n571), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n567), .A2(new_n573), .A3(new_n574), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  NOR2_X1   g657(.A1(new_n844), .A2(new_n858), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n840), .B(new_n843), .C1(new_n575), .C2(new_n576), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n856), .A2(new_n857), .A3(new_n661), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n859), .B1(new_n862), .B2(new_n707), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n833), .B1(new_n863), .B2(new_n720), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n864), .A2(new_n444), .ZN(new_n865));
  AND2_X1   g664(.A1(new_n462), .A2(new_n463), .ZN(new_n866));
  NOR2_X1   g665(.A1(new_n866), .A2(new_n440), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n869), .A2(new_n222), .A3(new_n705), .ZN(new_n870));
  AND2_X1   g669(.A1(new_n864), .A2(new_n335), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n445), .A2(new_n440), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n871), .A2(new_n408), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G113gat), .B1(new_n873), .B2(new_n577), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n870), .A2(new_n874), .ZN(new_n875));
  XNOR2_X1  g674(.A(new_n875), .B(KEYINPUT114), .ZN(G1340gat));
  OAI21_X1  g675(.A(G120gat), .B1(new_n873), .B2(new_n786), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n661), .A2(new_n225), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT115), .Z(new_n879));
  OAI21_X1  g678(.A(new_n877), .B1(new_n868), .B2(new_n879), .ZN(G1341gat));
  NAND3_X1  g679(.A1(new_n869), .A2(new_n597), .A3(new_n706), .ZN(new_n881));
  INV_X1    g680(.A(new_n720), .ZN(new_n882));
  OAI21_X1  g681(.A(G127gat), .B1(new_n873), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n881), .A2(new_n883), .ZN(G1342gat));
  OR3_X1    g683(.A1(new_n868), .A2(G134gat), .A3(new_n707), .ZN(new_n885));
  XNOR2_X1  g684(.A(KEYINPUT116), .B(KEYINPUT56), .ZN(new_n886));
  OR2_X1    g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  OAI21_X1  g687(.A(G134gat), .B1(new_n873), .B2(new_n707), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G1343gat));
  NAND2_X1  g689(.A1(new_n864), .A2(new_n694), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n475), .B(new_n872), .C1(new_n891), .C2(KEYINPUT57), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n894));
  XOR2_X1   g693(.A(KEYINPUT118), .B(KEYINPUT55), .Z(new_n895));
  OAI21_X1  g694(.A(new_n895), .B1(new_n842), .B2(new_n835), .ZN(new_n896));
  OAI211_X1 g695(.A(new_n840), .B(new_n896), .C1(new_n575), .C2(new_n576), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n898));
  NAND4_X1  g697(.A1(new_n856), .A2(new_n857), .A3(new_n661), .A4(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n894), .A2(new_n897), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n859), .B1(new_n900), .B2(new_n707), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n833), .B1(new_n901), .B2(new_n706), .ZN(new_n902));
  AOI21_X1  g701(.A(new_n893), .B1(new_n902), .B2(new_n694), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n892), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n205), .B1(new_n904), .B2(new_n705), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n755), .A2(new_n335), .A3(new_n440), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n865), .A2(new_n906), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n907), .A2(G141gat), .A3(new_n577), .ZN(new_n908));
  OR3_X1    g707(.A1(new_n905), .A2(KEYINPUT58), .A3(new_n908), .ZN(new_n909));
  OAI21_X1  g708(.A(KEYINPUT58), .B1(new_n905), .B2(new_n908), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n909), .A2(new_n910), .ZN(G1344gat));
  NAND2_X1  g710(.A1(new_n661), .A2(new_n206), .ZN(new_n912));
  NOR2_X1   g711(.A1(new_n907), .A2(new_n912), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT119), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n902), .A2(new_n893), .A3(new_n694), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n475), .A2(new_n661), .A3(new_n872), .ZN(new_n917));
  AND3_X1   g716(.A1(new_n915), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  NAND2_X1  g717(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n206), .B1(new_n904), .B2(new_n661), .ZN(new_n920));
  OAI221_X1 g719(.A(new_n914), .B1(new_n918), .B2(new_n919), .C1(new_n920), .C2(KEYINPUT59), .ZN(G1345gat));
  INV_X1    g720(.A(new_n907), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n922), .A2(new_n609), .A3(new_n706), .ZN(new_n923));
  NOR3_X1   g722(.A1(new_n892), .A2(new_n882), .A3(new_n903), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n923), .B1(new_n924), .B2(new_n609), .ZN(G1346gat));
  AOI21_X1  g724(.A(G162gat), .B1(new_n922), .B2(new_n679), .ZN(new_n926));
  AND2_X1   g725(.A1(new_n679), .A2(G162gat), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n926), .B1(new_n904), .B2(new_n927), .ZN(G1347gat));
  AND2_X1   g727(.A1(new_n864), .A2(new_n445), .ZN(new_n929));
  NOR2_X1   g728(.A1(new_n866), .A2(new_n446), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT120), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT120), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(new_n933), .A3(new_n930), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n577), .A2(G169gat), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n932), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  INV_X1    g735(.A(KEYINPUT121), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n936), .B(new_n937), .ZN(new_n938));
  NOR2_X1   g737(.A1(new_n446), .A2(new_n444), .ZN(new_n939));
  INV_X1    g738(.A(new_n939), .ZN(new_n940));
  NOR2_X1   g739(.A1(new_n940), .A2(new_n690), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT122), .B1(new_n871), .B2(new_n941), .ZN(new_n942));
  INV_X1    g741(.A(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n941), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI21_X1  g744(.A(G169gat), .B1(new_n945), .B2(new_n577), .ZN(new_n946));
  INV_X1    g745(.A(KEYINPUT123), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  OAI211_X1 g747(.A(KEYINPUT123), .B(G169gat), .C1(new_n945), .C2(new_n577), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n938), .A2(new_n948), .A3(new_n949), .ZN(G1348gat));
  AND3_X1   g749(.A1(new_n871), .A2(KEYINPUT122), .A3(new_n941), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n951), .A2(new_n942), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n786), .A2(new_n338), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n952), .A2(KEYINPUT124), .A3(new_n953), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n932), .A2(new_n661), .A3(new_n934), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n955), .A2(new_n338), .ZN(new_n956));
  AOI21_X1  g755(.A(KEYINPUT124), .B1(new_n952), .B2(new_n953), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n954), .A2(new_n956), .A3(new_n957), .ZN(G1349gat));
  AOI21_X1  g757(.A(new_n346), .B1(new_n952), .B2(new_n720), .ZN(new_n959));
  NAND4_X1  g758(.A1(new_n929), .A2(new_n353), .A3(new_n706), .A4(new_n930), .ZN(new_n960));
  INV_X1    g759(.A(new_n960), .ZN(new_n961));
  OAI21_X1  g760(.A(KEYINPUT60), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(G183gat), .B1(new_n945), .B2(new_n882), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n963), .A2(new_n964), .A3(new_n960), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n962), .A2(new_n965), .ZN(G1350gat));
  NOR2_X1   g765(.A1(new_n707), .A2(G190gat), .ZN(new_n967));
  NAND3_X1  g766(.A1(new_n932), .A2(new_n934), .A3(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT125), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n968), .B(new_n969), .ZN(new_n970));
  OAI21_X1  g769(.A(G190gat), .B1(new_n945), .B2(new_n707), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT61), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  OAI211_X1 g772(.A(KEYINPUT61), .B(G190gat), .C1(new_n945), .C2(new_n707), .ZN(new_n974));
  NAND3_X1  g773(.A1(new_n970), .A2(new_n973), .A3(new_n974), .ZN(G1351gat));
  NOR2_X1   g774(.A1(new_n755), .A2(new_n940), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n915), .A2(new_n916), .A3(new_n976), .ZN(new_n977));
  NOR3_X1   g776(.A1(new_n977), .A2(new_n289), .A3(new_n577), .ZN(new_n978));
  NOR3_X1   g777(.A1(new_n755), .A2(new_n335), .A3(new_n446), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n929), .A2(new_n979), .ZN(new_n980));
  INV_X1    g779(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g780(.A(G197gat), .B1(new_n981), .B2(new_n705), .ZN(new_n982));
  NOR2_X1   g781(.A1(new_n978), .A2(new_n982), .ZN(G1352gat));
  NOR3_X1   g782(.A1(new_n980), .A2(G204gat), .A3(new_n786), .ZN(new_n984));
  XNOR2_X1  g783(.A(new_n984), .B(KEYINPUT62), .ZN(new_n985));
  OAI21_X1  g784(.A(G204gat), .B1(new_n977), .B2(new_n786), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n985), .A2(new_n986), .ZN(G1353gat));
  OR3_X1    g786(.A1(new_n980), .A2(G211gat), .A3(new_n616), .ZN(new_n988));
  NAND4_X1  g787(.A1(new_n915), .A2(new_n706), .A3(new_n916), .A4(new_n976), .ZN(new_n989));
  AND3_X1   g788(.A1(new_n989), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n990));
  AOI21_X1  g789(.A(KEYINPUT63), .B1(new_n989), .B2(G211gat), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n988), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT126), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  OAI211_X1 g793(.A(KEYINPUT126), .B(new_n988), .C1(new_n990), .C2(new_n991), .ZN(new_n995));
  NAND2_X1  g794(.A1(new_n994), .A2(new_n995), .ZN(G1354gat));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n679), .ZN(new_n998));
  INV_X1    g797(.A(G218gat), .ZN(new_n999));
  AOI21_X1  g798(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI211_X1 g799(.A(KEYINPUT127), .B(G218gat), .C1(new_n981), .C2(new_n679), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n977), .A2(new_n999), .A3(new_n707), .ZN(new_n1002));
  NOR3_X1   g801(.A1(new_n1000), .A2(new_n1001), .A3(new_n1002), .ZN(G1355gat));
endmodule


