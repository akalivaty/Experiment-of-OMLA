//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 0 0 1 0 0 0 1 1 1 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 1 0 1 1 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 1 1 1 1 1 0 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:33 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n826, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n962, new_n963, new_n964, new_n965, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n990, new_n991, new_n992,
    new_n993, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1028, new_n1029, new_n1030, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(new_n187), .ZN(new_n188));
  INV_X1    g002(.A(G101), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT77), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n190), .A2(new_n191), .A3(new_n192), .A4(G104), .ZN(new_n193));
  INV_X1    g007(.A(G104), .ZN(new_n194));
  NOR3_X1   g008(.A1(new_n194), .A2(KEYINPUT77), .A3(G107), .ZN(new_n195));
  AOI21_X1  g009(.A(KEYINPUT3), .B1(new_n194), .B2(G107), .ZN(new_n196));
  OAI211_X1 g010(.A(new_n189), .B(new_n193), .C1(new_n195), .C2(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n192), .A2(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n194), .A2(G107), .ZN(new_n199));
  OAI21_X1  g013(.A(G101), .B1(new_n198), .B2(new_n199), .ZN(new_n200));
  AND2_X1   g014(.A1(new_n197), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G113), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT2), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n204), .A2(G113), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G116), .ZN(new_n208));
  INV_X1    g022(.A(G116), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G119), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n209), .A2(G119), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT5), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n208), .A2(new_n210), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n214), .B(G113), .C1(new_n215), .C2(new_n213), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n201), .A2(KEYINPUT84), .A3(new_n211), .A4(new_n216), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n216), .A2(new_n197), .A3(new_n211), .A4(new_n200), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT84), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(new_n191), .B1(new_n192), .B2(G104), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n190), .A2(new_n192), .A3(G104), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  AOI21_X1  g038(.A(new_n189), .B1(new_n224), .B2(new_n193), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT4), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n215), .A2(new_n203), .A3(new_n205), .ZN(new_n227));
  AOI22_X1  g041(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n211), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT83), .ZN(new_n229));
  OAI21_X1  g043(.A(new_n193), .B1(new_n195), .B2(new_n196), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n230), .A2(G101), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n231), .A2(KEYINPUT4), .A3(new_n197), .ZN(new_n232));
  AND3_X1   g046(.A1(new_n228), .A2(new_n229), .A3(new_n232), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n229), .B1(new_n228), .B2(new_n232), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n221), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(G110), .B(G122), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n235), .A2(new_n237), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n221), .B(new_n236), .C1(new_n233), .C2(new_n234), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT6), .ZN(new_n240));
  NOR2_X1   g054(.A1(new_n240), .A2(KEYINPUT85), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n238), .A2(new_n239), .A3(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G143), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT1), .B1(new_n243), .B2(G146), .ZN(new_n244));
  NOR2_X1   g058(.A1(new_n243), .A2(G146), .ZN(new_n245));
  INV_X1    g059(.A(G146), .ZN(new_n246));
  NOR2_X1   g060(.A1(new_n246), .A2(G143), .ZN(new_n247));
  OAI211_X1 g061(.A(G128), .B(new_n244), .C1(new_n245), .C2(new_n247), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n246), .A2(G143), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(G146), .ZN(new_n250));
  INV_X1    g064(.A(G128), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n249), .B(new_n250), .C1(KEYINPUT1), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n248), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(G125), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT0), .ZN(new_n256));
  OAI211_X1 g070(.A(new_n249), .B(new_n250), .C1(new_n256), .C2(new_n251), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n256), .A2(new_n251), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT0), .A2(G128), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G143), .B(G146), .ZN(new_n261));
  OAI211_X1 g075(.A(new_n257), .B(G125), .C1(new_n260), .C2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n255), .A2(new_n262), .ZN(new_n263));
  INV_X1    g077(.A(G224), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n264), .A2(G953), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n265), .B(KEYINPUT86), .ZN(new_n266));
  XNOR2_X1  g080(.A(new_n263), .B(new_n266), .ZN(new_n267));
  OAI211_X1 g081(.A(new_n235), .B(new_n237), .C1(KEYINPUT85), .C2(new_n240), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n242), .A2(new_n267), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g083(.A(KEYINPUT7), .B1(new_n264), .B2(G953), .ZN(new_n270));
  INV_X1    g084(.A(new_n262), .ZN(new_n271));
  AOI21_X1  g085(.A(G125), .B1(new_n248), .B2(new_n252), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n270), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n270), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n255), .A2(new_n262), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(G110), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n277), .A2(G122), .ZN(new_n278));
  INV_X1    g092(.A(G122), .ZN(new_n279));
  NOR2_X1   g093(.A1(new_n279), .A2(G110), .ZN(new_n280));
  NOR3_X1   g094(.A1(new_n278), .A2(new_n280), .A3(KEYINPUT87), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n279), .A2(G110), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n277), .A2(G122), .ZN(new_n284));
  AOI21_X1  g098(.A(new_n282), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(KEYINPUT8), .B1(new_n281), .B2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n236), .A2(new_n282), .ZN(new_n287));
  OAI21_X1  g101(.A(KEYINPUT87), .B1(new_n278), .B2(new_n280), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT8), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n287), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n286), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g105(.A1(new_n216), .A2(new_n211), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n197), .A2(new_n200), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n291), .B1(new_n294), .B2(new_n218), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n276), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n239), .A2(new_n296), .ZN(new_n297));
  INV_X1    g111(.A(G902), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(KEYINPUT88), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT88), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n297), .A2(new_n301), .A3(new_n298), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n269), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G210), .B1(G237), .B2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n307));
  AOI211_X1 g121(.A(KEYINPUT88), .B(G902), .C1(new_n239), .C2(new_n296), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n309), .A2(new_n304), .A3(new_n269), .ZN(new_n310));
  AOI21_X1  g124(.A(new_n188), .B1(new_n306), .B2(new_n310), .ZN(new_n311));
  INV_X1    g125(.A(G475), .ZN(new_n312));
  INV_X1    g126(.A(KEYINPUT89), .ZN(new_n313));
  INV_X1    g127(.A(G953), .ZN(new_n314));
  AND2_X1   g128(.A1(KEYINPUT65), .A2(G237), .ZN(new_n315));
  NOR2_X1   g129(.A1(KEYINPUT65), .A2(G237), .ZN(new_n316));
  OAI211_X1 g130(.A(G214), .B(new_n314), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n313), .B1(new_n317), .B2(new_n243), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT65), .ZN(new_n319));
  INV_X1    g133(.A(G237), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(KEYINPUT65), .A2(G237), .ZN(new_n322));
  AOI21_X1  g136(.A(G953), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(KEYINPUT89), .A3(G143), .A4(G214), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n318), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n317), .A2(new_n243), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n327), .A2(G131), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n329));
  AOI22_X1  g143(.A1(new_n318), .A2(new_n324), .B1(new_n243), .B2(new_n317), .ZN(new_n330));
  INV_X1    g144(.A(G131), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NAND3_X1  g146(.A1(new_n328), .A2(new_n329), .A3(new_n332), .ZN(new_n333));
  NOR3_X1   g147(.A1(new_n254), .A2(KEYINPUT16), .A3(G140), .ZN(new_n334));
  INV_X1    g148(.A(G140), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n335), .B1(new_n254), .B2(KEYINPUT72), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT72), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n337), .A2(G125), .A3(G140), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g153(.A(new_n334), .B1(new_n339), .B2(KEYINPUT16), .ZN(new_n340));
  XNOR2_X1  g154(.A(new_n340), .B(G146), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n331), .B1(new_n325), .B2(new_n326), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n341), .B1(new_n342), .B2(KEYINPUT17), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n333), .A2(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT91), .B(G104), .ZN(new_n346));
  XNOR2_X1  g160(.A(new_n345), .B(new_n346), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n327), .A2(KEYINPUT18), .A3(G131), .ZN(new_n348));
  NOR2_X1   g162(.A1(new_n339), .A2(new_n246), .ZN(new_n349));
  XNOR2_X1  g163(.A(G125), .B(G140), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n350), .A2(KEYINPUT74), .ZN(new_n351));
  INV_X1    g165(.A(KEYINPUT74), .ZN(new_n352));
  NOR2_X1   g166(.A1(new_n254), .A2(G140), .ZN(new_n353));
  NOR2_X1   g167(.A1(new_n335), .A2(G125), .ZN(new_n354));
  OAI21_X1  g168(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n351), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n349), .B1(new_n356), .B2(new_n246), .ZN(new_n357));
  NAND2_X1  g171(.A1(KEYINPUT18), .A2(G131), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n357), .B1(new_n330), .B2(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n348), .A2(new_n359), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n344), .A2(new_n347), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n347), .B1(new_n344), .B2(new_n360), .ZN(new_n362));
  OAI21_X1  g176(.A(new_n298), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(new_n312), .B1(new_n363), .B2(KEYINPUT92), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT92), .ZN(new_n365));
  OAI211_X1 g179(.A(new_n365), .B(new_n298), .C1(new_n361), .C2(new_n362), .ZN(new_n366));
  AND2_X1   g180(.A1(new_n340), .A2(G146), .ZN(new_n367));
  AND3_X1   g181(.A1(new_n336), .A2(KEYINPUT19), .A3(new_n338), .ZN(new_n368));
  XNOR2_X1  g182(.A(KEYINPUT90), .B(KEYINPUT19), .ZN(new_n369));
  AOI21_X1  g183(.A(new_n368), .B1(new_n356), .B2(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n367), .B1(new_n370), .B2(new_n246), .ZN(new_n371));
  AND3_X1   g185(.A1(new_n325), .A2(new_n331), .A3(new_n326), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(new_n342), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n347), .B1(new_n373), .B2(new_n360), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n333), .A2(new_n343), .B1(new_n348), .B2(new_n359), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n374), .B1(new_n347), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g190(.A1(G475), .A2(G902), .ZN(new_n377));
  INV_X1    g191(.A(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT20), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT20), .ZN(new_n380));
  OAI211_X1 g194(.A(new_n380), .B(new_n377), .C1(new_n361), .C2(new_n374), .ZN(new_n381));
  AOI22_X1  g195(.A1(new_n364), .A2(new_n366), .B1(new_n379), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g196(.A1(new_n314), .A2(G952), .ZN(new_n383));
  INV_X1    g197(.A(G234), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(new_n320), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI211_X1 g200(.A(new_n298), .B(new_n314), .C1(G234), .C2(G237), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT21), .B(G898), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n389), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n209), .A2(G122), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n209), .A2(G122), .ZN(new_n392));
  OAI21_X1  g206(.A(new_n391), .B1(new_n392), .B2(KEYINPUT14), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n393), .B1(KEYINPUT14), .B2(new_n391), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(G107), .ZN(new_n395));
  XNOR2_X1  g209(.A(G116), .B(G122), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n192), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n243), .A2(G128), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n251), .A2(G143), .ZN(new_n399));
  INV_X1    g213(.A(G134), .ZN(new_n400));
  AND3_X1   g214(.A1(new_n398), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n400), .B1(new_n398), .B2(new_n399), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n395), .B(new_n397), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n398), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n404), .B1(KEYINPUT13), .B2(new_n399), .ZN(new_n405));
  AND2_X1   g219(.A1(new_n404), .A2(KEYINPUT13), .ZN(new_n406));
  OAI21_X1  g220(.A(G134), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n401), .A2(KEYINPUT93), .ZN(new_n408));
  XNOR2_X1  g222(.A(new_n396), .B(new_n192), .ZN(new_n409));
  OR2_X1    g223(.A1(new_n401), .A2(KEYINPUT93), .ZN(new_n410));
  NAND4_X1  g224(.A1(new_n407), .A2(new_n408), .A3(new_n409), .A4(new_n410), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT9), .B(G234), .ZN(new_n412));
  INV_X1    g226(.A(G217), .ZN(new_n413));
  NOR3_X1   g227(.A1(new_n412), .A2(new_n413), .A3(G953), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n403), .A2(new_n411), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n414), .B1(new_n403), .B2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n298), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G478), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT15), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g234(.A1(new_n417), .A2(new_n419), .ZN(new_n421));
  OR3_X1    g235(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT94), .ZN(new_n422));
  OAI21_X1  g236(.A(KEYINPUT94), .B1(new_n420), .B2(new_n421), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND4_X1  g238(.A1(new_n311), .A2(new_n382), .A3(new_n390), .A4(new_n424), .ZN(new_n425));
  INV_X1    g239(.A(G221), .ZN(new_n426));
  INV_X1    g240(.A(new_n412), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n427), .B2(new_n298), .ZN(new_n428));
  INV_X1    g242(.A(new_n428), .ZN(new_n429));
  INV_X1    g243(.A(G469), .ZN(new_n430));
  XNOR2_X1  g244(.A(G110), .B(G140), .ZN(new_n431));
  AND2_X1   g245(.A1(new_n314), .A2(G227), .ZN(new_n432));
  XOR2_X1   g246(.A(new_n431), .B(new_n432), .Z(new_n433));
  NAND4_X1  g247(.A1(new_n197), .A2(new_n248), .A3(new_n252), .A4(new_n200), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n435), .A2(KEYINPUT10), .ZN(new_n436));
  OAI22_X1  g250(.A1(new_n245), .A2(new_n247), .B1(new_n258), .B2(new_n259), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n257), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n230), .A2(new_n226), .A3(G101), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n232), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  INV_X1    g254(.A(KEYINPUT79), .ZN(new_n441));
  XOR2_X1   g255(.A(KEYINPUT78), .B(KEYINPUT10), .Z(new_n442));
  AND3_X1   g256(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n441), .B1(new_n434), .B2(new_n442), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n436), .B(new_n440), .C1(new_n443), .C2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT11), .ZN(new_n446));
  OAI21_X1  g260(.A(new_n446), .B1(new_n400), .B2(G137), .ZN(new_n447));
  INV_X1    g261(.A(G137), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(KEYINPUT11), .A3(G134), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n400), .A2(G137), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n447), .A2(new_n449), .A3(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n451), .A2(G131), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n447), .A2(new_n449), .A3(new_n331), .A4(new_n450), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(KEYINPUT80), .B1(new_n445), .B2(new_n454), .ZN(new_n455));
  INV_X1    g269(.A(new_n444), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n434), .A2(new_n441), .A3(new_n442), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  AND2_X1   g272(.A1(new_n439), .A2(new_n438), .ZN(new_n459));
  AOI22_X1  g273(.A1(new_n459), .A2(new_n232), .B1(new_n435), .B2(KEYINPUT10), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n461));
  INV_X1    g275(.A(new_n454), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n458), .A2(new_n460), .A3(new_n461), .A4(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  INV_X1    g278(.A(KEYINPUT81), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n465), .B1(new_n452), .B2(new_n453), .ZN(new_n466));
  AOI22_X1  g280(.A1(new_n197), .A2(new_n200), .B1(new_n248), .B2(new_n252), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n466), .B1(new_n435), .B2(new_n467), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT12), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT12), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n470), .B(new_n466), .C1(new_n435), .C2(new_n467), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n433), .B1(new_n464), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n464), .A2(new_n433), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n445), .A2(new_n454), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(new_n433), .ZN(new_n479));
  AOI21_X1  g293(.A(new_n479), .B1(new_n455), .B2(new_n463), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT82), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n478), .B1(new_n480), .B2(new_n481), .ZN(new_n482));
  AOI211_X1 g296(.A(new_n430), .B(new_n474), .C1(new_n476), .C2(new_n482), .ZN(new_n483));
  AOI21_X1  g297(.A(new_n433), .B1(new_n464), .B2(new_n477), .ZN(new_n484));
  AOI211_X1 g298(.A(new_n479), .B(new_n472), .C1(new_n455), .C2(new_n463), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n430), .B(new_n298), .C1(new_n484), .C2(new_n485), .ZN(new_n486));
  NAND2_X1  g300(.A1(G469), .A2(G902), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n429), .B1(new_n483), .B2(new_n488), .ZN(new_n489));
  NOR2_X1   g303(.A1(new_n425), .A2(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(G472), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n454), .A2(new_n438), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n227), .A2(new_n211), .ZN(new_n494));
  INV_X1    g308(.A(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT64), .ZN(new_n496));
  XNOR2_X1  g310(.A(G134), .B(G137), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n496), .B1(new_n497), .B2(new_n331), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n400), .A2(G137), .ZN(new_n499));
  NOR2_X1   g313(.A1(new_n448), .A2(G134), .ZN(new_n500));
  OAI211_X1 g314(.A(KEYINPUT64), .B(G131), .C1(new_n499), .C2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n498), .A2(new_n453), .A3(new_n501), .ZN(new_n502));
  OAI211_X1 g316(.A(new_n493), .B(new_n495), .C1(new_n253), .C2(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT28), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NOR2_X1   g320(.A1(new_n502), .A2(new_n253), .ZN(new_n507));
  AOI22_X1  g321(.A1(new_n452), .A2(new_n453), .B1(new_n437), .B2(new_n257), .ZN(new_n508));
  OAI21_X1  g322(.A(new_n494), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n503), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n510), .A2(KEYINPUT28), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n506), .B1(new_n511), .B2(KEYINPUT69), .ZN(new_n512));
  AOI211_X1 g326(.A(KEYINPUT69), .B(new_n504), .C1(new_n509), .C2(new_n503), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n323), .A2(G210), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n515), .B(KEYINPUT67), .ZN(new_n516));
  XNOR2_X1  g330(.A(KEYINPUT26), .B(G101), .ZN(new_n517));
  OR2_X1    g331(.A1(new_n517), .A2(KEYINPUT68), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n517), .A2(KEYINPUT68), .ZN(new_n519));
  XOR2_X1   g333(.A(KEYINPUT66), .B(KEYINPUT27), .Z(new_n520));
  AND3_X1   g334(.A1(new_n518), .A2(new_n519), .A3(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(new_n520), .B1(new_n518), .B2(new_n519), .ZN(new_n522));
  OR3_X1    g336(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n516), .B1(new_n521), .B2(new_n522), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n512), .A2(new_n514), .A3(new_n525), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT29), .ZN(new_n527));
  INV_X1    g341(.A(KEYINPUT30), .ZN(new_n528));
  OR2_X1    g342(.A1(new_n502), .A2(new_n253), .ZN(new_n529));
  AOI21_X1  g343(.A(new_n528), .B1(new_n529), .B2(new_n493), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n507), .A2(new_n508), .A3(KEYINPUT30), .ZN(new_n531));
  OAI21_X1  g345(.A(new_n494), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(new_n503), .ZN(new_n533));
  INV_X1    g347(.A(new_n525), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n526), .A2(new_n527), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n534), .A2(new_n527), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n504), .B1(new_n509), .B2(new_n503), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n506), .A2(new_n538), .ZN(new_n539));
  AOI21_X1  g353(.A(G902), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n492), .B1(new_n536), .B2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT69), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n505), .B1(new_n538), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n534), .B1(new_n543), .B2(new_n513), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n544), .A2(KEYINPUT70), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT70), .ZN(new_n546));
  OAI211_X1 g360(.A(new_n546), .B(new_n534), .C1(new_n543), .C2(new_n513), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n532), .A2(new_n525), .A3(new_n503), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT31), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND4_X1  g364(.A1(new_n532), .A2(new_n525), .A3(KEYINPUT31), .A4(new_n503), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n545), .A2(new_n547), .A3(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n553), .A2(new_n492), .A3(new_n298), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT32), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT32), .ZN(new_n556));
  NAND4_X1  g370(.A1(new_n553), .A2(new_n556), .A3(new_n492), .A4(new_n298), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n541), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  XNOR2_X1  g372(.A(KEYINPUT22), .B(G137), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n426), .A2(new_n384), .A3(G953), .ZN(new_n560));
  XOR2_X1   g374(.A(new_n559), .B(new_n560), .Z(new_n561));
  INV_X1    g375(.A(new_n561), .ZN(new_n562));
  OAI21_X1  g376(.A(KEYINPUT71), .B1(new_n207), .B2(G128), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT23), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n207), .A2(G128), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n251), .A2(G119), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT23), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n566), .A2(KEYINPUT71), .A3(new_n567), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n564), .A2(new_n565), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(new_n277), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n566), .A2(new_n565), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT24), .B(G110), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  OR2_X1    g388(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(KEYINPUT73), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n367), .B1(new_n246), .B2(new_n356), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n575), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  OAI221_X1 g392(.A(new_n341), .B1(new_n277), .B2(new_n569), .C1(new_n571), .C2(new_n572), .ZN(new_n579));
  AOI21_X1  g393(.A(new_n562), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g394(.A(new_n580), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n578), .A2(new_n579), .A3(new_n562), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n413), .B1(G234), .B2(new_n298), .ZN(new_n584));
  NOR2_X1   g398(.A1(new_n584), .A2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n583), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n583), .A2(new_n298), .ZN(new_n587));
  NOR2_X1   g401(.A1(KEYINPUT75), .A2(KEYINPUT25), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n584), .B1(new_n587), .B2(new_n589), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n586), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n558), .A2(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT76), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  OAI21_X1  g410(.A(KEYINPUT76), .B1(new_n558), .B2(new_n593), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n491), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  XNOR2_X1  g412(.A(new_n598), .B(new_n189), .ZN(G3));
  AND3_X1   g413(.A1(new_n553), .A2(KEYINPUT95), .A3(new_n298), .ZN(new_n600));
  AOI21_X1  g414(.A(KEYINPUT95), .B1(new_n553), .B2(new_n298), .ZN(new_n601));
  OAI21_X1  g415(.A(G472), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n554), .A2(KEYINPUT96), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  OAI211_X1 g418(.A(KEYINPUT96), .B(G472), .C1(new_n600), .C2(new_n601), .ZN(new_n605));
  NOR2_X1   g419(.A1(new_n489), .A2(new_n593), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n604), .A2(new_n605), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n379), .A2(new_n381), .ZN(new_n609));
  NOR3_X1   g423(.A1(new_n372), .A2(new_n342), .A3(KEYINPUT17), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n327), .A2(KEYINPUT17), .A3(G131), .ZN(new_n611));
  INV_X1    g425(.A(new_n341), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g427(.A(new_n360), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n347), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n375), .A2(new_n347), .ZN(new_n617));
  AOI21_X1  g431(.A(G902), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  OAI21_X1  g432(.A(G475), .B1(new_n618), .B2(new_n365), .ZN(new_n619));
  INV_X1    g433(.A(new_n366), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n609), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  INV_X1    g435(.A(new_n417), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT98), .B(G478), .Z(new_n623));
  NOR2_X1   g437(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n625));
  AND2_X1   g439(.A1(KEYINPUT97), .A2(KEYINPUT33), .ZN(new_n626));
  OR4_X1    g440(.A1(new_n415), .A2(new_n416), .A3(new_n625), .A4(new_n626), .ZN(new_n627));
  OAI211_X1 g441(.A(KEYINPUT97), .B(KEYINPUT33), .C1(new_n415), .C2(new_n416), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n418), .A2(G902), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n624), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  INV_X1    g445(.A(new_n631), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n621), .A2(new_n632), .ZN(new_n633));
  AND4_X1   g447(.A1(new_n304), .A2(new_n269), .A3(new_n300), .A4(new_n302), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n304), .B1(new_n309), .B2(new_n269), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n390), .B(new_n187), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NOR2_X1   g450(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n608), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g452(.A(new_n638), .B(KEYINPUT99), .ZN(new_n639));
  XOR2_X1   g453(.A(KEYINPUT34), .B(G104), .Z(new_n640));
  XNOR2_X1  g454(.A(new_n639), .B(new_n640), .ZN(G6));
  INV_X1    g455(.A(new_n424), .ZN(new_n642));
  NAND2_X1  g456(.A1(new_n382), .A2(new_n642), .ZN(new_n643));
  NOR2_X1   g457(.A1(new_n643), .A2(new_n636), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n608), .A2(new_n644), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n645), .B(KEYINPUT100), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n646), .B(KEYINPUT35), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G107), .ZN(G9));
  INV_X1    g462(.A(new_n584), .ZN(new_n649));
  INV_X1    g463(.A(new_n582), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n650), .A2(new_n580), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n651), .A2(G902), .ZN(new_n652));
  AOI21_X1  g466(.A(new_n649), .B1(new_n652), .B2(new_n588), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n578), .A2(new_n579), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n562), .A2(KEYINPUT36), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  AOI22_X1  g470(.A1(new_n653), .A2(new_n590), .B1(new_n585), .B2(new_n656), .ZN(new_n657));
  NOR3_X1   g471(.A1(new_n425), .A2(new_n657), .A3(new_n489), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n605), .A3(new_n604), .ZN(new_n659));
  XOR2_X1   g473(.A(KEYINPUT37), .B(G110), .Z(new_n660));
  XNOR2_X1  g474(.A(new_n659), .B(new_n660), .ZN(G12));
  NAND2_X1  g475(.A1(new_n306), .A2(new_n310), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(new_n187), .ZN(new_n663));
  NOR3_X1   g477(.A1(new_n558), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  XOR2_X1   g478(.A(KEYINPUT101), .B(G900), .Z(new_n665));
  NAND2_X1  g479(.A1(new_n387), .A2(new_n665), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n667));
  NAND2_X1  g481(.A1(new_n666), .A2(KEYINPUT102), .ZN(new_n668));
  AND3_X1   g482(.A1(new_n667), .A2(new_n385), .A3(new_n668), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n489), .A2(new_n643), .A3(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n664), .A2(new_n670), .ZN(new_n671));
  XOR2_X1   g485(.A(KEYINPUT103), .B(G128), .Z(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(G30));
  NAND2_X1  g487(.A1(new_n657), .A2(new_n187), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n621), .A2(new_n642), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n555), .A2(new_n557), .ZN(new_n677));
  INV_X1    g491(.A(new_n548), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n510), .B2(new_n534), .ZN(new_n679));
  OAI21_X1  g493(.A(G472), .B1(new_n679), .B2(G902), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n662), .B(KEYINPUT38), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n676), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  INV_X1    g497(.A(new_n489), .ZN(new_n684));
  XOR2_X1   g498(.A(new_n669), .B(KEYINPUT39), .Z(new_n685));
  NAND2_X1  g499(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OR2_X1    g500(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n686), .A2(KEYINPUT40), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n683), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G143), .ZN(G45));
  INV_X1    g504(.A(KEYINPUT104), .ZN(new_n691));
  INV_X1    g505(.A(new_n669), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n621), .A2(new_n632), .A3(new_n692), .ZN(new_n693));
  OAI21_X1  g507(.A(new_n691), .B1(new_n693), .B2(new_n663), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n363), .A2(KEYINPUT92), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n695), .A2(G475), .A3(new_n366), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n631), .B1(new_n696), .B2(new_n609), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n697), .A2(KEYINPUT104), .A3(new_n311), .A4(new_n692), .ZN(new_n698));
  AND2_X1   g512(.A1(new_n694), .A2(new_n698), .ZN(new_n699));
  NOR3_X1   g513(.A1(new_n558), .A2(new_n489), .A3(new_n657), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n701), .B(G146), .ZN(G48));
  NOR2_X1   g516(.A1(new_n484), .A2(new_n485), .ZN(new_n703));
  OAI211_X1 g517(.A(KEYINPUT105), .B(G469), .C1(new_n703), .C2(G902), .ZN(new_n704));
  OR2_X1    g518(.A1(new_n484), .A2(new_n485), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n430), .B1(new_n705), .B2(new_n298), .ZN(new_n706));
  INV_X1    g520(.A(KEYINPUT105), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n486), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(new_n704), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n709), .A2(new_n429), .ZN(new_n710));
  INV_X1    g524(.A(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n709), .A2(KEYINPUT106), .A3(new_n429), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n594), .A2(new_n712), .A3(new_n637), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n594), .A2(new_n712), .A3(new_n644), .A4(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NOR3_X1   g532(.A1(new_n621), .A2(new_n642), .A3(new_n389), .ZN(new_n719));
  INV_X1    g533(.A(new_n710), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n664), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  AOI21_X1  g536(.A(new_n492), .B1(new_n553), .B2(new_n298), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT107), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n552), .B1(new_n525), .B2(new_n539), .ZN(new_n727));
  NOR2_X1   g541(.A1(G472), .A2(G902), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  OAI21_X1  g543(.A(new_n729), .B1(new_n723), .B2(new_n724), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n726), .A2(new_n730), .A3(new_n593), .ZN(new_n731));
  NOR3_X1   g545(.A1(new_n675), .A2(new_n663), .A3(new_n389), .ZN(new_n732));
  NAND4_X1  g546(.A1(new_n731), .A2(new_n712), .A3(new_n713), .A4(new_n732), .ZN(new_n733));
  XOR2_X1   g547(.A(KEYINPUT108), .B(G122), .Z(new_n734));
  XNOR2_X1  g548(.A(new_n733), .B(new_n734), .ZN(G24));
  AOI21_X1  g549(.A(new_n525), .B1(new_n512), .B2(new_n514), .ZN(new_n736));
  AOI22_X1  g550(.A1(new_n736), .A2(new_n546), .B1(new_n550), .B2(new_n551), .ZN(new_n737));
  AOI21_X1  g551(.A(G902), .B1(new_n737), .B2(new_n545), .ZN(new_n738));
  OAI21_X1  g552(.A(KEYINPUT107), .B1(new_n738), .B2(new_n492), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n656), .A2(new_n585), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n740), .B1(new_n591), .B2(new_n592), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n739), .A2(new_n741), .A3(new_n725), .A4(new_n729), .ZN(new_n742));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g558(.A(new_n730), .ZN(new_n745));
  NAND4_X1  g559(.A1(new_n745), .A2(KEYINPUT109), .A3(new_n741), .A4(new_n725), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n744), .A2(new_n746), .ZN(new_n747));
  NOR3_X1   g561(.A1(new_n710), .A2(new_n663), .A3(new_n693), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G125), .ZN(G27));
  NAND3_X1  g564(.A1(new_n306), .A2(new_n187), .A3(new_n310), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT111), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n306), .A2(KEYINPUT111), .A3(new_n187), .A4(new_n310), .ZN(new_n754));
  AND3_X1   g568(.A1(new_n753), .A2(new_n429), .A3(new_n754), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n756));
  AND2_X1   g570(.A1(new_n486), .A2(new_n487), .ZN(new_n757));
  INV_X1    g571(.A(new_n474), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n464), .A2(new_n481), .A3(new_n433), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n759), .A2(new_n477), .ZN(new_n760));
  NOR2_X1   g574(.A1(new_n480), .A2(new_n481), .ZN(new_n761));
  OAI211_X1 g575(.A(G469), .B(new_n758), .C1(new_n760), .C2(new_n761), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n756), .B1(new_n757), .B2(new_n762), .ZN(new_n763));
  AND4_X1   g577(.A1(new_n756), .A2(new_n762), .A3(new_n487), .A4(new_n486), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n755), .A2(new_n765), .A3(KEYINPUT112), .ZN(new_n766));
  INV_X1    g580(.A(KEYINPUT112), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n753), .A2(new_n429), .A3(new_n754), .ZN(new_n768));
  OAI21_X1  g582(.A(KEYINPUT110), .B1(new_n483), .B2(new_n488), .ZN(new_n769));
  NAND4_X1  g583(.A1(new_n762), .A2(new_n756), .A3(new_n487), .A4(new_n486), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n767), .B1(new_n768), .B2(new_n771), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n766), .A2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n693), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n594), .A3(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(KEYINPUT42), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(new_n558), .ZN(new_n778));
  INV_X1    g592(.A(new_n593), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n778), .A2(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n780), .B1(new_n766), .B2(new_n772), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(KEYINPUT42), .A3(new_n774), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n777), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  NOR2_X1   g598(.A1(new_n643), .A2(new_n669), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n773), .A2(new_n594), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G134), .ZN(G36));
  NAND2_X1  g601(.A1(new_n753), .A2(new_n754), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n382), .A2(new_n632), .ZN(new_n789));
  XOR2_X1   g603(.A(new_n789), .B(KEYINPUT43), .Z(new_n790));
  AND2_X1   g604(.A1(new_n790), .A2(new_n741), .ZN(new_n791));
  AND2_X1   g605(.A1(new_n604), .A2(new_n605), .ZN(new_n792));
  INV_X1    g606(.A(new_n792), .ZN(new_n793));
  NAND2_X1  g607(.A1(new_n791), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g608(.A1(new_n794), .A2(KEYINPUT44), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT44), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n791), .A2(new_n796), .A3(new_n793), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n788), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n476), .A2(new_n482), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n799), .A2(KEYINPUT45), .A3(new_n758), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n801));
  XNOR2_X1  g615(.A(new_n800), .B(new_n801), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT45), .B1(new_n799), .B2(new_n758), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n803), .A2(new_n430), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n802), .A2(new_n804), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT114), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT46), .B1(new_n806), .B2(new_n487), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n805), .A2(KEYINPUT114), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT114), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n809), .B1(new_n802), .B2(new_n804), .ZN(new_n810));
  OAI211_X1 g624(.A(KEYINPUT46), .B(new_n487), .C1(new_n808), .C2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n811), .A2(new_n486), .ZN(new_n812));
  OR2_X1    g626(.A1(new_n807), .A2(new_n812), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n798), .A2(new_n813), .A3(new_n429), .A4(new_n685), .ZN(new_n814));
  XNOR2_X1  g628(.A(new_n814), .B(G137), .ZN(G39));
  NAND3_X1  g629(.A1(new_n813), .A2(KEYINPUT47), .A3(new_n429), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n429), .B1(new_n807), .B2(new_n812), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT47), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n778), .A2(new_n788), .A3(new_n779), .A4(new_n693), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n822), .A2(KEYINPUT115), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT115), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n820), .A2(new_n824), .A3(new_n821), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n826), .B(G140), .ZN(G42));
  NAND3_X1  g641(.A1(new_n779), .A2(new_n429), .A3(new_n187), .ZN(new_n828));
  NOR4_X1   g642(.A1(new_n828), .A2(new_n681), .A3(new_n682), .A4(new_n789), .ZN(new_n829));
  XNOR2_X1  g643(.A(new_n709), .B(KEYINPUT49), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT116), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n832), .B1(new_n633), .B2(new_n636), .ZN(new_n833));
  NAND4_X1  g647(.A1(new_n697), .A2(KEYINPUT116), .A3(new_n311), .A4(new_n390), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(KEYINPUT118), .ZN(new_n836));
  OR3_X1    g650(.A1(new_n420), .A2(new_n421), .A3(KEYINPUT117), .ZN(new_n837));
  OAI21_X1  g651(.A(KEYINPUT117), .B1(new_n420), .B2(new_n421), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n837), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n836), .B1(new_n621), .B2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n382), .A2(KEYINPUT118), .A3(new_n839), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n636), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n835), .A2(new_n843), .ZN(new_n844));
  OAI21_X1  g658(.A(new_n659), .B1(new_n844), .B2(new_n607), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n598), .ZN(new_n846));
  INV_X1    g660(.A(new_n788), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n621), .A2(new_n669), .A3(new_n839), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n847), .A2(new_n684), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n778), .A2(new_n741), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n851), .B1(new_n781), .B2(new_n785), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n693), .B1(new_n744), .B2(new_n746), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n853), .A2(new_n773), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n846), .A2(new_n852), .A3(new_n854), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n699), .A2(new_n700), .B1(new_n664), .B2(new_n670), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n675), .A2(new_n663), .ZN(new_n857));
  AND4_X1   g671(.A1(new_n429), .A2(new_n857), .A3(new_n657), .A4(new_n692), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n858), .A2(new_n681), .A3(new_n765), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n856), .A2(new_n749), .A3(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n856), .A2(new_n749), .A3(new_n859), .A4(KEYINPUT52), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n855), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n714), .A2(new_n717), .A3(new_n721), .A4(new_n733), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n777), .B2(new_n782), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT119), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  AND4_X1   g682(.A1(new_n714), .A2(new_n717), .A3(new_n721), .A4(new_n733), .ZN(new_n869));
  AND4_X1   g683(.A1(KEYINPUT42), .A2(new_n773), .A3(new_n594), .A4(new_n774), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT42), .B1(new_n781), .B2(new_n774), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n869), .B1(new_n870), .B2(new_n871), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n873));
  NAND4_X1  g687(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n868), .A4(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT54), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n862), .A2(new_n863), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n596), .A2(new_n597), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n490), .ZN(new_n878));
  AOI21_X1  g692(.A(KEYINPUT118), .B1(new_n382), .B2(new_n839), .ZN(new_n879));
  AND4_X1   g693(.A1(KEYINPUT118), .A2(new_n696), .A3(new_n839), .A4(new_n609), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n833), .B(new_n834), .C1(new_n881), .C2(new_n636), .ZN(new_n882));
  AOI22_X1  g696(.A1(new_n608), .A2(new_n882), .B1(new_n792), .B2(new_n658), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n878), .A2(new_n883), .A3(new_n854), .ZN(new_n884));
  INV_X1    g698(.A(new_n851), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n786), .A2(new_n885), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n884), .A2(new_n886), .ZN(new_n887));
  NAND3_X1  g701(.A1(new_n876), .A2(new_n887), .A3(new_n866), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT53), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n888), .A2(new_n889), .ZN(new_n890));
  AND3_X1   g704(.A1(new_n874), .A2(new_n875), .A3(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n864), .A2(KEYINPUT53), .A3(new_n866), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n875), .B1(new_n892), .B2(new_n890), .ZN(new_n893));
  OAI21_X1  g707(.A(KEYINPUT120), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g708(.A(KEYINPUT120), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n874), .A2(new_n875), .A3(new_n890), .ZN(new_n896));
  AND2_X1   g710(.A1(new_n892), .A2(new_n890), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n895), .B(new_n896), .C1(new_n897), .C2(new_n875), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n894), .A2(new_n898), .ZN(new_n899));
  AND3_X1   g713(.A1(new_n790), .A2(new_n386), .A3(new_n731), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n900), .A2(new_n311), .A3(new_n720), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n755), .A2(new_n709), .ZN(new_n902));
  NOR4_X1   g716(.A1(new_n902), .A2(new_n593), .A3(new_n385), .A4(new_n681), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n697), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n901), .A2(new_n904), .A3(new_n383), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT122), .ZN(new_n907));
  AND4_X1   g721(.A1(new_n386), .A2(new_n790), .A3(new_n709), .A4(new_n755), .ZN(new_n908));
  NAND2_X1  g722(.A1(new_n908), .A2(new_n594), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(KEYINPUT48), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n906), .A2(new_n907), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT121), .ZN(new_n912));
  NOR3_X1   g726(.A1(new_n682), .A2(new_n710), .A3(new_n187), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n912), .B1(new_n900), .B2(new_n913), .ZN(new_n914));
  OR2_X1    g728(.A1(new_n914), .A2(KEYINPUT50), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n914), .A2(KEYINPUT50), .ZN(new_n916));
  NOR2_X1   g730(.A1(new_n621), .A2(new_n632), .ZN(new_n917));
  AOI22_X1  g731(.A1(new_n908), .A2(new_n747), .B1(new_n903), .B2(new_n917), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n916), .A3(new_n918), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n709), .A2(new_n428), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n816), .A2(new_n819), .A3(new_n920), .ZN(new_n921));
  AND2_X1   g735(.A1(new_n900), .A2(new_n847), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n919), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n911), .B1(new_n923), .B2(KEYINPUT51), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(KEYINPUT51), .B2(new_n923), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n899), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g740(.A1(G952), .A2(G953), .ZN(new_n927));
  OAI21_X1  g741(.A(new_n831), .B1(new_n926), .B2(new_n927), .ZN(G75));
  NAND2_X1  g742(.A1(new_n242), .A2(new_n268), .ZN(new_n929));
  XNOR2_X1  g743(.A(new_n929), .B(new_n267), .ZN(new_n930));
  INV_X1    g744(.A(new_n930), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n876), .A2(new_n887), .A3(KEYINPUT53), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n872), .A2(KEYINPUT119), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n867), .B1(new_n783), .B2(new_n869), .ZN(new_n934));
  NOR3_X1   g748(.A1(new_n932), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  AOI21_X1  g749(.A(KEYINPUT53), .B1(new_n864), .B2(new_n866), .ZN(new_n936));
  OAI211_X1 g750(.A(G210), .B(G902), .C1(new_n935), .C2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT55), .ZN(new_n938));
  NOR2_X1   g752(.A1(KEYINPUT123), .A2(KEYINPUT56), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n938), .B1(new_n937), .B2(new_n939), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n931), .B1(new_n940), .B2(new_n941), .ZN(new_n942));
  INV_X1    g756(.A(G210), .ZN(new_n943));
  AOI211_X1 g757(.A(new_n943), .B(new_n298), .C1(new_n874), .C2(new_n890), .ZN(new_n944));
  INV_X1    g758(.A(new_n939), .ZN(new_n945));
  OAI21_X1  g759(.A(KEYINPUT55), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n930), .A3(new_n947), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n314), .A2(G952), .ZN(new_n949));
  INV_X1    g763(.A(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n942), .A2(new_n948), .A3(new_n950), .ZN(G51));
  OAI21_X1  g765(.A(KEYINPUT54), .B1(new_n935), .B2(new_n936), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n952), .A2(new_n896), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n487), .B(KEYINPUT57), .Z(new_n954));
  NAND2_X1  g768(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  XNOR2_X1  g769(.A(new_n705), .B(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n874), .A2(new_n890), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n958), .A2(G902), .ZN(new_n959));
  OR2_X1    g773(.A1(new_n959), .A2(new_n806), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n949), .B1(new_n957), .B2(new_n960), .ZN(G54));
  NAND2_X1  g775(.A1(KEYINPUT58), .A2(G475), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n376), .B1(new_n959), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n963), .A2(new_n950), .ZN(new_n964));
  NOR3_X1   g778(.A1(new_n959), .A2(new_n376), .A3(new_n962), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n964), .A2(new_n965), .ZN(G60));
  INV_X1    g780(.A(KEYINPUT125), .ZN(new_n967));
  NAND2_X1  g781(.A1(G478), .A2(G902), .ZN(new_n968));
  XOR2_X1   g782(.A(new_n968), .B(KEYINPUT59), .Z(new_n969));
  INV_X1    g783(.A(new_n969), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n629), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n967), .B1(new_n953), .B2(new_n972), .ZN(new_n973));
  AOI211_X1 g787(.A(KEYINPUT125), .B(new_n971), .C1(new_n952), .C2(new_n896), .ZN(new_n974));
  OAI21_X1  g788(.A(new_n950), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n629), .B1(new_n899), .B2(new_n970), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n975), .A2(new_n976), .ZN(G63));
  NOR2_X1   g791(.A1(new_n933), .A2(new_n934), .ZN(new_n978));
  INV_X1    g792(.A(new_n932), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n978), .A2(new_n979), .B1(new_n889), .B2(new_n888), .ZN(new_n980));
  NAND2_X1  g794(.A1(G217), .A2(G902), .ZN(new_n981));
  XOR2_X1   g795(.A(new_n981), .B(KEYINPUT60), .Z(new_n982));
  INV_X1    g796(.A(new_n982), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n651), .B1(new_n980), .B2(new_n983), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n958), .A2(new_n656), .A3(new_n982), .ZN(new_n985));
  NAND3_X1  g799(.A1(new_n984), .A2(new_n950), .A3(new_n985), .ZN(new_n986));
  AND3_X1   g800(.A1(new_n986), .A2(KEYINPUT126), .A3(KEYINPUT61), .ZN(new_n987));
  AOI21_X1  g801(.A(KEYINPUT61), .B1(new_n986), .B2(KEYINPUT126), .ZN(new_n988));
  NOR2_X1   g802(.A1(new_n987), .A2(new_n988), .ZN(G66));
  NOR3_X1   g803(.A1(new_n388), .A2(new_n264), .A3(new_n314), .ZN(new_n990));
  NOR3_X1   g804(.A1(new_n865), .A2(new_n598), .A3(new_n845), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n990), .B1(new_n991), .B2(new_n314), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n929), .B1(G898), .B2(new_n314), .ZN(new_n993));
  XNOR2_X1  g807(.A(new_n992), .B(new_n993), .ZN(G69));
  NOR2_X1   g808(.A1(new_n530), .A2(new_n531), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n995), .B(new_n370), .ZN(new_n996));
  INV_X1    g810(.A(new_n996), .ZN(new_n997));
  AOI211_X1 g811(.A(new_n788), .B(new_n686), .C1(new_n633), .C2(new_n881), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n877), .ZN(new_n999));
  INV_X1    g813(.A(new_n689), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n856), .A2(new_n749), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g816(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1003));
  AND2_X1   g817(.A1(new_n1002), .A2(KEYINPUT62), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n814), .B(new_n999), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1005));
  INV_X1    g819(.A(new_n1005), .ZN(new_n1006));
  AND3_X1   g820(.A1(new_n820), .A2(new_n824), .A3(new_n821), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n824), .B1(new_n820), .B2(new_n821), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  AOI21_X1  g823(.A(new_n997), .B1(new_n1009), .B2(new_n314), .ZN(new_n1010));
  INV_X1    g824(.A(new_n1010), .ZN(new_n1011));
  AOI21_X1  g825(.A(new_n314), .B1(G227), .B2(G900), .ZN(new_n1012));
  INV_X1    g826(.A(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(new_n1001), .B1(new_n785), .B2(new_n781), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n798), .B1(new_n594), .B2(new_n857), .ZN(new_n1015));
  NAND3_X1  g829(.A1(new_n813), .A2(new_n429), .A3(new_n685), .ZN(new_n1016));
  OAI211_X1 g830(.A(new_n783), .B(new_n1014), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1017), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n826), .A2(new_n314), .A3(new_n1018), .ZN(new_n1019));
  AOI21_X1  g833(.A(new_n996), .B1(G900), .B2(G953), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  NAND3_X1  g835(.A1(new_n1011), .A2(new_n1013), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g836(.A(new_n1020), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1017), .B1(new_n823), .B2(new_n825), .ZN(new_n1024));
  AOI21_X1  g838(.A(new_n1023), .B1(new_n1024), .B2(new_n314), .ZN(new_n1025));
  OAI21_X1  g839(.A(new_n1012), .B1(new_n1025), .B2(new_n1010), .ZN(new_n1026));
  NAND2_X1  g840(.A1(new_n1022), .A2(new_n1026), .ZN(G72));
  NOR2_X1   g841(.A1(new_n533), .A2(new_n525), .ZN(new_n1028));
  XOR2_X1   g842(.A(new_n1028), .B(KEYINPUT127), .Z(new_n1029));
  NAND2_X1  g843(.A1(new_n1024), .A2(new_n991), .ZN(new_n1030));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  AOI21_X1  g846(.A(new_n1029), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  NAND2_X1  g847(.A1(new_n533), .A2(new_n525), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n826), .A2(new_n991), .A3(new_n1006), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1034), .B1(new_n1035), .B2(new_n1032), .ZN(new_n1036));
  INV_X1    g850(.A(new_n535), .ZN(new_n1037));
  OAI21_X1  g851(.A(new_n1032), .B1(new_n1037), .B2(new_n678), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n950), .B1(new_n897), .B2(new_n1038), .ZN(new_n1039));
  NOR3_X1   g853(.A1(new_n1033), .A2(new_n1036), .A3(new_n1039), .ZN(G57));
endmodule


