//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 0 1 1 1 1 1 1 1 0 0 1 1 0 1 1 0 1 0 0 0 1 0 0 0 1 0 0 1 0 0 0 1 0 1 1 1 1 1 1 0 0 1 0 0 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:47 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n205, new_n206, new_n207, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1277,
    new_n1278, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1287, new_n1288, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1351, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356, new_n1357;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  INV_X1    g0004(.A(G97), .ZN(new_n205));
  INV_X1    g0005(.A(G107), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n207), .A2(G87), .ZN(G355));
  INV_X1    g0008(.A(G1), .ZN(new_n209));
  INV_X1    g0009(.A(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g0011(.A(new_n211), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n212), .A2(G13), .ZN(new_n213));
  OAI211_X1 g0013(.A(new_n213), .B(G250), .C1(G257), .C2(G264), .ZN(new_n214));
  XNOR2_X1  g0014(.A(new_n214), .B(KEYINPUT0), .ZN(new_n215));
  AND2_X1   g0015(.A1(G1), .A2(G13), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n216), .A2(G20), .ZN(new_n217));
  INV_X1    g0017(.A(new_n201), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n218), .A2(G50), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT64), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G116), .B2(G270), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n212), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n215), .B1(new_n217), .B2(new_n219), .C1(new_n226), .C2(KEYINPUT1), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G250), .B(G257), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(KEYINPUT65), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G264), .B(G270), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  INV_X1    g0033(.A(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT2), .B(G226), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n232), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(KEYINPUT66), .Z(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G68), .ZN(new_n243));
  INV_X1    g0043(.A(G68), .ZN(new_n244));
  NAND2_X1  g0044(.A1(new_n244), .A2(G50), .ZN(new_n245));
  NAND2_X1  g0045(.A1(new_n243), .A2(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(G58), .B(G77), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(new_n242), .B(new_n248), .ZN(G351));
  INV_X1    g0049(.A(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n250), .A2(new_n244), .ZN(new_n251));
  OAI21_X1  g0051(.A(G20), .B1(new_n251), .B2(new_n201), .ZN(new_n252));
  NOR2_X1   g0052(.A1(G20), .A2(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(G159), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(KEYINPUT71), .ZN(new_n257));
  INV_X1    g0057(.A(KEYINPUT3), .ZN(new_n258));
  OAI21_X1  g0058(.A(new_n257), .B1(new_n258), .B2(G33), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(G33), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n261), .A2(KEYINPUT71), .A3(KEYINPUT3), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n259), .A2(new_n260), .A3(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(KEYINPUT7), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n263), .A2(new_n264), .A3(new_n210), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G68), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n264), .B1(new_n263), .B2(new_n210), .ZN(new_n267));
  OAI211_X1 g0067(.A(KEYINPUT16), .B(new_n256), .C1(new_n266), .C2(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT16), .ZN(new_n269));
  INV_X1    g0069(.A(KEYINPUT72), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT7), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n264), .A2(KEYINPUT72), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  OAI21_X1  g0074(.A(new_n273), .B1(new_n274), .B2(G20), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n260), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n277), .A2(new_n210), .A3(new_n272), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n244), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n269), .B1(new_n279), .B2(new_n255), .ZN(new_n280));
  NAND3_X1  g0080(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n281));
  NAND2_X1  g0081(.A1(G1), .A2(G13), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n268), .A2(new_n280), .A3(new_n283), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  AOI21_X1  g0085(.A(new_n285), .B1(new_n209), .B2(G20), .ZN(new_n286));
  NAND3_X1  g0086(.A1(new_n209), .A2(G13), .A3(G20), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NOR2_X1   g0088(.A1(new_n288), .A2(new_n283), .ZN(new_n289));
  AOI22_X1  g0089(.A1(new_n286), .A2(new_n289), .B1(new_n288), .B2(new_n285), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n284), .A2(new_n290), .ZN(new_n291));
  NAND2_X1  g0091(.A1(G33), .A2(G41), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G1), .A3(G13), .ZN(new_n293));
  NOR2_X1   g0093(.A1(G223), .A2(G1698), .ZN(new_n294));
  INV_X1    g0094(.A(G226), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n294), .B1(new_n295), .B2(G1698), .ZN(new_n296));
  NAND4_X1  g0096(.A1(new_n296), .A2(new_n260), .A3(new_n259), .A4(new_n262), .ZN(new_n297));
  NAND2_X1  g0097(.A1(G33), .A2(G87), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n293), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G41), .ZN(new_n300));
  INV_X1    g0100(.A(G45), .ZN(new_n301));
  AOI21_X1  g0101(.A(G1), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n302), .A2(new_n293), .A3(G274), .ZN(new_n303));
  OAI21_X1  g0103(.A(new_n209), .B1(G41), .B2(G45), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n293), .A2(G232), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  OAI21_X1  g0106(.A(G169), .B1(new_n299), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n295), .A2(G1698), .ZN(new_n308));
  OAI21_X1  g0108(.A(new_n308), .B1(G223), .B2(G1698), .ZN(new_n309));
  OAI21_X1  g0109(.A(new_n298), .B1(new_n263), .B2(new_n309), .ZN(new_n310));
  INV_X1    g0110(.A(new_n293), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n306), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n312), .A2(G179), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n307), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n291), .A2(new_n315), .A3(KEYINPUT18), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n291), .A2(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT18), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g0122(.A1(new_n319), .A2(new_n317), .A3(new_n320), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n284), .A2(new_n290), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT74), .ZN(new_n326));
  AOI211_X1 g0126(.A(G190), .B(new_n306), .C1(new_n311), .C2(new_n310), .ZN(new_n327));
  AOI21_X1  g0127(.A(G200), .B1(new_n312), .B2(new_n313), .ZN(new_n328));
  OAI21_X1  g0128(.A(new_n326), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G200), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n299), .B2(new_n306), .ZN(new_n331));
  INV_X1    g0131(.A(G190), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n312), .A2(new_n332), .A3(new_n313), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n331), .A2(KEYINPUT74), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n329), .A2(new_n334), .ZN(new_n335));
  AND3_X1   g0135(.A1(new_n325), .A2(new_n335), .A3(KEYINPUT17), .ZN(new_n336));
  AOI21_X1  g0136(.A(KEYINPUT17), .B1(new_n325), .B2(new_n335), .ZN(new_n337));
  INV_X1    g0137(.A(KEYINPUT75), .ZN(new_n338));
  NOR3_X1   g0138(.A1(new_n336), .A2(new_n337), .A3(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT17), .ZN(new_n340));
  NOR3_X1   g0140(.A1(new_n327), .A2(new_n328), .A3(new_n326), .ZN(new_n341));
  AOI21_X1  g0141(.A(KEYINPUT74), .B1(new_n331), .B2(new_n333), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n340), .B1(new_n343), .B2(new_n291), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n325), .A2(new_n335), .A3(KEYINPUT17), .ZN(new_n345));
  AOI21_X1  g0145(.A(KEYINPUT75), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n324), .B1(new_n339), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g0147(.A(new_n347), .B(KEYINPUT76), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n210), .A2(G33), .ZN(new_n349));
  INV_X1    g0149(.A(G150), .ZN(new_n350));
  INV_X1    g0150(.A(new_n253), .ZN(new_n351));
  OAI22_X1  g0151(.A1(new_n285), .A2(new_n349), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G20), .B2(new_n203), .ZN(new_n353));
  INV_X1    g0153(.A(new_n283), .ZN(new_n354));
  NOR2_X1   g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n202), .B1(new_n209), .B2(G20), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n289), .A2(new_n356), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n357), .B1(G50), .B2(new_n287), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(new_n359), .B(KEYINPUT9), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n293), .A2(new_n304), .ZN(new_n361));
  OAI21_X1  g0161(.A(new_n303), .B1(new_n295), .B2(new_n361), .ZN(new_n362));
  NOR2_X1   g0162(.A1(G222), .A2(G1698), .ZN(new_n363));
  INV_X1    g0163(.A(G1698), .ZN(new_n364));
  NOR2_X1   g0164(.A1(new_n364), .A2(G223), .ZN(new_n365));
  OAI21_X1  g0165(.A(new_n274), .B1(new_n363), .B2(new_n365), .ZN(new_n366));
  INV_X1    g0166(.A(G77), .ZN(new_n367));
  AOI21_X1  g0167(.A(new_n293), .B1(new_n277), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n362), .B1(new_n366), .B2(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(G190), .ZN(new_n370));
  OAI211_X1 g0170(.A(new_n370), .B(KEYINPUT68), .C1(new_n330), .C2(new_n369), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n360), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT10), .ZN(new_n373));
  XNOR2_X1  g0173(.A(new_n372), .B(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(G20), .A2(G77), .ZN(new_n375));
  XNOR2_X1  g0175(.A(KEYINPUT15), .B(G87), .ZN(new_n376));
  OAI221_X1 g0176(.A(new_n375), .B1(new_n285), .B2(new_n351), .C1(new_n349), .C2(new_n376), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n377), .A2(new_n283), .ZN(new_n378));
  INV_X1    g0178(.A(new_n289), .ZN(new_n379));
  OAI21_X1  g0179(.A(G77), .B1(new_n210), .B2(G1), .ZN(new_n380));
  OAI22_X1  g0180(.A1(new_n379), .A2(new_n380), .B1(G77), .B2(new_n287), .ZN(new_n381));
  NOR2_X1   g0181(.A1(new_n378), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n274), .A2(G232), .A3(new_n364), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n206), .B2(new_n274), .ZN(new_n384));
  INV_X1    g0184(.A(G238), .ZN(new_n385));
  NOR3_X1   g0185(.A1(new_n277), .A2(new_n385), .A3(new_n364), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n311), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n303), .ZN(new_n388));
  INV_X1    g0188(.A(new_n361), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n388), .B1(G244), .B2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n387), .A2(new_n390), .ZN(new_n391));
  INV_X1    g0191(.A(G169), .ZN(new_n392));
  AOI21_X1  g0192(.A(new_n382), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(G179), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n387), .A2(new_n394), .A3(new_n390), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n393), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(G200), .ZN(new_n397));
  OAI211_X1 g0197(.A(new_n397), .B(new_n382), .C1(new_n332), .C2(new_n391), .ZN(new_n398));
  AND2_X1   g0198(.A1(new_n396), .A2(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n399), .A2(KEYINPUT67), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n369), .A2(G169), .ZN(new_n401));
  AOI211_X1 g0201(.A(new_n401), .B(new_n359), .C1(new_n394), .C2(new_n369), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  OR2_X1    g0203(.A1(new_n399), .A2(KEYINPUT67), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n374), .A2(new_n400), .A3(new_n403), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n295), .A2(new_n364), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n234), .A2(G1698), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n274), .A2(new_n406), .A3(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n408), .B1(new_n261), .B2(new_n205), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n388), .B1(new_n409), .B2(new_n311), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT13), .ZN(new_n411));
  AOI21_X1  g0211(.A(KEYINPUT69), .B1(new_n293), .B2(new_n304), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n412), .A2(new_n385), .ZN(new_n413));
  INV_X1    g0213(.A(KEYINPUT69), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n413), .B1(new_n414), .B2(new_n361), .ZN(new_n415));
  NAND3_X1  g0215(.A1(new_n410), .A2(new_n411), .A3(new_n415), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n261), .A2(new_n205), .ZN(new_n417));
  AND2_X1   g0217(.A1(new_n406), .A2(new_n407), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n417), .B1(new_n418), .B2(new_n274), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n303), .B1(new_n419), .B2(new_n293), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n361), .A2(new_n414), .ZN(new_n421));
  NOR3_X1   g0221(.A1(new_n421), .A2(new_n385), .A3(new_n412), .ZN(new_n422));
  OAI21_X1  g0222(.A(KEYINPUT13), .B1(new_n420), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n416), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n424), .A2(G169), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(KEYINPUT14), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n416), .A2(new_n423), .A3(G179), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT14), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n424), .A2(new_n428), .A3(G169), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n426), .A2(new_n427), .A3(new_n429), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n288), .A2(new_n244), .ZN(new_n431));
  XNOR2_X1  g0231(.A(new_n431), .B(KEYINPUT12), .ZN(new_n432));
  AOI22_X1  g0232(.A1(new_n253), .A2(G50), .B1(G20), .B2(new_n244), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n367), .B2(new_n349), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n434), .A2(KEYINPUT11), .A3(new_n283), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n289), .B(G68), .C1(G1), .C2(new_n210), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(KEYINPUT11), .B1(new_n434), .B2(new_n283), .ZN(new_n438));
  NOR2_X1   g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g0239(.A(new_n439), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n416), .A2(new_n423), .A3(G190), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(new_n439), .ZN(new_n442));
  AOI21_X1  g0242(.A(new_n330), .B1(new_n416), .B2(new_n423), .ZN(new_n443));
  OAI21_X1  g0243(.A(KEYINPUT70), .B1(new_n442), .B2(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n424), .A2(G200), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT70), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n445), .A2(new_n446), .A3(new_n441), .A4(new_n439), .ZN(new_n447));
  AOI22_X1  g0247(.A1(new_n430), .A2(new_n440), .B1(new_n444), .B2(new_n447), .ZN(new_n448));
  INV_X1    g0248(.A(new_n448), .ZN(new_n449));
  NOR3_X1   g0249(.A1(new_n348), .A2(new_n405), .A3(new_n449), .ZN(new_n450));
  INV_X1    g0250(.A(G116), .ZN(new_n451));
  AOI22_X1  g0251(.A1(new_n281), .A2(new_n282), .B1(G20), .B2(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(G33), .A2(G283), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n453), .B(new_n210), .C1(G33), .C2(new_n205), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n452), .A2(new_n454), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n452), .A2(KEYINPUT20), .A3(new_n454), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n209), .A2(G33), .ZN(new_n460));
  AND3_X1   g0260(.A1(new_n354), .A2(new_n287), .A3(new_n460), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(G116), .ZN(new_n462));
  NAND2_X1  g0262(.A1(new_n288), .A2(new_n451), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  INV_X1    g0264(.A(KEYINPUT5), .ZN(new_n465));
  INV_X1    g0265(.A(KEYINPUT79), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n465), .B1(new_n466), .B2(G41), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n301), .A2(G1), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n300), .A2(KEYINPUT79), .A3(KEYINPUT5), .ZN(new_n469));
  NAND3_X1  g0269(.A1(new_n467), .A2(new_n468), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g0270(.A1(new_n470), .A2(G270), .A3(new_n293), .ZN(new_n471));
  INV_X1    g0271(.A(G274), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n472), .B1(new_n216), .B2(new_n292), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n473), .A2(new_n467), .A3(new_n468), .A4(new_n469), .ZN(new_n474));
  AND2_X1   g0274(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n277), .A2(G303), .ZN(new_n476));
  INV_X1    g0276(.A(G264), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n477), .A2(G1698), .ZN(new_n478));
  OAI21_X1  g0278(.A(new_n478), .B1(G257), .B2(G1698), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n476), .B1(new_n263), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n311), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n475), .A2(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n464), .A2(new_n482), .A3(G169), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT21), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  INV_X1    g0285(.A(new_n464), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n475), .A2(new_n481), .A3(G190), .ZN(new_n487));
  NOR2_X1   g0287(.A1(G257), .A2(G1698), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n488), .B1(new_n477), .B2(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n489), .A2(new_n260), .A3(new_n259), .A4(new_n262), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n293), .B1(new_n490), .B2(new_n476), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n471), .A2(new_n474), .ZN(new_n492));
  OAI21_X1  g0292(.A(G200), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n486), .A2(new_n487), .A3(new_n493), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n464), .A2(new_n482), .A3(KEYINPUT21), .A4(G169), .ZN(new_n495));
  NOR3_X1   g0295(.A1(new_n491), .A2(new_n492), .A3(new_n394), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n464), .ZN(new_n497));
  NAND4_X1  g0297(.A1(new_n485), .A2(new_n494), .A3(new_n495), .A4(new_n497), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  AND2_X1   g0300(.A1(new_n495), .A2(new_n497), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n501), .A2(KEYINPUT82), .A3(new_n485), .A4(new_n494), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(G33), .A2(G116), .ZN(new_n504));
  INV_X1    g0304(.A(G244), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G1698), .ZN(new_n506));
  OAI21_X1  g0306(.A(new_n506), .B1(G238), .B2(G1698), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n504), .B1(new_n263), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n508), .A2(KEYINPUT81), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT81), .ZN(new_n510));
  OAI211_X1 g0310(.A(new_n510), .B(new_n504), .C1(new_n263), .C2(new_n507), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n293), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n468), .ZN(new_n513));
  AND2_X1   g0313(.A1(new_n513), .A2(G250), .ZN(new_n514));
  AOI22_X1  g0314(.A1(new_n514), .A2(new_n293), .B1(new_n473), .B2(new_n468), .ZN(new_n515));
  INV_X1    g0315(.A(new_n515), .ZN(new_n516));
  NOR2_X1   g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(G190), .ZN(new_n518));
  OAI21_X1  g0318(.A(G200), .B1(new_n512), .B2(new_n516), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n349), .A2(KEYINPUT19), .A3(new_n205), .ZN(new_n520));
  OAI22_X1  g0320(.A1(new_n417), .A2(G20), .B1(new_n207), .B2(G87), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n520), .B1(new_n521), .B2(KEYINPUT19), .ZN(new_n522));
  NOR3_X1   g0322(.A1(new_n263), .A2(G20), .A3(new_n244), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n283), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n376), .A2(new_n288), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n461), .A2(G87), .ZN(new_n526));
  AND3_X1   g0326(.A1(new_n524), .A2(new_n525), .A3(new_n526), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n518), .A2(new_n519), .A3(new_n527), .ZN(new_n528));
  NOR2_X1   g0328(.A1(G238), .A2(G1698), .ZN(new_n529));
  AOI21_X1  g0329(.A(new_n529), .B1(new_n505), .B2(G1698), .ZN(new_n530));
  NAND4_X1  g0330(.A1(new_n530), .A2(new_n260), .A3(new_n259), .A4(new_n262), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n510), .B1(new_n531), .B2(new_n504), .ZN(new_n532));
  INV_X1    g0332(.A(new_n511), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n311), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n534), .A2(new_n394), .A3(new_n515), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n289), .A2(new_n460), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n524), .B(new_n525), .C1(new_n376), .C2(new_n536), .ZN(new_n537));
  OAI211_X1 g0337(.A(new_n535), .B(new_n537), .C1(new_n517), .C2(G169), .ZN(new_n538));
  AND2_X1   g0338(.A1(new_n528), .A2(new_n538), .ZN(new_n539));
  NOR2_X1   g0339(.A1(new_n505), .A2(G1698), .ZN(new_n540));
  NAND4_X1  g0340(.A1(new_n259), .A2(new_n262), .A3(new_n540), .A4(new_n260), .ZN(new_n541));
  INV_X1    g0341(.A(KEYINPUT4), .ZN(new_n542));
  AND2_X1   g0342(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n276), .A2(new_n260), .A3(G250), .A4(G1698), .ZN(new_n544));
  AND2_X1   g0344(.A1(KEYINPUT4), .A2(G244), .ZN(new_n545));
  NAND4_X1  g0345(.A1(new_n276), .A2(new_n260), .A3(new_n545), .A4(new_n364), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n546), .A3(new_n453), .ZN(new_n547));
  OAI21_X1  g0347(.A(new_n311), .B1(new_n543), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n470), .A2(G257), .A3(new_n293), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n549), .A2(new_n474), .ZN(new_n550));
  INV_X1    g0350(.A(new_n550), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(G169), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n541), .A2(new_n542), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n554), .A2(new_n453), .A3(new_n544), .A4(new_n546), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n550), .B1(new_n555), .B2(new_n311), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(G179), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n553), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n206), .A2(G97), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT77), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n560), .A2(KEYINPUT6), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n563));
  OAI21_X1  g0363(.A(new_n559), .B1(new_n561), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(KEYINPUT77), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n560), .A2(KEYINPUT6), .ZN(new_n566));
  NAND2_X1  g0366(.A1(G97), .A2(G107), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n207), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n564), .A2(new_n568), .A3(G20), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n253), .A2(G77), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n206), .B1(new_n275), .B2(new_n278), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n283), .B1(new_n571), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n287), .A2(G97), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n461), .B2(G97), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n558), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(KEYINPUT78), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n552), .A2(G200), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT78), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n573), .A2(new_n580), .A3(new_n575), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  INV_X1    g0382(.A(KEYINPUT80), .ZN(new_n583));
  OAI21_X1  g0383(.A(new_n583), .B1(new_n552), .B2(new_n332), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n556), .A2(KEYINPUT80), .A3(G190), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  OAI21_X1  g0386(.A(new_n577), .B1(new_n582), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(KEYINPUT22), .A2(G87), .ZN(new_n588));
  OR3_X1    g0388(.A1(new_n263), .A2(G20), .A3(new_n588), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT24), .ZN(new_n590));
  INV_X1    g0390(.A(KEYINPUT22), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n210), .A2(G87), .ZN(new_n592));
  OAI21_X1  g0392(.A(new_n591), .B1(new_n277), .B2(new_n592), .ZN(new_n593));
  NOR2_X1   g0393(.A1(new_n504), .A2(G20), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT23), .ZN(new_n595));
  OAI21_X1  g0395(.A(new_n595), .B1(new_n210), .B2(G107), .ZN(new_n596));
  NAND3_X1  g0396(.A1(new_n206), .A2(KEYINPUT23), .A3(G20), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n594), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n589), .A2(new_n590), .A3(new_n593), .A4(new_n598), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n593), .A2(new_n598), .ZN(new_n600));
  NOR3_X1   g0400(.A1(new_n263), .A2(G20), .A3(new_n588), .ZN(new_n601));
  OAI21_X1  g0401(.A(KEYINPUT24), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g0402(.A(new_n354), .B1(new_n599), .B2(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n287), .A2(G107), .ZN(new_n604));
  XNOR2_X1  g0404(.A(KEYINPUT83), .B(KEYINPUT25), .ZN(new_n605));
  XNOR2_X1  g0405(.A(new_n604), .B(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n206), .B2(new_n536), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  OR2_X1    g0408(.A1(G250), .A2(G1698), .ZN(new_n609));
  OAI21_X1  g0409(.A(new_n609), .B1(G257), .B2(new_n364), .ZN(new_n610));
  INV_X1    g0410(.A(G294), .ZN(new_n611));
  OAI22_X1  g0411(.A1(new_n263), .A2(new_n610), .B1(new_n261), .B2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n311), .ZN(new_n613));
  AND2_X1   g0413(.A1(new_n470), .A2(new_n293), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G264), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(new_n615), .A3(new_n474), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n616), .A2(new_n330), .ZN(new_n617));
  OAI21_X1  g0417(.A(new_n617), .B1(G190), .B2(new_n616), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n608), .A2(new_n618), .ZN(new_n619));
  AOI22_X1  g0419(.A1(new_n311), .A2(new_n612), .B1(new_n614), .B2(G264), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n620), .A2(new_n394), .A3(new_n474), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n616), .A2(new_n392), .ZN(new_n622));
  OAI211_X1 g0422(.A(new_n621), .B(new_n622), .C1(new_n603), .C2(new_n607), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n619), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n587), .A2(new_n624), .ZN(new_n625));
  AND4_X1   g0425(.A1(new_n450), .A2(new_n503), .A3(new_n539), .A4(new_n625), .ZN(G372));
  NAND2_X1  g0426(.A1(new_n519), .A2(new_n527), .ZN(new_n627));
  AOI22_X1  g0427(.A1(new_n627), .A2(KEYINPUT84), .B1(G190), .B2(new_n517), .ZN(new_n628));
  INV_X1    g0428(.A(KEYINPUT84), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n519), .A2(new_n629), .A3(new_n527), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n578), .A2(new_n581), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n632), .A2(new_n558), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT26), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n631), .A2(new_n633), .A3(new_n634), .A4(new_n538), .ZN(new_n635));
  INV_X1    g0435(.A(new_n538), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n553), .A2(new_n557), .B1(new_n573), .B2(new_n575), .ZN(new_n637));
  NAND3_X1  g0437(.A1(new_n528), .A2(new_n538), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n636), .B1(new_n638), .B2(KEYINPUT26), .ZN(new_n639));
  OR2_X1    g0439(.A1(new_n582), .A2(new_n586), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n501), .A2(new_n623), .A3(new_n485), .ZN(new_n641));
  NAND4_X1  g0441(.A1(new_n640), .A2(new_n619), .A3(new_n577), .A4(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n631), .A2(new_n538), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n635), .B(new_n639), .C1(new_n642), .C2(new_n643), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n450), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n321), .A2(new_n316), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n338), .B1(new_n336), .B2(new_n337), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n344), .A2(KEYINPUT75), .A3(new_n345), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n429), .A2(new_n427), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n428), .B1(new_n424), .B2(G169), .ZN(new_n652));
  OAI21_X1  g0452(.A(new_n440), .B1(new_n651), .B2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n444), .A2(new_n447), .ZN(new_n655));
  INV_X1    g0455(.A(new_n396), .ZN(new_n656));
  AOI21_X1  g0456(.A(new_n654), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  OAI21_X1  g0457(.A(new_n646), .B1(new_n650), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n402), .B1(new_n658), .B2(new_n374), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n645), .A2(new_n659), .ZN(G369));
  INV_X1    g0460(.A(KEYINPUT27), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n661), .A2(new_n209), .A3(new_n210), .A4(G13), .ZN(new_n662));
  XOR2_X1   g0462(.A(new_n662), .B(KEYINPUT85), .Z(new_n663));
  INV_X1    g0463(.A(G213), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n209), .A2(new_n210), .A3(G13), .ZN(new_n665));
  AOI21_X1  g0465(.A(new_n664), .B1(new_n665), .B2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n663), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT86), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND3_X1  g0469(.A1(new_n663), .A2(KEYINPUT86), .A3(new_n666), .ZN(new_n670));
  AND3_X1   g0470(.A1(new_n669), .A2(G343), .A3(new_n670), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n619), .B(new_n623), .C1(new_n608), .C2(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(new_n623), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n671), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n673), .A2(new_n675), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n671), .A2(new_n464), .ZN(new_n677));
  AND2_X1   g0477(.A1(new_n503), .A2(new_n677), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n501), .B2(new_n485), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n678), .A2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(KEYINPUT87), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NOR3_X1   g0482(.A1(new_n678), .A2(new_n679), .A3(KEYINPUT87), .ZN(new_n683));
  OAI211_X1 g0483(.A(G330), .B(new_n676), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n501), .A2(new_n485), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n685), .A2(new_n623), .A3(new_n619), .A4(new_n672), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n674), .A2(new_n672), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n686), .A2(KEYINPUT88), .A3(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  AOI21_X1  g0489(.A(KEYINPUT88), .B1(new_n686), .B2(new_n687), .ZN(new_n690));
  OR2_X1    g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n684), .A2(new_n691), .ZN(G399));
  INV_X1    g0492(.A(new_n213), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(G41), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n207), .A2(G87), .A3(G116), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n695), .A2(G1), .A3(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n697), .B1(new_n219), .B2(new_n695), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT28), .ZN(new_n699));
  OAI21_X1  g0499(.A(KEYINPUT92), .B1(new_n642), .B2(new_n643), .ZN(new_n700));
  NAND4_X1  g0500(.A1(new_n528), .A2(new_n634), .A3(new_n538), .A4(new_n637), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n701), .A2(new_n538), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n631), .A2(new_n633), .A3(new_n538), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n703), .B2(KEYINPUT26), .ZN(new_n704));
  OAI211_X1 g0504(.A(new_n619), .B(new_n577), .C1(new_n582), .C2(new_n586), .ZN(new_n705));
  INV_X1    g0505(.A(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n636), .B1(new_n628), .B2(new_n630), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT92), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n706), .A2(new_n707), .A3(new_n708), .A4(new_n641), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n700), .A2(new_n704), .A3(new_n709), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n710), .A2(new_n672), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(KEYINPUT29), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g0513(.A1(new_n644), .A2(new_n672), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(KEYINPUT29), .ZN(new_n715));
  INV_X1    g0515(.A(G330), .ZN(new_n716));
  XOR2_X1   g0516(.A(KEYINPUT90), .B(KEYINPUT30), .Z(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AND4_X1   g0518(.A1(new_n496), .A2(new_n534), .A3(new_n515), .A4(new_n620), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n718), .B1(new_n719), .B2(new_n556), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n496), .A2(new_n534), .A3(new_n515), .A4(new_n620), .ZN(new_n721));
  NAND2_X1  g0521(.A1(new_n556), .A2(KEYINPUT30), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n475), .B2(new_n481), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(new_n552), .A3(new_n616), .ZN(new_n724));
  OAI22_X1  g0524(.A1(new_n721), .A2(new_n722), .B1(new_n724), .B2(new_n517), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n720), .A2(new_n725), .ZN(new_n726));
  XNOR2_X1  g0526(.A(KEYINPUT89), .B(KEYINPUT31), .ZN(new_n727));
  NOR3_X1   g0527(.A1(new_n726), .A2(new_n672), .A3(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(KEYINPUT31), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT91), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(new_n720), .B2(new_n725), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n721), .A2(new_n722), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n717), .B1(new_n721), .B2(new_n552), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n534), .A2(new_n515), .ZN(new_n734));
  NAND4_X1  g0534(.A1(new_n734), .A2(new_n616), .A3(new_n552), .A4(new_n723), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n732), .A2(new_n733), .A3(KEYINPUT91), .A4(new_n735), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n731), .A2(new_n671), .A3(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n728), .B1(new_n729), .B2(new_n737), .ZN(new_n738));
  NAND4_X1  g0538(.A1(new_n625), .A2(new_n503), .A3(new_n539), .A4(new_n672), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n716), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NOR3_X1   g0540(.A1(new_n713), .A2(new_n715), .A3(new_n740), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n699), .B1(new_n741), .B2(G1), .ZN(G364));
  OR3_X1    g0542(.A1(new_n682), .A2(G330), .A3(new_n683), .ZN(new_n743));
  OAI21_X1  g0543(.A(G330), .B1(new_n682), .B2(new_n683), .ZN(new_n744));
  INV_X1    g0544(.A(G13), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n745), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n209), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n694), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n743), .A2(new_n744), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  AOI21_X1  g0554(.A(new_n282), .B1(G20), .B2(new_n392), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n248), .A2(new_n301), .ZN(new_n758));
  INV_X1    g0558(.A(new_n263), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n693), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n219), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n761), .B1(new_n301), .B2(new_n762), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n758), .B1(new_n763), .B2(KEYINPUT94), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(KEYINPUT94), .B2(new_n763), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n213), .A2(new_n274), .ZN(new_n766));
  INV_X1    g0566(.A(G355), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n766), .B1(KEYINPUT93), .B2(new_n767), .ZN(new_n768));
  OR2_X1    g0568(.A1(new_n767), .A2(KEYINPUT93), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n768), .A2(new_n769), .B1(new_n451), .B2(new_n693), .ZN(new_n770));
  AOI21_X1  g0570(.A(new_n757), .B1(new_n765), .B2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n755), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n332), .A2(G200), .ZN(new_n773));
  NAND2_X1  g0573(.A1(new_n773), .A2(new_n394), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(G20), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(G97), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n210), .A2(new_n394), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n777), .A2(G200), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n778), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n776), .B1(new_n780), .B2(new_n244), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  INV_X1    g0582(.A(KEYINPUT95), .ZN(new_n783));
  XNOR2_X1  g0583(.A(new_n777), .B(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(G190), .A2(G200), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n787), .A2(G77), .ZN(new_n788));
  NOR2_X1   g0588(.A1(new_n210), .A2(G179), .ZN(new_n789));
  NAND2_X1  g0589(.A1(new_n789), .A2(new_n785), .ZN(new_n790));
  INV_X1    g0590(.A(G159), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n790), .A2(KEYINPUT32), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n784), .A2(new_n773), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n277), .B(new_n792), .C1(new_n794), .C2(G58), .ZN(new_n795));
  OAI21_X1  g0595(.A(KEYINPUT32), .B1(new_n790), .B2(new_n791), .ZN(new_n796));
  NAND3_X1  g0596(.A1(new_n789), .A2(new_n332), .A3(G200), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n778), .A2(new_n332), .ZN(new_n798));
  INV_X1    g0598(.A(new_n798), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n796), .B1(new_n206), .B2(new_n797), .C1(new_n799), .C2(new_n202), .ZN(new_n800));
  NAND3_X1  g0600(.A1(new_n789), .A2(G190), .A3(G200), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT96), .ZN(new_n802));
  OR2_X1    g0602(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n801), .A2(new_n802), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g0605(.A(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n800), .B1(G87), .B2(new_n806), .ZN(new_n807));
  NAND4_X1  g0607(.A1(new_n782), .A2(new_n788), .A3(new_n795), .A4(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n798), .A2(G326), .B1(new_n775), .B2(G294), .ZN(new_n809));
  NOR2_X1   g0609(.A1(KEYINPUT33), .A2(G317), .ZN(new_n810));
  AND2_X1   g0610(.A1(KEYINPUT33), .A2(G317), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n779), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n813), .B1(G303), .B2(new_n806), .ZN(new_n814));
  INV_X1    g0614(.A(new_n790), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n274), .B1(new_n815), .B2(G329), .ZN(new_n816));
  INV_X1    g0616(.A(G283), .ZN(new_n817));
  OAI21_X1  g0617(.A(new_n816), .B1(new_n817), .B2(new_n797), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n818), .B1(new_n794), .B2(G322), .ZN(new_n819));
  INV_X1    g0619(.A(G311), .ZN(new_n820));
  OAI211_X1 g0620(.A(new_n814), .B(new_n819), .C1(new_n820), .C2(new_n786), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n772), .B1(new_n808), .B2(new_n821), .ZN(new_n822));
  NOR3_X1   g0622(.A1(new_n771), .A2(new_n822), .A3(new_n750), .ZN(new_n823));
  INV_X1    g0623(.A(new_n680), .ZN(new_n824));
  INV_X1    g0624(.A(new_n754), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n823), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  AND2_X1   g0626(.A1(new_n751), .A2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n827), .ZN(G396));
  NAND2_X1  g0628(.A1(new_n656), .A2(new_n672), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT99), .ZN(new_n830));
  OAI21_X1  g0630(.A(new_n671), .B1(new_n378), .B2(new_n381), .ZN(new_n831));
  AND2_X1   g0631(.A1(new_n831), .A2(new_n398), .ZN(new_n832));
  OAI211_X1 g0632(.A(new_n829), .B(new_n830), .C1(new_n656), .C2(new_n832), .ZN(new_n833));
  AOI22_X1  g0633(.A1(new_n831), .A2(new_n398), .B1(new_n395), .B2(new_n393), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n396), .A2(new_n671), .ZN(new_n835));
  OAI21_X1  g0635(.A(KEYINPUT99), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n833), .A2(new_n836), .ZN(new_n837));
  INV_X1    g0637(.A(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n714), .A2(new_n838), .ZN(new_n839));
  NAND3_X1  g0639(.A1(new_n644), .A2(new_n837), .A3(new_n672), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n740), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n841), .A2(new_n749), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n839), .A2(new_n740), .A3(new_n840), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n755), .A2(new_n752), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n750), .B1(new_n367), .B2(new_n845), .ZN(new_n846));
  AOI22_X1  g0646(.A1(G283), .A2(new_n779), .B1(new_n798), .B2(G303), .ZN(new_n847));
  OAI21_X1  g0647(.A(new_n847), .B1(new_n786), .B2(new_n451), .ZN(new_n848));
  XOR2_X1   g0648(.A(new_n848), .B(KEYINPUT98), .Z(new_n849));
  AOI21_X1  g0649(.A(new_n274), .B1(new_n815), .B2(G311), .ZN(new_n850));
  INV_X1    g0650(.A(new_n797), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n851), .A2(G87), .ZN(new_n852));
  AND3_X1   g0652(.A1(new_n850), .A2(new_n776), .A3(new_n852), .ZN(new_n853));
  OAI221_X1 g0653(.A(new_n853), .B1(new_n206), .B2(new_n805), .C1(new_n611), .C2(new_n793), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n849), .A2(new_n854), .ZN(new_n855));
  AOI22_X1  g0655(.A1(G137), .A2(new_n798), .B1(new_n779), .B2(G150), .ZN(new_n856));
  INV_X1    g0656(.A(G143), .ZN(new_n857));
  OAI221_X1 g0657(.A(new_n856), .B1(new_n786), .B2(new_n791), .C1(new_n857), .C2(new_n793), .ZN(new_n858));
  XNOR2_X1  g0658(.A(new_n858), .B(KEYINPUT34), .ZN(new_n859));
  AOI21_X1  g0659(.A(new_n263), .B1(new_n815), .B2(G132), .ZN(new_n860));
  INV_X1    g0660(.A(new_n775), .ZN(new_n861));
  OAI221_X1 g0661(.A(new_n860), .B1(new_n244), .B2(new_n797), .C1(new_n250), .C2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(new_n862), .B1(G50), .B2(new_n806), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n855), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n846), .B1(new_n772), .B2(new_n864), .C1(new_n837), .C2(new_n753), .ZN(new_n865));
  AND2_X1   g0665(.A1(new_n844), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(G384));
  NOR2_X1   g0667(.A1(new_n746), .A2(new_n209), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT40), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT38), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n256), .B1(new_n266), .B2(new_n267), .ZN(new_n871));
  AND2_X1   g0671(.A1(new_n871), .A2(new_n269), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n268), .A2(new_n283), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n290), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n669), .A2(new_n670), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g0677(.A(new_n877), .B1(new_n649), .B2(new_n324), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n325), .A2(new_n335), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n874), .A2(new_n315), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n879), .A2(new_n880), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n881), .A2(KEYINPUT37), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n291), .A2(new_n876), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n879), .A2(new_n319), .A3(new_n883), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n882), .B1(KEYINPUT37), .B2(new_n884), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n870), .B1(new_n878), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT101), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n647), .A2(new_n648), .B1(new_n322), .B2(new_n323), .ZN(new_n889));
  OAI211_X1 g0689(.A(KEYINPUT38), .B(new_n885), .C1(new_n889), .C2(new_n877), .ZN(new_n890));
  AND3_X1   g0690(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n891));
  AOI21_X1  g0691(.A(new_n888), .B1(new_n887), .B2(new_n890), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n430), .B1(new_n447), .B2(new_n444), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n440), .A2(new_n671), .ZN(new_n895));
  NOR2_X1   g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n655), .A2(new_n653), .A3(new_n895), .ZN(new_n897));
  INV_X1    g0697(.A(KEYINPUT100), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n448), .A2(KEYINPUT100), .A3(new_n895), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n896), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR2_X1   g0701(.A1(new_n901), .A2(new_n838), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n731), .A2(KEYINPUT31), .A3(new_n736), .A4(new_n671), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n739), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n737), .A2(KEYINPUT103), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT103), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n731), .A2(new_n906), .A3(new_n736), .A4(new_n671), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n905), .A2(new_n727), .A3(new_n907), .ZN(new_n908));
  INV_X1    g0708(.A(KEYINPUT104), .ZN(new_n909));
  AND3_X1   g0709(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n909), .B1(new_n904), .B2(new_n908), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n902), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n869), .B1(new_n893), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(KEYINPUT37), .ZN(new_n914));
  XNOR2_X1  g0714(.A(new_n884), .B(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n336), .A2(new_n337), .ZN(new_n916));
  AOI21_X1  g0716(.A(new_n883), .B1(new_n916), .B2(new_n646), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n870), .B1(new_n915), .B2(new_n917), .ZN(new_n918));
  AOI21_X1  g0718(.A(new_n869), .B1(new_n890), .B2(new_n918), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n919), .B(new_n902), .C1(new_n910), .C2(new_n911), .ZN(new_n920));
  AND2_X1   g0720(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n904), .A2(new_n908), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n922), .A2(KEYINPUT104), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n904), .A2(new_n908), .A3(new_n909), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n450), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n716), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n927), .B1(new_n921), .B2(new_n926), .ZN(new_n928));
  NAND2_X1  g0728(.A1(new_n840), .A2(new_n829), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n897), .A2(new_n898), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT100), .B1(new_n448), .B2(new_n895), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n930), .A2(new_n931), .B1(new_n895), .B2(new_n894), .ZN(new_n932));
  OAI211_X1 g0732(.A(new_n929), .B(new_n932), .C1(new_n891), .C2(new_n892), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n890), .A2(new_n918), .ZN(new_n934));
  INV_X1    g0734(.A(KEYINPUT39), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n887), .A2(KEYINPUT39), .A3(new_n890), .ZN(new_n937));
  NAND2_X1  g0737(.A1(new_n654), .A2(new_n672), .ZN(new_n938));
  XNOR2_X1  g0738(.A(new_n938), .B(KEYINPUT102), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n321), .A2(new_n316), .A3(new_n875), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n933), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n450), .B1(new_n713), .B2(new_n715), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n659), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n942), .B(new_n944), .ZN(new_n945));
  AOI21_X1  g0745(.A(new_n868), .B1(new_n928), .B2(new_n945), .ZN(new_n946));
  OAI21_X1  g0746(.A(new_n946), .B1(new_n945), .B2(new_n928), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n217), .A2(new_n451), .ZN(new_n948));
  NAND2_X1  g0748(.A1(new_n564), .A2(new_n568), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT35), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n951), .B1(new_n950), .B2(new_n949), .ZN(new_n952));
  XOR2_X1   g0752(.A(new_n952), .B(KEYINPUT36), .Z(new_n953));
  OAI21_X1  g0753(.A(G77), .B1(new_n250), .B2(new_n244), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n243), .B1(new_n219), .B2(new_n954), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n955), .A2(G1), .A3(new_n745), .ZN(new_n956));
  NAND3_X1  g0756(.A1(new_n947), .A2(new_n953), .A3(new_n956), .ZN(new_n957));
  XOR2_X1   g0757(.A(new_n957), .B(KEYINPUT105), .Z(G367));
  NAND2_X1  g0758(.A1(new_n633), .A2(new_n671), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n672), .B1(new_n578), .B2(new_n581), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n959), .B1(new_n587), .B2(new_n960), .ZN(new_n961));
  INV_X1    g0761(.A(new_n686), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT42), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  AND2_X1   g0765(.A1(new_n961), .A2(new_n674), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n672), .B1(new_n966), .B2(new_n637), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n965), .A2(new_n967), .ZN(new_n968));
  OR2_X1    g0768(.A1(new_n672), .A2(new_n527), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n707), .A2(new_n969), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n538), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  INV_X1    g0773(.A(KEYINPUT43), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n972), .A2(KEYINPUT43), .ZN(new_n976));
  NAND3_X1  g0776(.A1(new_n968), .A2(new_n975), .A3(new_n976), .ZN(new_n977));
  NAND4_X1  g0777(.A1(new_n965), .A2(new_n974), .A3(new_n973), .A4(new_n967), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  INV_X1    g0779(.A(KEYINPUT106), .ZN(new_n980));
  INV_X1    g0780(.A(new_n684), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n980), .B1(new_n981), .B2(new_n961), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n979), .A2(new_n982), .ZN(new_n983));
  AND2_X1   g0783(.A1(new_n981), .A2(new_n961), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n984), .A2(new_n980), .ZN(new_n985));
  XNOR2_X1  g0785(.A(new_n983), .B(new_n985), .ZN(new_n986));
  XOR2_X1   g0786(.A(new_n694), .B(KEYINPUT41), .Z(new_n987));
  INV_X1    g0787(.A(KEYINPUT44), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n691), .A2(new_n988), .A3(new_n961), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n988), .B1(new_n691), .B2(new_n961), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n989), .A2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n961), .B1(new_n689), .B2(new_n690), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(KEYINPUT107), .ZN(new_n993));
  INV_X1    g0793(.A(KEYINPUT107), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n994), .B(new_n961), .C1(new_n689), .C2(new_n690), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n993), .A2(KEYINPUT45), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n993), .A2(new_n995), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT45), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g0799(.A1(new_n991), .A2(new_n996), .A3(new_n999), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n1000), .A2(new_n981), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n685), .A2(new_n672), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n1002), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n686), .B1(new_n676), .B2(new_n1003), .ZN(new_n1004));
  XOR2_X1   g0804(.A(new_n744), .B(new_n1004), .Z(new_n1005));
  NAND4_X1  g0805(.A1(new_n991), .A2(new_n684), .A3(new_n996), .A4(new_n999), .ZN(new_n1006));
  NAND4_X1  g0806(.A1(new_n1001), .A2(new_n741), .A3(new_n1005), .A4(new_n1006), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n987), .B1(new_n1007), .B2(new_n741), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n986), .B1(new_n1008), .B2(new_n748), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n232), .A2(new_n761), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n756), .B1(new_n213), .B2(new_n376), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n749), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT108), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n805), .A2(new_n451), .ZN(new_n1014));
  XNOR2_X1  g0814(.A(new_n1014), .B(KEYINPUT46), .ZN(new_n1015));
  OAI22_X1  g0815(.A1(new_n780), .A2(new_n611), .B1(new_n205), .B2(new_n797), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n799), .A2(new_n820), .B1(new_n861), .B2(new_n206), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g0818(.A1(new_n787), .A2(G283), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n794), .A2(G303), .ZN(new_n1020));
  XOR2_X1   g0820(.A(KEYINPUT109), .B(G317), .Z(new_n1021));
  AOI21_X1  g0821(.A(new_n759), .B1(new_n815), .B2(new_n1021), .ZN(new_n1022));
  NAND4_X1  g0822(.A1(new_n1018), .A2(new_n1019), .A3(new_n1020), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g0823(.A(G137), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n274), .B1(new_n790), .B2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(G143), .B2(new_n798), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1026), .B1(new_n786), .B2(new_n202), .C1(new_n350), .C2(new_n793), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n797), .A2(new_n367), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(G68), .B2(new_n775), .ZN(new_n1029));
  OAI221_X1 g0829(.A(new_n1029), .B1(new_n791), .B2(new_n780), .C1(new_n805), .C2(new_n250), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n1015), .A2(new_n1023), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  INV_X1    g0831(.A(KEYINPUT47), .ZN(new_n1032));
  OR2_X1    g0832(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n772), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1034));
  AOI21_X1  g0834(.A(new_n1013), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  OAI21_X1  g0835(.A(new_n1035), .B1(new_n972), .B2(new_n825), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1009), .A2(new_n1036), .ZN(new_n1037));
  INV_X1    g0837(.A(KEYINPUT110), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1009), .A2(KEYINPUT110), .A3(new_n1036), .ZN(new_n1040));
  AND2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(G387));
  AOI21_X1  g0841(.A(new_n695), .B1(new_n1005), .B2(new_n741), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1042), .B1(new_n741), .B2(new_n1005), .ZN(new_n1043));
  NOR2_X1   g0843(.A1(new_n676), .A2(new_n825), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n766), .A2(new_n696), .B1(G107), .B2(new_n213), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n237), .A2(new_n301), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n696), .ZN(new_n1047));
  AOI211_X1 g0847(.A(G45), .B(new_n1047), .C1(G68), .C2(G77), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n285), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(KEYINPUT111), .B(KEYINPUT50), .ZN(new_n1050));
  XNOR2_X1  g0850(.A(new_n1049), .B(new_n1050), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n761), .B1(new_n1048), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1045), .B1(new_n1046), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n749), .B1(new_n1053), .B2(new_n757), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n805), .A2(new_n367), .ZN(new_n1055));
  OAI22_X1  g0855(.A1(new_n780), .A2(new_n285), .B1(new_n205), .B2(new_n797), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n799), .A2(new_n791), .B1(new_n861), .B2(new_n376), .ZN(new_n1057));
  NOR3_X1   g0857(.A1(new_n1055), .A2(new_n1056), .A3(new_n1057), .ZN(new_n1058));
  OAI21_X1  g0858(.A(new_n759), .B1(new_n350), .B2(new_n790), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1059), .B1(new_n794), .B2(G50), .ZN(new_n1060));
  OAI211_X1 g0860(.A(new_n1058), .B(new_n1060), .C1(new_n244), .C2(new_n786), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n759), .B1(G326), .B2(new_n815), .ZN(new_n1062));
  OAI22_X1  g0862(.A1(new_n805), .A2(new_n611), .B1(new_n817), .B2(new_n861), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n787), .A2(G303), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n794), .A2(new_n1021), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G311), .A2(new_n779), .B1(new_n798), .B2(G322), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1064), .A2(new_n1065), .A3(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1063), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1062), .B1(new_n451), .B2(new_n797), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1061), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI211_X1 g0874(.A(new_n1044), .B(new_n1054), .C1(new_n1074), .C2(new_n755), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n1075), .B1(new_n1005), .B2(new_n748), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1043), .A2(new_n1076), .ZN(G393));
  INV_X1    g0877(.A(new_n1001), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1006), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1078), .A2(new_n1079), .ZN(new_n1080));
  OR2_X1    g0880(.A1(new_n961), .A2(new_n825), .ZN(new_n1081));
  OAI22_X1  g0881(.A1(new_n793), .A2(new_n791), .B1(new_n350), .B2(new_n799), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT112), .Z(new_n1083));
  OR2_X1    g0883(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1083), .A2(KEYINPUT51), .ZN(new_n1085));
  OAI22_X1  g0885(.A1(new_n786), .A2(new_n285), .B1(new_n202), .B2(new_n780), .ZN(new_n1086));
  XOR2_X1   g0886(.A(new_n1086), .B(KEYINPUT113), .Z(new_n1087));
  AOI21_X1  g0887(.A(new_n263), .B1(new_n815), .B2(G143), .ZN(new_n1088));
  OAI211_X1 g0888(.A(new_n1088), .B(new_n852), .C1(new_n367), .C2(new_n861), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n1089), .B1(G68), .B2(new_n806), .ZN(new_n1090));
  NAND4_X1  g0890(.A1(new_n1084), .A2(new_n1085), .A3(new_n1087), .A4(new_n1090), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n794), .A2(G311), .B1(G317), .B2(new_n798), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT52), .Z(new_n1093));
  AOI21_X1  g0893(.A(new_n274), .B1(new_n815), .B2(G322), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n1094), .B1(new_n206), .B2(new_n797), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n779), .A2(G303), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n451), .B2(new_n861), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G294), .C2(new_n787), .ZN(new_n1098));
  OAI211_X1 g0898(.A(new_n1093), .B(new_n1098), .C1(new_n817), .C2(new_n805), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n772), .B1(new_n1091), .B2(new_n1099), .ZN(new_n1100));
  OR2_X1    g0900(.A1(new_n761), .A2(new_n241), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n757), .B1(G97), .B2(new_n693), .ZN(new_n1102));
  AOI211_X1 g0902(.A(new_n750), .B(new_n1100), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n1080), .A2(new_n748), .B1(new_n1081), .B2(new_n1104), .ZN(new_n1105));
  NAND2_X1  g0905(.A1(new_n1005), .A2(new_n741), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n1106), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1107), .A2(new_n694), .A3(new_n1007), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1105), .A2(new_n1108), .ZN(G390));
  NAND2_X1  g0909(.A1(new_n936), .A2(new_n937), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n929), .A2(new_n932), .ZN(new_n1111));
  INV_X1    g0911(.A(new_n939), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1111), .A2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1110), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n710), .A2(new_n672), .A3(new_n837), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1115), .A2(new_n829), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(new_n932), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n934), .A2(new_n1112), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1118), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1117), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n740), .A2(new_n837), .A3(new_n932), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(KEYINPUT115), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT115), .ZN(new_n1123));
  NAND4_X1  g0923(.A1(new_n740), .A2(new_n932), .A3(new_n1123), .A4(new_n837), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT116), .ZN(new_n1126));
  NAND4_X1  g0926(.A1(new_n1114), .A2(new_n1120), .A3(new_n1125), .A4(new_n1126), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n932), .A2(new_n837), .ZN(new_n1128));
  AOI211_X1 g0928(.A(new_n716), .B(new_n1128), .C1(new_n924), .C2(new_n923), .ZN(new_n1129));
  AOI22_X1  g0929(.A1(new_n936), .A2(new_n937), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1118), .B1(new_n932), .B2(new_n1116), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1129), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1127), .A2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n1110), .A2(new_n1113), .B1(new_n1117), .B2(new_n1119), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1126), .B1(new_n1134), .B2(new_n1125), .ZN(new_n1135));
  OR2_X1    g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  NAND3_X1  g0936(.A1(new_n925), .A2(G330), .A3(new_n837), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n901), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1116), .B1(new_n1122), .B2(new_n1124), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n932), .B1(new_n740), .B2(new_n837), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n929), .B1(new_n1129), .B2(new_n1141), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n716), .B1(new_n923), .B2(new_n924), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1144), .A2(new_n450), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1145), .A2(new_n943), .A3(new_n659), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n1146), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n695), .B1(new_n1136), .B2(new_n1148), .ZN(new_n1149));
  NOR2_X1   g0949(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1146), .B1(new_n1140), .B2(new_n1142), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n1150), .A2(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1149), .A2(new_n1152), .ZN(new_n1153));
  NAND2_X1  g0953(.A1(new_n1150), .A2(new_n748), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n750), .B1(new_n285), .B2(new_n845), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT117), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n277), .B1(new_n815), .B2(G125), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n202), .B2(new_n797), .ZN(new_n1158));
  XOR2_X1   g0958(.A(new_n1158), .B(KEYINPUT118), .Z(new_n1159));
  NAND2_X1  g0959(.A1(new_n779), .A2(G137), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n798), .A2(G128), .B1(new_n775), .B2(G159), .ZN(new_n1161));
  XOR2_X1   g0961(.A(KEYINPUT54), .B(G143), .Z(new_n1162));
  AOI22_X1  g0962(.A1(G132), .A2(new_n794), .B1(new_n787), .B2(new_n1162), .ZN(new_n1163));
  NAND4_X1  g0963(.A1(new_n1159), .A2(new_n1160), .A3(new_n1161), .A4(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n806), .A2(G150), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  OAI21_X1  g0966(.A(new_n277), .B1(new_n790), .B2(new_n611), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(G68), .B2(new_n851), .ZN(new_n1168));
  OAI221_X1 g0968(.A(new_n1168), .B1(new_n786), .B2(new_n205), .C1(new_n451), .C2(new_n793), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(new_n798), .A2(G283), .B1(new_n775), .B2(G77), .ZN(new_n1170));
  INV_X1    g0970(.A(G87), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1170), .B1(new_n206), .B2(new_n780), .C1(new_n805), .C2(new_n1171), .ZN(new_n1172));
  OAI22_X1  g0972(.A1(new_n1164), .A2(new_n1166), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1156), .B1(new_n1173), .B2(new_n755), .ZN(new_n1174));
  INV_X1    g0974(.A(new_n1110), .ZN(new_n1175));
  OAI21_X1  g0975(.A(new_n1174), .B1(new_n1175), .B2(new_n753), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1153), .A2(new_n1154), .A3(new_n1176), .ZN(G378));
  INV_X1    g0977(.A(KEYINPUT123), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n875), .A2(new_n359), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n374), .A2(new_n403), .A3(new_n1180), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n1181), .ZN(new_n1182));
  AOI21_X1  g0982(.A(new_n1180), .B1(new_n374), .B2(new_n403), .ZN(new_n1183));
  OAI21_X1  g0983(.A(KEYINPUT122), .B1(new_n1182), .B2(new_n1183), .ZN(new_n1184));
  INV_X1    g0984(.A(new_n1183), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT122), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1185), .A2(new_n1186), .A3(new_n1181), .ZN(new_n1187));
  XOR2_X1   g0987(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1188));
  NAND3_X1  g0988(.A1(new_n1184), .A2(new_n1187), .A3(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1184), .B2(new_n1187), .ZN(new_n1191));
  NOR2_X1   g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n877), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n347), .A2(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(KEYINPUT38), .B1(new_n1194), .B2(new_n885), .ZN(new_n1195));
  INV_X1    g0995(.A(new_n890), .ZN(new_n1196));
  OAI21_X1  g0996(.A(KEYINPUT101), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n887), .A2(new_n888), .A3(new_n890), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(new_n1198), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1128), .B1(new_n923), .B2(new_n924), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT40), .B1(new_n1199), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n920), .A2(G330), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1192), .B1(new_n1201), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n716), .B1(new_n1200), .B2(new_n919), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1184), .A2(new_n1187), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n1188), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1205), .A2(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1207), .A2(new_n1189), .ZN(new_n1208));
  AOI21_X1  g1008(.A(new_n912), .B1(new_n1197), .B2(new_n1198), .ZN(new_n1209));
  OAI211_X1 g1009(.A(new_n1204), .B(new_n1208), .C1(new_n1209), .C2(KEYINPUT40), .ZN(new_n1210));
  INV_X1    g1010(.A(new_n942), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1203), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1211), .B1(new_n1203), .B2(new_n1210), .ZN(new_n1213));
  OAI21_X1  g1013(.A(new_n1178), .B1(new_n1212), .B2(new_n1213), .ZN(new_n1214));
  NOR3_X1   g1014(.A1(new_n1201), .A2(new_n1192), .A3(new_n1202), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n1208), .B1(new_n913), .B2(new_n1204), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n942), .B1(new_n1215), .B2(new_n1216), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1203), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(KEYINPUT123), .A3(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1214), .A2(new_n1219), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1146), .B1(new_n1150), .B2(new_n1143), .ZN(new_n1221));
  INV_X1    g1021(.A(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(KEYINPUT57), .B1(new_n1220), .B2(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1217), .A2(new_n1218), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT57), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n694), .B1(new_n1225), .B2(new_n1221), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1223), .A2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n750), .B1(new_n202), .B2(new_n845), .ZN(new_n1229));
  AOI21_X1  g1029(.A(G41), .B1(new_n759), .B2(G33), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n1230), .A2(G50), .ZN(new_n1231));
  AOI211_X1 g1031(.A(G41), .B(new_n759), .C1(G283), .C2(new_n815), .ZN(new_n1232));
  OAI221_X1 g1032(.A(new_n1232), .B1(new_n786), .B2(new_n376), .C1(new_n206), .C2(new_n793), .ZN(new_n1233));
  AOI22_X1  g1033(.A1(G58), .A2(new_n851), .B1(new_n775), .B2(G68), .ZN(new_n1234));
  OAI221_X1 g1034(.A(new_n1234), .B1(new_n780), .B2(new_n205), .C1(new_n451), .C2(new_n799), .ZN(new_n1235));
  NOR3_X1   g1035(.A1(new_n1233), .A2(new_n1055), .A3(new_n1235), .ZN(new_n1236));
  XNOR2_X1  g1036(.A(KEYINPUT119), .B(KEYINPUT58), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1237), .ZN(new_n1238));
  AOI21_X1  g1038(.A(new_n1231), .B1(new_n1236), .B2(new_n1238), .ZN(new_n1239));
  OAI21_X1  g1039(.A(new_n1239), .B1(new_n1238), .B2(new_n1236), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n806), .A2(new_n1162), .ZN(new_n1241));
  OR2_X1    g1041(.A1(new_n1241), .A2(KEYINPUT120), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(KEYINPUT120), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n779), .A2(G132), .ZN(new_n1244));
  OAI21_X1  g1044(.A(new_n1244), .B1(new_n350), .B2(new_n861), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1245), .B1(G125), .B2(new_n798), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(G128), .A2(new_n794), .B1(new_n787), .B2(G137), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1243), .A3(new_n1246), .A4(new_n1247), .ZN(new_n1248));
  XNOR2_X1  g1048(.A(new_n1248), .B(KEYINPUT121), .ZN(new_n1249));
  OR2_X1    g1049(.A1(new_n1249), .A2(KEYINPUT59), .ZN(new_n1250));
  AOI211_X1 g1050(.A(G33), .B(G41), .C1(new_n815), .C2(G124), .ZN(new_n1251));
  OAI21_X1  g1051(.A(new_n1251), .B1(new_n791), .B2(new_n797), .ZN(new_n1252));
  AOI21_X1  g1052(.A(new_n1252), .B1(new_n1249), .B2(KEYINPUT59), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1240), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1254));
  OAI221_X1 g1054(.A(new_n1229), .B1(new_n772), .B2(new_n1254), .C1(new_n1208), .C2(new_n753), .ZN(new_n1255));
  INV_X1    g1055(.A(new_n1255), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1220), .B2(new_n748), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1228), .A2(new_n1257), .ZN(G375));
  NOR2_X1   g1058(.A1(new_n1143), .A2(new_n1147), .ZN(new_n1259));
  NOR3_X1   g1059(.A1(new_n1259), .A2(new_n987), .A3(new_n1151), .ZN(new_n1260));
  XNOR2_X1  g1060(.A(new_n1260), .B(KEYINPUT124), .ZN(new_n1261));
  AOI211_X1 g1061(.A(new_n274), .B(new_n1028), .C1(G303), .C2(new_n815), .ZN(new_n1262));
  OAI221_X1 g1062(.A(new_n1262), .B1(new_n206), .B2(new_n786), .C1(new_n817), .C2(new_n793), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n376), .ZN(new_n1264));
  AOI22_X1  g1064(.A1(new_n798), .A2(G294), .B1(new_n775), .B2(new_n1264), .ZN(new_n1265));
  OAI221_X1 g1065(.A(new_n1265), .B1(new_n451), .B2(new_n780), .C1(new_n805), .C2(new_n205), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n263), .B1(new_n815), .B2(G128), .ZN(new_n1267));
  OAI221_X1 g1067(.A(new_n1267), .B1(new_n786), .B2(new_n350), .C1(new_n1024), .C2(new_n793), .ZN(new_n1268));
  AOI22_X1  g1068(.A1(new_n798), .A2(G132), .B1(new_n851), .B2(G58), .ZN(new_n1269));
  AOI22_X1  g1069(.A1(new_n779), .A2(new_n1162), .B1(new_n775), .B2(G50), .ZN(new_n1270));
  OAI211_X1 g1070(.A(new_n1269), .B(new_n1270), .C1(new_n805), .C2(new_n791), .ZN(new_n1271));
  OAI22_X1  g1071(.A1(new_n1263), .A2(new_n1266), .B1(new_n1268), .B2(new_n1271), .ZN(new_n1272));
  NAND2_X1  g1072(.A1(new_n1272), .A2(new_n755), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n750), .B1(new_n244), .B2(new_n845), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n1273), .B(new_n1274), .C1(new_n932), .C2(new_n753), .ZN(new_n1275));
  AND2_X1   g1075(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1275), .B1(new_n1276), .B2(new_n747), .ZN(new_n1277));
  NOR2_X1   g1077(.A1(new_n1261), .A2(new_n1277), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1278), .ZN(G381));
  INV_X1    g1079(.A(G387), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1154), .A2(new_n1176), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1281), .B1(new_n1152), .B2(new_n1149), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(new_n1043), .A2(new_n827), .A3(new_n1076), .ZN(new_n1283));
  NOR3_X1   g1083(.A1(G390), .A2(G384), .A3(new_n1283), .ZN(new_n1284));
  NAND4_X1  g1084(.A1(new_n1280), .A2(new_n1282), .A3(new_n1278), .A4(new_n1284), .ZN(new_n1285));
  OR2_X1    g1085(.A1(new_n1285), .A2(G375), .ZN(G407));
  NOR2_X1   g1086(.A1(new_n664), .A2(G343), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1282), .A2(new_n1287), .ZN(new_n1288));
  OAI211_X1 g1088(.A(G407), .B(G213), .C1(G375), .C2(new_n1288), .ZN(G409));
  INV_X1    g1089(.A(G390), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1037), .A2(new_n1290), .ZN(new_n1291));
  NAND2_X1  g1091(.A1(new_n1291), .A2(KEYINPUT125), .ZN(new_n1292));
  INV_X1    g1092(.A(KEYINPUT125), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1037), .A2(new_n1290), .A3(new_n1293), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(G390), .A2(new_n1009), .A3(new_n1036), .ZN(new_n1295));
  NAND3_X1  g1095(.A1(new_n1292), .A2(new_n1294), .A3(new_n1295), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(G393), .A2(G396), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1297), .A2(new_n1283), .ZN(new_n1298));
  INV_X1    g1098(.A(new_n1298), .ZN(new_n1299));
  NAND3_X1  g1099(.A1(new_n1039), .A2(new_n1040), .A3(new_n1290), .ZN(new_n1300));
  AND2_X1   g1100(.A1(new_n1295), .A2(new_n1298), .ZN(new_n1301));
  AOI22_X1  g1101(.A1(new_n1296), .A2(new_n1299), .B1(new_n1300), .B2(new_n1301), .ZN(new_n1302));
  XNOR2_X1  g1102(.A(new_n1302), .B(KEYINPUT127), .ZN(new_n1303));
  OAI211_X1 g1103(.A(G378), .B(new_n1257), .C1(new_n1223), .C2(new_n1226), .ZN(new_n1304));
  AOI211_X1 g1104(.A(new_n987), .B(new_n1221), .C1(new_n1214), .C2(new_n1219), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1224), .A2(new_n748), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1306), .A2(new_n1255), .ZN(new_n1307));
  OAI21_X1  g1107(.A(new_n1282), .B1(new_n1305), .B2(new_n1307), .ZN(new_n1308));
  NAND2_X1  g1108(.A1(new_n1304), .A2(new_n1308), .ZN(new_n1309));
  INV_X1    g1109(.A(KEYINPUT62), .ZN(new_n1310));
  INV_X1    g1110(.A(new_n1287), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n1259), .B1(KEYINPUT60), .B2(new_n1148), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1276), .A2(KEYINPUT60), .A3(new_n1146), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(new_n694), .ZN(new_n1314));
  NOR2_X1   g1114(.A1(new_n1312), .A2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n866), .B1(new_n1315), .B2(new_n1277), .ZN(new_n1316));
  AND2_X1   g1116(.A1(new_n1313), .A2(new_n694), .ZN(new_n1317));
  NAND2_X1  g1117(.A1(new_n1148), .A2(KEYINPUT60), .ZN(new_n1318));
  INV_X1    g1118(.A(new_n1259), .ZN(new_n1319));
  NAND2_X1  g1119(.A1(new_n1318), .A2(new_n1319), .ZN(new_n1320));
  NAND2_X1  g1120(.A1(new_n1317), .A2(new_n1320), .ZN(new_n1321));
  INV_X1    g1121(.A(new_n1277), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1321), .A2(G384), .A3(new_n1322), .ZN(new_n1323));
  NAND2_X1  g1123(.A1(new_n1316), .A2(new_n1323), .ZN(new_n1324));
  INV_X1    g1124(.A(new_n1324), .ZN(new_n1325));
  NAND4_X1  g1125(.A1(new_n1309), .A2(new_n1310), .A3(new_n1311), .A4(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(KEYINPUT61), .ZN(new_n1327));
  AOI21_X1  g1127(.A(new_n1287), .B1(new_n1304), .B2(new_n1308), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1287), .A2(G2897), .ZN(new_n1329));
  INV_X1    g1129(.A(new_n1329), .ZN(new_n1330));
  AOI21_X1  g1130(.A(G384), .B1(new_n1321), .B2(new_n1322), .ZN(new_n1331));
  AOI211_X1 g1131(.A(new_n866), .B(new_n1277), .C1(new_n1317), .C2(new_n1320), .ZN(new_n1332));
  OAI21_X1  g1132(.A(new_n1330), .B1(new_n1331), .B2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1316), .A2(new_n1323), .A3(new_n1329), .ZN(new_n1334));
  NAND2_X1  g1134(.A1(new_n1333), .A2(new_n1334), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1326), .B(new_n1327), .C1(new_n1328), .C2(new_n1335), .ZN(new_n1336));
  AOI211_X1 g1136(.A(new_n1287), .B(new_n1324), .C1(new_n1304), .C2(new_n1308), .ZN(new_n1337));
  NOR2_X1   g1137(.A1(new_n1337), .A2(new_n1310), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1303), .B1(new_n1336), .B2(new_n1338), .ZN(new_n1339));
  OAI21_X1  g1139(.A(KEYINPUT63), .B1(new_n1328), .B2(new_n1335), .ZN(new_n1340));
  NAND2_X1  g1140(.A1(new_n1328), .A2(new_n1325), .ZN(new_n1341));
  NAND2_X1  g1141(.A1(new_n1340), .A2(new_n1341), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(new_n1337), .A2(KEYINPUT63), .ZN(new_n1343));
  INV_X1    g1143(.A(KEYINPUT126), .ZN(new_n1344));
  OAI21_X1  g1144(.A(new_n1344), .B1(new_n1302), .B2(KEYINPUT61), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1296), .A2(new_n1299), .ZN(new_n1346));
  AND2_X1   g1146(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1347));
  OAI211_X1 g1147(.A(KEYINPUT126), .B(new_n1327), .C1(new_n1346), .C2(new_n1347), .ZN(new_n1348));
  NAND4_X1  g1148(.A1(new_n1342), .A2(new_n1343), .A3(new_n1345), .A4(new_n1348), .ZN(new_n1349));
  NAND2_X1  g1149(.A1(new_n1339), .A2(new_n1349), .ZN(G405));
  NAND2_X1  g1150(.A1(G375), .A2(new_n1282), .ZN(new_n1351));
  NAND3_X1  g1151(.A1(new_n1351), .A2(new_n1304), .A3(new_n1324), .ZN(new_n1352));
  AOI21_X1  g1152(.A(G378), .B1(new_n1228), .B2(new_n1257), .ZN(new_n1353));
  INV_X1    g1153(.A(new_n1304), .ZN(new_n1354));
  OAI21_X1  g1154(.A(new_n1325), .B1(new_n1353), .B2(new_n1354), .ZN(new_n1355));
  AND3_X1   g1155(.A1(new_n1352), .A2(new_n1302), .A3(new_n1355), .ZN(new_n1356));
  AOI21_X1  g1156(.A(new_n1302), .B1(new_n1352), .B2(new_n1355), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1356), .A2(new_n1357), .ZN(G402));
endmodule


