//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:25 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n737, new_n738, new_n739, new_n740, new_n742,
    new_n743, new_n744, new_n745, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n757,
    new_n758, new_n759, new_n760, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n780,
    new_n781, new_n782, new_n783, new_n784, new_n785, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n822, new_n823, new_n824, new_n825, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n874, new_n875, new_n876, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n920, new_n921, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n964, new_n965,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n980, new_n981, new_n983,
    new_n984, new_n985, new_n986, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n994, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1004, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027;
  NAND2_X1  g000(.A1(KEYINPUT69), .A2(G127gat), .ZN(new_n202));
  INV_X1    g001(.A(G120gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G113gat), .ZN(new_n204));
  INV_X1    g003(.A(G113gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G120gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT1), .ZN(new_n208));
  AOI21_X1  g007(.A(new_n202), .B1(new_n207), .B2(new_n208), .ZN(new_n209));
  AOI211_X1 g008(.A(KEYINPUT1), .B(G127gat), .C1(new_n204), .C2(new_n206), .ZN(new_n210));
  OAI21_X1  g009(.A(G134gat), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n202), .ZN(new_n212));
  XNOR2_X1  g011(.A(G113gat), .B(G120gat), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n212), .B1(new_n213), .B2(KEYINPUT1), .ZN(new_n214));
  INV_X1    g013(.A(G134gat), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n205), .A2(G120gat), .ZN(new_n217));
  NOR2_X1   g016(.A1(new_n203), .A2(G113gat), .ZN(new_n218));
  OAI211_X1 g017(.A(new_n208), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n211), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT24), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT64), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(KEYINPUT64), .ZN(new_n228));
  INV_X1    g027(.A(G183gat), .ZN(new_n229));
  INV_X1    g028(.A(G190gat), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n229), .A2(new_n230), .ZN(new_n231));
  NAND3_X1  g030(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n226), .A2(new_n228), .A3(new_n231), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT23), .ZN(new_n234));
  NOR3_X1   g033(.A1(new_n234), .A2(G169gat), .A3(G176gat), .ZN(new_n235));
  INV_X1    g034(.A(G169gat), .ZN(new_n236));
  INV_X1    g035(.A(G176gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n236), .A2(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(G169gat), .A2(G176gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n239), .A2(KEYINPUT23), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n235), .B1(new_n238), .B2(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT25), .B1(new_n233), .B2(new_n241), .ZN(new_n242));
  INV_X1    g041(.A(KEYINPUT25), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n243), .B1(new_n240), .B2(new_n238), .ZN(new_n244));
  NAND3_X1  g043(.A1(new_n236), .A2(new_n237), .A3(KEYINPUT65), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT65), .ZN(new_n246));
  OAI21_X1  g045(.A(new_n246), .B1(G169gat), .B2(G176gat), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT23), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n244), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT67), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n232), .A2(KEYINPUT66), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT66), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n252), .A2(KEYINPUT24), .A3(G183gat), .A4(G190gat), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n251), .A2(new_n253), .A3(new_n224), .A4(new_n231), .ZN(new_n254));
  AOI21_X1  g053(.A(new_n249), .B1(new_n250), .B2(new_n254), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n227), .B1(new_n229), .B2(new_n230), .ZN(new_n256));
  NAND4_X1  g055(.A1(new_n256), .A2(KEYINPUT67), .A3(new_n253), .A4(new_n251), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n242), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(new_n229), .A2(KEYINPUT27), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT27), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(G183gat), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n259), .A2(new_n261), .A3(new_n230), .ZN(new_n262));
  NOR2_X1   g061(.A1(KEYINPUT68), .A2(KEYINPUT28), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT27), .B(G183gat), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(new_n230), .A3(new_n263), .ZN(new_n267));
  AND3_X1   g066(.A1(new_n265), .A2(new_n267), .A3(new_n222), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n238), .A2(KEYINPUT26), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n245), .A2(new_n247), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n239), .B(new_n269), .C1(new_n270), .C2(KEYINPUT26), .ZN(new_n271));
  AND2_X1   g070(.A1(new_n268), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n221), .B1(new_n258), .B2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G227gat), .ZN(new_n274));
  INV_X1    g073(.A(G233gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  AND2_X1   g075(.A1(new_n244), .A2(new_n248), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n254), .A2(new_n250), .ZN(new_n278));
  NAND3_X1  g077(.A1(new_n277), .A2(new_n257), .A3(new_n278), .ZN(new_n279));
  OAI211_X1 g078(.A(new_n231), .B(new_n232), .C1(new_n227), .C2(KEYINPUT64), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n224), .A2(new_n225), .ZN(new_n281));
  NOR2_X1   g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n240), .A2(new_n238), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n283), .B1(new_n234), .B2(new_n238), .ZN(new_n284));
  OAI21_X1  g083(.A(new_n243), .B1(new_n282), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n279), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n268), .A2(new_n271), .ZN(new_n287));
  NAND4_X1  g086(.A1(new_n286), .A2(new_n211), .A3(new_n220), .A4(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n273), .A2(new_n276), .A3(new_n288), .ZN(new_n289));
  INV_X1    g088(.A(KEYINPUT33), .ZN(new_n290));
  XNOR2_X1  g089(.A(G15gat), .B(G43gat), .ZN(new_n291));
  XNOR2_X1  g090(.A(new_n291), .B(KEYINPUT70), .ZN(new_n292));
  XNOR2_X1  g091(.A(G71gat), .B(G99gat), .ZN(new_n293));
  XNOR2_X1  g092(.A(new_n292), .B(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(new_n294), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n289), .B(KEYINPUT32), .C1(new_n290), .C2(new_n295), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n295), .B1(new_n289), .B2(KEYINPUT32), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n289), .A2(new_n290), .ZN(new_n298));
  AND3_X1   g097(.A1(new_n297), .A2(KEYINPUT71), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT71), .B1(new_n297), .B2(new_n298), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n296), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n273), .A2(new_n288), .ZN(new_n302));
  INV_X1    g101(.A(new_n276), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT72), .ZN(new_n305));
  XNOR2_X1  g104(.A(new_n305), .B(KEYINPUT34), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n289), .A2(KEYINPUT32), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n308), .A2(new_n298), .A3(new_n294), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT71), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n297), .A2(KEYINPUT71), .A3(new_n298), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n305), .A2(KEYINPUT34), .ZN(new_n314));
  INV_X1    g113(.A(KEYINPUT34), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n304), .B2(KEYINPUT72), .ZN(new_n316));
  NOR2_X1   g115(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n313), .A2(new_n317), .A3(new_n296), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n307), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT36), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n307), .A2(new_n318), .A3(KEYINPUT36), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(G228gat), .ZN(new_n324));
  NOR2_X1   g123(.A1(new_n324), .A2(new_n275), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  XOR2_X1   g125(.A(G141gat), .B(G148gat), .Z(new_n327));
  INV_X1    g126(.A(KEYINPUT2), .ZN(new_n328));
  AND2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(G155gat), .ZN(new_n330));
  INV_X1    g129(.A(G162gat), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(G155gat), .A2(G162gat), .ZN(new_n333));
  NOR3_X1   g132(.A1(new_n329), .A2(new_n332), .A3(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(G148gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT78), .B1(new_n335), .B2(G141gat), .ZN(new_n336));
  AND2_X1   g135(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n336), .B1(new_n339), .B2(G141gat), .ZN(new_n340));
  INV_X1    g139(.A(G141gat), .ZN(new_n341));
  NOR4_X1   g140(.A1(new_n337), .A2(new_n338), .A3(KEYINPUT78), .A4(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(KEYINPUT79), .B1(new_n340), .B2(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(KEYINPUT77), .A2(G148gat), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(G141gat), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(new_n336), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n349));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n350));
  NAND4_X1  g149(.A1(new_n344), .A2(new_n350), .A3(G141gat), .A4(new_n345), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n343), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g152(.A(new_n332), .B1(new_n328), .B2(new_n333), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n334), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT3), .ZN(new_n357));
  NAND2_X1  g156(.A1(G211gat), .A2(G218gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT22), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g159(.A1(new_n360), .A2(KEYINPUT73), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT73), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n358), .A2(new_n362), .A3(new_n359), .ZN(new_n363));
  XNOR2_X1  g162(.A(G197gat), .B(G204gat), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n361), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  XNOR2_X1  g164(.A(G211gat), .B(G218gat), .ZN(new_n366));
  INV_X1    g165(.A(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n361), .A2(new_n366), .A3(new_n364), .A4(new_n363), .ZN(new_n369));
  AOI21_X1  g168(.A(KEYINPUT29), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n357), .B1(new_n370), .B2(KEYINPUT83), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT83), .ZN(new_n373));
  AOI211_X1 g172(.A(new_n373), .B(KEYINPUT29), .C1(new_n368), .C2(new_n369), .ZN(new_n374));
  INV_X1    g173(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n356), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n368), .A2(new_n369), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT74), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(new_n368), .A2(KEYINPUT74), .A3(new_n369), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AND3_X1   g180(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n382));
  AOI21_X1  g181(.A(new_n349), .B1(new_n348), .B2(new_n351), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n355), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(new_n334), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n385), .A3(new_n357), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT29), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n381), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n326), .B1(new_n376), .B2(new_n388), .ZN(new_n389));
  AOI21_X1  g188(.A(new_n354), .B1(new_n343), .B2(new_n352), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT3), .B1(new_n390), .B2(new_n334), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n370), .B1(new_n390), .B2(new_n334), .ZN(new_n392));
  AND3_X1   g191(.A1(new_n391), .A2(new_n392), .A3(new_n325), .ZN(new_n393));
  INV_X1    g192(.A(new_n381), .ZN(new_n394));
  NOR3_X1   g193(.A1(new_n390), .A2(KEYINPUT3), .A3(new_n334), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(KEYINPUT29), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n393), .A2(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G22gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n389), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n399), .A2(KEYINPUT84), .ZN(new_n400));
  XNOR2_X1  g199(.A(G78gat), .B(G106gat), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT31), .B(G50gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n401), .B(new_n402), .Z(new_n403));
  OAI22_X1  g202(.A1(new_n371), .A2(new_n374), .B1(new_n390), .B2(new_n334), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n325), .B1(new_n396), .B2(new_n404), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n391), .A2(new_n392), .A3(new_n325), .ZN(new_n406));
  NOR2_X1   g205(.A1(new_n406), .A2(new_n388), .ZN(new_n407));
  OAI21_X1  g206(.A(G22gat), .B1(new_n405), .B2(new_n407), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n400), .A2(new_n403), .B1(new_n399), .B2(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT84), .ZN(new_n410));
  NAND4_X1  g209(.A1(new_n408), .A2(new_n399), .A3(new_n410), .A4(new_n403), .ZN(new_n411));
  INV_X1    g210(.A(new_n411), .ZN(new_n412));
  NOR2_X1   g211(.A1(new_n409), .A2(new_n412), .ZN(new_n413));
  AND3_X1   g212(.A1(new_n214), .A2(new_n215), .A3(new_n219), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n215), .B1(new_n214), .B2(new_n219), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT80), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT80), .B1(new_n211), .B2(new_n220), .ZN(new_n418));
  NOR2_X1   g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND3_X1  g218(.A1(new_n419), .A2(new_n391), .A3(new_n386), .ZN(new_n420));
  NAND2_X1  g219(.A1(G225gat), .A2(G233gat), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n384), .A2(new_n385), .A3(new_n221), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT4), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n356), .A2(KEYINPUT4), .A3(new_n221), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n420), .A2(new_n421), .A3(new_n424), .A4(new_n425), .ZN(new_n426));
  OR2_X1    g225(.A1(new_n426), .A2(KEYINPUT5), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT81), .ZN(new_n428));
  AND2_X1   g227(.A1(new_n426), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT5), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n416), .B1(new_n414), .B2(new_n415), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n211), .A2(KEYINPUT80), .A3(new_n220), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n422), .B1(new_n433), .B2(new_n356), .ZN(new_n434));
  INV_X1    g233(.A(new_n421), .ZN(new_n435));
  AOI21_X1  g234(.A(new_n430), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n436), .B1(new_n426), .B2(new_n428), .ZN(new_n437));
  OAI21_X1  g236(.A(new_n427), .B1(new_n429), .B2(new_n437), .ZN(new_n438));
  XOR2_X1   g237(.A(G1gat), .B(G29gat), .Z(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT0), .ZN(new_n440));
  XNOR2_X1  g239(.A(G57gat), .B(G85gat), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n440), .B(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XOR2_X1   g242(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n444));
  INV_X1    g243(.A(new_n444), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n438), .A2(new_n443), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n426), .A2(new_n428), .ZN(new_n447));
  AOI21_X1  g246(.A(KEYINPUT4), .B1(new_n356), .B2(new_n221), .ZN(new_n448));
  AND4_X1   g247(.A1(KEYINPUT4), .A2(new_n384), .A3(new_n385), .A4(new_n221), .ZN(new_n449));
  NOR2_X1   g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n450), .A2(KEYINPUT81), .A3(new_n421), .A4(new_n420), .ZN(new_n451));
  AND3_X1   g250(.A1(new_n447), .A2(new_n451), .A3(new_n436), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n442), .B1(new_n426), .B2(KEYINPUT5), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n444), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n447), .A2(new_n451), .A3(new_n436), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n442), .B1(new_n455), .B2(new_n427), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G8gat), .B(G36gat), .ZN(new_n458));
  XNOR2_X1  g257(.A(G64gat), .B(G92gat), .ZN(new_n459));
  XOR2_X1   g258(.A(new_n458), .B(new_n459), .Z(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n286), .A2(new_n287), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  INV_X1    g262(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g263(.A(KEYINPUT76), .B1(new_n462), .B2(new_n464), .ZN(new_n465));
  AOI22_X1  g264(.A1(new_n279), .A2(new_n285), .B1(new_n268), .B2(new_n271), .ZN(new_n466));
  INV_X1    g265(.A(KEYINPUT76), .ZN(new_n467));
  NOR3_X1   g266(.A1(new_n466), .A2(new_n467), .A3(new_n463), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AND3_X1   g268(.A1(new_n286), .A2(KEYINPUT75), .A3(new_n287), .ZN(new_n470));
  AOI21_X1  g269(.A(KEYINPUT75), .B1(new_n286), .B2(new_n287), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n470), .A2(new_n471), .A3(KEYINPUT29), .ZN(new_n472));
  OAI211_X1 g271(.A(new_n469), .B(new_n394), .C1(new_n472), .C2(new_n464), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n462), .A2(new_n387), .A3(new_n463), .ZN(new_n474));
  NOR2_X1   g273(.A1(new_n470), .A2(new_n471), .ZN(new_n475));
  OAI211_X1 g274(.A(new_n381), .B(new_n474), .C1(new_n475), .C2(new_n463), .ZN(new_n476));
  AOI21_X1  g275(.A(new_n461), .B1(new_n473), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g276(.A1(new_n477), .A2(KEYINPUT30), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT30), .ZN(new_n479));
  AOI211_X1 g278(.A(new_n479), .B(new_n461), .C1(new_n473), .C2(new_n476), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n473), .A2(new_n476), .A3(new_n461), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR3_X1   g281(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  AOI21_X1  g282(.A(new_n413), .B1(new_n457), .B2(new_n483), .ZN(new_n484));
  NOR2_X1   g283(.A1(new_n323), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n461), .A2(KEYINPUT37), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n481), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n473), .A2(KEYINPUT37), .A3(new_n476), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT38), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n442), .B(KEYINPUT85), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n438), .A2(new_n492), .ZN(new_n493));
  INV_X1    g292(.A(new_n453), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n445), .B1(new_n455), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n469), .B1(new_n472), .B2(new_n464), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(new_n381), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT37), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n474), .B1(new_n475), .B2(new_n463), .ZN(new_n500));
  AOI21_X1  g299(.A(new_n499), .B1(new_n500), .B2(new_n394), .ZN(new_n501));
  AOI21_X1  g300(.A(KEYINPUT38), .B1(new_n498), .B2(new_n501), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n477), .B1(new_n502), .B2(new_n487), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n490), .A2(new_n496), .A3(new_n446), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT40), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n420), .A2(new_n424), .A3(new_n425), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT39), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n506), .A2(new_n507), .A3(new_n435), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n508), .A2(new_n491), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT39), .B1(new_n434), .B2(new_n435), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n510), .B1(new_n435), .B2(new_n506), .ZN(new_n511));
  OAI21_X1  g310(.A(new_n505), .B1(new_n509), .B2(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT86), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  OAI211_X1 g313(.A(KEYINPUT86), .B(new_n505), .C1(new_n509), .C2(new_n511), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g315(.A1(new_n473), .A2(new_n476), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n479), .B1(new_n517), .B2(new_n461), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n477), .A2(KEYINPUT30), .ZN(new_n519));
  NAND3_X1  g318(.A1(new_n518), .A2(new_n481), .A3(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n509), .A2(new_n511), .ZN(new_n521));
  AOI22_X1  g320(.A1(KEYINPUT40), .A2(new_n521), .B1(new_n438), .B2(new_n492), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n520), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n504), .A2(new_n523), .A3(new_n413), .ZN(new_n524));
  NAND4_X1  g323(.A1(new_n457), .A2(new_n319), .A3(new_n413), .A4(new_n483), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n525), .A2(KEYINPUT35), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n408), .A2(new_n399), .ZN(new_n527));
  AOI21_X1  g326(.A(KEYINPUT29), .B1(new_n356), .B2(new_n357), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n404), .B1(new_n528), .B2(new_n381), .ZN(new_n529));
  AOI22_X1  g328(.A1(new_n529), .A2(new_n326), .B1(new_n393), .B2(new_n396), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n410), .B1(new_n530), .B2(new_n398), .ZN(new_n531));
  INV_X1    g330(.A(new_n403), .ZN(new_n532));
  OAI21_X1  g331(.A(new_n527), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(new_n411), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n534), .B1(new_n318), .B2(new_n307), .ZN(new_n535));
  AOI21_X1  g334(.A(KEYINPUT35), .B1(new_n496), .B2(new_n446), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n535), .A2(new_n536), .A3(new_n483), .ZN(new_n537));
  AOI22_X1  g336(.A1(new_n485), .A2(new_n524), .B1(new_n526), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT92), .ZN(new_n539));
  XOR2_X1   g338(.A(G15gat), .B(G22gat), .Z(new_n540));
  NAND2_X1  g339(.A1(new_n540), .A2(KEYINPUT89), .ZN(new_n541));
  XNOR2_X1  g340(.A(G15gat), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT89), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT16), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  AOI21_X1  g346(.A(KEYINPUT90), .B1(new_n541), .B2(new_n544), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(G1gat), .B2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT90), .ZN(new_n550));
  INV_X1    g349(.A(new_n544), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n542), .A2(new_n543), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n550), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(G1gat), .ZN(new_n554));
  NOR2_X1   g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NOR3_X1   g354(.A1(new_n549), .A2(new_n555), .A3(G8gat), .ZN(new_n556));
  INV_X1    g355(.A(G8gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n553), .A2(new_n554), .B1(new_n546), .B2(new_n545), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n548), .A2(G1gat), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n539), .B1(new_n556), .B2(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(G29gat), .ZN(new_n562));
  INV_X1    g361(.A(G36gat), .ZN(new_n563));
  NAND3_X1  g362(.A1(new_n562), .A2(new_n563), .A3(KEYINPUT14), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT14), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n565), .B1(G29gat), .B2(G36gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(G29gat), .A2(G36gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT15), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n564), .A2(new_n566), .A3(KEYINPUT15), .A4(new_n567), .ZN(new_n571));
  XNOR2_X1  g370(.A(G43gat), .B(G50gat), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n570), .A2(new_n571), .A3(new_n572), .ZN(new_n573));
  OR2_X1    g372(.A1(new_n571), .A2(new_n572), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(KEYINPUT88), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(KEYINPUT88), .B1(new_n573), .B2(new_n574), .ZN(new_n577));
  NOR2_X1   g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  OAI21_X1  g377(.A(G8gat), .B1(new_n549), .B2(new_n555), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n558), .A2(new_n557), .A3(new_n559), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT92), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n561), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(KEYINPUT91), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n583), .B1(new_n556), .B2(new_n560), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT17), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n585), .B1(new_n576), .B2(new_n577), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n573), .A2(new_n574), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n587), .A2(KEYINPUT17), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n586), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n579), .A2(new_n580), .A3(KEYINPUT91), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n584), .A2(new_n589), .A3(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G229gat), .A2(G233gat), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n591), .A3(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT93), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT18), .ZN(new_n596));
  NAND4_X1  g395(.A1(new_n582), .A2(new_n591), .A3(KEYINPUT93), .A4(new_n592), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g397(.A(new_n592), .B(KEYINPUT13), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n561), .A2(new_n581), .ZN(new_n601));
  OR2_X1    g400(.A1(new_n576), .A2(new_n577), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n600), .B1(new_n603), .B2(new_n582), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n598), .A2(new_n605), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n582), .A2(new_n591), .A3(KEYINPUT18), .A4(new_n592), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT94), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XNOR2_X1  g408(.A(G113gat), .B(G141gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(G169gat), .B(G197gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(KEYINPUT87), .B(KEYINPUT11), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n612), .B(new_n613), .ZN(new_n614));
  XOR2_X1   g413(.A(new_n614), .B(KEYINPUT12), .Z(new_n615));
  NOR3_X1   g414(.A1(new_n606), .A2(new_n609), .A3(new_n615), .ZN(new_n616));
  INV_X1    g415(.A(new_n615), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT18), .B1(new_n593), .B2(new_n594), .ZN(new_n618));
  AOI21_X1  g417(.A(new_n604), .B1(new_n618), .B2(new_n597), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n607), .B(KEYINPUT94), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n617), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(G71gat), .A2(G78gat), .ZN(new_n623));
  OR2_X1    g422(.A1(G71gat), .A2(G78gat), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT9), .ZN(new_n625));
  OAI21_X1  g424(.A(new_n623), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(G57gat), .ZN(new_n627));
  OAI21_X1  g426(.A(G64gat), .B1(new_n627), .B2(KEYINPUT95), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT95), .ZN(new_n629));
  INV_X1    g428(.A(G64gat), .ZN(new_n630));
  NAND3_X1  g429(.A1(new_n629), .A2(new_n630), .A3(G57gat), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  NOR2_X1   g432(.A1(new_n627), .A2(new_n630), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n623), .B(new_n624), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  AND2_X1   g435(.A1(new_n633), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n601), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n637), .A2(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g439(.A1(G231gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G127gat), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n639), .A2(new_n643), .ZN(new_n644));
  INV_X1    g443(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n639), .A2(new_n643), .ZN(new_n646));
  XNOR2_X1  g445(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n647), .B(new_n330), .ZN(new_n648));
  XOR2_X1   g447(.A(G183gat), .B(G211gat), .Z(new_n649));
  XNOR2_X1  g448(.A(new_n648), .B(new_n649), .ZN(new_n650));
  INV_X1    g449(.A(new_n650), .ZN(new_n651));
  OR3_X1    g450(.A1(new_n645), .A2(new_n646), .A3(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n651), .B1(new_n645), .B2(new_n646), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(G134gat), .B(G162gat), .Z(new_n655));
  INV_X1    g454(.A(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT96), .ZN(new_n657));
  XNOR2_X1  g456(.A(G99gat), .B(G106gat), .ZN(new_n658));
  INV_X1    g457(.A(KEYINPUT97), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n658), .B(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(G85gat), .A2(G92gat), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(KEYINPUT7), .ZN(new_n662));
  NAND2_X1  g461(.A1(G99gat), .A2(G106gat), .ZN(new_n663));
  INV_X1    g462(.A(G85gat), .ZN(new_n664));
  INV_X1    g463(.A(G92gat), .ZN(new_n665));
  AOI22_X1  g464(.A1(KEYINPUT8), .A2(new_n663), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n660), .A2(new_n662), .A3(new_n666), .ZN(new_n667));
  XNOR2_X1  g466(.A(new_n658), .B(KEYINPUT97), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n662), .A2(new_n666), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n589), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n671), .ZN(new_n673));
  AND2_X1   g472(.A1(G232gat), .A2(G233gat), .ZN(new_n674));
  AOI22_X1  g473(.A1(new_n578), .A2(new_n673), .B1(KEYINPUT41), .B2(new_n674), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n672), .A2(new_n230), .A3(new_n675), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n674), .A2(KEYINPUT41), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n602), .B2(new_n671), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n673), .B1(new_n586), .B2(new_n588), .ZN(new_n679));
  OAI21_X1  g478(.A(G190gat), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n676), .A2(new_n680), .ZN(new_n681));
  INV_X1    g480(.A(G218gat), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n657), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n674), .A2(KEYINPUT41), .ZN(new_n684));
  INV_X1    g483(.A(new_n684), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n676), .A2(new_n680), .A3(G218gat), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n683), .A2(new_n685), .A3(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  AOI21_X1  g487(.A(new_n685), .B1(new_n683), .B2(new_n686), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n656), .B1(new_n688), .B2(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n683), .A2(new_n686), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n684), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n692), .A2(new_n655), .A3(new_n687), .ZN(new_n693));
  AOI21_X1  g492(.A(new_n637), .B1(new_n667), .B2(new_n670), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT99), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT98), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n696), .B1(new_n662), .B2(new_n666), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n637), .B1(new_n668), .B2(new_n697), .ZN(new_n698));
  AND3_X1   g497(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n695), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  OR2_X1    g499(.A1(new_n668), .A2(new_n697), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n668), .A2(KEYINPUT98), .A3(new_n669), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n701), .A2(new_n702), .A3(KEYINPUT99), .A4(new_n637), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n694), .B1(new_n700), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(G230gat), .A2(G233gat), .ZN(new_n705));
  OR3_X1    g504(.A1(new_n704), .A2(KEYINPUT100), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(KEYINPUT100), .B1(new_n704), .B2(new_n705), .ZN(new_n707));
  XNOR2_X1  g506(.A(G120gat), .B(G148gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(G176gat), .B(G204gat), .ZN(new_n709));
  XOR2_X1   g508(.A(new_n708), .B(new_n709), .Z(new_n710));
  NAND3_X1  g509(.A1(new_n706), .A2(new_n707), .A3(new_n710), .ZN(new_n711));
  AOI211_X1 g510(.A(KEYINPUT10), .B(new_n694), .C1(new_n700), .C2(new_n703), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n673), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n713));
  INV_X1    g512(.A(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n705), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n711), .A2(new_n716), .ZN(new_n717));
  INV_X1    g516(.A(new_n717), .ZN(new_n718));
  INV_X1    g517(.A(new_n710), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n705), .B(KEYINPUT101), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n700), .A2(new_n703), .ZN(new_n721));
  INV_X1    g520(.A(KEYINPUT10), .ZN(new_n722));
  INV_X1    g521(.A(new_n694), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n721), .A2(new_n722), .A3(new_n723), .ZN(new_n724));
  AOI21_X1  g523(.A(new_n720), .B1(new_n724), .B2(new_n713), .ZN(new_n725));
  NOR2_X1   g524(.A1(new_n704), .A2(new_n705), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n719), .B1(new_n725), .B2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n718), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  AND4_X1   g528(.A1(new_n654), .A2(new_n690), .A3(new_n693), .A4(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NOR3_X1   g530(.A1(new_n538), .A2(new_n622), .A3(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(new_n457), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  XOR2_X1   g533(.A(KEYINPUT102), .B(G1gat), .Z(new_n735));
  XNOR2_X1  g534(.A(new_n734), .B(new_n735), .ZN(G1324gat));
  NAND2_X1  g535(.A1(new_n732), .A2(new_n520), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT16), .B(G8gat), .ZN(new_n738));
  OAI21_X1  g537(.A(KEYINPUT103), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n739), .A2(KEYINPUT42), .B1(G8gat), .B2(new_n737), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT42), .B2(new_n739), .ZN(G1325gat));
  NAND2_X1  g540(.A1(new_n732), .A2(new_n323), .ZN(new_n742));
  INV_X1    g541(.A(new_n319), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(G15gat), .ZN(new_n744));
  AOI22_X1  g543(.A1(new_n742), .A2(G15gat), .B1(new_n732), .B2(new_n744), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(KEYINPUT104), .ZN(G1326gat));
  NAND2_X1  g545(.A1(new_n457), .A2(new_n483), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n747), .A2(new_n534), .ZN(new_n748));
  INV_X1    g547(.A(new_n322), .ZN(new_n749));
  AOI21_X1  g548(.A(KEYINPUT36), .B1(new_n307), .B2(new_n318), .ZN(new_n750));
  NOR2_X1   g549(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n524), .A2(new_n748), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n526), .A2(new_n537), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(new_n615), .B1(new_n606), .B2(new_n609), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n619), .A2(new_n620), .A3(new_n617), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n754), .A2(new_n534), .A3(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n758), .A2(new_n731), .ZN(new_n759));
  XOR2_X1   g558(.A(KEYINPUT43), .B(G22gat), .Z(new_n760));
  XNOR2_X1  g559(.A(new_n759), .B(new_n760), .ZN(G1327gat));
  NAND2_X1  g560(.A1(new_n690), .A2(new_n693), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n754), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n654), .A2(new_n728), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(new_n757), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n766), .A2(new_n562), .A3(new_n733), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT45), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT44), .ZN(new_n769));
  NOR3_X1   g568(.A1(new_n688), .A2(new_n689), .A3(new_n656), .ZN(new_n770));
  AOI21_X1  g569(.A(new_n655), .B1(new_n692), .B2(new_n687), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n769), .B1(new_n538), .B2(new_n772), .ZN(new_n773));
  NAND3_X1  g572(.A1(new_n754), .A2(KEYINPUT44), .A3(new_n762), .ZN(new_n774));
  AND2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n765), .B(KEYINPUT105), .ZN(new_n776));
  AND2_X1   g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  AND2_X1   g576(.A1(new_n777), .A2(new_n733), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n768), .B1(new_n562), .B2(new_n778), .ZN(G1328gat));
  NAND3_X1  g578(.A1(new_n766), .A2(new_n563), .A3(new_n520), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT46), .Z(new_n781));
  NAND3_X1  g580(.A1(new_n775), .A2(new_n520), .A3(new_n776), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n782), .A2(KEYINPUT106), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(G36gat), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n782), .A2(KEYINPUT106), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n781), .B1(new_n784), .B2(new_n785), .ZN(G1329gat));
  NAND3_X1  g585(.A1(new_n775), .A2(new_n323), .A3(new_n776), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n743), .A2(G43gat), .ZN(new_n788));
  AOI22_X1  g587(.A1(new_n787), .A2(G43gat), .B1(new_n766), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g588(.A(new_n789), .B(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n534), .A4(new_n776), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(G50gat), .ZN(new_n792));
  INV_X1    g591(.A(KEYINPUT108), .ZN(new_n793));
  INV_X1    g592(.A(G50gat), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n762), .A2(new_n764), .A3(new_n794), .ZN(new_n795));
  OR2_X1    g594(.A1(new_n758), .A2(new_n795), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n792), .A2(new_n793), .A3(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g597(.A(new_n793), .B1(new_n792), .B2(new_n796), .ZN(new_n799));
  AOI21_X1  g598(.A(KEYINPUT107), .B1(new_n791), .B2(G50gat), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n798), .A2(new_n799), .B1(KEYINPUT48), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(new_n799), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n800), .A2(KEYINPUT48), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n802), .A2(new_n803), .A3(new_n797), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n801), .A2(new_n804), .ZN(G1331gat));
  NAND4_X1  g604(.A1(new_n772), .A2(new_n622), .A3(new_n654), .A4(new_n728), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT109), .ZN(new_n807));
  XNOR2_X1  g606(.A(new_n806), .B(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n754), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n809), .A2(new_n457), .ZN(new_n810));
  XNOR2_X1  g609(.A(KEYINPUT110), .B(G57gat), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n810), .B(new_n811), .ZN(G1332gat));
  INV_X1    g611(.A(KEYINPUT111), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n809), .A2(new_n813), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n808), .A2(KEYINPUT111), .A3(new_n754), .ZN(new_n815));
  AND2_X1   g614(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n816), .A2(new_n520), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n818));
  XNOR2_X1  g617(.A(KEYINPUT49), .B(G64gat), .ZN(new_n819));
  NAND3_X1  g618(.A1(new_n816), .A2(new_n520), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g619(.A1(new_n818), .A2(new_n820), .ZN(G1333gat));
  NAND4_X1  g620(.A1(new_n814), .A2(G71gat), .A3(new_n323), .A4(new_n815), .ZN(new_n822));
  INV_X1    g621(.A(G71gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n823), .B1(new_n809), .B2(new_n743), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n822), .A2(new_n824), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g625(.A1(new_n816), .A2(new_n534), .ZN(new_n827));
  XNOR2_X1  g626(.A(KEYINPUT112), .B(G78gat), .ZN(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n827), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g629(.A1(new_n816), .A2(new_n534), .A3(new_n828), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(G1335gat));
  NOR2_X1   g631(.A1(new_n757), .A2(new_n654), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n729), .ZN(new_n835));
  AND2_X1   g634(.A1(new_n775), .A2(new_n835), .ZN(new_n836));
  AND2_X1   g635(.A1(new_n836), .A2(new_n733), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n772), .B1(new_n752), .B2(new_n753), .ZN(new_n838));
  XNOR2_X1  g637(.A(KEYINPUT113), .B(KEYINPUT51), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n833), .A3(new_n840), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n763), .A2(new_n834), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n843), .A2(KEYINPUT113), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n841), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n733), .A2(new_n664), .A3(new_n728), .ZN(new_n847));
  OAI22_X1  g646(.A1(new_n837), .A2(new_n664), .B1(new_n846), .B2(new_n847), .ZN(G1336gat));
  INV_X1    g647(.A(KEYINPUT116), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n729), .A2(new_n483), .A3(G92gat), .ZN(new_n850));
  NOR4_X1   g649(.A1(new_n538), .A2(new_n772), .A3(new_n834), .A4(new_n839), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n844), .B1(new_n838), .B2(new_n833), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n850), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT52), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n773), .A2(new_n774), .A3(new_n520), .A4(new_n835), .ZN(new_n856));
  INV_X1    g655(.A(KEYINPUT115), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n665), .B1(new_n856), .B2(new_n857), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n855), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n856), .A2(G92gat), .ZN(new_n861));
  XOR2_X1   g660(.A(new_n850), .B(KEYINPUT114), .Z(new_n862));
  OAI21_X1  g661(.A(new_n862), .B1(new_n851), .B2(new_n852), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n854), .B1(new_n861), .B2(new_n863), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n849), .B1(new_n860), .B2(new_n864), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(new_n845), .B2(new_n850), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n856), .A2(new_n857), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(G92gat), .ZN(new_n868));
  NOR2_X1   g667(.A1(new_n856), .A2(new_n857), .ZN(new_n869));
  OAI21_X1  g668(.A(new_n866), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(new_n864), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n870), .A2(KEYINPUT116), .A3(new_n871), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n865), .A2(new_n872), .ZN(G1337gat));
  INV_X1    g672(.A(G99gat), .ZN(new_n874));
  NAND4_X1  g673(.A1(new_n845), .A2(new_n874), .A3(new_n319), .A4(new_n728), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n836), .A2(new_n323), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n876), .B2(new_n874), .ZN(G1338gat));
  NAND3_X1  g676(.A1(new_n775), .A2(new_n534), .A3(new_n835), .ZN(new_n878));
  XNOR2_X1  g677(.A(KEYINPUT117), .B(G106gat), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n729), .A2(new_n413), .A3(G106gat), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT118), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n845), .A2(new_n881), .B1(new_n882), .B2(KEYINPUT53), .ZN(new_n883));
  OR2_X1    g682(.A1(new_n882), .A2(KEYINPUT53), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n880), .B2(new_n883), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(G1339gat));
  INV_X1    g686(.A(KEYINPUT54), .ZN(new_n888));
  AOI21_X1  g687(.A(new_n710), .B1(new_n725), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g688(.A1(new_n724), .A2(new_n720), .A3(new_n713), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n715), .A2(KEYINPUT54), .A3(new_n890), .ZN(new_n891));
  AND3_X1   g690(.A1(new_n889), .A2(new_n891), .A3(KEYINPUT55), .ZN(new_n892));
  AOI21_X1  g691(.A(KEYINPUT55), .B1(new_n889), .B2(new_n891), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n892), .A2(new_n893), .A3(new_n717), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n894), .B1(new_n616), .B2(new_n621), .ZN(new_n895));
  AND3_X1   g694(.A1(new_n603), .A2(new_n582), .A3(new_n600), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n592), .B1(new_n582), .B2(new_n591), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n614), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n756), .A2(new_n728), .A3(new_n898), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n772), .A2(new_n895), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n756), .A2(new_n894), .A3(new_n898), .ZN(new_n901));
  AOI21_X1  g700(.A(new_n654), .B1(new_n762), .B2(new_n901), .ZN(new_n902));
  AOI22_X1  g701(.A1(new_n900), .A2(new_n902), .B1(new_n730), .B2(new_n622), .ZN(new_n903));
  INV_X1    g702(.A(new_n535), .ZN(new_n904));
  NOR4_X1   g703(.A1(new_n903), .A2(new_n457), .A3(new_n520), .A4(new_n904), .ZN(new_n905));
  AOI21_X1  g704(.A(G113gat), .B1(new_n905), .B2(new_n757), .ZN(new_n906));
  OAI21_X1  g705(.A(new_n901), .B1(new_n770), .B2(new_n771), .ZN(new_n907));
  INV_X1    g706(.A(new_n654), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n899), .A2(new_n693), .A3(new_n690), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n892), .A2(new_n893), .A3(new_n717), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n910), .B1(new_n755), .B2(new_n756), .ZN(new_n911));
  OAI211_X1 g710(.A(new_n907), .B(new_n908), .C1(new_n909), .C2(new_n911), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n730), .A2(new_n622), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n457), .A2(new_n520), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n914), .A2(new_n535), .A3(new_n915), .ZN(new_n916));
  XOR2_X1   g715(.A(new_n916), .B(KEYINPUT119), .Z(new_n917));
  NOR2_X1   g716(.A1(new_n622), .A2(new_n205), .ZN(new_n918));
  AOI21_X1  g717(.A(new_n906), .B1(new_n917), .B2(new_n918), .ZN(G1340gat));
  AOI21_X1  g718(.A(G120gat), .B1(new_n905), .B2(new_n728), .ZN(new_n920));
  NOR2_X1   g719(.A1(new_n729), .A2(new_n203), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n920), .B1(new_n917), .B2(new_n921), .ZN(G1341gat));
  AND3_X1   g721(.A1(new_n905), .A2(KEYINPUT120), .A3(new_n654), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT120), .B1(new_n905), .B2(new_n654), .ZN(new_n924));
  NOR3_X1   g723(.A1(new_n923), .A2(G127gat), .A3(new_n924), .ZN(new_n925));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n216), .ZN(new_n926));
  AOI21_X1  g725(.A(new_n925), .B1(new_n917), .B2(new_n926), .ZN(G1342gat));
  XOR2_X1   g726(.A(KEYINPUT69), .B(G134gat), .Z(new_n928));
  NAND3_X1  g727(.A1(new_n905), .A2(new_n762), .A3(new_n928), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT56), .Z(new_n930));
  AND2_X1   g729(.A1(new_n917), .A2(new_n762), .ZN(new_n931));
  OAI21_X1  g730(.A(new_n930), .B1(new_n931), .B2(new_n215), .ZN(G1343gat));
  NAND2_X1  g731(.A1(new_n751), .A2(new_n915), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT57), .ZN(new_n934));
  AOI211_X1 g733(.A(new_n934), .B(new_n413), .C1(new_n912), .C2(new_n913), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n933), .B1(new_n935), .B2(KEYINPUT121), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n934), .B1(new_n903), .B2(new_n413), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n914), .A2(KEYINPUT57), .A3(new_n534), .ZN(new_n938));
  INV_X1    g737(.A(KEYINPUT121), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n937), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n936), .A2(new_n940), .A3(new_n757), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n941), .A2(G141gat), .ZN(new_n942));
  NOR2_X1   g741(.A1(new_n323), .A2(new_n413), .ZN(new_n943));
  AND4_X1   g742(.A1(new_n733), .A2(new_n914), .A3(new_n483), .A4(new_n943), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n341), .A3(new_n757), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n946), .A2(KEYINPUT58), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT58), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n942), .A2(new_n948), .A3(new_n945), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n947), .A2(new_n949), .ZN(G1344gat));
  NOR2_X1   g749(.A1(new_n339), .A2(KEYINPUT59), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n940), .ZN(new_n952));
  OAI21_X1  g751(.A(new_n951), .B1(new_n952), .B2(new_n729), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT59), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n937), .A2(new_n938), .ZN(new_n955));
  AND2_X1   g754(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n956));
  NOR2_X1   g755(.A1(new_n933), .A2(KEYINPUT123), .ZN(new_n957));
  NOR3_X1   g756(.A1(new_n956), .A2(new_n957), .A3(new_n729), .ZN(new_n958));
  AOI21_X1  g757(.A(new_n335), .B1(new_n955), .B2(new_n958), .ZN(new_n959));
  OAI21_X1  g758(.A(new_n953), .B1(new_n954), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g759(.A1(new_n944), .A2(new_n339), .A3(new_n728), .ZN(new_n961));
  XNOR2_X1  g760(.A(new_n961), .B(KEYINPUT122), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1345gat));
  OAI21_X1  g762(.A(G155gat), .B1(new_n952), .B2(new_n908), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n944), .A2(new_n330), .A3(new_n654), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n964), .A2(new_n965), .ZN(G1346gat));
  NOR3_X1   g765(.A1(new_n952), .A2(new_n331), .A3(new_n772), .ZN(new_n967));
  AOI21_X1  g766(.A(G162gat), .B1(new_n944), .B2(new_n762), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n967), .A2(new_n968), .ZN(G1347gat));
  NOR2_X1   g768(.A1(new_n903), .A2(new_n733), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n904), .A2(new_n483), .ZN(new_n971));
  NAND2_X1  g770(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G169gat), .B1(new_n973), .B2(new_n757), .ZN(new_n974));
  NOR2_X1   g773(.A1(new_n733), .A2(new_n483), .ZN(new_n975));
  INV_X1    g774(.A(new_n975), .ZN(new_n976));
  NOR3_X1   g775(.A1(new_n903), .A2(new_n904), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g776(.A1(new_n622), .A2(new_n236), .ZN(new_n978));
  AOI21_X1  g777(.A(new_n974), .B1(new_n977), .B2(new_n978), .ZN(G1348gat));
  NAND3_X1  g778(.A1(new_n973), .A2(new_n237), .A3(new_n728), .ZN(new_n980));
  AND2_X1   g779(.A1(new_n977), .A2(new_n728), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n981), .B2(new_n237), .ZN(G1349gat));
  AOI21_X1  g781(.A(new_n229), .B1(new_n977), .B2(new_n654), .ZN(new_n983));
  INV_X1    g782(.A(new_n266), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n908), .A2(new_n984), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n983), .B1(new_n973), .B2(new_n985), .ZN(new_n986));
  XOR2_X1   g785(.A(new_n986), .B(KEYINPUT60), .Z(G1350gat));
  NAND3_X1  g786(.A1(new_n973), .A2(new_n230), .A3(new_n762), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n977), .A2(new_n762), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n989), .A2(G190gat), .ZN(new_n990));
  AND2_X1   g789(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n990), .A2(KEYINPUT61), .ZN(new_n992));
  OAI21_X1  g791(.A(new_n988), .B1(new_n991), .B2(new_n992), .ZN(G1351gat));
  INV_X1    g792(.A(G197gat), .ZN(new_n994));
  NOR2_X1   g793(.A1(new_n976), .A2(new_n323), .ZN(new_n995));
  INV_X1    g794(.A(new_n995), .ZN(new_n996));
  AOI21_X1  g795(.A(new_n996), .B1(new_n937), .B2(new_n938), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n994), .B1(new_n997), .B2(new_n757), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n943), .A2(new_n520), .ZN(new_n999));
  XNOR2_X1  g798(.A(new_n999), .B(KEYINPUT124), .ZN(new_n1000));
  NAND2_X1  g799(.A1(new_n970), .A2(new_n1000), .ZN(new_n1001));
  NOR3_X1   g800(.A1(new_n1001), .A2(G197gat), .A3(new_n622), .ZN(new_n1002));
  OR3_X1    g801(.A1(new_n998), .A2(KEYINPUT125), .A3(new_n1002), .ZN(new_n1003));
  OAI21_X1  g802(.A(KEYINPUT125), .B1(new_n998), .B2(new_n1002), .ZN(new_n1004));
  NAND2_X1  g803(.A1(new_n1003), .A2(new_n1004), .ZN(G1352gat));
  INV_X1    g804(.A(KEYINPUT127), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n970), .A2(new_n1000), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n729), .A2(G204gat), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1007), .A2(KEYINPUT126), .A3(new_n1008), .ZN(new_n1009));
  INV_X1    g808(.A(KEYINPUT126), .ZN(new_n1010));
  INV_X1    g809(.A(new_n1008), .ZN(new_n1011));
  OAI21_X1  g810(.A(new_n1010), .B1(new_n1001), .B2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g811(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  OAI21_X1  g812(.A(new_n1006), .B1(new_n1013), .B2(KEYINPUT62), .ZN(new_n1014));
  NAND2_X1  g813(.A1(new_n1013), .A2(KEYINPUT62), .ZN(new_n1015));
  INV_X1    g814(.A(KEYINPUT62), .ZN(new_n1016));
  NAND4_X1  g815(.A1(new_n1009), .A2(new_n1012), .A3(KEYINPUT127), .A4(new_n1016), .ZN(new_n1017));
  INV_X1    g816(.A(new_n997), .ZN(new_n1018));
  OAI21_X1  g817(.A(G204gat), .B1(new_n1018), .B2(new_n729), .ZN(new_n1019));
  NAND4_X1  g818(.A1(new_n1014), .A2(new_n1015), .A3(new_n1017), .A4(new_n1019), .ZN(G1353gat));
  OR3_X1    g819(.A1(new_n1001), .A2(G211gat), .A3(new_n908), .ZN(new_n1021));
  NAND2_X1  g820(.A1(new_n997), .A2(new_n654), .ZN(new_n1022));
  AND3_X1   g821(.A1(new_n1022), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1023));
  AOI21_X1  g822(.A(KEYINPUT63), .B1(new_n1022), .B2(G211gat), .ZN(new_n1024));
  OAI21_X1  g823(.A(new_n1021), .B1(new_n1023), .B2(new_n1024), .ZN(G1354gat));
  OAI21_X1  g824(.A(G218gat), .B1(new_n1018), .B2(new_n772), .ZN(new_n1026));
  NAND3_X1  g825(.A1(new_n1007), .A2(new_n682), .A3(new_n762), .ZN(new_n1027));
  NAND2_X1  g826(.A1(new_n1026), .A2(new_n1027), .ZN(G1355gat));
endmodule


