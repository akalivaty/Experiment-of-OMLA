

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803;

  AND2_X1 U382 ( .A1(n507), .A2(n506), .ZN(n396) );
  XNOR2_X1 U383 ( .A(n618), .B(n366), .ZN(n372) );
  XNOR2_X1 U384 ( .A(n468), .B(n467), .ZN(n687) );
  OR2_X1 U385 ( .A1(n587), .A2(n724), .ZN(n600) );
  INV_X1 U386 ( .A(n436), .ZN(n438) );
  XOR2_X1 U387 ( .A(KEYINPUT67), .B(G101), .Z(n553) );
  XNOR2_X1 U388 ( .A(n516), .B(n515), .ZN(n555) );
  XNOR2_X1 U389 ( .A(n367), .B(n419), .ZN(n445) );
  XNOR2_X1 U390 ( .A(n651), .B(KEYINPUT109), .ZN(n652) );
  NOR2_X1 U391 ( .A1(n653), .A2(n652), .ZN(n704) );
  AND2_X1 U392 ( .A1(n438), .A2(n437), .ZN(n360) );
  XOR2_X1 U393 ( .A(n561), .B(KEYINPUT62), .Z(n361) );
  AND2_X1 U394 ( .A1(n390), .A2(n387), .ZN(n362) );
  INV_X1 U395 ( .A(n649), .ZN(n683) );
  NAND2_X4 U396 ( .A1(n461), .A2(n474), .ZN(n507) );
  AND2_X2 U397 ( .A1(n472), .A2(n470), .ZN(n461) );
  XNOR2_X1 U398 ( .A(n392), .B(n552), .ZN(n367) );
  XNOR2_X1 U399 ( .A(n393), .B(n553), .ZN(n392) );
  XNOR2_X1 U400 ( .A(n551), .B(n462), .ZN(n393) );
  NOR2_X2 U401 ( .A1(n743), .A2(n729), .ZN(n595) );
  XNOR2_X2 U402 ( .A(n594), .B(KEYINPUT100), .ZN(n743) );
  INV_X1 U403 ( .A(n721), .ZN(n506) );
  NOR2_X2 U404 ( .A1(n721), .A2(n720), .ZN(n722) );
  NAND2_X2 U405 ( .A1(n452), .A2(n595), .ZN(n596) );
  NAND2_X2 U406 ( .A1(n687), .A2(n686), .ZN(n791) );
  OR2_X2 U407 ( .A1(n561), .A2(G902), .ZN(n420) );
  NOR2_X1 U408 ( .A1(n791), .A2(n371), .ZN(n370) );
  NAND2_X1 U409 ( .A1(n603), .A2(n602), .ZN(n594) );
  OR2_X1 U410 ( .A1(n763), .A2(n423), .ZN(n422) );
  XNOR2_X1 U411 ( .A(G113), .B(G143), .ZN(n536) );
  INV_X1 U412 ( .A(KEYINPUT69), .ZN(n418) );
  INV_X1 U413 ( .A(KEYINPUT22), .ZN(n364) );
  INV_X1 U414 ( .A(KEYINPUT2), .ZN(n371) );
  AND2_X1 U415 ( .A1(n383), .A2(n389), .ZN(n382) );
  NAND2_X1 U416 ( .A1(n475), .A2(KEYINPUT81), .ZN(n474) );
  NAND2_X1 U417 ( .A1(n372), .A2(n370), .ZN(n691) );
  OR2_X1 U418 ( .A1(n372), .A2(KEYINPUT2), .ZN(n718) );
  NOR2_X1 U419 ( .A1(n471), .A2(n412), .ZN(n470) );
  NOR2_X1 U420 ( .A1(n377), .A2(n599), .ZN(n380) );
  OR2_X1 U421 ( .A1(n607), .A2(n608), .ZN(n606) );
  OR2_X1 U422 ( .A1(n592), .A2(n591), .ZN(n599) );
  XNOR2_X1 U423 ( .A(n612), .B(KEYINPUT32), .ZN(n801) );
  XNOR2_X1 U424 ( .A(n369), .B(KEYINPUT31), .ZN(n710) );
  XNOR2_X1 U425 ( .A(n373), .B(KEYINPUT42), .ZN(n803) );
  AND2_X1 U426 ( .A1(n482), .A2(n405), .ZN(n481) );
  INV_X1 U427 ( .A(n670), .ZN(n705) );
  AND2_X1 U428 ( .A1(n723), .A2(n655), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n368), .B(n636), .ZN(n723) );
  NAND2_X1 U430 ( .A1(n435), .A2(n439), .ZN(n436) );
  NOR2_X1 U431 ( .A1(n633), .A2(n632), .ZN(n655) );
  NOR2_X1 U432 ( .A1(n657), .A2(n626), .ZN(n627) );
  XNOR2_X1 U433 ( .A(n762), .B(n761), .ZN(n409) );
  NAND2_X2 U434 ( .A1(n425), .A2(n422), .ZN(n631) );
  XNOR2_X1 U435 ( .A(n593), .B(G475), .ZN(n603) );
  INV_X1 U436 ( .A(n660), .ZN(n363) );
  AND2_X1 U437 ( .A1(n427), .A2(n426), .ZN(n425) );
  XOR2_X1 U438 ( .A(n765), .B(n764), .Z(n411) );
  OR2_X1 U439 ( .A1(n767), .A2(G902), .ZN(n414) );
  XOR2_X1 U440 ( .A(n767), .B(n766), .Z(n410) );
  XNOR2_X1 U441 ( .A(n586), .B(n585), .ZN(n763) );
  XNOR2_X1 U442 ( .A(n586), .B(n522), .ZN(n561) );
  XNOR2_X1 U443 ( .A(n541), .B(n540), .ZN(n767) );
  XNOR2_X1 U444 ( .A(n458), .B(n565), .ZN(n541) );
  XNOR2_X1 U445 ( .A(n416), .B(n415), .ZN(n458) );
  XNOR2_X1 U446 ( .A(n478), .B(n582), .ZN(n419) );
  XNOR2_X1 U447 ( .A(n555), .B(KEYINPUT16), .ZN(n477) );
  XNOR2_X1 U448 ( .A(n417), .B(n536), .ZN(n416) );
  XNOR2_X1 U449 ( .A(n499), .B(n498), .ZN(n497) );
  AND2_X1 U450 ( .A1(KEYINPUT122), .A2(n464), .ZN(n384) );
  XNOR2_X1 U451 ( .A(n421), .B(G110), .ZN(n582) );
  XNOR2_X1 U452 ( .A(n418), .B(G131), .ZN(n535) );
  XNOR2_X1 U453 ( .A(n550), .B(KEYINPUT10), .ZN(n565) );
  INV_X1 U454 ( .A(n617), .ZN(n366) );
  INV_X1 U455 ( .A(n374), .ZN(n365) );
  XNOR2_X1 U456 ( .A(G125), .B(G146), .ZN(n550) );
  XNOR2_X1 U457 ( .A(KEYINPUT3), .B(G119), .ZN(n515) );
  NOR2_X2 U458 ( .A1(G953), .A2(G237), .ZN(n534) );
  INV_X1 U459 ( .A(G475), .ZN(n399) );
  XOR2_X1 U460 ( .A(G113), .B(G116), .Z(n516) );
  BUF_X1 U461 ( .A(G953), .Z(n374) );
  XNOR2_X1 U462 ( .A(KEYINPUT96), .B(KEYINPUT95), .ZN(n498) );
  XNOR2_X1 U463 ( .A(G119), .B(G110), .ZN(n569) );
  XNOR2_X1 U464 ( .A(G137), .B(KEYINPUT5), .ZN(n517) );
  XOR2_X1 U465 ( .A(G902), .B(KEYINPUT15), .Z(n562) );
  XOR2_X1 U466 ( .A(KEYINPUT45), .B(KEYINPUT64), .Z(n617) );
  XNOR2_X1 U467 ( .A(G128), .B(KEYINPUT24), .ZN(n566) );
  XNOR2_X1 U468 ( .A(KEYINPUT30), .B(KEYINPUT108), .ZN(n500) );
  AND2_X1 U469 ( .A1(n510), .A2(n363), .ZN(n611) );
  XNOR2_X1 U470 ( .A(n596), .B(n364), .ZN(n510) );
  NAND2_X1 U471 ( .A1(n372), .A2(n365), .ZN(n779) );
  XNOR2_X1 U472 ( .A(n619), .B(KEYINPUT82), .ZN(n476) );
  NAND2_X1 U473 ( .A1(n469), .A2(n648), .ZN(n605) );
  NAND2_X1 U474 ( .A1(n360), .A2(n430), .ZN(n434) );
  INV_X2 U475 ( .A(G143), .ZN(n503) );
  XNOR2_X2 U476 ( .A(n504), .B(n450), .ZN(n452) );
  XNOR2_X1 U477 ( .A(n609), .B(KEYINPUT102), .ZN(n641) );
  NAND2_X1 U478 ( .A1(n738), .A2(n635), .ZN(n368) );
  XNOR2_X2 U479 ( .A(n683), .B(KEYINPUT38), .ZN(n741) );
  NAND2_X1 U480 ( .A1(n430), .A2(n734), .ZN(n369) );
  XNOR2_X2 U481 ( .A(n605), .B(KEYINPUT35), .ZN(n607) );
  NAND2_X1 U482 ( .A1(n375), .A2(KEYINPUT44), .ZN(n381) );
  NAND2_X1 U483 ( .A1(n615), .A2(n613), .ZN(n375) );
  NAND2_X1 U484 ( .A1(n376), .A2(n616), .ZN(n378) );
  XNOR2_X1 U485 ( .A(n615), .B(KEYINPUT86), .ZN(n376) );
  NAND2_X1 U486 ( .A1(n606), .A2(n465), .ZN(n377) );
  NAND2_X2 U487 ( .A1(n379), .A2(n378), .ZN(n618) );
  AND2_X2 U488 ( .A1(n381), .A2(n380), .ZN(n379) );
  NAND2_X1 U489 ( .A1(n382), .A2(n386), .ZN(G75) );
  NAND2_X1 U490 ( .A1(n388), .A2(n464), .ZN(n383) );
  NAND2_X1 U491 ( .A1(n385), .A2(KEYINPUT122), .ZN(n391) );
  NAND2_X1 U492 ( .A1(n385), .A2(n384), .ZN(n389) );
  INV_X1 U493 ( .A(n449), .ZN(n385) );
  NAND2_X1 U494 ( .A1(n391), .A2(n362), .ZN(n386) );
  AND2_X1 U495 ( .A1(n447), .A2(KEYINPUT53), .ZN(n387) );
  NAND2_X1 U496 ( .A1(n390), .A2(n447), .ZN(n388) );
  NAND2_X1 U497 ( .A1(n449), .A2(n406), .ZN(n390) );
  BUF_X1 U498 ( .A(n728), .Z(n394) );
  BUF_X1 U499 ( .A(n772), .Z(n395) );
  XNOR2_X1 U500 ( .A(n578), .B(n577), .ZN(n728) );
  AND2_X1 U501 ( .A1(n506), .A2(G472), .ZN(n397) );
  NAND2_X1 U502 ( .A1(n507), .A2(n398), .ZN(n486) );
  NOR2_X1 U503 ( .A1(n721), .A2(n399), .ZN(n398) );
  NAND2_X1 U504 ( .A1(n400), .A2(n507), .ZN(n494) );
  AND2_X1 U505 ( .A1(n506), .A2(G469), .ZN(n400) );
  INV_X4 U506 ( .A(G953), .ZN(n792) );
  NAND2_X1 U507 ( .A1(n363), .A2(n408), .ZN(n439) );
  NAND2_X1 U508 ( .A1(n429), .A2(n428), .ZN(n437) );
  INV_X1 U509 ( .A(n600), .ZN(n429) );
  NOR2_X1 U510 ( .A1(n363), .A2(n408), .ZN(n428) );
  XNOR2_X1 U511 ( .A(n535), .B(n520), .ZN(n502) );
  INV_X1 U512 ( .A(G134), .ZN(n520) );
  NAND2_X1 U513 ( .A1(n557), .A2(G214), .ZN(n740) );
  XOR2_X1 U514 ( .A(G137), .B(G140), .Z(n580) );
  XNOR2_X1 U515 ( .A(n581), .B(n460), .ZN(n459) );
  INV_X1 U516 ( .A(KEYINPUT77), .ZN(n460) );
  XNOR2_X1 U517 ( .A(G107), .B(KEYINPUT70), .ZN(n421) );
  NAND2_X1 U518 ( .A1(G469), .A2(n424), .ZN(n423) );
  INV_X1 U519 ( .A(KEYINPUT6), .ZN(n495) );
  XNOR2_X1 U520 ( .A(n497), .B(n496), .ZN(n518) );
  XNOR2_X1 U521 ( .A(n517), .B(KEYINPUT73), .ZN(n496) );
  XOR2_X1 U522 ( .A(KEYINPUT68), .B(KEYINPUT8), .Z(n528) );
  XNOR2_X1 U523 ( .A(G134), .B(KEYINPUT7), .ZN(n526) );
  XNOR2_X1 U524 ( .A(n539), .B(n514), .ZN(n540) );
  XNOR2_X1 U525 ( .A(n576), .B(n513), .ZN(n577) );
  NOR2_X1 U526 ( .A1(n448), .A2(n374), .ZN(n447) );
  NOR2_X1 U527 ( .A1(n403), .A2(n759), .ZN(n448) );
  NAND2_X1 U528 ( .A1(G234), .A2(G237), .ZN(n543) );
  NOR2_X1 U529 ( .A1(G237), .A2(G902), .ZN(n549) );
  INV_X1 U530 ( .A(G902), .ZN(n424) );
  NAND2_X1 U531 ( .A1(n446), .A2(G902), .ZN(n426) );
  INV_X1 U532 ( .A(KEYINPUT48), .ZN(n467) );
  XNOR2_X1 U533 ( .A(G140), .B(KEYINPUT98), .ZN(n537) );
  XOR2_X1 U534 ( .A(KEYINPUT12), .B(KEYINPUT97), .Z(n538) );
  NOR2_X1 U535 ( .A1(n689), .A2(n487), .ZN(n471) );
  NAND2_X1 U536 ( .A1(n792), .A2(G224), .ZN(n551) );
  INV_X1 U537 ( .A(KEYINPUT4), .ZN(n519) );
  XNOR2_X1 U538 ( .A(n550), .B(KEYINPUT88), .ZN(n478) );
  INV_X1 U539 ( .A(KEYINPUT111), .ZN(n628) );
  XNOR2_X1 U540 ( .A(n569), .B(n568), .ZN(n570) );
  INV_X1 U541 ( .A(n580), .ZN(n463) );
  XNOR2_X1 U542 ( .A(n459), .B(n580), .ZN(n584) );
  INV_X1 U543 ( .A(KEYINPUT122), .ZN(n759) );
  INV_X1 U544 ( .A(KEYINPUT0), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n501), .B(n500), .ZN(n642) );
  NOR2_X1 U546 ( .A1(n681), .A2(n511), .ZN(n509) );
  XOR2_X1 U547 ( .A(G122), .B(KEYINPUT9), .Z(n530) );
  XNOR2_X1 U548 ( .A(n598), .B(KEYINPUT101), .ZN(n800) );
  INV_X1 U549 ( .A(KEYINPUT60), .ZN(n483) );
  INV_X1 U550 ( .A(KEYINPUT124), .ZN(n491) );
  INV_X1 U551 ( .A(KEYINPUT56), .ZN(n453) );
  INV_X1 U552 ( .A(KEYINPUT53), .ZN(n464) );
  AND2_X1 U553 ( .A1(n437), .A2(KEYINPUT34), .ZN(n401) );
  XOR2_X1 U554 ( .A(KEYINPUT13), .B(KEYINPUT99), .Z(n402) );
  XOR2_X1 U555 ( .A(KEYINPUT121), .B(n758), .Z(n403) );
  AND2_X1 U556 ( .A1(n506), .A2(G210), .ZN(n404) );
  INV_X1 U557 ( .A(G469), .ZN(n446) );
  AND2_X1 U558 ( .A1(n508), .A2(n626), .ZN(n405) );
  AND2_X1 U559 ( .A1(n403), .A2(n759), .ZN(n406) );
  NOR2_X1 U560 ( .A1(n724), .A2(n620), .ZN(n407) );
  XOR2_X1 U561 ( .A(KEYINPUT104), .B(KEYINPUT33), .Z(n408) );
  INV_X1 U562 ( .A(KEYINPUT34), .ZN(n440) );
  NOR2_X1 U563 ( .A1(n690), .A2(n371), .ZN(n412) );
  NOR2_X1 U564 ( .A1(G952), .A2(n792), .ZN(n774) );
  INV_X1 U565 ( .A(n774), .ZN(n455) );
  XOR2_X1 U566 ( .A(KEYINPUT63), .B(KEYINPUT89), .Z(n413) );
  INV_X1 U567 ( .A(KEYINPUT81), .ZN(n487) );
  XNOR2_X2 U568 ( .A(n414), .B(n402), .ZN(n593) );
  INV_X1 U569 ( .A(n535), .ZN(n415) );
  NAND2_X1 U570 ( .A1(n534), .A2(G214), .ZN(n417) );
  XNOR2_X2 U571 ( .A(n523), .B(n519), .ZN(n552) );
  XNOR2_X2 U572 ( .A(n503), .B(G128), .ZN(n523) );
  XNOR2_X2 U573 ( .A(n420), .B(G472), .ZN(n609) );
  NAND2_X1 U574 ( .A1(n763), .A2(n446), .ZN(n427) );
  XNOR2_X2 U575 ( .A(n631), .B(KEYINPUT1), .ZN(n724) );
  INV_X1 U576 ( .A(n601), .ZN(n430) );
  NAND2_X1 U577 ( .A1(n433), .A2(n431), .ZN(n469) );
  NAND2_X1 U578 ( .A1(n401), .A2(n432), .ZN(n431) );
  NOR2_X1 U579 ( .A1(n436), .A2(n601), .ZN(n432) );
  NAND2_X1 U580 ( .A1(n434), .A2(n440), .ZN(n433) );
  NAND2_X1 U581 ( .A1(n600), .A2(n408), .ZN(n435) );
  NAND2_X1 U582 ( .A1(n438), .A2(n437), .ZN(n755) );
  XNOR2_X1 U583 ( .A(n596), .B(KEYINPUT22), .ZN(n610) );
  BUF_X1 U584 ( .A(n760), .Z(n441) );
  XNOR2_X1 U585 ( .A(n571), .B(n570), .ZN(n573) );
  XNOR2_X1 U586 ( .A(G110), .B(G107), .ZN(n442) );
  XNOR2_X1 U587 ( .A(n618), .B(n617), .ZN(n775) );
  NAND2_X1 U588 ( .A1(n534), .A2(G210), .ZN(n499) );
  NAND2_X1 U589 ( .A1(n456), .A2(n455), .ZN(n454) );
  NOR2_X1 U590 ( .A1(n802), .A2(n803), .ZN(n647) );
  NAND2_X1 U591 ( .A1(n641), .A2(n740), .ZN(n501) );
  XNOR2_X1 U592 ( .A(n609), .B(n495), .ZN(n660) );
  BUF_X1 U593 ( .A(n654), .Z(n443) );
  XNOR2_X1 U594 ( .A(n505), .B(KEYINPUT19), .ZN(n654) );
  XNOR2_X1 U595 ( .A(n457), .B(n409), .ZN(n456) );
  BUF_X1 U596 ( .A(n699), .Z(n444) );
  NAND2_X1 U597 ( .A1(n481), .A2(n480), .ZN(n479) );
  XNOR2_X2 U598 ( .A(n445), .B(n780), .ZN(n760) );
  NAND2_X1 U599 ( .A1(n404), .A2(n507), .ZN(n457) );
  NAND2_X1 U600 ( .A1(n397), .A2(n507), .ZN(n490) );
  NAND2_X1 U601 ( .A1(n396), .A2(G478), .ZN(n768) );
  NAND2_X1 U602 ( .A1(n396), .A2(G217), .ZN(n771) );
  XNOR2_X2 U603 ( .A(n789), .B(n521), .ZN(n586) );
  INV_X1 U604 ( .A(n724), .ZN(n681) );
  XNOR2_X1 U605 ( .A(n722), .B(KEYINPUT83), .ZN(n449) );
  INV_X1 U606 ( .A(n452), .ZN(n601) );
  OR2_X1 U607 ( .A1(n601), .A2(n451), .ZN(n588) );
  INV_X1 U608 ( .A(n637), .ZN(n451) );
  XNOR2_X1 U609 ( .A(n454), .B(n453), .ZN(G51) );
  AND2_X1 U610 ( .A1(n611), .A2(n407), .ZN(n612) );
  XNOR2_X1 U611 ( .A(n479), .B(KEYINPUT65), .ZN(n466) );
  INV_X1 U612 ( .A(n800), .ZN(n465) );
  XNOR2_X2 U613 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n462) );
  AND2_X2 U614 ( .A1(n466), .A2(n394), .ZN(n699) );
  XNOR2_X1 U615 ( .A(n574), .B(n790), .ZN(n772) );
  XNOR2_X1 U616 ( .A(n565), .B(n463), .ZN(n790) );
  NOR2_X2 U617 ( .A1(n699), .A2(n801), .ZN(n615) );
  NAND2_X1 U618 ( .A1(n610), .A2(n511), .ZN(n482) );
  XNOR2_X1 U619 ( .A(n791), .B(n688), .ZN(n689) );
  NAND2_X1 U620 ( .A1(n676), .A2(n677), .ZN(n468) );
  NAND2_X1 U621 ( .A1(n476), .A2(n473), .ZN(n472) );
  AND2_X1 U622 ( .A1(n689), .A2(n487), .ZN(n473) );
  INV_X1 U623 ( .A(n476), .ZN(n475) );
  XNOR2_X2 U624 ( .A(n556), .B(n477), .ZN(n780) );
  NAND2_X1 U625 ( .A1(n510), .A2(n509), .ZN(n480) );
  XNOR2_X1 U626 ( .A(n484), .B(n483), .ZN(G60) );
  NAND2_X1 U627 ( .A1(n485), .A2(n455), .ZN(n484) );
  XNOR2_X1 U628 ( .A(n486), .B(n410), .ZN(n485) );
  XNOR2_X1 U629 ( .A(n488), .B(n413), .ZN(G57) );
  NAND2_X1 U630 ( .A1(n489), .A2(n455), .ZN(n488) );
  XNOR2_X1 U631 ( .A(n490), .B(n361), .ZN(n489) );
  XNOR2_X1 U632 ( .A(n492), .B(n491), .ZN(G54) );
  NAND2_X1 U633 ( .A1(n493), .A2(n455), .ZN(n492) );
  XNOR2_X1 U634 ( .A(n494), .B(n411), .ZN(n493) );
  XNOR2_X2 U635 ( .A(n552), .B(n502), .ZN(n789) );
  NAND2_X1 U636 ( .A1(n654), .A2(n560), .ZN(n504) );
  NAND2_X1 U637 ( .A1(n649), .A2(n740), .ZN(n505) );
  XNOR2_X2 U638 ( .A(n691), .B(KEYINPUT75), .ZN(n721) );
  NAND2_X1 U639 ( .A1(n681), .A2(n511), .ZN(n508) );
  INV_X1 U640 ( .A(KEYINPUT103), .ZN(n511) );
  NOR2_X2 U641 ( .A1(n760), .A2(n562), .ZN(n559) );
  NOR2_X2 U642 ( .A1(n643), .A2(n642), .ZN(n650) );
  AND2_X1 U643 ( .A1(n572), .A2(G221), .ZN(n512) );
  XOR2_X1 U644 ( .A(KEYINPUT25), .B(KEYINPUT94), .Z(n513) );
  XOR2_X1 U645 ( .A(n538), .B(n537), .Z(n514) );
  INV_X1 U646 ( .A(KEYINPUT74), .ZN(n688) );
  INV_X1 U647 ( .A(KEYINPUT92), .ZN(n568) );
  INV_X1 U648 ( .A(KEYINPUT76), .ZN(n639) );
  XNOR2_X1 U649 ( .A(n628), .B(KEYINPUT28), .ZN(n629) );
  XNOR2_X1 U650 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U651 ( .A1(n715), .A2(n685), .ZN(n686) );
  XNOR2_X1 U652 ( .A(n630), .B(n629), .ZN(n633) );
  XNOR2_X1 U653 ( .A(n573), .B(n512), .ZN(n574) );
  XOR2_X1 U654 ( .A(n555), .B(n518), .Z(n522) );
  XOR2_X1 U655 ( .A(n553), .B(G146), .Z(n521) );
  XNOR2_X1 U656 ( .A(n523), .B(G116), .ZN(n524) );
  XNOR2_X1 U657 ( .A(n524), .B(G107), .ZN(n525) );
  XNOR2_X1 U658 ( .A(n526), .B(n525), .ZN(n532) );
  NAND2_X1 U659 ( .A1(G234), .A2(n792), .ZN(n527) );
  XNOR2_X1 U660 ( .A(n528), .B(n527), .ZN(n572) );
  NAND2_X1 U661 ( .A1(G217), .A2(n572), .ZN(n529) );
  XNOR2_X1 U662 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U663 ( .A(n532), .B(n531), .ZN(n769) );
  NOR2_X1 U664 ( .A1(G902), .A2(n769), .ZN(n533) );
  XNOR2_X1 U665 ( .A(G478), .B(n533), .ZN(n602) );
  XOR2_X1 U666 ( .A(G122), .B(G104), .Z(n554) );
  XNOR2_X1 U667 ( .A(n554), .B(KEYINPUT11), .ZN(n539) );
  XOR2_X1 U668 ( .A(G475), .B(n593), .Z(n542) );
  NAND2_X1 U669 ( .A1(n602), .A2(n542), .ZN(n692) );
  NOR2_X1 U670 ( .A1(n542), .A2(n602), .ZN(n709) );
  INV_X1 U671 ( .A(n709), .ZN(n678) );
  NAND2_X1 U672 ( .A1(n692), .A2(n678), .ZN(n737) );
  XOR2_X1 U673 ( .A(n737), .B(KEYINPUT78), .Z(n590) );
  XNOR2_X1 U674 ( .A(KEYINPUT14), .B(n543), .ZN(n546) );
  AND2_X1 U675 ( .A1(n374), .A2(n546), .ZN(n544) );
  NAND2_X1 U676 ( .A1(G902), .A2(n544), .ZN(n621) );
  NOR2_X1 U677 ( .A1(G898), .A2(n621), .ZN(n545) );
  XNOR2_X1 U678 ( .A(KEYINPUT91), .B(n545), .ZN(n548) );
  NAND2_X1 U679 ( .A1(G952), .A2(n546), .ZN(n753) );
  NOR2_X1 U680 ( .A1(n374), .A2(n753), .ZN(n547) );
  XOR2_X1 U681 ( .A(KEYINPUT90), .B(n547), .Z(n623) );
  NAND2_X1 U682 ( .A1(n548), .A2(n623), .ZN(n560) );
  XOR2_X1 U683 ( .A(KEYINPUT72), .B(n549), .Z(n557) );
  XOR2_X1 U684 ( .A(n554), .B(KEYINPUT71), .Z(n556) );
  NAND2_X1 U685 ( .A1(n557), .A2(G210), .ZN(n558) );
  XNOR2_X2 U686 ( .A(n559), .B(n558), .ZN(n649) );
  INV_X1 U687 ( .A(n609), .ZN(n726) );
  INV_X1 U688 ( .A(n562), .ZN(n690) );
  NAND2_X1 U689 ( .A1(n690), .A2(G234), .ZN(n563) );
  XNOR2_X1 U690 ( .A(n563), .B(KEYINPUT20), .ZN(n575) );
  NAND2_X1 U691 ( .A1(n575), .A2(G221), .ZN(n564) );
  XNOR2_X1 U692 ( .A(KEYINPUT21), .B(n564), .ZN(n729) );
  XOR2_X1 U693 ( .A(KEYINPUT93), .B(KEYINPUT23), .Z(n567) );
  XNOR2_X1 U694 ( .A(n567), .B(n566), .ZN(n571) );
  NOR2_X1 U695 ( .A1(n772), .A2(G902), .ZN(n578) );
  NAND2_X1 U696 ( .A1(n575), .A2(G217), .ZN(n576) );
  NOR2_X1 U697 ( .A1(n729), .A2(n728), .ZN(n579) );
  INV_X1 U698 ( .A(n579), .ZN(n587) );
  NAND2_X1 U699 ( .A1(n792), .A2(G227), .ZN(n581) );
  XNOR2_X1 U700 ( .A(n582), .B(G104), .ZN(n583) );
  XNOR2_X1 U701 ( .A(n584), .B(n583), .ZN(n585) );
  NOR2_X1 U702 ( .A1(n726), .A2(n600), .ZN(n734) );
  NOR2_X2 U703 ( .A1(n587), .A2(n631), .ZN(n637) );
  NOR2_X1 U704 ( .A1(n609), .A2(n588), .ZN(n694) );
  NOR2_X1 U705 ( .A1(n710), .A2(n694), .ZN(n589) );
  NOR2_X1 U706 ( .A1(n590), .A2(n589), .ZN(n592) );
  INV_X1 U707 ( .A(KEYINPUT85), .ZN(n608) );
  NOR2_X1 U708 ( .A1(KEYINPUT44), .A2(n608), .ZN(n591) );
  NOR2_X1 U709 ( .A1(n681), .A2(n394), .ZN(n597) );
  NAND2_X1 U710 ( .A1(n611), .A2(n597), .ZN(n598) );
  OR2_X1 U711 ( .A1(n603), .A2(n602), .ZN(n604) );
  XNOR2_X1 U712 ( .A(KEYINPUT105), .B(n604), .ZN(n648) );
  NAND2_X1 U713 ( .A1(n608), .A2(n607), .ZN(n613) );
  INV_X1 U714 ( .A(n394), .ZN(n620) );
  INV_X1 U715 ( .A(KEYINPUT44), .ZN(n614) );
  INV_X1 U716 ( .A(n607), .ZN(n799) );
  AND2_X1 U717 ( .A1(n614), .A2(n799), .ZN(n616) );
  NOR2_X2 U718 ( .A1(n775), .A2(n690), .ZN(n619) );
  NOR2_X1 U719 ( .A1(n729), .A2(n620), .ZN(n663) );
  XNOR2_X1 U720 ( .A(KEYINPUT106), .B(n621), .ZN(n622) );
  NOR2_X1 U721 ( .A1(G900), .A2(n622), .ZN(n625) );
  INV_X1 U722 ( .A(n623), .ZN(n624) );
  NOR2_X1 U723 ( .A1(n625), .A2(n624), .ZN(n657) );
  INV_X1 U724 ( .A(n641), .ZN(n626) );
  NAND2_X1 U725 ( .A1(n663), .A2(n627), .ZN(n630) );
  XNOR2_X1 U726 ( .A(n631), .B(KEYINPUT110), .ZN(n632) );
  XOR2_X1 U727 ( .A(KEYINPUT113), .B(KEYINPUT41), .Z(n636) );
  INV_X1 U728 ( .A(n743), .ZN(n635) );
  NAND2_X1 U729 ( .A1(n741), .A2(n740), .ZN(n634) );
  XOR2_X1 U730 ( .A(KEYINPUT112), .B(n634), .Z(n738) );
  XNOR2_X1 U731 ( .A(n637), .B(KEYINPUT107), .ZN(n638) );
  NOR2_X1 U732 ( .A1(n638), .A2(n657), .ZN(n640) );
  NAND2_X1 U733 ( .A1(n650), .A2(n741), .ZN(n645) );
  XOR2_X1 U734 ( .A(KEYINPUT39), .B(KEYINPUT84), .Z(n644) );
  XNOR2_X1 U735 ( .A(n645), .B(n644), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n679), .A2(n692), .ZN(n646) );
  XNOR2_X1 U737 ( .A(n646), .B(KEYINPUT40), .ZN(n802) );
  XNOR2_X1 U738 ( .A(n647), .B(KEYINPUT46), .ZN(n677) );
  INV_X1 U739 ( .A(n648), .ZN(n653) );
  AND2_X1 U740 ( .A1(n649), .A2(n650), .ZN(n651) );
  XOR2_X1 U741 ( .A(KEYINPUT79), .B(n704), .Z(n675) );
  NAND2_X1 U742 ( .A1(n655), .A2(n443), .ZN(n670) );
  NAND2_X1 U743 ( .A1(n737), .A2(n705), .ZN(n656) );
  NAND2_X1 U744 ( .A1(n656), .A2(KEYINPUT47), .ZN(n673) );
  INV_X1 U745 ( .A(n740), .ZN(n658) );
  NOR2_X1 U746 ( .A1(n658), .A2(n657), .ZN(n659) );
  NAND2_X1 U747 ( .A1(n660), .A2(n659), .ZN(n661) );
  NOR2_X1 U748 ( .A1(n692), .A2(n661), .ZN(n662) );
  NAND2_X1 U749 ( .A1(n663), .A2(n662), .ZN(n680) );
  NOR2_X1 U750 ( .A1(n683), .A2(n680), .ZN(n664) );
  XOR2_X1 U751 ( .A(KEYINPUT36), .B(n664), .Z(n665) );
  NOR2_X1 U752 ( .A1(n724), .A2(n665), .ZN(n713) );
  NOR2_X1 U753 ( .A1(KEYINPUT78), .A2(n737), .ZN(n668) );
  NAND2_X1 U754 ( .A1(KEYINPUT78), .A2(n737), .ZN(n666) );
  NOR2_X1 U755 ( .A1(KEYINPUT47), .A2(n666), .ZN(n667) );
  NOR2_X1 U756 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U757 ( .A1(n670), .A2(n669), .ZN(n671) );
  NOR2_X1 U758 ( .A1(n713), .A2(n671), .ZN(n672) );
  NAND2_X1 U759 ( .A1(n673), .A2(n672), .ZN(n674) );
  NOR2_X1 U760 ( .A1(n675), .A2(n674), .ZN(n676) );
  NOR2_X1 U761 ( .A1(n679), .A2(n678), .ZN(n715) );
  OR2_X1 U762 ( .A1(n681), .A2(n680), .ZN(n682) );
  XNOR2_X1 U763 ( .A(n682), .B(KEYINPUT43), .ZN(n684) );
  NAND2_X1 U764 ( .A1(n684), .A2(n683), .ZN(n716) );
  INV_X1 U765 ( .A(n716), .ZN(n685) );
  INV_X1 U766 ( .A(n692), .ZN(n707) );
  NAND2_X1 U767 ( .A1(n694), .A2(n707), .ZN(n693) );
  XNOR2_X1 U768 ( .A(n693), .B(G104), .ZN(G6) );
  XNOR2_X1 U769 ( .A(G107), .B(KEYINPUT27), .ZN(n698) );
  XOR2_X1 U770 ( .A(KEYINPUT114), .B(KEYINPUT26), .Z(n696) );
  NAND2_X1 U771 ( .A1(n694), .A2(n709), .ZN(n695) );
  XNOR2_X1 U772 ( .A(n696), .B(n695), .ZN(n697) );
  XNOR2_X1 U773 ( .A(n698), .B(n697), .ZN(G9) );
  XNOR2_X1 U774 ( .A(n444), .B(G110), .ZN(n700) );
  XNOR2_X1 U775 ( .A(n700), .B(KEYINPUT115), .ZN(G12) );
  XOR2_X1 U776 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n702) );
  NAND2_X1 U777 ( .A1(n705), .A2(n709), .ZN(n701) );
  XNOR2_X1 U778 ( .A(n702), .B(n701), .ZN(n703) );
  XNOR2_X1 U779 ( .A(G128), .B(n703), .ZN(G30) );
  XOR2_X1 U780 ( .A(G143), .B(n704), .Z(G45) );
  NAND2_X1 U781 ( .A1(n705), .A2(n707), .ZN(n706) );
  XNOR2_X1 U782 ( .A(n706), .B(G146), .ZN(G48) );
  NAND2_X1 U783 ( .A1(n710), .A2(n707), .ZN(n708) );
  XNOR2_X1 U784 ( .A(n708), .B(G113), .ZN(G15) );
  XOR2_X1 U785 ( .A(G116), .B(KEYINPUT117), .Z(n712) );
  NAND2_X1 U786 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U787 ( .A(n712), .B(n711), .ZN(G18) );
  XNOR2_X1 U788 ( .A(G125), .B(n713), .ZN(n714) );
  XNOR2_X1 U789 ( .A(n714), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U790 ( .A(G134), .B(n715), .Z(G36) );
  XNOR2_X1 U791 ( .A(G140), .B(n716), .ZN(G42) );
  NAND2_X1 U792 ( .A1(n791), .A2(n371), .ZN(n717) );
  XNOR2_X1 U793 ( .A(n717), .B(KEYINPUT80), .ZN(n719) );
  NAND2_X1 U794 ( .A1(n719), .A2(n718), .ZN(n720) );
  INV_X1 U795 ( .A(n723), .ZN(n754) );
  NAND2_X1 U796 ( .A1(n724), .A2(n587), .ZN(n725) );
  XNOR2_X1 U797 ( .A(n725), .B(KEYINPUT50), .ZN(n727) );
  NAND2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n732) );
  NAND2_X1 U799 ( .A1(n729), .A2(n394), .ZN(n730) );
  XNOR2_X1 U800 ( .A(KEYINPUT49), .B(n730), .ZN(n731) );
  NOR2_X1 U801 ( .A1(n732), .A2(n731), .ZN(n733) );
  NOR2_X1 U802 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U803 ( .A(KEYINPUT51), .B(n735), .Z(n736) );
  NOR2_X1 U804 ( .A1(n754), .A2(n736), .ZN(n749) );
  NAND2_X1 U805 ( .A1(n738), .A2(n737), .ZN(n739) );
  XNOR2_X1 U806 ( .A(KEYINPUT119), .B(n739), .ZN(n746) );
  NOR2_X1 U807 ( .A1(n741), .A2(n740), .ZN(n742) );
  NOR2_X1 U808 ( .A1(n743), .A2(n742), .ZN(n744) );
  XNOR2_X1 U809 ( .A(n744), .B(KEYINPUT118), .ZN(n745) );
  NOR2_X1 U810 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U811 ( .A1(n755), .A2(n747), .ZN(n748) );
  NOR2_X1 U812 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U813 ( .A(n750), .B(KEYINPUT52), .ZN(n751) );
  XNOR2_X1 U814 ( .A(KEYINPUT120), .B(n751), .ZN(n752) );
  NOR2_X1 U815 ( .A1(n753), .A2(n752), .ZN(n757) );
  NOR2_X1 U816 ( .A1(n755), .A2(n754), .ZN(n756) );
  NOR2_X1 U817 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U818 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n762) );
  XNOR2_X1 U819 ( .A(n441), .B(KEYINPUT87), .ZN(n761) );
  XNOR2_X1 U820 ( .A(KEYINPUT58), .B(KEYINPUT123), .ZN(n765) );
  XNOR2_X1 U821 ( .A(n763), .B(KEYINPUT57), .ZN(n764) );
  XOR2_X1 U822 ( .A(KEYINPUT59), .B(KEYINPUT66), .Z(n766) );
  XNOR2_X1 U823 ( .A(n769), .B(n768), .ZN(n770) );
  NOR2_X1 U824 ( .A1(n770), .A2(n774), .ZN(G63) );
  XNOR2_X1 U825 ( .A(n395), .B(n771), .ZN(n773) );
  NOR2_X1 U826 ( .A1(n773), .A2(n774), .ZN(G66) );
  XNOR2_X1 U827 ( .A(KEYINPUT125), .B(KEYINPUT127), .ZN(n788) );
  NAND2_X1 U828 ( .A1(n374), .A2(G224), .ZN(n776) );
  XNOR2_X1 U829 ( .A(KEYINPUT61), .B(n776), .ZN(n777) );
  NAND2_X1 U830 ( .A1(n777), .A2(G898), .ZN(n778) );
  NAND2_X1 U831 ( .A1(n779), .A2(n778), .ZN(n786) );
  XNOR2_X1 U832 ( .A(n442), .B(KEYINPUT126), .ZN(n782) );
  XNOR2_X1 U833 ( .A(G101), .B(n780), .ZN(n781) );
  XNOR2_X1 U834 ( .A(n782), .B(n781), .ZN(n784) );
  NOR2_X1 U835 ( .A1(G898), .A2(n792), .ZN(n783) );
  NOR2_X1 U836 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U837 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U838 ( .A(n788), .B(n787), .ZN(G69) );
  XNOR2_X1 U839 ( .A(n789), .B(n790), .ZN(n794) );
  XNOR2_X1 U840 ( .A(n791), .B(n794), .ZN(n793) );
  NAND2_X1 U841 ( .A1(n793), .A2(n792), .ZN(n798) );
  XNOR2_X1 U842 ( .A(G227), .B(n794), .ZN(n795) );
  NAND2_X1 U843 ( .A1(n795), .A2(G900), .ZN(n796) );
  NAND2_X1 U844 ( .A1(n796), .A2(n374), .ZN(n797) );
  NAND2_X1 U845 ( .A1(n798), .A2(n797), .ZN(G72) );
  XNOR2_X1 U846 ( .A(G122), .B(n799), .ZN(G24) );
  XOR2_X1 U847 ( .A(G101), .B(n800), .Z(G3) );
  XOR2_X1 U848 ( .A(G119), .B(n801), .Z(G21) );
  XOR2_X1 U849 ( .A(n802), .B(G131), .Z(G33) );
  XOR2_X1 U850 ( .A(n803), .B(G137), .Z(G39) );
endmodule

