//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 1 1 1 1 0 1 1 1 1 0 0 0 1 0 0 0 1 0 0 0 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 1 0 0 0 1 1 1 0 0 0 0 0 1 1 0 1 1 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:33 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1217, new_n1218,
    new_n1219, new_n1221, new_n1222, new_n1223, new_n1224, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1288, new_n1289, new_n1290;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  NOR2_X1   g0005(.A1(new_n205), .A2(G13), .ZN(new_n206));
  OAI211_X1 g0006(.A(new_n206), .B(G250), .C1(G257), .C2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT0), .ZN(new_n208));
  NAND2_X1  g0008(.A1(new_n202), .A2(G50), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NAND2_X1  g0010(.A1(G1), .A2(G13), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n210), .A2(new_n213), .ZN(new_n214));
  AOI22_X1  g0014(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n215));
  INV_X1    g0015(.A(G68), .ZN(new_n216));
  INV_X1    g0016(.A(G238), .ZN(new_n217));
  INV_X1    g0017(.A(G87), .ZN(new_n218));
  INV_X1    g0018(.A(G250), .ZN(new_n219));
  OAI221_X1 g0019(.A(new_n215), .B1(new_n216), .B2(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  INV_X1    g0021(.A(G77), .ZN(new_n222));
  INV_X1    g0022(.A(G244), .ZN(new_n223));
  INV_X1    g0023(.A(G107), .ZN(new_n224));
  INV_X1    g0024(.A(G264), .ZN(new_n225));
  OAI221_X1 g0025(.A(new_n221), .B1(new_n222), .B2(new_n223), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n205), .B1(new_n220), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n208), .B(new_n214), .C1(KEYINPUT1), .C2(new_n227), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XOR2_X1   g0029(.A(G238), .B(G244), .Z(new_n230));
  XNOR2_X1  g0030(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(G226), .B(G232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XOR2_X1   g0034(.A(G264), .B(G270), .Z(new_n235));
  XNOR2_X1  g0035(.A(G250), .B(G257), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XNOR2_X1  g0038(.A(G50), .B(G68), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G58), .B(G77), .ZN(new_n240));
  XOR2_X1   g0040(.A(new_n239), .B(new_n240), .Z(new_n241));
  XOR2_X1   g0041(.A(G87), .B(G97), .Z(new_n242));
  XNOR2_X1  g0042(.A(G107), .B(G116), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n241), .B(new_n244), .ZN(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n211), .ZN(new_n247));
  OR2_X1    g0047(.A1(KEYINPUT8), .A2(G58), .ZN(new_n248));
  AND2_X1   g0048(.A1(KEYINPUT66), .A2(G58), .ZN(new_n249));
  NOR2_X1   g0049(.A1(KEYINPUT66), .A2(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g0051(.A(KEYINPUT8), .ZN(new_n252));
  OAI21_X1  g0052(.A(new_n248), .B1(new_n251), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n212), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  NOR2_X1   g0055(.A1(G20), .A2(G33), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT67), .ZN(new_n259));
  AND2_X1   g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n261), .B1(new_n258), .B2(new_n259), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n247), .B1(new_n260), .B2(new_n262), .ZN(new_n263));
  INV_X1    g0063(.A(G13), .ZN(new_n264));
  NOR3_X1   g0064(.A1(new_n264), .A2(new_n212), .A3(G1), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(G50), .ZN(new_n267));
  INV_X1    g0067(.A(G1), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n247), .B1(new_n268), .B2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n267), .B1(new_n269), .B2(G50), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n263), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n211), .ZN(new_n273));
  INV_X1    g0073(.A(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(G33), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT3), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n277), .A2(G33), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n276), .A2(new_n278), .ZN(new_n279));
  AOI21_X1  g0079(.A(new_n274), .B1(new_n222), .B2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(G222), .A2(G1698), .ZN(new_n281));
  INV_X1    g0081(.A(G223), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n281), .B1(new_n282), .B2(G1698), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n280), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT65), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n285), .B1(new_n272), .B2(new_n211), .ZN(new_n286));
  OAI21_X1  g0086(.A(new_n268), .B1(G41), .B2(G45), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(G33), .A2(G41), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n289), .A2(KEYINPUT65), .A3(G1), .A4(G13), .ZN(new_n290));
  NAND4_X1  g0090(.A1(new_n286), .A2(new_n288), .A3(G274), .A4(new_n290), .ZN(new_n291));
  AND2_X1   g0091(.A1(new_n286), .A2(new_n290), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n287), .ZN(new_n293));
  INV_X1    g0093(.A(G226), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n284), .B(new_n291), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  OAI211_X1 g0097(.A(new_n271), .B(new_n297), .C1(G179), .C2(new_n295), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  XNOR2_X1  g0099(.A(new_n271), .B(KEYINPUT9), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n295), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n302), .B1(G200), .B2(new_n295), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n300), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n304), .A2(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT10), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n300), .A2(new_n306), .A3(new_n303), .ZN(new_n307));
  AOI21_X1  g0107(.A(new_n299), .B1(new_n305), .B2(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n293), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(G238), .ZN(new_n310));
  MUX2_X1   g0110(.A(G226), .B(G232), .S(G1698), .Z(new_n311));
  XNOR2_X1  g0111(.A(KEYINPUT3), .B(G33), .ZN(new_n312));
  AOI22_X1  g0112(.A1(new_n311), .A2(new_n312), .B1(G33), .B2(G97), .ZN(new_n313));
  OR2_X1    g0113(.A1(new_n313), .A2(new_n274), .ZN(new_n314));
  NAND3_X1  g0114(.A1(new_n310), .A2(new_n291), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT13), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  NAND4_X1  g0117(.A1(new_n310), .A2(new_n317), .A3(new_n291), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  INV_X1    g0120(.A(G200), .ZN(new_n321));
  NOR2_X1   g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(G50), .ZN(new_n323));
  OAI22_X1  g0123(.A1(new_n257), .A2(new_n323), .B1(new_n212), .B2(G68), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n254), .A2(new_n222), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n247), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n269), .A2(G68), .ZN(new_n330));
  NOR3_X1   g0130(.A1(new_n266), .A2(KEYINPUT12), .A3(G68), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT12), .ZN(new_n332));
  AOI21_X1  g0132(.A(new_n332), .B1(new_n265), .B2(new_n216), .ZN(new_n333));
  OAI21_X1  g0133(.A(new_n330), .B1(new_n331), .B2(new_n333), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n326), .A2(new_n327), .ZN(new_n335));
  NOR3_X1   g0135(.A1(new_n329), .A2(new_n334), .A3(new_n335), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n336), .B1(new_n319), .B2(new_n301), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n322), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n319), .A2(G169), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n339), .A2(KEYINPUT14), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n320), .A2(G179), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT14), .ZN(new_n342));
  NAND3_X1  g0142(.A1(new_n319), .A2(new_n342), .A3(G169), .ZN(new_n343));
  NAND3_X1  g0143(.A1(new_n340), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n336), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n338), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(new_n291), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n347), .B1(new_n309), .B2(G244), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n312), .A2(G232), .A3(new_n349), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT68), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n279), .A2(new_n217), .A3(new_n349), .ZN(new_n352));
  AOI21_X1  g0152(.A(new_n352), .B1(G107), .B2(new_n279), .ZN(new_n353));
  AND2_X1   g0153(.A1(new_n351), .A2(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n348), .B1(new_n354), .B2(new_n274), .ZN(new_n355));
  OR2_X1    g0155(.A1(new_n355), .A2(G179), .ZN(new_n356));
  XOR2_X1   g0156(.A(KEYINPUT8), .B(G58), .Z(new_n357));
  AOI22_X1  g0157(.A1(new_n357), .A2(new_n256), .B1(G20), .B2(G77), .ZN(new_n358));
  XNOR2_X1  g0158(.A(KEYINPUT15), .B(G87), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n358), .B1(new_n254), .B2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(new_n247), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n269), .A2(G77), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n361), .B(new_n362), .C1(G77), .C2(new_n266), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n355), .A2(new_n296), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n363), .B1(new_n355), .B2(G200), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n366), .B1(new_n301), .B2(new_n355), .ZN(new_n367));
  AND2_X1   g0167(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g0168(.A1(new_n308), .A2(new_n346), .A3(new_n368), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  NAND4_X1  g0170(.A1(new_n286), .A2(G232), .A3(new_n287), .A4(new_n290), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n291), .A2(new_n371), .ZN(new_n372));
  INV_X1    g0172(.A(KEYINPUT72), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT69), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n374), .B1(new_n277), .B2(G33), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n275), .A2(KEYINPUT69), .A3(KEYINPUT3), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n375), .A2(new_n278), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n349), .A2(G223), .ZN(new_n378));
  OAI21_X1  g0178(.A(new_n373), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  OAI22_X1  g0179(.A1(new_n378), .A2(new_n373), .B1(new_n294), .B2(new_n349), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n380), .A2(new_n375), .A3(new_n278), .A4(new_n376), .ZN(new_n381));
  NAND2_X1  g0181(.A1(G33), .A2(G87), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n379), .A2(new_n381), .A3(new_n382), .ZN(new_n383));
  AOI211_X1 g0183(.A(new_n301), .B(new_n372), .C1(new_n383), .C2(new_n273), .ZN(new_n384));
  AND3_X1   g0184(.A1(new_n375), .A2(new_n278), .A3(new_n376), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n282), .A2(G1698), .ZN(new_n386));
  AOI21_X1  g0186(.A(KEYINPUT72), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  AOI22_X1  g0187(.A1(new_n386), .A2(KEYINPUT72), .B1(G226), .B2(G1698), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n382), .B1(new_n388), .B2(new_n377), .ZN(new_n389));
  OAI21_X1  g0189(.A(new_n273), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n372), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n321), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NOR2_X1   g0192(.A1(new_n384), .A2(new_n392), .ZN(new_n393));
  INV_X1    g0193(.A(KEYINPUT16), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT66), .B(G58), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n201), .B1(new_n395), .B2(G68), .ZN(new_n396));
  INV_X1    g0196(.A(G159), .ZN(new_n397));
  OAI22_X1  g0197(.A1(new_n396), .A2(new_n212), .B1(new_n397), .B2(new_n257), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT7), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n399), .B1(new_n312), .B2(G20), .ZN(new_n400));
  NOR2_X1   g0200(.A1(new_n277), .A2(G33), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n275), .A2(KEYINPUT3), .ZN(new_n402));
  OAI211_X1 g0202(.A(KEYINPUT7), .B(new_n212), .C1(new_n401), .C2(new_n402), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n216), .B1(new_n400), .B2(new_n403), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n394), .B1(new_n398), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(KEYINPUT70), .ZN(new_n406));
  INV_X1    g0206(.A(new_n247), .ZN(new_n407));
  OAI21_X1  g0207(.A(KEYINPUT7), .B1(new_n385), .B2(G20), .ZN(new_n408));
  NAND3_X1  g0208(.A1(new_n377), .A2(new_n399), .A3(new_n212), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n408), .A2(G68), .A3(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G68), .B1(new_n249), .B2(new_n250), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n212), .B1(new_n411), .B2(new_n202), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n257), .A2(new_n397), .ZN(new_n413));
  NOR3_X1   g0213(.A1(new_n412), .A2(new_n394), .A3(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n407), .B1(new_n410), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT70), .ZN(new_n416));
  OAI211_X1 g0216(.A(new_n416), .B(new_n394), .C1(new_n398), .C2(new_n404), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n406), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n253), .A2(new_n266), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n419), .B1(new_n253), .B2(new_n269), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n393), .A2(new_n418), .A3(KEYINPUT73), .A4(new_n420), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n421), .B(KEYINPUT17), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n418), .A2(new_n420), .ZN(new_n423));
  INV_X1    g0223(.A(KEYINPUT71), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n418), .A2(KEYINPUT71), .A3(new_n420), .ZN(new_n426));
  INV_X1    g0226(.A(new_n389), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n274), .B1(new_n427), .B2(new_n379), .ZN(new_n428));
  OAI21_X1  g0228(.A(G169), .B1(new_n428), .B2(new_n372), .ZN(new_n429));
  NAND3_X1  g0229(.A1(new_n390), .A2(G179), .A3(new_n391), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g0231(.A1(new_n425), .A2(new_n426), .A3(new_n431), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n432), .A2(KEYINPUT18), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT18), .ZN(new_n434));
  NAND4_X1  g0234(.A1(new_n425), .A2(new_n434), .A3(new_n426), .A4(new_n431), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n422), .A2(new_n433), .A3(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n370), .A2(new_n437), .A3(KEYINPUT74), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT74), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n369), .B2(new_n436), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n440), .ZN(new_n441));
  XNOR2_X1  g0241(.A(G97), .B(G107), .ZN(new_n442));
  INV_X1    g0242(.A(KEYINPUT75), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n442), .B1(new_n443), .B2(KEYINPUT6), .ZN(new_n444));
  MUX2_X1   g0244(.A(new_n443), .B(G97), .S(KEYINPUT6), .Z(new_n445));
  OAI21_X1  g0245(.A(new_n444), .B1(new_n442), .B2(new_n445), .ZN(new_n446));
  OAI22_X1  g0246(.A1(new_n446), .A2(new_n212), .B1(new_n222), .B2(new_n257), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n224), .B1(new_n400), .B2(new_n403), .ZN(new_n448));
  OAI21_X1  g0248(.A(new_n247), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n266), .A2(G97), .ZN(new_n450));
  OAI211_X1 g0250(.A(new_n266), .B(new_n407), .C1(G1), .C2(new_n275), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n450), .B1(new_n452), .B2(G97), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G41), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n455), .A2(KEYINPUT5), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n268), .A2(G45), .ZN(new_n457));
  OAI21_X1  g0257(.A(KEYINPUT78), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(KEYINPUT5), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n459), .A2(G41), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT78), .ZN(new_n461));
  NAND4_X1  g0261(.A1(new_n460), .A2(new_n461), .A3(new_n268), .A4(G45), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n458), .B(new_n462), .C1(new_n459), .C2(G41), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n286), .A2(G274), .A3(new_n290), .ZN(new_n464));
  OR3_X1    g0264(.A1(new_n463), .A2(KEYINPUT79), .A3(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT79), .B1(new_n463), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT77), .ZN(new_n468));
  NOR2_X1   g0268(.A1(new_n223), .A2(G1698), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n469), .A2(KEYINPUT4), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n468), .B1(new_n470), .B2(new_n279), .ZN(new_n471));
  NAND2_X1  g0271(.A1(G33), .A2(G283), .ZN(new_n472));
  NAND4_X1  g0272(.A1(new_n312), .A2(KEYINPUT77), .A3(KEYINPUT4), .A4(new_n469), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n312), .A2(G250), .A3(G1698), .ZN(new_n474));
  NAND4_X1  g0274(.A1(new_n471), .A2(new_n472), .A3(new_n473), .A4(new_n474), .ZN(new_n475));
  XOR2_X1   g0275(.A(KEYINPUT76), .B(KEYINPUT4), .Z(new_n476));
  AOI21_X1  g0276(.A(new_n476), .B1(new_n385), .B2(new_n469), .ZN(new_n477));
  OAI21_X1  g0277(.A(new_n273), .B1(new_n475), .B2(new_n477), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n463), .A2(new_n292), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n479), .A2(G257), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n467), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n454), .B1(G200), .B2(new_n481), .ZN(new_n482));
  AOI22_X1  g0282(.A1(new_n465), .A2(new_n466), .B1(new_n479), .B2(G257), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n483), .A2(KEYINPUT80), .A3(G190), .A4(new_n478), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT80), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n481), .B2(new_n301), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n482), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n481), .A2(new_n296), .ZN(new_n488));
  INV_X1    g0288(.A(G179), .ZN(new_n489));
  NAND3_X1  g0289(.A1(new_n483), .A2(new_n489), .A3(new_n478), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n488), .A2(new_n490), .A3(new_n454), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n265), .A2(KEYINPUT25), .A3(new_n224), .ZN(new_n493));
  INV_X1    g0293(.A(new_n493), .ZN(new_n494));
  AOI21_X1  g0294(.A(KEYINPUT25), .B1(new_n265), .B2(new_n224), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n451), .A2(new_n224), .B1(new_n494), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n312), .A2(new_n212), .A3(G87), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT22), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT82), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G116), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n499), .B1(new_n500), .B2(G20), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n212), .A2(KEYINPUT82), .A3(G33), .A4(G116), .ZN(new_n502));
  AOI22_X1  g0302(.A1(new_n497), .A2(new_n498), .B1(new_n501), .B2(new_n502), .ZN(new_n503));
  NAND4_X1  g0303(.A1(new_n385), .A2(KEYINPUT22), .A3(new_n212), .A4(G87), .ZN(new_n504));
  OAI21_X1  g0304(.A(KEYINPUT23), .B1(new_n212), .B2(G107), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(KEYINPUT83), .ZN(new_n506));
  INV_X1    g0306(.A(KEYINPUT83), .ZN(new_n507));
  OAI211_X1 g0307(.A(new_n507), .B(KEYINPUT23), .C1(new_n212), .C2(G107), .ZN(new_n508));
  OR3_X1    g0308(.A1(new_n212), .A2(KEYINPUT23), .A3(G107), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n506), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n503), .A2(new_n504), .A3(new_n510), .ZN(new_n511));
  XNOR2_X1  g0311(.A(new_n511), .B(KEYINPUT24), .ZN(new_n512));
  AOI21_X1  g0312(.A(new_n496), .B1(new_n512), .B2(new_n247), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(KEYINPUT84), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n463), .A2(G264), .A3(new_n292), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(KEYINPUT85), .ZN(new_n517));
  AND2_X1   g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n219), .A2(new_n349), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n519), .B1(G257), .B2(new_n349), .ZN(new_n520));
  INV_X1    g0320(.A(G294), .ZN(new_n521));
  OAI22_X1  g0321(.A1(new_n520), .A2(new_n377), .B1(new_n275), .B2(new_n521), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n465), .A2(new_n466), .B1(new_n273), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n518), .A2(G179), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n522), .A2(new_n273), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n467), .A2(new_n515), .A3(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n526), .A2(G169), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n524), .A2(new_n527), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT84), .ZN(new_n529));
  OR2_X1    g0329(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n511), .A2(KEYINPUT24), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n407), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n529), .B1(new_n532), .B2(new_n496), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n514), .A2(new_n528), .A3(new_n533), .ZN(new_n534));
  AOI21_X1  g0334(.A(G200), .B1(new_n518), .B2(new_n523), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n526), .A2(G190), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n513), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G97), .ZN(new_n539));
  OAI211_X1 g0339(.A(new_n472), .B(new_n212), .C1(G33), .C2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n540), .B(new_n247), .C1(new_n212), .C2(G116), .ZN(new_n541));
  XOR2_X1   g0341(.A(new_n541), .B(KEYINPUT20), .Z(new_n542));
  NAND2_X1  g0342(.A1(new_n452), .A2(G116), .ZN(new_n543));
  OAI211_X1 g0343(.A(new_n542), .B(new_n543), .C1(G116), .C2(new_n266), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n225), .A2(G1698), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G257), .B2(G1698), .ZN(new_n546));
  INV_X1    g0346(.A(G303), .ZN(new_n547));
  OAI22_X1  g0347(.A1(new_n377), .A2(new_n546), .B1(new_n547), .B2(new_n312), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n479), .A2(G270), .B1(new_n273), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n467), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n544), .B1(new_n550), .B2(G200), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n551), .B1(new_n301), .B2(new_n550), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n544), .A3(G169), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT21), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND4_X1  g0355(.A1(new_n550), .A2(new_n544), .A3(KEYINPUT21), .A4(G169), .ZN(new_n556));
  NAND4_X1  g0356(.A1(new_n544), .A2(G179), .A3(new_n467), .A4(new_n549), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n552), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NOR2_X1   g0358(.A1(new_n216), .A2(G20), .ZN(new_n559));
  NOR3_X1   g0359(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n560));
  AOI21_X1  g0360(.A(G20), .B1(G33), .B2(G97), .ZN(new_n561));
  OAI21_X1  g0361(.A(KEYINPUT19), .B1(new_n560), .B2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT19), .ZN(new_n563));
  NAND4_X1  g0363(.A1(new_n563), .A2(new_n212), .A3(G33), .A4(G97), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n385), .A2(new_n559), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g0365(.A(new_n359), .ZN(new_n566));
  OAI22_X1  g0366(.A1(new_n565), .A2(new_n407), .B1(new_n266), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n452), .A2(new_n566), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n223), .A2(G1698), .ZN(new_n571));
  OAI21_X1  g0371(.A(new_n571), .B1(G238), .B2(G1698), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n500), .B1(new_n377), .B2(new_n572), .ZN(new_n573));
  NOR2_X1   g0373(.A1(new_n457), .A2(G274), .ZN(new_n574));
  AOI21_X1  g0374(.A(new_n574), .B1(new_n219), .B2(new_n457), .ZN(new_n575));
  AOI22_X1  g0375(.A1(new_n273), .A2(new_n573), .B1(new_n575), .B2(new_n292), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n576), .A2(new_n296), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n573), .A2(new_n273), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n575), .A2(new_n292), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g0380(.A1(new_n580), .A2(new_n489), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n570), .B1(new_n577), .B2(new_n581), .ZN(new_n582));
  AOI21_X1  g0382(.A(new_n567), .B1(G87), .B2(new_n452), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(G200), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n576), .A2(G190), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n583), .A2(new_n584), .A3(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  INV_X1    g0387(.A(KEYINPUT81), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n582), .A2(new_n586), .A3(KEYINPUT81), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NOR2_X1   g0391(.A1(new_n558), .A2(new_n591), .ZN(new_n592));
  AND4_X1   g0392(.A1(new_n441), .A2(new_n492), .A3(new_n538), .A4(new_n592), .ZN(G372));
  INV_X1    g0393(.A(KEYINPUT86), .ZN(new_n594));
  OAI21_X1  g0394(.A(new_n594), .B1(new_n581), .B2(new_n577), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n576), .A2(G179), .ZN(new_n596));
  OAI211_X1 g0396(.A(new_n596), .B(KEYINPUT86), .C1(new_n296), .C2(new_n576), .ZN(new_n597));
  AOI22_X1  g0397(.A1(new_n595), .A2(new_n597), .B1(new_n568), .B2(new_n569), .ZN(new_n598));
  INV_X1    g0398(.A(new_n586), .ZN(new_n599));
  NOR3_X1   g0399(.A1(new_n491), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT26), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n598), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g0402(.A(KEYINPUT26), .B1(new_n591), .B2(new_n491), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n555), .A2(new_n556), .A3(new_n557), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n513), .B1(new_n527), .B2(new_n524), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NOR2_X1   g0406(.A1(new_n598), .A2(new_n599), .ZN(new_n607));
  NAND4_X1  g0407(.A1(new_n607), .A2(new_n537), .A3(new_n487), .A4(new_n491), .ZN(new_n608));
  OAI211_X1 g0408(.A(new_n602), .B(new_n603), .C1(new_n606), .C2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n441), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n423), .A2(new_n431), .ZN(new_n611));
  XNOR2_X1  g0411(.A(new_n611), .B(new_n434), .ZN(new_n612));
  INV_X1    g0412(.A(new_n338), .ZN(new_n613));
  INV_X1    g0413(.A(new_n365), .ZN(new_n614));
  AOI22_X1  g0414(.A1(new_n613), .A2(new_n614), .B1(new_n344), .B2(new_n345), .ZN(new_n615));
  INV_X1    g0415(.A(new_n422), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n612), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n305), .A2(new_n307), .ZN(new_n618));
  AOI21_X1  g0418(.A(new_n299), .B1(new_n617), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n610), .A2(new_n619), .ZN(G369));
  INV_X1    g0420(.A(G330), .ZN(new_n621));
  INV_X1    g0421(.A(new_n604), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n268), .A2(new_n212), .A3(G13), .ZN(new_n623));
  OR2_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n623), .A2(KEYINPUT27), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n544), .A2(new_n628), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n622), .A2(new_n552), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n604), .A2(new_n544), .A3(new_n628), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n621), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  INV_X1    g0432(.A(new_n534), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(new_n628), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n514), .A2(new_n533), .A3(new_n628), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n534), .A2(new_n635), .A3(new_n537), .ZN(new_n636));
  NAND2_X1  g0436(.A1(new_n634), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g0437(.A1(new_n632), .A2(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n628), .ZN(new_n639));
  NAND4_X1  g0439(.A1(new_n534), .A2(new_n537), .A3(new_n604), .A4(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n605), .A2(new_n639), .ZN(new_n641));
  AND2_X1   g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NAND2_X1  g0442(.A1(new_n638), .A2(new_n642), .ZN(G399));
  INV_X1    g0443(.A(new_n206), .ZN(new_n644));
  NOR2_X1   g0444(.A1(new_n644), .A2(G41), .ZN(new_n645));
  INV_X1    g0445(.A(G116), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n560), .A2(new_n646), .ZN(new_n647));
  NOR3_X1   g0447(.A1(new_n645), .A2(new_n647), .A3(new_n268), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n648), .B1(new_n210), .B2(new_n645), .ZN(new_n649));
  XOR2_X1   g0449(.A(new_n649), .B(KEYINPUT28), .Z(new_n650));
  AND3_X1   g0450(.A1(new_n488), .A2(new_n454), .A3(new_n490), .ZN(new_n651));
  NAND4_X1  g0451(.A1(new_n589), .A2(new_n651), .A3(new_n601), .A4(new_n590), .ZN(new_n652));
  INV_X1    g0452(.A(new_n598), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n600), .A2(new_n601), .ZN(new_n655));
  NOR2_X1   g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n622), .A2(new_n534), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n657), .A2(new_n492), .A3(new_n537), .A4(new_n607), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n628), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(KEYINPUT88), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n660), .A3(KEYINPUT29), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n516), .A2(new_n525), .A3(new_n517), .A4(new_n576), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n662), .A2(new_n481), .ZN(new_n663));
  INV_X1    g0463(.A(KEYINPUT87), .ZN(new_n664));
  OAI21_X1  g0464(.A(new_n664), .B1(new_n550), .B2(new_n489), .ZN(new_n665));
  NAND4_X1  g0465(.A1(new_n467), .A2(new_n549), .A3(KEYINPUT87), .A4(G179), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n663), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT30), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n663), .A2(new_n665), .A3(KEYINPUT30), .A4(new_n666), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n518), .A2(new_n523), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n576), .A2(G179), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n671), .A2(new_n481), .A3(new_n550), .A4(new_n672), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n669), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n674), .A2(new_n628), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT31), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n592), .A2(new_n538), .A3(new_n492), .A4(new_n639), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n674), .A2(KEYINPUT31), .A3(new_n628), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(G330), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n608), .B1(new_n534), .B2(new_n622), .ZN(new_n682));
  OAI211_X1 g0482(.A(new_n652), .B(new_n653), .C1(new_n601), .C2(new_n600), .ZN(new_n683));
  OAI211_X1 g0483(.A(KEYINPUT29), .B(new_n639), .C1(new_n682), .C2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n684), .A2(KEYINPUT88), .ZN(new_n685));
  AOI21_X1  g0485(.A(KEYINPUT29), .B1(new_n609), .B2(new_n639), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n661), .B(new_n681), .C1(new_n685), .C2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n650), .B1(new_n688), .B2(G1), .ZN(G364));
  NAND2_X1  g0489(.A1(new_n630), .A2(new_n631), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n690), .A2(G330), .ZN(new_n691));
  XNOR2_X1  g0491(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  INV_X1    g0492(.A(new_n632), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n264), .A2(G20), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n268), .B1(new_n694), .B2(G45), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n645), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n692), .A2(new_n693), .A3(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n312), .A2(G355), .A3(new_n206), .ZN(new_n700));
  OAI21_X1  g0500(.A(new_n700), .B1(G116), .B2(new_n206), .ZN(new_n701));
  INV_X1    g0501(.A(G45), .ZN(new_n702));
  OR2_X1    g0502(.A1(new_n241), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n385), .A2(new_n644), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n702), .B2(new_n210), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n701), .B1(new_n703), .B2(new_n706), .ZN(new_n707));
  NOR2_X1   g0507(.A1(G13), .A2(G33), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n709), .A2(G20), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n211), .B1(G20), .B2(new_n296), .ZN(new_n711));
  NOR2_X1   g0511(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  OAI21_X1  g0513(.A(new_n697), .B1(new_n707), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n212), .A2(G179), .ZN(new_n715));
  NAND3_X1  g0515(.A1(new_n715), .A2(new_n301), .A3(G200), .ZN(new_n716));
  INV_X1    g0516(.A(G283), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n301), .A2(G200), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n719), .A2(new_n489), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G20), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n715), .A2(G190), .A3(G200), .ZN(new_n723));
  OAI22_X1  g0523(.A1(new_n722), .A2(new_n521), .B1(new_n723), .B2(new_n547), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n212), .A2(new_n489), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n725), .A2(G200), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(new_n301), .ZN(new_n727));
  AOI211_X1 g0527(.A(new_n718), .B(new_n724), .C1(G326), .C2(new_n727), .ZN(new_n728));
  XNOR2_X1  g0528(.A(KEYINPUT33), .B(G317), .ZN(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n726), .A2(G190), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n730), .A2(KEYINPUT93), .ZN(new_n733));
  NAND3_X1  g0533(.A1(new_n731), .A2(new_n732), .A3(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT90), .ZN(new_n735));
  AND3_X1   g0535(.A1(new_n725), .A2(new_n735), .A3(new_n719), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n735), .B1(new_n725), .B2(new_n719), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n739), .A2(G322), .ZN(new_n740));
  NOR2_X1   g0540(.A1(G190), .A2(G200), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n725), .A2(new_n741), .ZN(new_n742));
  INV_X1    g0542(.A(G311), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n715), .A2(new_n741), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  AOI211_X1 g0546(.A(new_n312), .B(new_n744), .C1(G329), .C2(new_n746), .ZN(new_n747));
  NAND4_X1  g0547(.A1(new_n728), .A2(new_n734), .A3(new_n740), .A4(new_n747), .ZN(new_n748));
  AOI22_X1  g0548(.A1(new_n732), .A2(G68), .B1(new_n721), .B2(G97), .ZN(new_n749));
  XNOR2_X1  g0549(.A(new_n749), .B(KEYINPUT92), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT91), .B(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n745), .A2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(KEYINPUT32), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  INV_X1    g0554(.A(new_n727), .ZN(new_n755));
  OAI21_X1  g0555(.A(new_n754), .B1(new_n755), .B2(new_n323), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n738), .A2(new_n251), .ZN(new_n757));
  OAI22_X1  g0557(.A1(new_n752), .A2(new_n753), .B1(new_n224), .B2(new_n716), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n312), .B1(new_n742), .B2(new_n222), .C1(new_n218), .C2(new_n723), .ZN(new_n759));
  OR4_X1    g0559(.A1(new_n756), .A2(new_n757), .A3(new_n758), .A4(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n748), .B1(new_n750), .B2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n714), .B1(new_n761), .B2(new_n711), .ZN(new_n762));
  INV_X1    g0562(.A(new_n710), .ZN(new_n763));
  OAI21_X1  g0563(.A(new_n762), .B1(new_n690), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n699), .A2(new_n764), .ZN(G396));
  NAND2_X1  g0565(.A1(new_n363), .A2(new_n628), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n365), .A2(new_n367), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n767), .A2(KEYINPUT94), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n614), .A2(new_n628), .ZN(new_n769));
  INV_X1    g0569(.A(KEYINPUT94), .ZN(new_n770));
  NAND4_X1  g0570(.A1(new_n365), .A2(new_n367), .A3(new_n770), .A4(new_n766), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n768), .A2(new_n769), .A3(new_n771), .ZN(new_n772));
  XNOR2_X1  g0572(.A(new_n772), .B(KEYINPUT95), .ZN(new_n773));
  INV_X1    g0573(.A(new_n609), .ZN(new_n774));
  OAI21_X1  g0574(.A(new_n773), .B1(new_n774), .B2(new_n628), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n768), .A2(new_n771), .ZN(new_n776));
  NAND3_X1  g0576(.A1(new_n609), .A2(new_n639), .A3(new_n776), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n697), .B1(new_n778), .B2(new_n681), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n779), .B1(new_n681), .B2(new_n778), .ZN(new_n780));
  INV_X1    g0580(.A(new_n711), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n781), .A2(new_n709), .ZN(new_n782));
  OAI21_X1  g0582(.A(new_n697), .B1(new_n782), .B2(G77), .ZN(new_n783));
  INV_X1    g0583(.A(new_n732), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n784), .A2(new_n717), .B1(new_n224), .B2(new_n723), .ZN(new_n785));
  AOI21_X1  g0585(.A(new_n785), .B1(G303), .B2(new_n727), .ZN(new_n786));
  NAND2_X1  g0586(.A1(new_n739), .A2(G294), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n279), .B1(new_n742), .B2(new_n646), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n788), .B1(G311), .B2(new_n746), .ZN(new_n789));
  INV_X1    g0589(.A(new_n716), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n790), .A2(G87), .B1(new_n721), .B2(G97), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n786), .A2(new_n787), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(new_n742), .ZN(new_n793));
  INV_X1    g0593(.A(new_n751), .ZN(new_n794));
  AOI22_X1  g0594(.A1(new_n727), .A2(G137), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n795), .B1(new_n255), .B2(new_n784), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n796), .B1(G143), .B2(new_n739), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n798));
  INV_X1    g0598(.A(G132), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n385), .B1(new_n799), .B2(new_n745), .ZN(new_n800));
  OAI22_X1  g0600(.A1(new_n722), .A2(new_n251), .B1(new_n716), .B2(new_n216), .ZN(new_n801));
  INV_X1    g0601(.A(new_n723), .ZN(new_n802));
  AOI211_X1 g0602(.A(new_n800), .B(new_n801), .C1(G50), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n797), .A2(KEYINPUT34), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n792), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n783), .B1(new_n806), .B2(new_n711), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n807), .B1(new_n772), .B2(new_n709), .ZN(new_n808));
  AND2_X1   g0608(.A1(new_n780), .A2(new_n808), .ZN(new_n809));
  INV_X1    g0609(.A(new_n809), .ZN(G384));
  INV_X1    g0610(.A(KEYINPUT97), .ZN(new_n811));
  NAND3_X1  g0611(.A1(new_n393), .A2(new_n418), .A3(new_n420), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n409), .A2(G68), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n399), .B1(new_n377), .B2(new_n212), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OAI221_X1 g0615(.A(KEYINPUT16), .B1(new_n397), .B2(new_n257), .C1(new_n396), .C2(new_n212), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n247), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n398), .ZN(new_n818));
  AOI21_X1  g0618(.A(KEYINPUT16), .B1(new_n410), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g0619(.A(new_n420), .B1(new_n817), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n820), .A2(new_n431), .ZN(new_n821));
  INV_X1    g0621(.A(new_n626), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g0623(.A1(new_n812), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  AND2_X1   g0624(.A1(new_n824), .A2(KEYINPUT37), .ZN(new_n825));
  INV_X1    g0625(.A(KEYINPUT37), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n812), .A2(new_n826), .ZN(new_n827));
  AND3_X1   g0627(.A1(new_n418), .A2(KEYINPUT71), .A3(new_n420), .ZN(new_n828));
  AOI21_X1  g0628(.A(KEYINPUT71), .B1(new_n418), .B2(new_n420), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n827), .B1(new_n830), .B2(new_n431), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n425), .A2(new_n426), .A3(new_n822), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n825), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT96), .ZN(new_n834));
  INV_X1    g0634(.A(new_n823), .ZN(new_n835));
  AOI22_X1  g0635(.A1(new_n833), .A2(new_n834), .B1(new_n436), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n827), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n432), .A2(new_n832), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n824), .A2(KEYINPUT37), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n840), .A2(KEYINPUT96), .ZN(new_n841));
  AOI21_X1  g0641(.A(KEYINPUT38), .B1(new_n836), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n436), .A2(new_n835), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n838), .A2(new_n834), .A3(new_n839), .ZN(new_n844));
  AND4_X1   g0644(.A1(KEYINPUT38), .A2(new_n841), .A3(new_n843), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n811), .B1(new_n842), .B2(new_n845), .ZN(new_n846));
  NAND3_X1  g0646(.A1(new_n841), .A2(new_n843), .A3(new_n844), .ZN(new_n847));
  INV_X1    g0647(.A(KEYINPUT38), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n836), .A2(KEYINPUT38), .A3(new_n841), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT97), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(new_n772), .ZN(new_n853));
  OAI21_X1  g0653(.A(new_n346), .B1(new_n336), .B2(new_n639), .ZN(new_n854));
  OAI211_X1 g0654(.A(new_n345), .B(new_n628), .C1(new_n344), .C2(new_n338), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n853), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n856), .A2(new_n680), .ZN(new_n857));
  INV_X1    g0657(.A(new_n857), .ZN(new_n858));
  AOI21_X1  g0658(.A(KEYINPUT40), .B1(new_n852), .B2(new_n858), .ZN(new_n859));
  NOR3_X1   g0659(.A1(new_n828), .A2(new_n829), .A3(new_n626), .ZN(new_n860));
  NAND2_X1  g0660(.A1(new_n611), .A2(new_n812), .ZN(new_n861));
  OAI21_X1  g0661(.A(KEYINPUT37), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  AOI21_X1  g0662(.A(KEYINPUT98), .B1(new_n862), .B2(new_n838), .ZN(new_n863));
  AOI21_X1  g0663(.A(new_n832), .B1(new_n612), .B2(new_n422), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(KEYINPUT98), .A3(new_n838), .ZN(new_n866));
  AND2_X1   g0666(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n850), .B1(new_n867), .B2(KEYINPUT38), .ZN(new_n868));
  AND3_X1   g0668(.A1(new_n856), .A2(KEYINPUT40), .A3(new_n680), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n859), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  AND2_X1   g0670(.A1(new_n441), .A2(new_n680), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n870), .A2(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n872), .ZN(new_n873));
  NOR2_X1   g0673(.A1(new_n870), .A2(new_n871), .ZN(new_n874));
  NOR3_X1   g0674(.A1(new_n873), .A2(new_n621), .A3(new_n874), .ZN(new_n875));
  NOR2_X1   g0675(.A1(new_n365), .A2(new_n628), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n777), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n854), .A2(new_n855), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  INV_X1    g0680(.A(new_n880), .ZN(new_n881));
  INV_X1    g0681(.A(new_n851), .ZN(new_n882));
  AOI21_X1  g0682(.A(KEYINPUT97), .B1(new_n849), .B2(new_n850), .ZN(new_n883));
  OAI21_X1  g0683(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT39), .ZN(new_n885));
  AOI21_X1  g0685(.A(KEYINPUT38), .B1(new_n865), .B2(new_n866), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n885), .B1(new_n886), .B2(new_n845), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n344), .A2(new_n345), .A3(new_n639), .ZN(new_n888));
  INV_X1    g0688(.A(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n849), .A2(new_n850), .A3(KEYINPUT39), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n887), .A2(new_n889), .A3(new_n890), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n612), .A2(new_n822), .ZN(new_n892));
  AND3_X1   g0692(.A1(new_n884), .A2(new_n891), .A3(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n661), .B1(new_n685), .B2(new_n686), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT99), .ZN(new_n895));
  AND3_X1   g0695(.A1(new_n441), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n895), .B1(new_n441), .B2(new_n894), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n619), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  XNOR2_X1  g0698(.A(new_n893), .B(new_n898), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n875), .A2(new_n899), .B1(new_n268), .B2(new_n694), .ZN(new_n900));
  AOI21_X1  g0700(.A(new_n900), .B1(new_n899), .B2(new_n875), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  OAI211_X1 g0702(.A(G116), .B(new_n213), .C1(new_n446), .C2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n446), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n904), .B(KEYINPUT36), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n210), .A2(G77), .A3(new_n411), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n323), .A2(G68), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n268), .B(G13), .C1(new_n906), .C2(new_n907), .ZN(new_n908));
  OR3_X1    g0708(.A1(new_n901), .A2(new_n905), .A3(new_n908), .ZN(G367));
  OR2_X1    g0709(.A1(new_n583), .A2(new_n639), .ZN(new_n910));
  OR2_X1    g0710(.A1(new_n653), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n607), .A2(new_n910), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n454), .A2(new_n628), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n492), .A2(new_n916), .B1(new_n651), .B2(new_n628), .ZN(new_n917));
  NOR2_X1   g0717(.A1(new_n917), .A2(KEYINPUT102), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n487), .A2(new_n491), .A3(new_n916), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n491), .B2(new_n639), .ZN(new_n920));
  INV_X1    g0720(.A(KEYINPUT102), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n633), .B1(new_n918), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n628), .B1(new_n923), .B2(new_n491), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n917), .A2(new_n640), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT42), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n925), .B(new_n926), .ZN(new_n927));
  OAI21_X1  g0727(.A(new_n915), .B1(new_n924), .B2(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(KEYINPUT100), .B(KEYINPUT43), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n913), .A2(new_n929), .ZN(new_n930));
  XOR2_X1   g0730(.A(new_n930), .B(KEYINPUT101), .Z(new_n931));
  NAND2_X1  g0731(.A1(new_n928), .A2(new_n931), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n918), .A2(new_n922), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n933), .A2(new_n638), .ZN(new_n934));
  INV_X1    g0734(.A(new_n931), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n935), .B(new_n915), .C1(new_n924), .C2(new_n927), .ZN(new_n936));
  AND3_X1   g0736(.A1(new_n932), .A2(new_n934), .A3(new_n936), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n934), .B1(new_n932), .B2(new_n936), .ZN(new_n938));
  NOR2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  XOR2_X1   g0739(.A(new_n645), .B(KEYINPUT41), .Z(new_n940));
  NOR2_X1   g0740(.A1(new_n684), .A2(KEYINPUT88), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n660), .B1(new_n659), .B2(KEYINPUT29), .ZN(new_n942));
  INV_X1    g0742(.A(new_n686), .ZN(new_n943));
  AOI21_X1  g0743(.A(new_n941), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n634), .B(new_n636), .C1(new_n622), .C2(new_n628), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n640), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n632), .A2(KEYINPUT104), .ZN(new_n947));
  INV_X1    g0747(.A(KEYINPUT104), .ZN(new_n948));
  AOI211_X1 g0748(.A(new_n948), .B(new_n621), .C1(new_n630), .C2(new_n631), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n946), .B1(new_n947), .B2(new_n949), .ZN(new_n950));
  OAI211_X1 g0750(.A(new_n945), .B(new_n640), .C1(new_n632), .C2(KEYINPUT104), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NAND4_X1  g0752(.A1(new_n944), .A2(new_n952), .A3(KEYINPUT105), .A4(new_n681), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n950), .A2(new_n951), .ZN(new_n955));
  OAI21_X1  g0755(.A(new_n954), .B1(new_n687), .B2(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT45), .ZN(new_n957));
  INV_X1    g0757(.A(KEYINPUT103), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n958), .B1(new_n642), .B2(new_n920), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n640), .A2(new_n641), .ZN(new_n960));
  NOR3_X1   g0760(.A1(new_n960), .A2(new_n917), .A3(KEYINPUT103), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n957), .B1(new_n959), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n917), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT44), .ZN(new_n964));
  XNOR2_X1  g0764(.A(new_n963), .B(new_n964), .ZN(new_n965));
  NAND3_X1  g0765(.A1(new_n642), .A2(new_n958), .A3(new_n920), .ZN(new_n966));
  OAI21_X1  g0766(.A(KEYINPUT103), .B1(new_n917), .B2(new_n960), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n966), .A2(new_n967), .A3(KEYINPUT45), .ZN(new_n968));
  NAND4_X1  g0768(.A1(new_n962), .A2(new_n965), .A3(new_n638), .A4(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n962), .A2(new_n965), .A3(new_n968), .ZN(new_n970));
  INV_X1    g0770(.A(new_n638), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n953), .A2(new_n956), .A3(new_n969), .A4(new_n972), .ZN(new_n973));
  AOI21_X1  g0773(.A(new_n940), .B1(new_n973), .B2(new_n688), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n939), .B1(new_n974), .B2(new_n696), .ZN(new_n975));
  OAI221_X1 g0775(.A(new_n712), .B1(new_n206), .B2(new_n359), .C1(new_n705), .C2(new_n237), .ZN(new_n976));
  AND2_X1   g0776(.A1(new_n976), .A2(new_n697), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT106), .B1(new_n802), .B2(G116), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT46), .ZN(new_n979));
  AOI22_X1  g0779(.A1(new_n732), .A2(G294), .B1(new_n721), .B2(G107), .ZN(new_n980));
  NOR2_X1   g0780(.A1(new_n716), .A2(new_n539), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n981), .B1(G311), .B2(new_n727), .ZN(new_n982));
  INV_X1    g0782(.A(G317), .ZN(new_n983));
  OAI221_X1 g0783(.A(new_n377), .B1(new_n745), .B2(new_n983), .C1(new_n717), .C2(new_n742), .ZN(new_n984));
  AOI21_X1  g0784(.A(new_n984), .B1(new_n739), .B2(G303), .ZN(new_n985));
  NAND4_X1  g0785(.A1(new_n979), .A2(new_n980), .A3(new_n982), .A4(new_n985), .ZN(new_n986));
  XNOR2_X1  g0786(.A(new_n986), .B(KEYINPUT107), .ZN(new_n987));
  OAI22_X1  g0787(.A1(new_n738), .A2(new_n255), .B1(new_n722), .B2(new_n216), .ZN(new_n988));
  XOR2_X1   g0788(.A(new_n988), .B(KEYINPUT108), .Z(new_n989));
  XNOR2_X1  g0789(.A(KEYINPUT109), .B(G137), .ZN(new_n990));
  OAI221_X1 g0790(.A(new_n312), .B1(new_n745), .B2(new_n990), .C1(new_n323), .C2(new_n742), .ZN(new_n991));
  INV_X1    g0791(.A(new_n991), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n732), .A2(new_n794), .B1(new_n802), .B2(new_n395), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n716), .A2(new_n222), .ZN(new_n994));
  AOI21_X1  g0794(.A(new_n994), .B1(G143), .B2(new_n727), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n992), .A2(new_n993), .A3(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n987), .B1(new_n989), .B2(new_n996), .ZN(new_n997));
  XOR2_X1   g0797(.A(new_n997), .B(KEYINPUT47), .Z(new_n998));
  OAI221_X1 g0798(.A(new_n977), .B1(new_n914), .B2(new_n763), .C1(new_n998), .C2(new_n781), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n975), .A2(new_n999), .ZN(G387));
  NAND2_X1  g0800(.A1(new_n688), .A2(new_n952), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n687), .A2(new_n955), .ZN(new_n1002));
  XNOR2_X1  g0802(.A(new_n645), .B(KEYINPUT113), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n634), .A2(new_n636), .A3(new_n710), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n732), .A2(G311), .B1(new_n793), .B2(G303), .ZN(new_n1006));
  INV_X1    g0806(.A(G322), .ZN(new_n1007));
  OAI221_X1 g0807(.A(new_n1006), .B1(new_n1007), .B2(new_n755), .C1(new_n738), .C2(new_n983), .ZN(new_n1008));
  INV_X1    g0808(.A(KEYINPUT48), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n802), .A2(G294), .B1(new_n721), .B2(G283), .ZN(new_n1012));
  NAND3_X1  g0812(.A1(new_n1010), .A2(new_n1011), .A3(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT49), .ZN(new_n1014));
  OR2_X1    g0814(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n716), .A2(new_n646), .ZN(new_n1017));
  AOI211_X1 g0817(.A(new_n385), .B(new_n1017), .C1(G326), .C2(new_n746), .ZN(new_n1018));
  NAND3_X1  g0818(.A1(new_n1015), .A2(new_n1016), .A3(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n727), .A2(G159), .ZN(new_n1020));
  XOR2_X1   g0820(.A(new_n1020), .B(KEYINPUT112), .Z(new_n1021));
  NOR2_X1   g0821(.A1(new_n723), .A2(new_n222), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n722), .A2(new_n359), .ZN(new_n1023));
  NOR4_X1   g0823(.A1(new_n1021), .A2(new_n981), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n385), .B1(new_n216), .B2(new_n742), .C1(new_n255), .C2(new_n745), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n1025), .B1(new_n739), .B2(G50), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n1024), .B(new_n1026), .C1(new_n253), .C2(new_n784), .ZN(new_n1027));
  AOI21_X1  g0827(.A(new_n781), .B1(new_n1019), .B2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g0828(.A1(new_n647), .A2(new_n206), .A3(new_n312), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(G107), .B2(new_n206), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT110), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n357), .A2(new_n323), .ZN(new_n1032));
  XNOR2_X1  g0832(.A(new_n1032), .B(KEYINPUT50), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  AOI211_X1 g0834(.A(G45), .B(new_n647), .C1(G68), .C2(G77), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n705), .B1(new_n1034), .B2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT111), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  OAI21_X1  g0838(.A(new_n1038), .B1(new_n702), .B2(new_n234), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1040));
  OAI21_X1  g0840(.A(new_n1031), .B1(new_n1039), .B2(new_n1040), .ZN(new_n1041));
  AOI211_X1 g0841(.A(new_n698), .B(new_n1028), .C1(new_n712), .C2(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n952), .A2(new_n696), .B1(new_n1005), .B2(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1004), .A2(new_n1043), .ZN(G393));
  INV_X1    g0844(.A(KEYINPUT114), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n972), .A2(new_n1045), .A3(new_n969), .ZN(new_n1046));
  OR3_X1    g0846(.A1(new_n970), .A2(new_n1045), .A3(new_n971), .ZN(new_n1047));
  NAND3_X1  g0847(.A1(new_n1046), .A2(new_n1047), .A3(new_n1001), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1048), .A2(new_n973), .A3(new_n1003), .ZN(new_n1049));
  OAI221_X1 g0849(.A(new_n712), .B1(new_n539), .B2(new_n206), .C1(new_n705), .C2(new_n244), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n397), .A2(new_n738), .B1(new_n755), .B2(new_n255), .ZN(new_n1051));
  XNOR2_X1  g0851(.A(new_n1051), .B(KEYINPUT51), .ZN(new_n1052));
  NOR2_X1   g0852(.A1(new_n722), .A2(new_n222), .ZN(new_n1053));
  AOI21_X1  g0853(.A(new_n1053), .B1(G50), .B2(new_n732), .ZN(new_n1054));
  AOI22_X1  g0854(.A1(new_n357), .A2(new_n793), .B1(new_n746), .B2(G143), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n802), .A2(G68), .B1(new_n790), .B2(G87), .ZN(new_n1056));
  AND4_X1   g0856(.A1(new_n385), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  OAI221_X1 g0857(.A(new_n279), .B1(new_n742), .B2(new_n521), .C1(new_n224), .C2(new_n716), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n784), .A2(new_n547), .B1(new_n722), .B2(new_n646), .ZN(new_n1059));
  OAI22_X1  g0859(.A1(new_n723), .A2(new_n717), .B1(new_n745), .B2(new_n1007), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(KEYINPUT116), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1058), .B(new_n1059), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  OAI22_X1  g0863(.A1(new_n743), .A2(new_n738), .B1(new_n755), .B2(new_n983), .ZN(new_n1064));
  XOR2_X1   g0864(.A(KEYINPUT115), .B(KEYINPUT52), .Z(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  AOI22_X1  g0866(.A1(new_n1052), .A2(new_n1057), .B1(new_n1063), .B2(new_n1066), .ZN(new_n1067));
  OAI211_X1 g0867(.A(new_n697), .B(new_n1050), .C1(new_n1067), .C2(new_n781), .ZN(new_n1068));
  XOR2_X1   g0868(.A(new_n1068), .B(KEYINPUT117), .Z(new_n1069));
  AOI21_X1  g0869(.A(new_n1069), .B1(new_n933), .B2(new_n710), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1046), .A2(new_n1047), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n1070), .B1(new_n1071), .B2(new_n696), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1049), .A2(new_n1072), .ZN(G390));
  INV_X1    g0873(.A(new_n1003), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n887), .A2(new_n890), .B1(new_n880), .B2(new_n888), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1075), .ZN(new_n1076));
  NAND4_X1  g0876(.A1(new_n680), .A2(new_n879), .A3(G330), .A4(new_n772), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n776), .B(new_n639), .C1(new_n682), .C2(new_n683), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1078), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n879), .B1(new_n1079), .B2(new_n876), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n868), .A2(new_n888), .A3(new_n1080), .ZN(new_n1081));
  NAND3_X1  g0881(.A1(new_n1076), .A2(new_n1077), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1077), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1081), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1083), .B1(new_n1084), .B2(new_n1075), .ZN(new_n1085));
  AND2_X1   g0885(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n441), .A2(G330), .A3(new_n680), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n619), .B(new_n1087), .C1(new_n896), .C2(new_n897), .ZN(new_n1088));
  NOR3_X1   g0888(.A1(new_n1083), .A2(new_n876), .A3(new_n1079), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n879), .ZN(new_n1090));
  OAI21_X1  g0890(.A(new_n1090), .B1(new_n681), .B2(new_n773), .ZN(new_n1091));
  OAI21_X1  g0891(.A(new_n1090), .B1(new_n681), .B2(new_n853), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1077), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1089), .A2(new_n1091), .B1(new_n1093), .B2(new_n878), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g0895(.A(new_n1074), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n1096), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n887), .A2(new_n890), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1098), .A2(new_n708), .ZN(new_n1099));
  NAND3_X1  g0899(.A1(new_n253), .A2(new_n709), .A3(new_n781), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n697), .A2(new_n1100), .ZN(new_n1101));
  AOI21_X1  g0901(.A(new_n1053), .B1(G283), .B2(new_n727), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1102), .B1(new_n224), .B2(new_n784), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n738), .A2(new_n646), .ZN(new_n1104));
  OAI221_X1 g0904(.A(new_n279), .B1(new_n745), .B2(new_n521), .C1(new_n539), .C2(new_n742), .ZN(new_n1105));
  OAI22_X1  g0905(.A1(new_n216), .A2(new_n716), .B1(new_n723), .B2(new_n218), .ZN(new_n1106));
  OR4_X1    g0906(.A1(new_n1103), .A2(new_n1104), .A3(new_n1105), .A4(new_n1106), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n723), .A2(new_n255), .ZN(new_n1108));
  XNOR2_X1  g0908(.A(KEYINPUT118), .B(KEYINPUT53), .ZN(new_n1109));
  XNOR2_X1  g0909(.A(new_n1108), .B(new_n1109), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  XNOR2_X1  g0911(.A(KEYINPUT54), .B(G143), .ZN(new_n1112));
  OAI221_X1 g0912(.A(new_n312), .B1(new_n745), .B2(new_n1111), .C1(new_n742), .C2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(new_n1113), .B1(new_n739), .B2(G132), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n990), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n732), .A2(new_n1115), .B1(new_n790), .B2(G50), .ZN(new_n1116));
  AOI22_X1  g0916(.A1(new_n727), .A2(G128), .B1(new_n721), .B2(G159), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1107), .B1(new_n1110), .B2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1101), .B1(new_n1119), .B2(new_n711), .ZN(new_n1120));
  AOI22_X1  g0920(.A1(new_n1086), .A2(new_n696), .B1(new_n1099), .B2(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1097), .A2(new_n1121), .ZN(G378));
  NAND2_X1  g0922(.A1(new_n271), .A2(new_n822), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n308), .B(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n708), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n697), .B1(new_n782), .B2(G50), .ZN(new_n1128));
  NOR2_X1   g0928(.A1(new_n385), .A2(G41), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(G33), .A2(G41), .ZN(new_n1130));
  NOR3_X1   g0930(.A1(new_n1129), .A2(G50), .A3(new_n1130), .ZN(new_n1131));
  OAI22_X1  g0931(.A1(new_n784), .A2(new_n539), .B1(new_n251), .B2(new_n716), .ZN(new_n1132));
  AOI211_X1 g0932(.A(new_n1022), .B(new_n1132), .C1(G116), .C2(new_n727), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n739), .A2(G107), .ZN(new_n1134));
  OAI22_X1  g0934(.A1(new_n742), .A2(new_n359), .B1(new_n745), .B2(new_n717), .ZN(new_n1135));
  AOI21_X1  g0935(.A(new_n1135), .B1(G68), .B2(new_n721), .ZN(new_n1136));
  NAND4_X1  g0936(.A1(new_n1133), .A2(new_n1129), .A3(new_n1134), .A4(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT58), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1131), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT119), .ZN(new_n1140));
  INV_X1    g0940(.A(G124), .ZN(new_n1141));
  OAI221_X1 g0941(.A(new_n1130), .B1(new_n745), .B2(new_n1141), .C1(new_n716), .C2(new_n751), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n793), .A2(G137), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n1143), .B1(new_n784), .B2(new_n799), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1144), .B1(new_n739), .B2(G128), .ZN(new_n1145));
  INV_X1    g0945(.A(new_n1112), .ZN(new_n1146));
  AOI22_X1  g0946(.A1(new_n802), .A2(new_n1146), .B1(new_n721), .B2(G150), .ZN(new_n1147));
  OAI211_X1 g0947(.A(new_n1145), .B(new_n1147), .C1(new_n1111), .C2(new_n755), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n1142), .B1(new_n1148), .B2(KEYINPUT59), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(KEYINPUT59), .B2(new_n1148), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1140), .B(new_n1150), .C1(new_n1138), .C2(new_n1137), .ZN(new_n1151));
  INV_X1    g0951(.A(KEYINPUT120), .ZN(new_n1152));
  OR2_X1    g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n781), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1154));
  AOI21_X1  g0954(.A(new_n1128), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1127), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  INV_X1    g0957(.A(KEYINPUT121), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n868), .A2(new_n869), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1159), .A2(G330), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1126), .B1(new_n859), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n621), .B1(new_n868), .B2(new_n869), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1126), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n857), .B1(new_n846), .B2(new_n851), .ZN(new_n1164));
  OAI211_X1 g0964(.A(new_n1162), .B(new_n1163), .C1(new_n1164), .C2(KEYINPUT40), .ZN(new_n1165));
  AND3_X1   g0965(.A1(new_n1161), .A2(new_n893), .A3(new_n1165), .ZN(new_n1166));
  AOI21_X1  g0966(.A(new_n893), .B1(new_n1161), .B2(new_n1165), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1158), .B1(new_n1166), .B2(new_n1167), .ZN(new_n1168));
  INV_X1    g0968(.A(new_n893), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n858), .B1(new_n882), .B2(new_n883), .ZN(new_n1170));
  INV_X1    g0970(.A(KEYINPUT40), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1163), .B1(new_n1172), .B2(new_n1162), .ZN(new_n1173));
  INV_X1    g0973(.A(new_n1165), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1169), .B1(new_n1173), .B2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g0975(.A1(new_n1161), .A2(new_n893), .A3(new_n1165), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n1175), .A2(KEYINPUT121), .A3(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1168), .A2(new_n1177), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1157), .B1(new_n1178), .B2(new_n696), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n1088), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1082), .A2(new_n1085), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n1180), .B1(new_n1181), .B2(new_n1094), .ZN(new_n1182));
  AOI21_X1  g0982(.A(KEYINPUT57), .B1(new_n1178), .B2(new_n1182), .ZN(new_n1183));
  NAND2_X1  g0983(.A1(new_n1182), .A2(KEYINPUT57), .ZN(new_n1184));
  NOR2_X1   g0984(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1185));
  OAI21_X1  g0985(.A(new_n1003), .B1(new_n1184), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1179), .B1(new_n1183), .B2(new_n1186), .ZN(G375));
  OR2_X1    g0987(.A1(new_n1094), .A2(new_n695), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n697), .B1(new_n782), .B2(G68), .ZN(new_n1189));
  OAI22_X1  g0989(.A1(new_n722), .A2(new_n323), .B1(new_n723), .B2(new_n397), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1190), .B1(G132), .B2(new_n727), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n739), .A2(new_n1115), .ZN(new_n1192));
  NOR2_X1   g0992(.A1(new_n742), .A2(new_n255), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n377), .B(new_n1193), .C1(G128), .C2(new_n746), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n732), .A2(new_n1146), .B1(new_n790), .B2(new_n395), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1191), .A2(new_n1192), .A3(new_n1194), .A4(new_n1195), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1023), .B1(G294), .B2(new_n727), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n802), .A2(G97), .ZN(new_n1198));
  AOI211_X1 g0998(.A(new_n312), .B(new_n994), .C1(G303), .C2(new_n746), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n739), .A2(G283), .ZN(new_n1200));
  NAND4_X1  g1000(.A1(new_n1197), .A2(new_n1198), .A3(new_n1199), .A4(new_n1200), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(new_n732), .A2(G116), .B1(new_n793), .B2(G107), .ZN(new_n1202));
  XOR2_X1   g1002(.A(new_n1202), .B(KEYINPUT123), .Z(new_n1203));
  OAI21_X1  g1003(.A(new_n1196), .B1(new_n1201), .B2(new_n1203), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n1189), .B1(new_n1204), .B2(new_n711), .ZN(new_n1205));
  OAI21_X1  g1005(.A(new_n1205), .B1(new_n879), .B2(new_n709), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1188), .A2(new_n1206), .ZN(new_n1207));
  INV_X1    g1007(.A(new_n1207), .ZN(new_n1208));
  AND2_X1   g1008(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1209), .A2(KEYINPUT122), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1088), .A2(new_n1094), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT122), .ZN(new_n1212));
  NAND2_X1  g1012(.A1(new_n1211), .A2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1210), .A2(new_n1213), .ZN(new_n1214));
  OR2_X1    g1014(.A1(new_n1095), .A2(new_n940), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1208), .B1(new_n1214), .B2(new_n1215), .ZN(G381));
  INV_X1    g1016(.A(G396), .ZN(new_n1217));
  NAND3_X1  g1017(.A1(new_n1004), .A2(new_n1217), .A3(new_n1043), .ZN(new_n1218));
  OR4_X1    g1018(.A1(G384), .A2(G387), .A3(G390), .A4(new_n1218), .ZN(new_n1219));
  OR4_X1    g1019(.A1(G378), .A2(G375), .A3(G381), .A4(new_n1219), .ZN(G407));
  INV_X1    g1020(.A(G378), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n627), .A2(G213), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1221), .A2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(G407), .B(G213), .C1(G375), .C2(new_n1224), .ZN(G409));
  INV_X1    g1025(.A(KEYINPUT127), .ZN(new_n1226));
  AND3_X1   g1026(.A1(new_n1004), .A2(new_n1217), .A3(new_n1043), .ZN(new_n1227));
  AOI21_X1  g1027(.A(new_n1217), .B1(new_n1004), .B2(new_n1043), .ZN(new_n1228));
  OAI21_X1  g1028(.A(KEYINPUT124), .B1(new_n1227), .B2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(G393), .A2(G396), .ZN(new_n1230));
  INV_X1    g1030(.A(KEYINPUT124), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1230), .A2(new_n1231), .A3(new_n1218), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1233));
  NAND3_X1  g1033(.A1(new_n975), .A2(G390), .A3(new_n999), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(G390), .B1(new_n975), .B2(new_n999), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1233), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  INV_X1    g1037(.A(G390), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(G387), .A2(new_n1238), .ZN(new_n1239));
  AND2_X1   g1039(.A1(new_n1229), .A2(new_n1232), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(new_n1234), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1237), .A2(new_n1241), .ZN(new_n1242));
  XOR2_X1   g1042(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1243));
  OAI211_X1 g1043(.A(G378), .B(new_n1179), .C1(new_n1183), .C2(new_n1186), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1088), .B1(new_n1086), .B2(new_n1095), .ZN(new_n1245));
  AOI211_X1 g1045(.A(new_n940), .B(new_n1245), .C1(new_n1168), .C2(new_n1177), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1156), .B1(new_n1185), .B2(new_n695), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1221), .B1(new_n1246), .B2(new_n1247), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n1223), .B1(new_n1244), .B2(new_n1248), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT60), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1210), .A2(new_n1250), .A3(new_n1213), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1074), .B1(new_n1209), .B2(KEYINPUT60), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1251), .A2(new_n1252), .ZN(new_n1253));
  AOI21_X1  g1053(.A(G384), .B1(new_n1253), .B2(new_n1208), .ZN(new_n1254));
  AOI211_X1 g1054(.A(new_n809), .B(new_n1207), .C1(new_n1251), .C2(new_n1252), .ZN(new_n1255));
  OAI211_X1 g1055(.A(G2897), .B(new_n1223), .C1(new_n1254), .C2(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1253), .A2(new_n1208), .ZN(new_n1257));
  NAND2_X1  g1057(.A1(new_n1257), .A2(new_n809), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1253), .A2(G384), .A3(new_n1208), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1223), .A2(G2897), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1258), .A2(new_n1259), .A3(new_n1260), .ZN(new_n1261));
  NAND2_X1  g1061(.A1(new_n1256), .A2(new_n1261), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1243), .B1(new_n1249), .B2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(KEYINPUT62), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1254), .A2(new_n1255), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1264), .B1(new_n1249), .B2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1263), .A2(new_n1266), .ZN(new_n1267));
  NAND3_X1  g1067(.A1(new_n1249), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1268));
  AOI21_X1  g1068(.A(new_n1242), .B1(new_n1267), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT125), .ZN(new_n1270));
  INV_X1    g1070(.A(KEYINPUT61), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1270), .B1(new_n1242), .B2(new_n1271), .ZN(new_n1272));
  AOI211_X1 g1072(.A(KEYINPUT125), .B(KEYINPUT61), .C1(new_n1237), .C2(new_n1241), .ZN(new_n1273));
  NOR2_X1   g1073(.A1(new_n1272), .A2(new_n1273), .ZN(new_n1274));
  OAI21_X1  g1074(.A(new_n1274), .B1(new_n1249), .B2(new_n1262), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(new_n1249), .A2(KEYINPUT63), .A3(new_n1265), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1276), .ZN(new_n1277));
  AOI21_X1  g1077(.A(KEYINPUT63), .B1(new_n1249), .B2(new_n1265), .ZN(new_n1278));
  NOR3_X1   g1078(.A1(new_n1275), .A2(new_n1277), .A3(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1226), .B1(new_n1269), .B2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1278), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1249), .A2(new_n1262), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1281), .A2(new_n1282), .A3(new_n1276), .A4(new_n1274), .ZN(new_n1283));
  INV_X1    g1083(.A(new_n1268), .ZN(new_n1284));
  NOR3_X1   g1084(.A1(new_n1284), .A2(new_n1263), .A3(new_n1266), .ZN(new_n1285));
  OAI211_X1 g1085(.A(KEYINPUT127), .B(new_n1283), .C1(new_n1285), .C2(new_n1242), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1280), .A2(new_n1286), .ZN(G405));
  NAND2_X1  g1087(.A1(G375), .A2(new_n1221), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(new_n1244), .ZN(new_n1289));
  XNOR2_X1  g1089(.A(new_n1289), .B(new_n1265), .ZN(new_n1290));
  XOR2_X1   g1090(.A(new_n1290), .B(new_n1242), .Z(G402));
endmodule


