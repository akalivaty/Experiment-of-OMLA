//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 0 0 0 1 1 0 1 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 1 1 1 1 1 0 1 0 0 1 1 0 0 1 1 1 0 1 1 0 0 0 1 0 0 0 0 1 1 0 0 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:10 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n796, new_n798, new_n799, new_n800, new_n801,
    new_n802, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n825, new_n826, new_n827, new_n828, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n883,
    new_n885, new_n886, new_n888, new_n889, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n895, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n965, new_n966, new_n967,
    new_n969, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n985,
    new_n986, new_n987, new_n988, new_n989, new_n990, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1010, new_n1011, new_n1012;
  INV_X1    g000(.A(KEYINPUT18), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT15), .ZN(new_n203));
  XNOR2_X1  g002(.A(G43gat), .B(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT89), .ZN(new_n205));
  AOI21_X1  g004(.A(new_n203), .B1(new_n204), .B2(new_n205), .ZN(new_n206));
  OR2_X1    g005(.A1(G43gat), .A2(G50gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  NAND3_X1  g007(.A1(new_n207), .A2(KEYINPUT89), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n206), .A2(new_n209), .ZN(new_n210));
  INV_X1    g009(.A(KEYINPUT90), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n211), .B1(new_n204), .B2(KEYINPUT15), .ZN(new_n212));
  INV_X1    g011(.A(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n214), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  XNOR2_X1  g015(.A(KEYINPUT14), .B(G29gat), .ZN(new_n217));
  INV_X1    g016(.A(G36gat), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI21_X1  g018(.A(new_n210), .B1(new_n213), .B2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT17), .ZN(new_n221));
  NOR2_X1   g020(.A1(new_n204), .A2(KEYINPUT15), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n206), .A2(new_n209), .B1(new_n222), .B2(KEYINPUT90), .ZN(new_n223));
  OAI211_X1 g022(.A(new_n220), .B(new_n221), .C1(new_n219), .C2(new_n223), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n222), .A2(KEYINPUT90), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n219), .B1(new_n210), .B2(new_n225), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n217), .A2(new_n218), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(new_n215), .ZN(new_n228));
  AOI22_X1  g027(.A1(new_n228), .A2(new_n212), .B1(new_n206), .B2(new_n209), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT17), .B1(new_n226), .B2(new_n229), .ZN(new_n230));
  XNOR2_X1  g029(.A(G15gat), .B(G22gat), .ZN(new_n231));
  OR2_X1    g030(.A1(new_n231), .A2(G1gat), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT16), .ZN(new_n233));
  OAI21_X1  g032(.A(new_n231), .B1(new_n233), .B2(G1gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT91), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G8gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n232), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(G8gat), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(new_n238), .ZN(new_n240));
  NAND4_X1  g039(.A1(new_n232), .A2(new_n234), .A3(new_n240), .A4(new_n236), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n239), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n224), .A2(new_n230), .A3(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(G229gat), .A2(G233gat), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n239), .A2(new_n241), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n226), .A2(new_n229), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n243), .A2(new_n244), .A3(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n245), .B(new_n246), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n244), .B(KEYINPUT13), .Z(new_n250));
  AOI22_X1  g049(.A1(new_n202), .A2(new_n248), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n243), .A2(KEYINPUT18), .A3(new_n247), .A4(new_n244), .ZN(new_n252));
  AND2_X1   g051(.A1(new_n252), .A2(KEYINPUT92), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n252), .A2(KEYINPUT92), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n251), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  XNOR2_X1  g054(.A(G113gat), .B(G141gat), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G197gat), .ZN(new_n257));
  XOR2_X1   g056(.A(KEYINPUT11), .B(G169gat), .Z(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  XNOR2_X1  g058(.A(new_n259), .B(KEYINPUT12), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n261), .ZN(new_n262));
  OAI211_X1 g061(.A(new_n251), .B(new_n260), .C1(new_n253), .C2(new_n254), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(G134gat), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n266), .A2(G127gat), .ZN(new_n267));
  INV_X1    g066(.A(G127gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(G134gat), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  XNOR2_X1  g069(.A(G113gat), .B(G120gat), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n270), .B1(new_n271), .B2(KEYINPUT1), .ZN(new_n272));
  INV_X1    g071(.A(G120gat), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(G113gat), .ZN(new_n274));
  INV_X1    g073(.A(G113gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n275), .A2(G120gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n274), .A2(new_n276), .ZN(new_n277));
  XNOR2_X1  g076(.A(G127gat), .B(G134gat), .ZN(new_n278));
  INV_X1    g077(.A(KEYINPUT1), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  AND2_X1   g079(.A1(new_n272), .A2(new_n280), .ZN(new_n281));
  OR2_X1    g080(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n282));
  NAND2_X1  g081(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(G148gat), .A3(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G148gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G141gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(G155gat), .A2(G162gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(G155gat), .A2(G162gat), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT2), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n288), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n284), .A2(new_n286), .B1(new_n287), .B2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G155gat), .B(G162gat), .ZN(new_n292));
  INV_X1    g091(.A(G141gat), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(G148gat), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n286), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(KEYINPUT76), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT76), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT2), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n296), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n292), .B1(new_n295), .B2(new_n299), .ZN(new_n300));
  NOR2_X1   g099(.A1(new_n291), .A2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(KEYINPUT3), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n281), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  OAI21_X1  g102(.A(KEYINPUT78), .B1(new_n291), .B2(new_n300), .ZN(new_n304));
  INV_X1    g103(.A(new_n287), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n305), .A2(new_n288), .ZN(new_n306));
  XNOR2_X1  g105(.A(G141gat), .B(G148gat), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT76), .B(KEYINPUT2), .ZN(new_n308));
  OAI21_X1  g107(.A(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT78), .ZN(new_n310));
  INV_X1    g109(.A(new_n286), .ZN(new_n311));
  AND2_X1   g110(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(KEYINPUT77), .A2(G141gat), .ZN(new_n313));
  NOR2_X1   g112(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n311), .B1(new_n314), .B2(G148gat), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n305), .B1(new_n289), .B2(new_n288), .ZN(new_n316));
  OAI211_X1 g115(.A(new_n309), .B(new_n310), .C1(new_n315), .C2(new_n316), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n304), .A2(new_n317), .A3(KEYINPUT3), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n303), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT79), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n303), .A2(new_n318), .A3(KEYINPUT79), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT5), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT4), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n309), .B1(new_n315), .B2(new_n316), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n272), .A2(new_n280), .ZN(new_n327));
  OAI21_X1  g126(.A(new_n325), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n301), .A2(new_n281), .A3(KEYINPUT4), .ZN(new_n329));
  NAND2_X1  g128(.A1(G225gat), .A2(G233gat), .ZN(new_n330));
  AND3_X1   g129(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n323), .A2(new_n324), .A3(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT80), .ZN(new_n333));
  AND3_X1   g132(.A1(new_n303), .A2(new_n318), .A3(KEYINPUT79), .ZN(new_n334));
  AOI21_X1  g133(.A(KEYINPUT79), .B1(new_n303), .B2(new_n318), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n331), .C1(new_n334), .C2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT81), .ZN(new_n337));
  NAND3_X1  g136(.A1(new_n304), .A2(new_n317), .A3(new_n327), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n301), .A2(new_n281), .ZN(new_n339));
  AOI21_X1  g138(.A(new_n330), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n337), .B1(new_n340), .B2(new_n324), .ZN(new_n341));
  AND2_X1   g140(.A1(new_n338), .A2(new_n339), .ZN(new_n342));
  OAI211_X1 g141(.A(KEYINPUT81), .B(KEYINPUT5), .C1(new_n342), .C2(new_n330), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n336), .A2(new_n341), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(new_n333), .B1(new_n323), .B2(new_n331), .ZN(new_n345));
  OAI21_X1  g144(.A(new_n332), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  XOR2_X1   g145(.A(G1gat), .B(G29gat), .Z(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G85gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT6), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n331), .B1(new_n334), .B2(new_n335), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT80), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n355), .A2(new_n336), .A3(new_n341), .A4(new_n343), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n356), .A2(new_n351), .A3(new_n332), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n353), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n351), .B1(new_n356), .B2(new_n332), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT83), .B1(new_n359), .B2(KEYINPUT6), .ZN(new_n360));
  AND4_X1   g159(.A1(KEYINPUT83), .A2(new_n346), .A3(KEYINPUT6), .A4(new_n352), .ZN(new_n361));
  OAI21_X1  g160(.A(new_n358), .B1(new_n360), .B2(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(G211gat), .A2(G218gat), .ZN(new_n363));
  INV_X1    g162(.A(G211gat), .ZN(new_n364));
  INV_X1    g163(.A(G218gat), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g165(.A1(G197gat), .A2(G204gat), .ZN(new_n367));
  NOR2_X1   g166(.A1(G197gat), .A2(G204gat), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT22), .ZN(new_n370));
  OAI211_X1 g169(.A(new_n363), .B(new_n366), .C1(new_n369), .C2(new_n370), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n366), .A2(new_n363), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n363), .A2(new_n370), .ZN(new_n373));
  OAI211_X1 g172(.A(new_n372), .B(new_n373), .C1(new_n368), .C2(new_n367), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n377));
  NAND2_X1  g176(.A1(G183gat), .A2(G190gat), .ZN(new_n378));
  NAND2_X1  g177(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  NAND3_X1  g178(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT23), .ZN(new_n382));
  OAI21_X1  g181(.A(new_n382), .B1(G169gat), .B2(G176gat), .ZN(new_n383));
  NAND2_X1  g182(.A1(G169gat), .A2(G176gat), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n383), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G169gat), .ZN(new_n386));
  INV_X1    g185(.A(G176gat), .ZN(new_n387));
  NAND3_X1  g186(.A1(new_n386), .A2(new_n387), .A3(KEYINPUT23), .ZN(new_n388));
  NAND3_X1  g187(.A1(new_n381), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT25), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT64), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n378), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393));
  NAND3_X1  g192(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n393), .A3(new_n394), .ZN(new_n395));
  OR2_X1    g194(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n396));
  INV_X1    g195(.A(G183gat), .ZN(new_n397));
  NAND2_X1  g196(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n396), .A2(new_n397), .A3(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n395), .A2(new_n399), .A3(new_n380), .ZN(new_n400));
  AND4_X1   g199(.A1(KEYINPUT25), .A2(new_n388), .A3(new_n383), .A4(new_n384), .ZN(new_n401));
  AOI22_X1  g200(.A1(new_n389), .A2(new_n390), .B1(new_n400), .B2(new_n401), .ZN(new_n402));
  NOR2_X1   g201(.A1(G169gat), .A2(G176gat), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n403), .A2(KEYINPUT26), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT26), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n384), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n404), .B(new_n378), .C1(new_n406), .C2(new_n403), .ZN(new_n407));
  AND2_X1   g206(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n408));
  NOR2_X1   g207(.A1(KEYINPUT65), .A2(G190gat), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n408), .A2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(KEYINPUT27), .B(G183gat), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT28), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT28), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n407), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(KEYINPUT71), .B1(new_n402), .B2(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT29), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n400), .A2(new_n401), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n393), .A2(new_n397), .ZN(new_n420));
  AOI22_X1  g219(.A1(new_n420), .A2(G190gat), .B1(new_n377), .B2(new_n378), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n388), .A2(new_n383), .A3(new_n384), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n390), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n419), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  INV_X1    g224(.A(new_n407), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n410), .A2(new_n411), .A3(KEYINPUT28), .ZN(new_n427));
  AOI21_X1  g226(.A(KEYINPUT28), .B1(new_n410), .B2(new_n411), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n424), .A2(new_n425), .A3(new_n429), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n417), .A2(new_n418), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(G226gat), .A2(G233gat), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n431), .A2(KEYINPUT72), .A3(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n424), .A2(new_n429), .ZN(new_n435));
  INV_X1    g234(.A(new_n432), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AOI22_X1  g236(.A1(new_n431), .A2(new_n432), .B1(KEYINPUT72), .B2(new_n437), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n376), .B1(new_n434), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n417), .A2(new_n430), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n440), .A2(new_n436), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n435), .A2(new_n418), .A3(new_n432), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n376), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  XOR2_X1   g243(.A(G8gat), .B(G36gat), .Z(new_n445));
  XNOR2_X1  g244(.A(new_n445), .B(KEYINPUT73), .ZN(new_n446));
  XNOR2_X1  g245(.A(G64gat), .B(G92gat), .ZN(new_n447));
  XNOR2_X1  g246(.A(new_n446), .B(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n439), .A2(new_n444), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(KEYINPUT30), .ZN(new_n450));
  AND3_X1   g249(.A1(new_n449), .A2(KEYINPUT75), .A3(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n450), .B1(new_n449), .B2(KEYINPUT75), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n448), .B(KEYINPUT74), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n431), .A2(new_n432), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n437), .A2(KEYINPUT72), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n375), .B1(new_n456), .B2(new_n433), .ZN(new_n457));
  OAI21_X1  g256(.A(new_n453), .B1(new_n457), .B2(new_n443), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR3_X1   g258(.A1(new_n451), .A2(new_n452), .A3(new_n459), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n418), .B1(new_n326), .B2(KEYINPUT3), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(new_n376), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT29), .B1(new_n371), .B2(new_n374), .ZN(new_n463));
  OAI211_X1 g262(.A(new_n304), .B(new_n317), .C1(new_n463), .C2(KEYINPUT3), .ZN(new_n464));
  AND4_X1   g263(.A1(G228gat), .A2(new_n462), .A3(G233gat), .A4(new_n464), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n302), .B1(new_n463), .B2(KEYINPUT85), .ZN(new_n466));
  AND3_X1   g265(.A1(new_n375), .A2(KEYINPUT85), .A3(new_n418), .ZN(new_n467));
  OAI21_X1  g266(.A(new_n326), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT86), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  OAI211_X1 g269(.A(KEYINPUT86), .B(new_n326), .C1(new_n466), .C2(new_n467), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n470), .A2(new_n471), .A3(new_n462), .ZN(new_n472));
  NAND2_X1  g271(.A1(G228gat), .A2(G233gat), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n465), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(G22gat), .ZN(new_n475));
  AOI21_X1  g274(.A(KEYINPUT87), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n477));
  INV_X1    g276(.A(G50gat), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n477), .B(new_n478), .ZN(new_n479));
  XOR2_X1   g278(.A(G78gat), .B(G106gat), .Z(new_n480));
  XOR2_X1   g279(.A(new_n479), .B(new_n480), .Z(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n474), .A2(new_n475), .ZN(new_n483));
  AOI211_X1 g282(.A(G22gat), .B(new_n465), .C1(new_n472), .C2(new_n473), .ZN(new_n484));
  OAI22_X1  g283(.A1(new_n476), .A2(new_n482), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n472), .A2(new_n473), .ZN(new_n486));
  OAI21_X1  g285(.A(G22gat), .B1(new_n486), .B2(new_n465), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n474), .A2(new_n475), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n487), .A2(new_n488), .A3(KEYINPUT87), .A4(new_n481), .ZN(new_n489));
  AND2_X1   g288(.A1(new_n485), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n281), .B1(new_n424), .B2(new_n429), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT66), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n424), .A2(new_n281), .A3(new_n429), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n491), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n424), .A2(KEYINPUT66), .A3(new_n281), .A4(new_n429), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  XOR2_X1   g296(.A(new_n497), .B(KEYINPUT34), .Z(new_n498));
  INV_X1    g297(.A(KEYINPUT67), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n495), .B1(new_n494), .B2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT32), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n493), .A2(new_n492), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n435), .A2(new_n327), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n503), .A2(new_n496), .A3(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(new_n495), .ZN(new_n506));
  AOI21_X1  g305(.A(new_n501), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n507), .A2(KEYINPUT67), .ZN(new_n508));
  XOR2_X1   g307(.A(G15gat), .B(G43gat), .Z(new_n509));
  XNOR2_X1  g308(.A(new_n509), .B(KEYINPUT68), .ZN(new_n510));
  XOR2_X1   g309(.A(G71gat), .B(G99gat), .Z(new_n511));
  XNOR2_X1  g310(.A(new_n510), .B(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n505), .A2(new_n506), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT33), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n502), .A2(new_n508), .A3(new_n515), .ZN(new_n516));
  OR2_X1    g315(.A1(new_n512), .A2(new_n514), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n507), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(KEYINPUT69), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT69), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n507), .A2(new_n520), .A3(new_n517), .ZN(new_n521));
  AND4_X1   g320(.A1(new_n498), .A2(new_n516), .A3(new_n519), .A4(new_n521), .ZN(new_n522));
  AND3_X1   g321(.A1(new_n507), .A2(new_n520), .A3(new_n517), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n520), .B1(new_n507), .B2(new_n517), .ZN(new_n524));
  NOR2_X1   g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n498), .B1(new_n525), .B2(new_n516), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n522), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n362), .A2(new_n460), .A3(new_n490), .A4(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n528), .A2(KEYINPUT35), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n485), .A2(new_n489), .ZN(new_n530));
  NOR3_X1   g329(.A1(new_n530), .A2(new_n526), .A3(new_n522), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT35), .ZN(new_n532));
  NAND4_X1  g331(.A1(new_n531), .A2(new_n532), .A3(new_n362), .A4(new_n460), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n529), .A2(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n448), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n457), .A2(new_n443), .A3(new_n535), .ZN(new_n536));
  NAND3_X1  g335(.A1(new_n456), .A2(new_n375), .A3(new_n433), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n537), .A2(KEYINPUT88), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT88), .ZN(new_n539));
  NAND4_X1  g338(.A1(new_n456), .A2(new_n539), .A3(new_n375), .A4(new_n433), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n441), .A2(new_n376), .A3(new_n442), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n538), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(new_n542), .A2(KEYINPUT37), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n439), .A2(new_n444), .A3(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(new_n453), .ZN(new_n546));
  NOR2_X1   g345(.A1(new_n546), .A2(KEYINPUT38), .ZN(new_n547));
  AND2_X1   g346(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  AOI21_X1  g347(.A(new_n536), .B1(new_n543), .B2(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n346), .A2(KEYINPUT6), .A3(new_n352), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT83), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n359), .A2(KEYINPUT83), .A3(KEYINPUT6), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n545), .A2(new_n535), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n544), .B1(new_n439), .B2(new_n444), .ZN(new_n556));
  OAI21_X1  g355(.A(KEYINPUT38), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n549), .A2(new_n554), .A3(new_n358), .A4(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT75), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT30), .B1(new_n536), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n449), .A2(KEYINPUT75), .A3(new_n450), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n561), .A3(new_n458), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n342), .A2(new_n330), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT39), .ZN(new_n564));
  OAI211_X1 g363(.A(new_n328), .B(new_n329), .C1(new_n334), .C2(new_n335), .ZN(new_n565));
  INV_X1    g364(.A(new_n330), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n564), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(KEYINPUT39), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n565), .A2(new_n569), .A3(new_n566), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n568), .A2(KEYINPUT40), .A3(new_n351), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n346), .A2(new_n352), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT40), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n570), .A2(new_n351), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n567), .ZN(new_n575));
  AND3_X1   g374(.A1(new_n571), .A2(new_n572), .A3(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n530), .B1(new_n562), .B2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n558), .A2(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n552), .A2(new_n553), .B1(new_n357), .B2(new_n353), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n530), .B1(new_n579), .B2(new_n562), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT70), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT36), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n584));
  OAI211_X1 g383(.A(new_n583), .B(new_n584), .C1(new_n522), .C2(new_n526), .ZN(new_n585));
  INV_X1    g384(.A(new_n498), .ZN(new_n586));
  INV_X1    g385(.A(new_n516), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n519), .A2(new_n521), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n587), .B2(new_n588), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n525), .A2(new_n498), .A3(new_n516), .ZN(new_n590));
  NAND4_X1  g389(.A1(new_n589), .A2(new_n581), .A3(new_n582), .A4(new_n590), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n585), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n578), .A2(new_n580), .A3(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n265), .B1(new_n534), .B2(new_n593), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(G71gat), .A2(G78gat), .ZN(new_n596));
  INV_X1    g395(.A(KEYINPUT93), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(G71gat), .ZN(new_n599));
  INV_X1    g398(.A(G78gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n599), .A2(new_n600), .A3(KEYINPUT94), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT94), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n602), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g403(.A(KEYINPUT95), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n596), .B(KEYINPUT93), .ZN(new_n606));
  INV_X1    g405(.A(KEYINPUT95), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n606), .A2(new_n607), .A3(new_n603), .A4(new_n601), .ZN(new_n608));
  INV_X1    g407(.A(G57gat), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n609), .A2(G64gat), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NOR2_X1   g410(.A1(new_n609), .A2(G64gat), .ZN(new_n612));
  INV_X1    g411(.A(new_n596), .ZN(new_n613));
  OAI22_X1  g412(.A1(new_n611), .A2(new_n612), .B1(new_n613), .B2(KEYINPUT9), .ZN(new_n614));
  NAND3_X1  g413(.A1(new_n605), .A2(new_n608), .A3(new_n614), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n612), .B1(KEYINPUT96), .B2(new_n610), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n616), .B1(KEYINPUT96), .B2(new_n610), .ZN(new_n617));
  INV_X1    g416(.A(KEYINPUT9), .ZN(new_n618));
  NOR3_X1   g417(.A1(new_n618), .A2(G71gat), .A3(G78gat), .ZN(new_n619));
  OAI21_X1  g418(.A(new_n617), .B1(new_n613), .B2(new_n619), .ZN(new_n620));
  AND2_X1   g419(.A1(new_n615), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n595), .B1(new_n621), .B2(KEYINPUT21), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n615), .A2(new_n620), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT21), .ZN(new_n624));
  INV_X1    g423(.A(new_n595), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  AND2_X1   g425(.A1(new_n622), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT98), .ZN(new_n629));
  AND3_X1   g428(.A1(new_n628), .A2(new_n629), .A3(new_n242), .ZN(new_n630));
  AOI21_X1  g429(.A(new_n629), .B1(new_n628), .B2(new_n242), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n627), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n628), .A2(new_n242), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(KEYINPUT98), .ZN(new_n634));
  NAND2_X1  g433(.A1(new_n622), .A2(new_n626), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n628), .A2(new_n629), .A3(new_n242), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n634), .A2(new_n635), .A3(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(G231gat), .A2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(KEYINPUT97), .ZN(new_n639));
  XOR2_X1   g438(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g440(.A(G183gat), .B(G211gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(new_n643));
  AND3_X1   g442(.A1(new_n632), .A2(new_n637), .A3(new_n643), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n643), .B1(new_n632), .B2(new_n637), .ZN(new_n645));
  NOR2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(KEYINPUT101), .ZN(new_n647));
  XNOR2_X1  g446(.A(G190gat), .B(G218gat), .ZN(new_n648));
  NAND2_X1  g447(.A1(G85gat), .A2(G92gat), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT7), .ZN(new_n650));
  XNOR2_X1  g449(.A(G99gat), .B(G106gat), .ZN(new_n651));
  NAND2_X1  g450(.A1(G99gat), .A2(G106gat), .ZN(new_n652));
  INV_X1    g451(.A(G85gat), .ZN(new_n653));
  INV_X1    g452(.A(G92gat), .ZN(new_n654));
  AOI22_X1  g453(.A1(KEYINPUT8), .A2(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  AND3_X1   g454(.A1(new_n650), .A2(new_n651), .A3(new_n655), .ZN(new_n656));
  AOI21_X1  g455(.A(new_n651), .B1(new_n650), .B2(new_n655), .ZN(new_n657));
  NOR2_X1   g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n224), .A2(new_n230), .A3(new_n659), .ZN(new_n660));
  AND2_X1   g459(.A1(G232gat), .A2(G233gat), .ZN(new_n661));
  AOI22_X1  g460(.A1(new_n246), .A2(new_n658), .B1(KEYINPUT41), .B2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT99), .ZN(new_n663));
  NAND3_X1  g462(.A1(new_n660), .A2(new_n662), .A3(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n663), .B1(new_n660), .B2(new_n662), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n648), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  XOR2_X1   g466(.A(G134gat), .B(G162gat), .Z(new_n668));
  NOR2_X1   g467(.A1(new_n661), .A2(KEYINPUT41), .ZN(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT100), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n660), .A2(new_n662), .ZN(new_n673));
  NAND2_X1  g472(.A1(new_n673), .A2(KEYINPUT99), .ZN(new_n674));
  INV_X1    g473(.A(new_n648), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n664), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n667), .A2(new_n672), .A3(new_n676), .ZN(new_n677));
  INV_X1    g476(.A(new_n677), .ZN(new_n678));
  XNOR2_X1  g477(.A(new_n670), .B(KEYINPUT100), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  AOI21_X1  g479(.A(new_n680), .B1(new_n667), .B2(new_n676), .ZN(new_n681));
  OAI211_X1 g480(.A(new_n646), .B(new_n647), .C1(new_n678), .C2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NOR3_X1   g482(.A1(new_n665), .A2(new_n648), .A3(new_n666), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n675), .B1(new_n674), .B2(new_n664), .ZN(new_n685));
  NOR2_X1   g484(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n677), .B1(new_n686), .B2(new_n680), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n647), .B1(new_n687), .B2(new_n646), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n623), .A2(new_n659), .ZN(new_n690));
  INV_X1    g489(.A(KEYINPUT10), .ZN(new_n691));
  NAND3_X1  g490(.A1(new_n658), .A2(new_n615), .A3(new_n620), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n690), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n621), .A2(KEYINPUT10), .A3(new_n658), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(KEYINPUT102), .ZN(new_n696));
  NAND2_X1  g495(.A1(G230gat), .A2(G233gat), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT102), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n693), .A2(new_n698), .A3(new_n694), .ZN(new_n699));
  NAND3_X1  g498(.A1(new_n696), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n697), .B1(new_n690), .B2(new_n692), .ZN(new_n701));
  XOR2_X1   g500(.A(G120gat), .B(G148gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT103), .ZN(new_n703));
  XOR2_X1   g502(.A(G176gat), .B(G204gat), .Z(new_n704));
  XNOR2_X1  g503(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n701), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n700), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n697), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n693), .B2(new_n694), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n706), .B1(new_n710), .B2(new_n701), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n689), .A2(new_n713), .ZN(new_n714));
  INV_X1    g513(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n594), .A2(new_n715), .ZN(new_n716));
  OR2_X1    g515(.A1(new_n362), .A2(KEYINPUT104), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n362), .A2(KEYINPUT104), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g518(.A1(new_n716), .A2(new_n719), .ZN(new_n720));
  XOR2_X1   g519(.A(KEYINPUT105), .B(G1gat), .Z(new_n721));
  XNOR2_X1  g520(.A(new_n720), .B(new_n721), .ZN(G1324gat));
  NOR2_X1   g521(.A1(new_n716), .A2(new_n460), .ZN(new_n723));
  XOR2_X1   g522(.A(KEYINPUT16), .B(G8gat), .Z(new_n724));
  NAND2_X1  g523(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(G8gat), .ZN(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(new_n723), .ZN(new_n727));
  MUX2_X1   g526(.A(new_n725), .B(new_n727), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g527(.A1(new_n585), .A2(new_n591), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT106), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND3_X1  g530(.A1(new_n585), .A2(new_n591), .A3(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(G15gat), .B1(new_n716), .B2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n527), .ZN(new_n735));
  OR2_X1    g534(.A1(new_n735), .A2(G15gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n716), .B2(new_n736), .ZN(G1326gat));
  NOR2_X1   g536(.A1(new_n716), .A2(new_n490), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(KEYINPUT107), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT43), .B(G22gat), .ZN(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  NOR3_X1   g540(.A1(new_n687), .A2(new_n646), .A3(new_n712), .ZN(new_n742));
  XNOR2_X1  g541(.A(new_n742), .B(KEYINPUT108), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n594), .A2(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n719), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n745), .A2(new_n214), .A3(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT45), .ZN(new_n748));
  INV_X1    g547(.A(new_n646), .ZN(new_n749));
  NAND3_X1  g548(.A1(new_n749), .A2(new_n264), .A3(new_n713), .ZN(new_n750));
  XOR2_X1   g549(.A(new_n750), .B(KEYINPUT109), .Z(new_n751));
  INV_X1    g550(.A(KEYINPUT44), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n534), .A2(new_n593), .ZN(new_n753));
  INV_X1    g552(.A(new_n687), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n754), .A2(new_n752), .ZN(new_n756));
  AND3_X1   g555(.A1(new_n585), .A2(new_n591), .A3(KEYINPUT106), .ZN(new_n757));
  AOI21_X1  g556(.A(KEYINPUT106), .B1(new_n585), .B2(new_n591), .ZN(new_n758));
  OAI211_X1 g557(.A(new_n578), .B(new_n580), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n756), .B1(new_n759), .B2(new_n534), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n751), .B1(new_n755), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G29gat), .B1(new_n761), .B2(new_n719), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n748), .A2(new_n762), .ZN(G1328gat));
  NOR3_X1   g562(.A1(new_n744), .A2(G36gat), .A3(new_n460), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT46), .ZN(new_n765));
  OAI21_X1  g564(.A(G36gat), .B1(new_n761), .B2(new_n460), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(G1329gat));
  OAI21_X1  g566(.A(G43gat), .B1(new_n761), .B2(new_n733), .ZN(new_n768));
  INV_X1    g567(.A(G43gat), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n745), .A2(new_n769), .A3(new_n527), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  AOI21_X1  g570(.A(KEYINPUT47), .B1(new_n770), .B2(KEYINPUT110), .ZN(new_n772));
  XNOR2_X1  g571(.A(new_n771), .B(new_n772), .ZN(G1330gat));
  OAI21_X1  g572(.A(G50gat), .B1(new_n761), .B2(new_n490), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n530), .A2(new_n478), .ZN(new_n775));
  XNOR2_X1  g574(.A(new_n775), .B(KEYINPUT111), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n745), .A2(new_n776), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n774), .A2(new_n777), .ZN(new_n778));
  XNOR2_X1  g577(.A(KEYINPUT112), .B(KEYINPUT48), .ZN(new_n779));
  XNOR2_X1  g578(.A(new_n778), .B(new_n779), .ZN(G1331gat));
  NAND2_X1  g579(.A1(new_n759), .A2(new_n534), .ZN(new_n781));
  NOR4_X1   g580(.A1(new_n683), .A2(new_n688), .A3(new_n264), .A4(new_n713), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NOR2_X1   g582(.A1(new_n783), .A2(new_n719), .ZN(new_n784));
  XOR2_X1   g583(.A(KEYINPUT113), .B(G57gat), .Z(new_n785));
  XNOR2_X1  g584(.A(new_n784), .B(new_n785), .ZN(G1332gat));
  NOR2_X1   g585(.A1(new_n783), .A2(new_n460), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  OAI21_X1  g590(.A(G71gat), .B1(new_n783), .B2(new_n733), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n527), .A2(new_n599), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n792), .B1(new_n783), .B2(new_n793), .ZN(new_n794));
  XOR2_X1   g593(.A(new_n794), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g594(.A1(new_n783), .A2(new_n490), .ZN(new_n796));
  XNOR2_X1  g595(.A(new_n796), .B(new_n600), .ZN(G1335gat));
  NOR3_X1   g596(.A1(new_n264), .A2(new_n713), .A3(new_n646), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n755), .B2(new_n760), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT114), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  OAI211_X1 g600(.A(KEYINPUT114), .B(new_n798), .C1(new_n755), .C2(new_n760), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n801), .A2(new_n746), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(G85gat), .ZN(new_n804));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n362), .A2(new_n460), .ZN(new_n806));
  AOI22_X1  g605(.A1(new_n558), .A2(new_n577), .B1(new_n806), .B2(new_n530), .ZN(new_n807));
  AOI22_X1  g606(.A1(new_n733), .A2(new_n807), .B1(new_n529), .B2(new_n533), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n264), .A2(new_n646), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n754), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(new_n811));
  NAND4_X1  g610(.A1(new_n781), .A2(KEYINPUT51), .A3(new_n754), .A4(new_n809), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n713), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n653), .A3(new_n746), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n804), .A2(new_n814), .ZN(G1336gat));
  NAND3_X1  g614(.A1(new_n813), .A2(new_n654), .A3(new_n562), .ZN(new_n816));
  OAI21_X1  g615(.A(G92gat), .B1(new_n799), .B2(new_n460), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT52), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n816), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n811), .A2(new_n812), .ZN(new_n820));
  AND4_X1   g619(.A1(new_n654), .A2(new_n820), .A3(new_n562), .A4(new_n712), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n801), .A2(new_n562), .A3(new_n802), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(G92gat), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n819), .B1(new_n823), .B2(new_n818), .ZN(G1337gat));
  AOI21_X1  g623(.A(G99gat), .B1(new_n813), .B2(new_n527), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n801), .A2(new_n802), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n757), .A2(new_n758), .ZN(new_n827));
  AND2_X1   g626(.A1(new_n827), .A2(G99gat), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n826), .B2(new_n828), .ZN(G1338gat));
  NOR3_X1   g628(.A1(new_n490), .A2(G106gat), .A3(new_n713), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n820), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n801), .A2(new_n530), .A3(new_n802), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n831), .B1(new_n832), .B2(G106gat), .ZN(new_n833));
  INV_X1    g632(.A(KEYINPUT53), .ZN(new_n834));
  AOI21_X1  g633(.A(KEYINPUT53), .B1(new_n820), .B2(new_n830), .ZN(new_n835));
  OAI211_X1 g634(.A(new_n530), .B(new_n798), .C1(new_n755), .C2(new_n760), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n836), .A2(G106gat), .ZN(new_n837));
  AOI21_X1  g636(.A(KEYINPUT115), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n835), .A2(new_n837), .A3(KEYINPUT115), .ZN(new_n839));
  OAI22_X1  g638(.A1(new_n833), .A2(new_n834), .B1(new_n838), .B2(new_n839), .ZN(G1339gat));
  INV_X1    g639(.A(new_n531), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT116), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n693), .A2(new_n709), .A3(new_n694), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(KEYINPUT54), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n709), .B1(new_n695), .B2(KEYINPUT102), .ZN(new_n845));
  AOI21_X1  g644(.A(new_n844), .B1(new_n845), .B2(new_n699), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n695), .A2(new_n847), .A3(new_n697), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n848), .A2(KEYINPUT55), .A3(new_n706), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n842), .B1(new_n846), .B2(new_n849), .ZN(new_n850));
  INV_X1    g649(.A(new_n844), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n700), .A2(new_n851), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT55), .ZN(new_n853));
  AOI211_X1 g652(.A(new_n853), .B(new_n705), .C1(new_n710), .C2(new_n847), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n852), .A2(new_n854), .A3(KEYINPUT116), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n850), .A2(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n708), .ZN(new_n857));
  INV_X1    g656(.A(KEYINPUT117), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(new_n708), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n860), .B1(new_n850), .B2(new_n855), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n861), .A2(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n848), .A2(new_n706), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n853), .B1(new_n846), .B2(new_n863), .ZN(new_n864));
  NAND4_X1  g663(.A1(new_n859), .A2(new_n264), .A3(new_n862), .A4(new_n864), .ZN(new_n865));
  NOR2_X1   g664(.A1(new_n249), .A2(new_n250), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n244), .B1(new_n243), .B2(new_n247), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n259), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n712), .A2(new_n263), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n754), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n263), .A2(new_n868), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n687), .A2(new_n871), .ZN(new_n872));
  NAND4_X1  g671(.A1(new_n859), .A2(new_n862), .A3(new_n864), .A4(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n749), .B1(new_n870), .B2(new_n874), .ZN(new_n875));
  INV_X1    g674(.A(new_n688), .ZN(new_n876));
  NAND4_X1  g675(.A1(new_n876), .A2(new_n265), .A3(new_n682), .A4(new_n713), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n841), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n719), .A2(new_n562), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n880), .A2(new_n265), .ZN(new_n881));
  XNOR2_X1  g680(.A(new_n881), .B(new_n275), .ZN(G1340gat));
  NOR2_X1   g681(.A1(new_n880), .A2(new_n713), .ZN(new_n883));
  XNOR2_X1  g682(.A(new_n883), .B(new_n273), .ZN(G1341gat));
  NOR2_X1   g683(.A1(new_n880), .A2(new_n749), .ZN(new_n885));
  XOR2_X1   g684(.A(KEYINPUT118), .B(G127gat), .Z(new_n886));
  XNOR2_X1  g685(.A(new_n885), .B(new_n886), .ZN(G1342gat));
  NAND4_X1  g686(.A1(new_n878), .A2(new_n266), .A3(new_n754), .A4(new_n879), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT56), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT120), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n889), .B(new_n890), .ZN(new_n891));
  OR3_X1    g690(.A1(new_n888), .A2(KEYINPUT119), .A3(KEYINPUT56), .ZN(new_n892));
  OAI21_X1  g691(.A(KEYINPUT119), .B1(new_n888), .B2(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  OAI21_X1  g693(.A(G134gat), .B1(new_n880), .B2(new_n687), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n891), .A2(new_n894), .A3(new_n895), .ZN(G1343gat));
  NOR3_X1   g695(.A1(new_n827), .A2(new_n719), .A3(new_n562), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n875), .A2(new_n877), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n898), .B2(new_n530), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n490), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n864), .A2(KEYINPUT121), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT121), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n903), .B(new_n853), .C1(new_n846), .C2(new_n863), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n902), .A2(new_n264), .A3(new_n904), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n869), .B1(new_n905), .B2(new_n857), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n687), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n646), .B1(new_n907), .B2(new_n873), .ZN(new_n908));
  INV_X1    g707(.A(new_n877), .ZN(new_n909));
  OAI21_X1  g708(.A(new_n901), .B1(new_n908), .B2(new_n909), .ZN(new_n910));
  INV_X1    g709(.A(KEYINPUT122), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI211_X1 g711(.A(KEYINPUT122), .B(new_n901), .C1(new_n908), .C2(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  OAI211_X1 g713(.A(new_n264), .B(new_n897), .C1(new_n899), .C2(new_n914), .ZN(new_n915));
  INV_X1    g714(.A(new_n314), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n490), .B1(new_n875), .B2(new_n877), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n265), .A2(G141gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n918), .A2(new_n897), .A3(new_n919), .ZN(new_n920));
  OR2_X1    g719(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT58), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n920), .A2(KEYINPUT123), .ZN(new_n923));
  NAND3_X1  g722(.A1(new_n921), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n898), .A2(new_n530), .ZN(new_n925));
  INV_X1    g724(.A(new_n897), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g726(.A1(new_n915), .A2(new_n916), .B1(new_n927), .B2(new_n919), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n917), .A2(new_n924), .B1(new_n928), .B2(new_n922), .ZN(G1344gat));
  NAND4_X1  g728(.A1(new_n918), .A2(new_n285), .A3(new_n712), .A4(new_n897), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT59), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n897), .A2(new_n712), .ZN(new_n932));
  OAI21_X1  g731(.A(new_n864), .B1(new_n861), .B2(KEYINPUT117), .ZN(new_n933));
  AOI211_X1 g732(.A(new_n858), .B(new_n860), .C1(new_n850), .C2(new_n855), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n933), .A2(new_n265), .A3(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n869), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n687), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  AOI21_X1  g736(.A(new_n646), .B1(new_n937), .B2(new_n873), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n901), .B1(new_n938), .B2(new_n909), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n877), .A2(KEYINPUT124), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT124), .ZN(new_n941));
  NAND4_X1  g740(.A1(new_n689), .A2(new_n941), .A3(new_n265), .A4(new_n713), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n940), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g742(.A(new_n530), .B1(new_n943), .B2(new_n908), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n944), .A2(new_n900), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n932), .B1(new_n939), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g745(.A(new_n285), .B1(new_n946), .B2(KEYINPUT125), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT125), .ZN(new_n948));
  AOI22_X1  g747(.A1(new_n898), .A2(new_n901), .B1(new_n944), .B2(new_n900), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n932), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n931), .B1(new_n947), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g750(.A1(new_n931), .A2(G148gat), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n925), .A2(new_n900), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n912), .A2(new_n913), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n926), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n952), .B1(new_n955), .B2(new_n712), .ZN(new_n956));
  OAI21_X1  g755(.A(new_n930), .B1(new_n951), .B2(new_n956), .ZN(G1345gat));
  AOI21_X1  g756(.A(G155gat), .B1(new_n927), .B2(new_n646), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n646), .A2(G155gat), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n955), .B2(new_n959), .ZN(G1346gat));
  INV_X1    g759(.A(G162gat), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n961), .B1(new_n955), .B2(new_n754), .ZN(new_n962));
  NOR4_X1   g761(.A1(new_n925), .A2(G162gat), .A3(new_n687), .A4(new_n926), .ZN(new_n963));
  OR2_X1    g762(.A1(new_n962), .A2(new_n963), .ZN(G1347gat));
  NAND2_X1  g763(.A1(new_n719), .A2(new_n562), .ZN(new_n965));
  AOI211_X1 g764(.A(new_n841), .B(new_n965), .C1(new_n875), .C2(new_n877), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(new_n264), .ZN(new_n967));
  XNOR2_X1  g766(.A(new_n967), .B(G169gat), .ZN(G1348gat));
  NAND2_X1  g767(.A1(new_n966), .A2(new_n712), .ZN(new_n969));
  XNOR2_X1  g768(.A(new_n969), .B(G176gat), .ZN(G1349gat));
  INV_X1    g769(.A(KEYINPUT126), .ZN(new_n971));
  AOI21_X1  g770(.A(new_n411), .B1(new_n971), .B2(G183gat), .ZN(new_n972));
  AND3_X1   g771(.A1(new_n966), .A2(new_n646), .A3(new_n972), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n966), .A2(new_n646), .B1(KEYINPUT126), .B2(G183gat), .ZN(new_n974));
  INV_X1    g773(.A(KEYINPUT60), .ZN(new_n975));
  OR3_X1    g774(.A1(new_n973), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g775(.A(new_n975), .B1(new_n973), .B2(new_n974), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(G1350gat));
  AND3_X1   g777(.A1(new_n966), .A2(new_n410), .A3(new_n754), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n966), .A2(new_n754), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n980), .A2(G190gat), .ZN(new_n981));
  INV_X1    g780(.A(KEYINPUT61), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n979), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  OAI21_X1  g782(.A(new_n983), .B1(new_n982), .B2(new_n981), .ZN(G1351gat));
  NAND3_X1  g783(.A1(new_n733), .A2(new_n562), .A3(new_n719), .ZN(new_n985));
  AOI21_X1  g784(.A(new_n985), .B1(new_n939), .B2(new_n945), .ZN(new_n986));
  INV_X1    g785(.A(G197gat), .ZN(new_n987));
  NOR2_X1   g786(.A1(new_n265), .A2(new_n987), .ZN(new_n988));
  NOR3_X1   g787(.A1(new_n965), .A2(new_n490), .A3(new_n827), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n898), .A2(new_n264), .A3(new_n989), .ZN(new_n990));
  AOI22_X1  g789(.A1(new_n986), .A2(new_n988), .B1(new_n987), .B2(new_n990), .ZN(G1352gat));
  INV_X1    g790(.A(KEYINPUT127), .ZN(new_n992));
  INV_X1    g791(.A(G204gat), .ZN(new_n993));
  NAND4_X1  g792(.A1(new_n898), .A2(new_n993), .A3(new_n712), .A4(new_n989), .ZN(new_n994));
  XNOR2_X1  g793(.A(new_n994), .B(KEYINPUT62), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n993), .B1(new_n986), .B2(new_n712), .ZN(new_n996));
  OAI21_X1  g795(.A(new_n992), .B1(new_n995), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n986), .A2(new_n712), .ZN(new_n998));
  NAND2_X1  g797(.A1(new_n998), .A2(G204gat), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n1000));
  XNOR2_X1  g799(.A(new_n994), .B(new_n1000), .ZN(new_n1001));
  NAND3_X1  g800(.A1(new_n999), .A2(new_n1001), .A3(KEYINPUT127), .ZN(new_n1002));
  NAND2_X1  g801(.A1(new_n997), .A2(new_n1002), .ZN(G1353gat));
  NAND2_X1  g802(.A1(new_n986), .A2(new_n646), .ZN(new_n1004));
  AND3_X1   g803(.A1(new_n1004), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1005));
  AOI21_X1  g804(.A(KEYINPUT63), .B1(new_n1004), .B2(G211gat), .ZN(new_n1006));
  NAND2_X1  g805(.A1(new_n898), .A2(new_n989), .ZN(new_n1007));
  NAND2_X1  g806(.A1(new_n646), .A2(new_n364), .ZN(new_n1008));
  OAI22_X1  g807(.A1(new_n1005), .A2(new_n1006), .B1(new_n1007), .B2(new_n1008), .ZN(G1354gat));
  NAND2_X1  g808(.A1(new_n986), .A2(new_n754), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1010), .A2(G218gat), .ZN(new_n1011));
  NAND2_X1  g810(.A1(new_n754), .A2(new_n365), .ZN(new_n1012));
  OAI21_X1  g811(.A(new_n1011), .B1(new_n1007), .B2(new_n1012), .ZN(G1355gat));
endmodule


