//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 1 0 1 1 0 0 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:00 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n235, new_n236, new_n237,
    new_n238, new_n240, new_n241, new_n242, new_n243, new_n244, new_n245,
    new_n246, new_n248, new_n249, new_n250, new_n251, new_n252, new_n253,
    new_n254, new_n255, new_n256, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1168, new_n1169,
    new_n1170, new_n1171, new_n1172, new_n1173, new_n1174, new_n1175,
    new_n1176, new_n1177, new_n1178, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1191, new_n1192, new_n1193, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1251,
    new_n1252, new_n1253, new_n1254, new_n1255, new_n1256, new_n1257;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(G13), .ZN(new_n206));
  NAND2_X1  g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT64), .ZN(new_n208));
  OAI211_X1 g0008(.A(new_n208), .B(G250), .C1(G257), .C2(G264), .ZN(new_n209));
  XOR2_X1   g0009(.A(new_n209), .B(KEYINPUT0), .Z(new_n210));
  INV_X1    g0010(.A(new_n205), .ZN(new_n211));
  INV_X1    g0011(.A(G68), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  INV_X1    g0014(.A(G87), .ZN(new_n215));
  INV_X1    g0015(.A(G250), .ZN(new_n216));
  INV_X1    g0016(.A(G97), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  OAI22_X1  g0018(.A1(new_n215), .A2(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n214), .B(new_n219), .C1(G107), .C2(G264), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G50), .A2(G226), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G77), .A2(G244), .ZN(new_n222));
  NAND2_X1  g0022(.A1(G116), .A2(G270), .ZN(new_n223));
  NAND4_X1  g0023(.A1(new_n220), .A2(new_n221), .A3(new_n222), .A4(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G58), .ZN(new_n225));
  INV_X1    g0025(.A(G232), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n211), .B1(new_n224), .B2(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  INV_X1    g0030(.A(KEYINPUT65), .ZN(new_n231));
  NAND2_X1  g0031(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g0032(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n233));
  NAND2_X1  g0033(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  INV_X1    g0034(.A(new_n234), .ZN(new_n235));
  NOR2_X1   g0035(.A1(new_n235), .A2(new_n204), .ZN(new_n236));
  OAI21_X1  g0036(.A(G50), .B1(G58), .B2(G68), .ZN(new_n237));
  XOR2_X1   g0037(.A(new_n237), .B(KEYINPUT66), .Z(new_n238));
  AOI211_X1 g0038(.A(new_n210), .B(new_n229), .C1(new_n236), .C2(new_n238), .ZN(G361));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n240), .B(G264), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n241), .B(G270), .Z(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT2), .B(G226), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(new_n226), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G238), .B(G244), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(new_n242), .B(new_n246), .Z(G358));
  XOR2_X1   g0047(.A(G68), .B(G77), .Z(new_n248));
  XNOR2_X1  g0048(.A(new_n248), .B(KEYINPUT67), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G50), .B(G58), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(G87), .B(G97), .ZN(new_n252));
  INV_X1    g0052(.A(G107), .ZN(new_n253));
  XNOR2_X1  g0053(.A(new_n252), .B(new_n253), .ZN(new_n254));
  INV_X1    g0054(.A(G116), .ZN(new_n255));
  XNOR2_X1  g0055(.A(new_n254), .B(new_n255), .ZN(new_n256));
  XNOR2_X1  g0056(.A(new_n251), .B(new_n256), .ZN(G351));
  NAND3_X1  g0057(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n232), .A2(new_n233), .A3(new_n258), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  NOR2_X1   g0060(.A1(G58), .A2(G68), .ZN(new_n261));
  INV_X1    g0061(.A(G50), .ZN(new_n262));
  AOI21_X1  g0062(.A(new_n204), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(G20), .A2(G33), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n263), .B1(G150), .B2(new_n264), .ZN(new_n265));
  XOR2_X1   g0065(.A(KEYINPUT8), .B(G58), .Z(new_n266));
  NAND3_X1  g0066(.A1(new_n266), .A2(new_n204), .A3(G33), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n260), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AOI21_X1  g0068(.A(new_n259), .B1(new_n203), .B2(G20), .ZN(new_n269));
  AOI21_X1  g0069(.A(new_n268), .B1(G50), .B2(new_n269), .ZN(new_n270));
  NAND3_X1  g0070(.A1(new_n203), .A2(G13), .A3(G20), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  NAND2_X1  g0072(.A1(new_n272), .A2(new_n262), .ZN(new_n273));
  NAND2_X1  g0073(.A1(new_n270), .A2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(new_n274), .B(KEYINPUT9), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(G33), .ZN(new_n279));
  INV_X1    g0079(.A(G41), .ZN(new_n280));
  OAI211_X1 g0080(.A(G1), .B(G13), .C1(new_n279), .C2(new_n280), .ZN(new_n281));
  AND2_X1   g0081(.A1(new_n281), .A2(new_n276), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n278), .B1(new_n282), .B2(G226), .ZN(new_n283));
  AND2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(KEYINPUT3), .A2(G33), .ZN(new_n285));
  NOR2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  XNOR2_X1  g0086(.A(KEYINPUT68), .B(G1698), .ZN(new_n287));
  AOI21_X1  g0087(.A(new_n286), .B1(G222), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(G223), .ZN(new_n289));
  INV_X1    g0089(.A(G1698), .ZN(new_n290));
  OAI21_X1  g0090(.A(new_n288), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OR2_X1    g0091(.A1(KEYINPUT3), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(KEYINPUT3), .A2(G33), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n291), .B1(G77), .B2(new_n294), .ZN(new_n295));
  AOI22_X1  g0095(.A1(new_n232), .A2(new_n233), .B1(G33), .B2(G41), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n283), .B1(new_n295), .B2(new_n297), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n275), .B(new_n299), .C1(new_n300), .C2(new_n298), .ZN(new_n301));
  OAI21_X1  g0101(.A(new_n301), .B1(KEYINPUT71), .B2(KEYINPUT10), .ZN(new_n302));
  NAND2_X1  g0102(.A1(KEYINPUT71), .A2(KEYINPUT10), .ZN(new_n303));
  XNOR2_X1  g0103(.A(new_n302), .B(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n298), .A2(G179), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(new_n298), .ZN(new_n307));
  AND2_X1   g0107(.A1(new_n307), .A2(new_n274), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n304), .A2(new_n309), .ZN(new_n310));
  XOR2_X1   g0110(.A(KEYINPUT15), .B(G87), .Z(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  NOR3_X1   g0112(.A1(new_n312), .A2(G20), .A3(new_n279), .ZN(new_n313));
  INV_X1    g0113(.A(new_n266), .ZN(new_n314));
  INV_X1    g0114(.A(new_n264), .ZN(new_n315));
  INV_X1    g0115(.A(G77), .ZN(new_n316));
  OAI22_X1  g0116(.A1(new_n314), .A2(new_n315), .B1(new_n204), .B2(new_n316), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n259), .B1(new_n313), .B2(new_n317), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n269), .A2(G77), .ZN(new_n319));
  OAI211_X1 g0119(.A(new_n318), .B(new_n319), .C1(G77), .C2(new_n271), .ZN(new_n320));
  XNOR2_X1  g0120(.A(new_n320), .B(KEYINPUT70), .ZN(new_n321));
  AND2_X1   g0121(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n322));
  NOR2_X1   g0122(.A1(KEYINPUT68), .A2(G1698), .ZN(new_n323));
  NOR2_X1   g0123(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI221_X1 g0124(.A(new_n294), .B1(new_n213), .B2(new_n290), .C1(new_n324), .C2(new_n226), .ZN(new_n325));
  XNOR2_X1  g0125(.A(KEYINPUT69), .B(G107), .ZN(new_n326));
  INV_X1    g0126(.A(new_n326), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n325), .B(new_n296), .C1(new_n294), .C2(new_n327), .ZN(new_n328));
  INV_X1    g0128(.A(new_n278), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n282), .A2(G244), .ZN(new_n330));
  NAND3_X1  g0130(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n331), .A2(new_n306), .ZN(new_n332));
  INV_X1    g0132(.A(new_n331), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n321), .A2(new_n332), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n310), .A2(new_n337), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n204), .A2(G33), .A3(G77), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n339), .B1(new_n204), .B2(G68), .ZN(new_n340));
  XNOR2_X1  g0140(.A(new_n340), .B(KEYINPUT74), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n315), .A2(new_n262), .ZN(new_n342));
  INV_X1    g0142(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n341), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n344), .A2(new_n259), .ZN(new_n345));
  XOR2_X1   g0145(.A(KEYINPUT75), .B(KEYINPUT11), .Z(new_n346));
  INV_X1    g0146(.A(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n344), .A2(new_n259), .A3(new_n346), .ZN(new_n349));
  NOR2_X1   g0149(.A1(new_n271), .A2(G68), .ZN(new_n350));
  XNOR2_X1  g0150(.A(new_n350), .B(KEYINPUT12), .ZN(new_n351));
  AOI21_X1  g0151(.A(new_n351), .B1(G68), .B2(new_n269), .ZN(new_n352));
  NAND3_X1  g0152(.A1(new_n348), .A2(new_n349), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT76), .ZN(new_n354));
  OR2_X1    g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n353), .A2(new_n354), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g0157(.A1(G33), .A2(G97), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n294), .A2(new_n287), .A3(G226), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n290), .B1(new_n292), .B2(new_n293), .ZN(new_n360));
  AOI21_X1  g0160(.A(KEYINPUT72), .B1(new_n360), .B2(G232), .ZN(new_n361));
  OAI211_X1 g0161(.A(G232), .B(G1698), .C1(new_n284), .C2(new_n285), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT72), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  OAI211_X1 g0164(.A(new_n358), .B(new_n359), .C1(new_n361), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n296), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n282), .A2(G238), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n366), .A2(new_n329), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT13), .ZN(new_n369));
  INV_X1    g0169(.A(KEYINPUT73), .ZN(new_n370));
  INV_X1    g0170(.A(KEYINPUT13), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n366), .A2(new_n371), .A3(new_n329), .A4(new_n367), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n369), .A2(new_n370), .A3(new_n372), .ZN(new_n373));
  OR3_X1    g0173(.A1(new_n368), .A2(new_n370), .A3(KEYINPUT13), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(G200), .ZN(new_n375));
  NAND3_X1  g0175(.A1(new_n369), .A2(G190), .A3(new_n372), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n357), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n377), .A2(KEYINPUT77), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT77), .ZN(new_n379));
  NAND4_X1  g0179(.A1(new_n357), .A2(new_n375), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND3_X1  g0181(.A1(new_n373), .A2(new_n374), .A3(G169), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(KEYINPUT14), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT14), .ZN(new_n384));
  NAND4_X1  g0184(.A1(new_n373), .A2(new_n374), .A3(new_n384), .A4(G169), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n369), .A2(G179), .A3(new_n372), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n383), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AND2_X1   g0187(.A1(new_n355), .A2(new_n356), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n381), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n292), .A2(new_n204), .A3(new_n293), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT7), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n292), .A2(KEYINPUT7), .A3(new_n204), .A4(new_n293), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n212), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NOR2_X1   g0196(.A1(new_n225), .A2(new_n212), .ZN(new_n397));
  OAI21_X1  g0197(.A(G20), .B1(new_n397), .B2(new_n261), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n264), .A2(G159), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n391), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g0201(.A(KEYINPUT7), .B1(new_n286), .B2(new_n204), .ZN(new_n402));
  NOR4_X1   g0202(.A1(new_n284), .A2(new_n285), .A3(new_n393), .A4(G20), .ZN(new_n403));
  OAI21_X1  g0203(.A(G68), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(new_n400), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(KEYINPUT16), .A3(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n401), .A2(new_n406), .A3(new_n259), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n266), .A2(new_n271), .ZN(new_n408));
  AOI21_X1  g0208(.A(new_n408), .B1(new_n269), .B2(new_n266), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G223), .B1(new_n322), .B2(new_n323), .ZN(new_n411));
  NAND2_X1  g0211(.A1(G226), .A2(G1698), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n286), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n279), .A2(new_n215), .ZN(new_n414));
  OAI21_X1  g0214(.A(new_n296), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  AOI21_X1  g0215(.A(new_n278), .B1(new_n282), .B2(G232), .ZN(new_n416));
  AOI21_X1  g0216(.A(G169), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n416), .ZN(new_n418));
  INV_X1    g0218(.A(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n417), .B1(new_n419), .B2(new_n334), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n410), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT18), .ZN(new_n422));
  XNOR2_X1  g0222(.A(new_n421), .B(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n418), .A2(G200), .ZN(new_n424));
  XNOR2_X1  g0224(.A(KEYINPUT78), .B(G190), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n415), .A2(new_n416), .A3(new_n425), .ZN(new_n426));
  NAND4_X1  g0226(.A1(new_n407), .A2(new_n424), .A3(new_n426), .A4(new_n409), .ZN(new_n427));
  XNOR2_X1  g0227(.A(new_n427), .B(KEYINPUT17), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n423), .A2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n321), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n331), .A2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n333), .A2(G190), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n433), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n390), .A2(new_n429), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g0235(.A1(new_n338), .A2(new_n435), .ZN(new_n436));
  INV_X1    g0236(.A(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n294), .A2(new_n287), .A3(G257), .ZN(new_n438));
  INV_X1    g0238(.A(KEYINPUT82), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  AOI22_X1  g0240(.A1(new_n360), .A2(G264), .B1(new_n286), .B2(G303), .ZN(new_n441));
  NAND4_X1  g0241(.A1(new_n294), .A2(new_n287), .A3(KEYINPUT82), .A4(G257), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(G45), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n444), .A2(G1), .ZN(new_n445));
  AND2_X1   g0245(.A1(KEYINPUT5), .A2(G41), .ZN(new_n446));
  NOR2_X1   g0246(.A1(KEYINPUT5), .A2(G41), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n445), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  AND2_X1   g0248(.A1(new_n448), .A2(new_n281), .ZN(new_n449));
  AOI22_X1  g0249(.A1(new_n443), .A2(new_n296), .B1(G270), .B2(new_n449), .ZN(new_n450));
  OR2_X1    g0250(.A1(new_n448), .A2(new_n277), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT85), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT84), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(KEYINPUT20), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n255), .A2(G20), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n259), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT83), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g0259(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  AOI21_X1  g0261(.A(G20), .B1(G33), .B2(G283), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n462), .B1(G33), .B2(new_n217), .ZN(new_n463));
  AOI21_X1  g0263(.A(new_n455), .B1(new_n461), .B2(new_n463), .ZN(new_n464));
  AND3_X1   g0264(.A1(new_n259), .A2(KEYINPUT83), .A3(new_n456), .ZN(new_n465));
  AOI21_X1  g0265(.A(KEYINPUT83), .B1(new_n259), .B2(new_n456), .ZN(new_n466));
  OAI211_X1 g0266(.A(new_n455), .B(new_n463), .C1(new_n465), .C2(new_n466), .ZN(new_n467));
  INV_X1    g0267(.A(new_n467), .ZN(new_n468));
  OAI22_X1  g0268(.A1(new_n464), .A2(new_n468), .B1(new_n454), .B2(KEYINPUT20), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n272), .A2(G116), .ZN(new_n470));
  NOR2_X1   g0270(.A1(new_n279), .A2(G1), .ZN(new_n471));
  OR3_X1    g0271(.A1(new_n259), .A2(new_n272), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n472), .B2(G116), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n453), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  NOR2_X1   g0275(.A1(new_n454), .A2(KEYINPUT20), .ZN(new_n476));
  OAI21_X1  g0276(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n477));
  INV_X1    g0277(.A(new_n455), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n476), .B1(new_n479), .B2(new_n467), .ZN(new_n480));
  NOR3_X1   g0280(.A1(new_n480), .A2(KEYINPUT85), .A3(new_n473), .ZN(new_n481));
  OAI211_X1 g0281(.A(G169), .B(new_n452), .C1(new_n475), .C2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT21), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n469), .A2(new_n453), .A3(new_n474), .ZN(new_n485));
  OAI21_X1  g0285(.A(KEYINPUT85), .B1(new_n480), .B2(new_n473), .ZN(new_n486));
  AOI21_X1  g0286(.A(new_n306), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n487), .A2(KEYINPUT21), .A3(new_n452), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n449), .A2(G264), .ZN(new_n489));
  OAI22_X1  g0289(.A1(new_n324), .A2(new_n216), .B1(new_n218), .B2(new_n290), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n490), .A2(new_n294), .B1(G33), .B2(G294), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n489), .B(new_n451), .C1(new_n491), .C2(new_n297), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(KEYINPUT88), .ZN(new_n493));
  AOI22_X1  g0293(.A1(new_n287), .A2(G250), .B1(G257), .B2(G1698), .ZN(new_n494));
  INV_X1    g0294(.A(G294), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n494), .A2(new_n286), .B1(new_n279), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n496), .A2(new_n296), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT88), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n497), .A2(new_n498), .A3(new_n489), .A4(new_n451), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n493), .A2(new_n499), .ZN(new_n500));
  OAI22_X1  g0300(.A1(new_n500), .A2(new_n306), .B1(new_n334), .B2(new_n492), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n294), .A2(new_n204), .A3(G87), .ZN(new_n502));
  XOR2_X1   g0302(.A(KEYINPUT86), .B(KEYINPUT22), .Z(new_n503));
  INV_X1    g0303(.A(new_n503), .ZN(new_n504));
  XNOR2_X1  g0304(.A(new_n502), .B(new_n504), .ZN(new_n505));
  OR3_X1    g0305(.A1(new_n204), .A2(KEYINPUT23), .A3(G107), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n507), .A2(G20), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n326), .A2(G20), .ZN(new_n509));
  XNOR2_X1  g0309(.A(KEYINPUT87), .B(KEYINPUT23), .ZN(new_n510));
  AOI21_X1  g0310(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NAND4_X1  g0311(.A1(new_n505), .A2(KEYINPUT24), .A3(new_n506), .A4(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  XNOR2_X1  g0313(.A(new_n502), .B(new_n503), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n511), .A2(new_n506), .ZN(new_n515));
  OAI21_X1  g0315(.A(new_n513), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n512), .A2(new_n516), .A3(new_n259), .ZN(new_n517));
  OR2_X1    g0317(.A1(new_n472), .A2(new_n253), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n271), .A2(G107), .ZN(new_n519));
  XNOR2_X1  g0319(.A(new_n519), .B(KEYINPUT25), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n517), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n501), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n485), .A2(new_n486), .ZN(new_n523));
  NOR2_X1   g0323(.A1(new_n452), .A2(new_n334), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n484), .A2(new_n488), .A3(new_n522), .A4(new_n525), .ZN(new_n526));
  NAND2_X1  g0326(.A1(G250), .A2(G1698), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT79), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n287), .B1(new_n528), .B2(KEYINPUT4), .ZN(new_n529));
  INV_X1    g0329(.A(G244), .ZN(new_n530));
  OAI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(new_n294), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n294), .A2(new_n287), .A3(G244), .ZN(new_n533));
  NOR2_X1   g0333(.A1(new_n528), .A2(KEYINPUT4), .ZN(new_n534));
  AOI22_X1  g0334(.A1(new_n533), .A2(new_n534), .B1(G33), .B2(G283), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n297), .B1(new_n532), .B2(new_n535), .ZN(new_n536));
  INV_X1    g0336(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n449), .A2(G257), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n537), .A2(new_n451), .A3(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(KEYINPUT80), .ZN(new_n540));
  NAND3_X1  g0340(.A1(new_n539), .A2(new_n540), .A3(G200), .ZN(new_n541));
  INV_X1    g0341(.A(new_n451), .ZN(new_n542));
  INV_X1    g0342(.A(new_n538), .ZN(new_n543));
  NOR3_X1   g0343(.A1(new_n536), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(G200), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT80), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT6), .ZN(new_n547));
  NOR3_X1   g0347(.A1(new_n547), .A2(new_n217), .A3(G107), .ZN(new_n548));
  XNOR2_X1  g0348(.A(G97), .B(G107), .ZN(new_n549));
  AOI21_X1  g0349(.A(new_n548), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  OAI22_X1  g0350(.A1(new_n550), .A2(new_n204), .B1(new_n316), .B2(new_n315), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n326), .B1(new_n394), .B2(new_n395), .ZN(new_n552));
  OAI21_X1  g0352(.A(new_n259), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n272), .A2(new_n217), .ZN(new_n554));
  OAI211_X1 g0354(.A(new_n553), .B(new_n554), .C1(new_n217), .C2(new_n472), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n555), .B1(new_n544), .B2(G190), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n541), .A2(new_n546), .A3(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n521), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n493), .A2(new_n300), .A3(new_n499), .ZN(new_n559));
  INV_X1    g0359(.A(new_n492), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n559), .B1(G200), .B2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n558), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g0362(.A1(new_n358), .A2(G20), .ZN(new_n563));
  NOR2_X1   g0363(.A1(new_n563), .A2(KEYINPUT19), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n286), .A2(G20), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n564), .B1(new_n565), .B2(G68), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n326), .A2(new_n215), .A3(new_n217), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n358), .A2(new_n204), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n567), .A2(KEYINPUT19), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n259), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n311), .A2(new_n271), .ZN(new_n572));
  INV_X1    g0372(.A(new_n572), .ZN(new_n573));
  OAI211_X1 g0373(.A(new_n571), .B(new_n573), .C1(new_n312), .C2(new_n472), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n445), .A2(new_n277), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n575), .B(new_n281), .C1(G250), .C2(new_n445), .ZN(new_n576));
  OAI22_X1  g0376(.A1(new_n324), .A2(new_n213), .B1(new_n530), .B2(new_n290), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n577), .A2(new_n294), .B1(G33), .B2(G116), .ZN(new_n578));
  OAI21_X1  g0378(.A(new_n576), .B1(new_n578), .B2(new_n297), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n579), .A2(new_n306), .ZN(new_n580));
  OAI211_X1 g0380(.A(new_n574), .B(new_n580), .C1(G179), .C2(new_n579), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT81), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n582), .B1(new_n579), .B2(new_n300), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n577), .A2(new_n294), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n507), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n296), .ZN(new_n586));
  NAND4_X1  g0386(.A1(new_n586), .A2(KEYINPUT81), .A3(G190), .A4(new_n576), .ZN(new_n587));
  NOR4_X1   g0387(.A1(new_n259), .A2(new_n272), .A3(new_n215), .A4(new_n471), .ZN(new_n588));
  AOI211_X1 g0388(.A(new_n572), .B(new_n588), .C1(new_n570), .C2(new_n259), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n579), .A2(G200), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n583), .A2(new_n587), .A3(new_n589), .A4(new_n590), .ZN(new_n591));
  AND2_X1   g0391(.A1(new_n581), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n544), .A2(new_n334), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n593), .B(new_n555), .C1(G169), .C2(new_n544), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n557), .A2(new_n562), .A3(new_n592), .A4(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(new_n452), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n596), .A2(new_n425), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n597), .B1(new_n545), .B2(new_n596), .ZN(new_n598));
  NOR2_X1   g0398(.A1(new_n598), .A2(new_n523), .ZN(new_n599));
  NOR4_X1   g0399(.A1(new_n437), .A2(new_n526), .A3(new_n595), .A4(new_n599), .ZN(G372));
  INV_X1    g0400(.A(new_n389), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n601), .B1(new_n377), .B2(new_n337), .ZN(new_n602));
  INV_X1    g0402(.A(new_n428), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n423), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n308), .B1(new_n604), .B2(new_n304), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n482), .A2(new_n483), .ZN(new_n606));
  AOI21_X1  g0406(.A(KEYINPUT21), .B1(new_n487), .B2(new_n452), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND4_X1  g0408(.A1(new_n608), .A2(KEYINPUT89), .A3(new_n522), .A4(new_n525), .ZN(new_n609));
  INV_X1    g0409(.A(new_n595), .ZN(new_n610));
  INV_X1    g0410(.A(KEYINPUT89), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n526), .A2(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n609), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n581), .A2(new_n591), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n594), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g0415(.A(new_n615), .B(KEYINPUT26), .ZN(new_n616));
  AND2_X1   g0416(.A1(new_n616), .A2(new_n581), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  INV_X1    g0418(.A(new_n618), .ZN(new_n619));
  OAI21_X1  g0419(.A(new_n605), .B1(new_n437), .B2(new_n619), .ZN(G369));
  NAND3_X1  g0420(.A1(new_n484), .A2(new_n525), .A3(new_n488), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n206), .A2(G20), .ZN(new_n622));
  INV_X1    g0422(.A(new_n622), .ZN(new_n623));
  OR3_X1    g0423(.A1(new_n623), .A2(KEYINPUT27), .A3(G1), .ZN(new_n624));
  OAI21_X1  g0424(.A(KEYINPUT27), .B1(new_n623), .B2(G1), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n624), .A2(G213), .A3(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(G343), .ZN(new_n627));
  NOR2_X1   g0427(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g0428(.A1(new_n621), .A2(new_n523), .A3(new_n628), .ZN(new_n629));
  INV_X1    g0429(.A(KEYINPUT90), .ZN(new_n630));
  NOR2_X1   g0430(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  AND3_X1   g0431(.A1(new_n484), .A2(new_n525), .A3(new_n488), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n523), .A2(new_n628), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  OAI21_X1  g0434(.A(KEYINPUT90), .B1(new_n634), .B2(new_n599), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n631), .B1(new_n635), .B2(new_n629), .ZN(new_n636));
  INV_X1    g0436(.A(G330), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n521), .B1(new_n501), .B2(new_n628), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n638), .A2(new_n562), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(KEYINPUT91), .ZN(new_n640));
  INV_X1    g0440(.A(KEYINPUT91), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n638), .B2(new_n562), .ZN(new_n642));
  INV_X1    g0442(.A(new_n628), .ZN(new_n643));
  OAI22_X1  g0443(.A1(new_n640), .A2(new_n642), .B1(new_n522), .B2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  NOR3_X1   g0445(.A1(new_n636), .A2(new_n637), .A3(new_n645), .ZN(new_n646));
  INV_X1    g0446(.A(KEYINPUT92), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n621), .A2(new_n647), .A3(new_n643), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  AOI21_X1  g0449(.A(new_n647), .B1(new_n621), .B2(new_n643), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n644), .B1(new_n649), .B2(new_n650), .ZN(new_n651));
  INV_X1    g0451(.A(new_n522), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n652), .A2(new_n643), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n646), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g0455(.A(new_n655), .B(KEYINPUT93), .ZN(G399));
  NAND2_X1  g0456(.A1(new_n208), .A2(new_n280), .ZN(new_n657));
  INV_X1    g0457(.A(new_n657), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n567), .A2(G116), .ZN(new_n659));
  NOR3_X1   g0459(.A1(new_n658), .A2(new_n203), .A3(new_n659), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n660), .B1(new_n238), .B2(new_n658), .ZN(new_n661));
  XNOR2_X1  g0461(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n662));
  XNOR2_X1  g0462(.A(new_n661), .B(new_n662), .ZN(new_n663));
  NAND2_X1  g0463(.A1(new_n526), .A2(new_n610), .ZN(new_n664));
  AOI21_X1  g0464(.A(new_n628), .B1(new_n617), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(KEYINPUT29), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n628), .B1(new_n613), .B2(new_n617), .ZN(new_n667));
  OAI21_X1  g0467(.A(new_n666), .B1(new_n667), .B2(KEYINPUT29), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n595), .A2(new_n599), .ZN(new_n669));
  NAND4_X1  g0469(.A1(new_n632), .A2(new_n669), .A3(new_n522), .A4(new_n643), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n536), .A2(new_n543), .ZN(new_n671));
  NOR2_X1   g0471(.A1(new_n492), .A2(new_n579), .ZN(new_n672));
  NAND3_X1  g0472(.A1(new_n524), .A2(new_n671), .A3(new_n672), .ZN(new_n673));
  INV_X1    g0473(.A(KEYINPUT30), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NOR2_X1   g0475(.A1(new_n596), .A2(G179), .ZN(new_n676));
  NAND4_X1  g0476(.A1(new_n676), .A2(new_n492), .A3(new_n539), .A4(new_n579), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n524), .A2(KEYINPUT30), .A3(new_n671), .A4(new_n672), .ZN(new_n678));
  NAND3_X1  g0478(.A1(new_n675), .A2(new_n677), .A3(new_n678), .ZN(new_n679));
  NAND2_X1  g0479(.A1(new_n679), .A2(new_n628), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n680), .A2(KEYINPUT31), .ZN(new_n681));
  INV_X1    g0481(.A(KEYINPUT31), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n679), .A2(new_n682), .A3(new_n628), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n681), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n670), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n685), .A2(G330), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n668), .A2(new_n686), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n663), .B1(new_n688), .B2(G1), .ZN(G364));
  AOI21_X1  g0489(.A(new_n203), .B1(new_n622), .B2(G45), .ZN(new_n690));
  INV_X1    g0490(.A(new_n690), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n658), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g0493(.A1(G13), .A2(G33), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NOR2_X1   g0495(.A1(new_n695), .A2(G20), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n693), .B1(new_n636), .B2(new_n696), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n235), .B1(G20), .B2(new_n306), .ZN(new_n698));
  NOR2_X1   g0498(.A1(new_n204), .A2(G190), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G179), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(new_n701), .ZN(new_n702));
  AND2_X1   g0502(.A1(new_n702), .A2(G329), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n204), .A2(new_n334), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n425), .A2(new_n704), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(G200), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n705), .A2(new_n545), .ZN(new_n707));
  AOI22_X1  g0507(.A1(G322), .A2(new_n706), .B1(new_n707), .B2(G326), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n204), .B1(new_n700), .B2(G190), .ZN(new_n709));
  INV_X1    g0509(.A(G311), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n704), .A2(new_n300), .A3(new_n545), .ZN(new_n711));
  OAI221_X1 g0511(.A(new_n708), .B1(new_n495), .B2(new_n709), .C1(new_n710), .C2(new_n711), .ZN(new_n712));
  INV_X1    g0512(.A(new_n699), .ZN(new_n713));
  NOR3_X1   g0513(.A1(new_n713), .A2(new_n334), .A3(new_n545), .ZN(new_n714));
  XNOR2_X1  g0514(.A(KEYINPUT33), .B(G317), .ZN(new_n715));
  AOI211_X1 g0515(.A(new_n703), .B(new_n712), .C1(new_n714), .C2(new_n715), .ZN(new_n716));
  INV_X1    g0516(.A(G283), .ZN(new_n717));
  NOR2_X1   g0517(.A1(new_n545), .A2(G179), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n699), .A2(new_n718), .ZN(new_n719));
  OAI211_X1 g0519(.A(new_n716), .B(new_n286), .C1(new_n717), .C2(new_n719), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n718), .A2(G20), .A3(G190), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  AOI21_X1  g0522(.A(new_n720), .B1(G303), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n709), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n725));
  NOR2_X1   g0525(.A1(new_n724), .A2(KEYINPUT96), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(new_n217), .ZN(new_n728));
  NAND2_X1  g0528(.A1(new_n702), .A2(G159), .ZN(new_n729));
  XNOR2_X1  g0529(.A(new_n729), .B(KEYINPUT32), .ZN(new_n730));
  INV_X1    g0530(.A(new_n706), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n731), .A2(new_n225), .ZN(new_n732));
  INV_X1    g0532(.A(new_n714), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n733), .A2(new_n212), .ZN(new_n734));
  NOR4_X1   g0534(.A1(new_n728), .A2(new_n730), .A3(new_n732), .A4(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n719), .ZN(new_n736));
  AOI22_X1  g0536(.A1(new_n722), .A2(G87), .B1(new_n736), .B2(G107), .ZN(new_n737));
  XOR2_X1   g0537(.A(new_n711), .B(KEYINPUT95), .Z(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  AOI21_X1  g0539(.A(new_n286), .B1(new_n739), .B2(G77), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n735), .A2(new_n737), .A3(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(G50), .B2(new_n707), .ZN(new_n742));
  OAI21_X1  g0542(.A(new_n698), .B1(new_n723), .B2(new_n742), .ZN(new_n743));
  AND2_X1   g0543(.A1(new_n697), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n698), .A2(new_n696), .ZN(new_n745));
  OR2_X1    g0545(.A1(new_n251), .A2(new_n444), .ZN(new_n746));
  INV_X1    g0546(.A(new_n238), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(new_n444), .ZN(new_n748));
  AOI21_X1  g0548(.A(new_n294), .B1(new_n746), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(G355), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n208), .B1(new_n750), .B2(new_n286), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n745), .B1(new_n255), .B2(new_n208), .C1(new_n749), .C2(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n636), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  INV_X1    g0554(.A(new_n754), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n692), .B1(new_n753), .B2(G330), .ZN(new_n756));
  AOI22_X1  g0556(.A1(new_n744), .A2(new_n752), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(G396));
  OAI21_X1  g0558(.A(new_n433), .B1(new_n430), .B2(new_n643), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n759), .A2(new_n336), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n336), .A2(new_n628), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n667), .A2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n628), .B(new_n763), .C1(new_n613), .C2(new_n617), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(new_n686), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n768), .A2(new_n693), .ZN(new_n769));
  AOI22_X1  g0569(.A1(new_n706), .A2(G294), .B1(G283), .B2(new_n714), .ZN(new_n770));
  OAI21_X1  g0570(.A(new_n770), .B1(new_n215), .B2(new_n719), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n286), .B1(new_n701), .B2(new_n710), .ZN(new_n772));
  INV_X1    g0572(.A(new_n707), .ZN(new_n773));
  INV_X1    g0573(.A(G303), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  NOR4_X1   g0575(.A1(new_n771), .A2(new_n728), .A3(new_n772), .A4(new_n775), .ZN(new_n776));
  OAI221_X1 g0576(.A(new_n776), .B1(new_n253), .B2(new_n721), .C1(new_n255), .C2(new_n738), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n706), .A2(G143), .B1(G150), .B2(new_n714), .ZN(new_n778));
  INV_X1    g0578(.A(G137), .ZN(new_n779));
  INV_X1    g0579(.A(G159), .ZN(new_n780));
  OAI221_X1 g0580(.A(new_n778), .B1(new_n779), .B2(new_n773), .C1(new_n738), .C2(new_n780), .ZN(new_n781));
  XOR2_X1   g0581(.A(new_n781), .B(KEYINPUT97), .Z(new_n782));
  XNOR2_X1  g0582(.A(new_n782), .B(KEYINPUT34), .ZN(new_n783));
  INV_X1    g0583(.A(G132), .ZN(new_n784));
  OAI211_X1 g0584(.A(new_n783), .B(new_n294), .C1(new_n784), .C2(new_n701), .ZN(new_n785));
  AOI22_X1  g0585(.A1(new_n722), .A2(G50), .B1(new_n736), .B2(G68), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n786), .B1(new_n225), .B2(new_n709), .ZN(new_n787));
  OAI21_X1  g0587(.A(new_n777), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n693), .B1(new_n788), .B2(new_n698), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n698), .A2(new_n694), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI221_X1 g0591(.A(new_n789), .B1(G77), .B2(new_n791), .C1(new_n695), .C2(new_n764), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n769), .A2(new_n792), .ZN(G384));
  AOI21_X1  g0593(.A(new_n763), .B1(new_n670), .B2(new_n684), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n388), .A2(new_n628), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n795), .A2(KEYINPUT99), .ZN(new_n796));
  OR3_X1    g0596(.A1(new_n357), .A2(KEYINPUT99), .A3(new_n643), .ZN(new_n797));
  NAND4_X1  g0597(.A1(new_n389), .A2(new_n377), .A3(new_n796), .A4(new_n797), .ZN(new_n798));
  AOI22_X1  g0598(.A1(new_n378), .A2(new_n380), .B1(new_n387), .B2(new_n388), .ZN(new_n799));
  OAI21_X1  g0599(.A(new_n798), .B1(new_n799), .B2(new_n795), .ZN(new_n800));
  AND2_X1   g0600(.A1(new_n794), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(KEYINPUT101), .ZN(new_n802));
  INV_X1    g0602(.A(KEYINPUT37), .ZN(new_n803));
  INV_X1    g0603(.A(new_n626), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n410), .A2(new_n804), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n805), .A2(KEYINPUT100), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n626), .B1(new_n407), .B2(new_n409), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT100), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n806), .A2(new_n809), .ZN(new_n810));
  AND2_X1   g0610(.A1(new_n421), .A2(new_n427), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n803), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g0612(.A1(new_n421), .A2(new_n427), .ZN(new_n813));
  NOR3_X1   g0613(.A1(new_n813), .A2(new_n807), .A3(KEYINPUT37), .ZN(new_n814));
  OAI21_X1  g0614(.A(new_n802), .B1(new_n812), .B2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n810), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n429), .A2(new_n816), .ZN(new_n817));
  NAND3_X1  g0617(.A1(new_n811), .A2(new_n803), .A3(new_n805), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n813), .B1(new_n806), .B2(new_n809), .ZN(new_n819));
  OAI211_X1 g0619(.A(new_n818), .B(KEYINPUT101), .C1(new_n819), .C2(new_n803), .ZN(new_n820));
  NAND4_X1  g0620(.A1(new_n815), .A2(KEYINPUT38), .A3(new_n817), .A4(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT38), .ZN(new_n822));
  AOI21_X1  g0622(.A(new_n803), .B1(new_n811), .B2(new_n805), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n823), .A2(new_n814), .ZN(new_n824));
  AOI21_X1  g0624(.A(new_n805), .B1(new_n423), .B2(new_n428), .ZN(new_n825));
  OAI21_X1  g0625(.A(new_n822), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n821), .A2(new_n826), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n801), .A2(KEYINPUT40), .A3(new_n827), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n829), .A2(new_n822), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n830), .A2(KEYINPUT102), .A3(new_n821), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT102), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n829), .A2(new_n832), .A3(new_n822), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n831), .A2(new_n794), .A3(new_n833), .A4(new_n800), .ZN(new_n834));
  INV_X1    g0634(.A(KEYINPUT106), .ZN(new_n835));
  INV_X1    g0635(.A(KEYINPUT40), .ZN(new_n836));
  AND3_X1   g0636(.A1(new_n834), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n835), .B1(new_n834), .B2(new_n836), .ZN(new_n838));
  OAI21_X1  g0638(.A(new_n828), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  XOR2_X1   g0639(.A(new_n839), .B(KEYINPUT107), .Z(new_n840));
  INV_X1    g0640(.A(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(new_n685), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n841), .B1(new_n437), .B2(new_n842), .ZN(new_n843));
  NAND3_X1  g0643(.A1(new_n840), .A2(new_n436), .A3(new_n685), .ZN(new_n844));
  NAND3_X1  g0644(.A1(new_n843), .A2(G330), .A3(new_n844), .ZN(new_n845));
  OAI211_X1 g0645(.A(new_n436), .B(new_n666), .C1(KEYINPUT29), .C2(new_n667), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n605), .ZN(new_n847));
  XOR2_X1   g0647(.A(new_n847), .B(KEYINPUT105), .Z(new_n848));
  XNOR2_X1  g0648(.A(new_n845), .B(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n821), .A2(KEYINPUT102), .ZN(new_n850));
  XNOR2_X1  g0650(.A(new_n850), .B(new_n830), .ZN(new_n851));
  OAI211_X1 g0651(.A(new_n851), .B(new_n800), .C1(new_n766), .C2(new_n761), .ZN(new_n852));
  INV_X1    g0652(.A(new_n423), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n853), .A2(new_n626), .ZN(new_n854));
  AND2_X1   g0654(.A1(new_n852), .A2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n601), .A2(new_n643), .ZN(new_n856));
  XNOR2_X1  g0656(.A(new_n856), .B(KEYINPUT103), .ZN(new_n857));
  NAND3_X1  g0657(.A1(new_n831), .A2(KEYINPUT39), .A3(new_n833), .ZN(new_n858));
  OAI21_X1  g0658(.A(KEYINPUT104), .B1(new_n827), .B2(KEYINPUT39), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n858), .A2(new_n859), .ZN(new_n860));
  NAND4_X1  g0660(.A1(new_n831), .A2(KEYINPUT104), .A3(KEYINPUT39), .A4(new_n833), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n857), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND2_X1  g0663(.A1(new_n855), .A2(new_n863), .ZN(new_n864));
  OR2_X1    g0664(.A1(new_n849), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n849), .A2(new_n864), .ZN(new_n866));
  OAI211_X1 g0666(.A(new_n865), .B(new_n866), .C1(new_n203), .C2(new_n622), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT35), .ZN(new_n868));
  AOI211_X1 g0668(.A(new_n204), .B(new_n235), .C1(new_n550), .C2(new_n868), .ZN(new_n869));
  OAI211_X1 g0669(.A(new_n869), .B(G116), .C1(new_n868), .C2(new_n550), .ZN(new_n870));
  XNOR2_X1  g0670(.A(new_n870), .B(KEYINPUT36), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n747), .A2(new_n316), .A3(new_n397), .ZN(new_n872));
  AOI21_X1  g0672(.A(new_n872), .B1(new_n262), .B2(G68), .ZN(new_n873));
  NOR3_X1   g0673(.A1(new_n873), .A2(new_n203), .A3(G13), .ZN(new_n874));
  XOR2_X1   g0674(.A(new_n874), .B(KEYINPUT98), .Z(new_n875));
  NAND3_X1  g0675(.A1(new_n867), .A2(new_n871), .A3(new_n875), .ZN(G367));
  NOR2_X1   g0676(.A1(new_n721), .A2(new_n255), .ZN(new_n877));
  XNOR2_X1  g0677(.A(new_n877), .B(KEYINPUT46), .ZN(new_n878));
  AOI22_X1  g0678(.A1(new_n739), .A2(G283), .B1(new_n327), .B2(new_n724), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  NOR2_X1   g0680(.A1(new_n880), .A2(KEYINPUT115), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n736), .A2(G97), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n882), .B1(new_n773), .B2(new_n710), .C1(new_n774), .C2(new_n731), .ZN(new_n883));
  INV_X1    g0683(.A(G317), .ZN(new_n884));
  OAI21_X1  g0684(.A(new_n286), .B1(new_n701), .B2(new_n884), .ZN(new_n885));
  NOR3_X1   g0685(.A1(new_n881), .A2(new_n883), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n886), .B1(new_n495), .B2(new_n733), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n878), .B(new_n887), .C1(KEYINPUT115), .C2(new_n880), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n706), .A2(G150), .B1(G58), .B2(new_n722), .ZN(new_n889));
  OAI21_X1  g0689(.A(new_n889), .B1(new_n779), .B2(new_n701), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n727), .A2(new_n212), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n719), .A2(new_n316), .ZN(new_n892));
  AND2_X1   g0692(.A1(new_n707), .A2(G143), .ZN(new_n893));
  NOR4_X1   g0693(.A1(new_n890), .A2(new_n891), .A3(new_n892), .A4(new_n893), .ZN(new_n894));
  OAI211_X1 g0694(.A(new_n894), .B(new_n294), .C1(new_n262), .C2(new_n738), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n895), .B1(G159), .B2(new_n714), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n888), .A2(new_n896), .ZN(new_n897));
  XOR2_X1   g0697(.A(new_n897), .B(KEYINPUT47), .Z(new_n898));
  NAND2_X1  g0698(.A1(new_n898), .A2(new_n698), .ZN(new_n899));
  OR2_X1    g0699(.A1(new_n589), .A2(new_n643), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n592), .A2(new_n900), .ZN(new_n901));
  OR2_X1    g0701(.A1(new_n581), .A2(new_n900), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n901), .A2(new_n696), .A3(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n208), .A2(new_n286), .ZN(new_n904));
  OAI221_X1 g0704(.A(new_n745), .B1(new_n208), .B2(new_n312), .C1(new_n242), .C2(new_n904), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n899), .A2(new_n692), .A3(new_n903), .A4(new_n905), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  OAI21_X1  g0707(.A(KEYINPUT92), .B1(new_n632), .B2(new_n628), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(new_n648), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g0710(.A(new_n645), .B1(new_n636), .B2(new_n637), .ZN(new_n911));
  INV_X1    g0711(.A(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n910), .B1(new_n912), .B2(new_n646), .ZN(new_n913));
  INV_X1    g0713(.A(new_n646), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n914), .A2(new_n909), .A3(new_n911), .ZN(new_n915));
  NAND3_X1  g0715(.A1(new_n688), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  XNOR2_X1  g0716(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n917));
  INV_X1    g0717(.A(new_n917), .ZN(new_n918));
  AND2_X1   g0718(.A1(new_n557), .A2(new_n594), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n555), .A2(new_n628), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  OR2_X1    g0721(.A1(new_n594), .A2(new_n643), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n918), .B1(new_n654), .B2(new_n924), .ZN(new_n925));
  AOI211_X1 g0725(.A(new_n923), .B(new_n917), .C1(new_n651), .C2(new_n653), .ZN(new_n926));
  NOR2_X1   g0726(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  AOI22_X1  g0727(.A1(new_n909), .A2(new_n644), .B1(new_n652), .B2(new_n643), .ZN(new_n928));
  XNOR2_X1  g0728(.A(KEYINPUT112), .B(KEYINPUT45), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n928), .A2(new_n923), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n651), .A2(new_n653), .A3(new_n923), .ZN(new_n931));
  INV_X1    g0731(.A(new_n929), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n646), .B1(new_n927), .B2(new_n934), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n930), .A2(new_n933), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n917), .B1(new_n928), .B2(new_n923), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n654), .A2(new_n924), .A3(new_n918), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND3_X1  g0739(.A1(new_n936), .A2(new_n914), .A3(new_n939), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n940), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n916), .B1(new_n941), .B2(KEYINPUT114), .ZN(new_n942));
  NOR2_X1   g0742(.A1(new_n646), .A2(KEYINPUT114), .ZN(new_n943));
  INV_X1    g0743(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n687), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  XOR2_X1   g0745(.A(new_n657), .B(KEYINPUT41), .Z(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n690), .B1(new_n945), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n914), .A2(new_n924), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n901), .A2(new_n902), .ZN(new_n950));
  AOI22_X1  g0750(.A1(new_n949), .A2(KEYINPUT111), .B1(KEYINPUT43), .B2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT110), .ZN(new_n952));
  OAI211_X1 g0752(.A(new_n644), .B(new_n923), .C1(new_n649), .C2(new_n650), .ZN(new_n953));
  OAI21_X1  g0753(.A(new_n952), .B1(new_n953), .B2(KEYINPUT42), .ZN(new_n954));
  OR3_X1    g0754(.A1(new_n953), .A2(new_n952), .A3(KEYINPUT42), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT109), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n953), .A2(KEYINPUT42), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n919), .A2(new_n652), .A3(new_n920), .ZN(new_n958));
  AOI21_X1  g0758(.A(new_n628), .B1(new_n958), .B2(new_n594), .ZN(new_n959));
  INV_X1    g0759(.A(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n956), .B1(new_n957), .B2(new_n960), .ZN(new_n961));
  AOI211_X1 g0761(.A(KEYINPUT109), .B(new_n959), .C1(new_n953), .C2(KEYINPUT42), .ZN(new_n962));
  OAI211_X1 g0762(.A(new_n954), .B(new_n955), .C1(new_n961), .C2(new_n962), .ZN(new_n963));
  INV_X1    g0763(.A(KEYINPUT108), .ZN(new_n964));
  OR2_X1    g0764(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n964), .A2(KEYINPUT43), .ZN(new_n966));
  AOI21_X1  g0766(.A(new_n950), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g0767(.A(new_n967), .ZN(new_n968));
  AND2_X1   g0768(.A1(new_n963), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g0769(.A1(new_n963), .A2(new_n968), .ZN(new_n970));
  OAI21_X1  g0770(.A(new_n951), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n949), .A2(KEYINPUT111), .ZN(new_n972));
  INV_X1    g0772(.A(new_n972), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n971), .A2(new_n973), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n972), .B(new_n951), .C1(new_n969), .C2(new_n970), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(new_n976), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n907), .B1(new_n948), .B2(new_n977), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(G387));
  NOR3_X1   g0779(.A1(new_n912), .A2(new_n646), .A3(new_n910), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n909), .B1(new_n914), .B2(new_n911), .ZN(new_n981));
  OAI21_X1  g0781(.A(new_n687), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g0782(.A1(new_n982), .A2(new_n658), .A3(new_n916), .ZN(new_n983));
  AOI21_X1  g0783(.A(new_n286), .B1(new_n702), .B2(G150), .ZN(new_n984));
  OAI211_X1 g0784(.A(new_n984), .B(new_n882), .C1(new_n316), .C2(new_n721), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT116), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n985), .A2(new_n986), .B1(new_n266), .B2(new_n714), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n727), .A2(new_n312), .ZN(new_n988));
  INV_X1    g0788(.A(new_n988), .ZN(new_n989));
  AOI22_X1  g0789(.A1(G50), .A2(new_n706), .B1(new_n707), .B2(G159), .ZN(new_n990));
  AND3_X1   g0790(.A1(new_n987), .A2(new_n989), .A3(new_n990), .ZN(new_n991));
  OAI221_X1 g0791(.A(new_n991), .B1(new_n986), .B2(new_n985), .C1(new_n212), .C2(new_n711), .ZN(new_n992));
  AOI22_X1  g0792(.A1(new_n706), .A2(G317), .B1(G311), .B2(new_n714), .ZN(new_n993));
  INV_X1    g0793(.A(G322), .ZN(new_n994));
  OAI221_X1 g0794(.A(new_n993), .B1(new_n994), .B2(new_n773), .C1(new_n738), .C2(new_n774), .ZN(new_n995));
  XNOR2_X1  g0795(.A(new_n995), .B(KEYINPUT48), .ZN(new_n996));
  OAI221_X1 g0796(.A(new_n996), .B1(new_n717), .B2(new_n709), .C1(new_n495), .C2(new_n721), .ZN(new_n997));
  INV_X1    g0797(.A(KEYINPUT49), .ZN(new_n998));
  OR2_X1    g0798(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n736), .A2(G116), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n702), .A2(G326), .ZN(new_n1001));
  NAND4_X1  g0801(.A1(new_n999), .A2(new_n286), .A3(new_n1000), .A4(new_n1001), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n997), .A2(new_n998), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n992), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n693), .B1(new_n1004), .B2(new_n698), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n696), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n1005), .B1(new_n644), .B2(new_n1006), .ZN(new_n1007));
  NOR2_X1   g0807(.A1(new_n208), .A2(new_n253), .ZN(new_n1008));
  NAND3_X1  g0808(.A1(new_n246), .A2(G45), .A3(new_n286), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n314), .A2(G50), .ZN(new_n1010));
  INV_X1    g0810(.A(new_n1010), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(new_n1011), .A2(KEYINPUT50), .B1(G68), .B2(G77), .ZN(new_n1012));
  INV_X1    g0812(.A(KEYINPUT50), .ZN(new_n1013));
  AOI21_X1  g0813(.A(G45), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n294), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1009), .B1(new_n1015), .B2(new_n659), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n1008), .B1(new_n1016), .B2(new_n208), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1007), .B1(new_n745), .B2(new_n1017), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n980), .A2(new_n981), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1018), .B1(new_n1019), .B2(new_n691), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n983), .A2(new_n1020), .ZN(G393));
  AND2_X1   g0821(.A1(new_n935), .A2(new_n940), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1022), .A2(new_n691), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n256), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n745), .B1(new_n217), .B2(new_n208), .C1(new_n1024), .C2(new_n904), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n1025), .A2(new_n692), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G311), .A2(new_n706), .B1(new_n707), .B2(G317), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT52), .ZN(new_n1028));
  NOR2_X1   g0828(.A1(new_n719), .A2(new_n253), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n286), .B1(new_n709), .B2(new_n255), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n733), .A2(new_n774), .B1(new_n701), .B2(new_n994), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1028), .A2(new_n1029), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  OAI221_X1 g0832(.A(new_n1032), .B1(new_n717), .B2(new_n721), .C1(new_n495), .C2(new_n711), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n721), .A2(new_n212), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n727), .A2(new_n316), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n286), .B(new_n1035), .C1(new_n266), .C2(new_n739), .ZN(new_n1036));
  AOI22_X1  g0836(.A1(G150), .A2(new_n707), .B1(new_n706), .B2(G159), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(KEYINPUT51), .ZN(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(G87), .B2(new_n736), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n702), .A2(G143), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n1037), .A2(KEYINPUT51), .B1(G50), .B2(new_n714), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1036), .A2(new_n1039), .A3(new_n1040), .A4(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1033), .B1(new_n1034), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1026), .B1(new_n1043), .B2(new_n698), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n1044), .B1(new_n923), .B2(new_n1006), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1023), .A2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g0846(.A1(new_n942), .A2(new_n944), .B1(new_n916), .B2(new_n941), .ZN(new_n1047));
  AOI21_X1  g0847(.A(new_n1046), .B1(new_n1047), .B2(new_n658), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1048), .ZN(G390));
  NAND3_X1  g0849(.A1(new_n860), .A2(new_n694), .A3(new_n861), .ZN(new_n1050));
  OAI22_X1  g0850(.A1(new_n738), .A2(new_n217), .B1(new_n326), .B2(new_n733), .ZN(new_n1051));
  XOR2_X1   g0851(.A(new_n1051), .B(KEYINPUT120), .Z(new_n1052));
  AOI21_X1  g0852(.A(new_n1035), .B1(G116), .B2(new_n706), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1053), .B1(new_n495), .B2(new_n701), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n773), .A2(new_n717), .ZN(new_n1055));
  OAI221_X1 g0855(.A(new_n286), .B1(new_n719), .B2(new_n212), .C1(new_n215), .C2(new_n721), .ZN(new_n1056));
  NOR4_X1   g0856(.A1(new_n1052), .A2(new_n1054), .A3(new_n1055), .A4(new_n1056), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n727), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1058), .A2(G159), .B1(G125), .B2(new_n702), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n722), .A2(G150), .ZN(new_n1060));
  XOR2_X1   g0860(.A(new_n1060), .B(KEYINPUT53), .Z(new_n1061));
  NAND2_X1  g0861(.A1(new_n714), .A2(G137), .ZN(new_n1062));
  NAND4_X1  g0862(.A1(new_n1059), .A2(new_n1061), .A3(new_n294), .A4(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n731), .A2(new_n784), .ZN(new_n1064));
  INV_X1    g0864(.A(G128), .ZN(new_n1065));
  NOR2_X1   g0865(.A1(new_n773), .A2(new_n1065), .ZN(new_n1066));
  XOR2_X1   g0866(.A(KEYINPUT54), .B(G143), .Z(new_n1067));
  INV_X1    g0867(.A(new_n1067), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n738), .A2(new_n1068), .B1(new_n262), .B2(new_n719), .ZN(new_n1069));
  NOR4_X1   g0869(.A1(new_n1063), .A2(new_n1064), .A3(new_n1066), .A4(new_n1069), .ZN(new_n1070));
  OAI21_X1  g0870(.A(new_n698), .B1(new_n1057), .B2(new_n1070), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n692), .B1(new_n266), .B2(new_n791), .ZN(new_n1072));
  XNOR2_X1  g0872(.A(new_n1072), .B(KEYINPUT119), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n1050), .A2(new_n1071), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g0874(.A(new_n1074), .ZN(new_n1075));
  AOI21_X1  g0875(.A(new_n761), .B1(new_n665), .B2(new_n760), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n800), .ZN(new_n1077));
  OAI211_X1 g0877(.A(new_n857), .B(new_n827), .C1(new_n1076), .C2(new_n1077), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n857), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n618), .A2(new_n643), .A3(new_n764), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1080), .A2(new_n762), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1079), .B1(new_n1081), .B2(new_n800), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n860), .A2(new_n861), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n1078), .B1(new_n1082), .B2(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n801), .A2(G330), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  OAI211_X1 g0887(.A(new_n1078), .B(new_n1085), .C1(new_n1082), .C2(new_n1083), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1087), .A2(new_n1088), .ZN(new_n1089));
  OAI221_X1 g0889(.A(new_n798), .B1(KEYINPUT117), .B2(new_n763), .C1(new_n799), .C2(new_n795), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n794), .A2(G330), .ZN(new_n1091));
  XNOR2_X1  g0891(.A(new_n1090), .B(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1076), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1091), .A2(new_n1077), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n1085), .A2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1095), .A2(new_n1081), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n436), .A2(G330), .A3(new_n685), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n846), .A2(new_n605), .A3(new_n1098), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n1099), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  AND2_X1   g0901(.A1(new_n1101), .A2(KEYINPUT118), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1089), .B1(new_n1102), .B2(new_n657), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1101), .A2(KEYINPUT118), .A3(new_n658), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1104), .A2(new_n690), .A3(new_n1087), .A4(new_n1088), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1075), .B1(new_n1103), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g0906(.A(new_n1106), .ZN(G378));
  NAND3_X1  g0907(.A1(new_n1087), .A2(new_n1088), .A3(new_n1097), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1108), .A2(new_n1100), .ZN(new_n1109));
  XOR2_X1   g0909(.A(KEYINPUT55), .B(KEYINPUT56), .Z(new_n1110));
  XNOR2_X1  g0910(.A(new_n310), .B(new_n1110), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n626), .B1(new_n270), .B2(new_n273), .ZN(new_n1112));
  XNOR2_X1  g0912(.A(new_n1111), .B(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OAI211_X1 g0914(.A(G330), .B(new_n828), .C1(new_n837), .C2(new_n838), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1115), .A2(new_n863), .A3(new_n855), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n852), .A2(new_n854), .ZN(new_n1117));
  NOR2_X1   g0917(.A1(new_n1117), .A2(new_n862), .ZN(new_n1118));
  NOR2_X1   g0918(.A1(new_n1118), .A2(new_n1115), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1114), .B1(new_n1116), .B2(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1115), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1121), .A2(new_n864), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1118), .A2(new_n1115), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1122), .A2(new_n1113), .A3(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1109), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT57), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1127));
  NAND4_X1  g0927(.A1(new_n1109), .A2(new_n1120), .A3(KEYINPUT57), .A4(new_n1124), .ZN(new_n1128));
  NAND3_X1  g0928(.A1(new_n1127), .A2(new_n658), .A3(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n1120), .A2(new_n691), .A3(new_n1124), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(new_n719), .A2(new_n225), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n891), .B1(G97), .B2(new_n714), .ZN(new_n1132));
  OAI221_X1 g0932(.A(new_n1132), .B1(new_n255), .B2(new_n773), .C1(new_n717), .C2(new_n701), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n711), .ZN(new_n1134));
  AOI211_X1 g0934(.A(new_n1131), .B(new_n1133), .C1(new_n311), .C2(new_n1134), .ZN(new_n1135));
  OAI211_X1 g0935(.A(new_n280), .B(new_n286), .C1(new_n721), .C2(new_n316), .ZN(new_n1136));
  XNOR2_X1  g0936(.A(new_n1136), .B(KEYINPUT121), .ZN(new_n1137));
  OAI211_X1 g0937(.A(new_n1135), .B(new_n1137), .C1(new_n253), .C2(new_n731), .ZN(new_n1138));
  XOR2_X1   g0938(.A(new_n1138), .B(KEYINPUT58), .Z(new_n1139));
  OAI21_X1  g0939(.A(new_n262), .B1(new_n284), .B2(G41), .ZN(new_n1140));
  OAI22_X1  g0940(.A1(new_n1068), .A2(new_n721), .B1(new_n779), .B2(new_n711), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n731), .A2(new_n1065), .ZN(new_n1142));
  AOI211_X1 g0942(.A(new_n1141), .B(new_n1142), .C1(G150), .C2(new_n1058), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n707), .A2(G125), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1143), .B(new_n1144), .C1(new_n784), .C2(new_n733), .ZN(new_n1145));
  XOR2_X1   g0945(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n1146));
  XOR2_X1   g0946(.A(new_n1145), .B(new_n1146), .Z(new_n1147));
  AOI211_X1 g0947(.A(G33), .B(G41), .C1(new_n702), .C2(G124), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n780), .B2(new_n719), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1140), .B1(new_n1147), .B2(new_n1149), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n698), .B1(new_n1139), .B2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g0951(.A(new_n692), .B1(G50), .B2(new_n791), .ZN(new_n1152));
  XNOR2_X1  g0952(.A(new_n1152), .B(KEYINPUT123), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1151), .B(new_n1153), .C1(new_n1113), .C2(new_n695), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1130), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1129), .A2(new_n1156), .ZN(G375));
  AOI22_X1  g0957(.A1(new_n1092), .A2(new_n1076), .B1(new_n1095), .B2(new_n1081), .ZN(new_n1158));
  NAND2_X1  g0958(.A1(new_n1158), .A2(new_n1099), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1101), .A2(new_n946), .A3(new_n1159), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n988), .A2(new_n892), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n706), .A2(G283), .B1(G116), .B2(new_n714), .ZN(new_n1162));
  OAI211_X1 g0962(.A(new_n1161), .B(new_n1162), .C1(new_n217), .C2(new_n721), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n701), .A2(new_n774), .ZN(new_n1164));
  NOR2_X1   g0964(.A1(new_n738), .A2(new_n326), .ZN(new_n1165));
  OAI21_X1  g0965(.A(new_n286), .B1(new_n773), .B2(new_n495), .ZN(new_n1166));
  NOR4_X1   g0966(.A1(new_n1163), .A2(new_n1164), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1058), .A2(G50), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n719), .A2(new_n225), .B1(new_n701), .B2(new_n1065), .ZN(new_n1169));
  AOI211_X1 g0969(.A(new_n286), .B(new_n1169), .C1(G150), .C2(new_n1134), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n706), .A2(G137), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n707), .A2(G132), .B1(new_n714), .B2(new_n1067), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1170), .A3(new_n1171), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n1173), .B1(G159), .B2(new_n722), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n698), .B1(new_n1167), .B2(new_n1174), .ZN(new_n1175));
  OAI211_X1 g0975(.A(new_n1175), .B(new_n692), .C1(G68), .C2(new_n791), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1077), .B2(new_n694), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n1097), .B2(new_n691), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1160), .A2(new_n1178), .ZN(G381));
  INV_X1    g0979(.A(new_n916), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT114), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n944), .B(new_n1180), .C1(new_n1022), .C2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1182), .A2(new_n688), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n691), .B1(new_n1183), .B2(new_n946), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n906), .B(new_n1048), .C1(new_n1184), .C2(new_n976), .ZN(new_n1185));
  NOR3_X1   g0985(.A1(new_n1185), .A2(G384), .A3(G381), .ZN(new_n1186));
  AOI21_X1  g0986(.A(new_n657), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1155), .B1(new_n1187), .B2(new_n1128), .ZN(new_n1188));
  NOR2_X1   g0988(.A1(G393), .A2(G396), .ZN(new_n1189));
  NAND4_X1  g0989(.A1(new_n1186), .A2(new_n1106), .A3(new_n1188), .A4(new_n1189), .ZN(G407));
  NAND2_X1  g0990(.A1(new_n1188), .A2(new_n1106), .ZN(new_n1191));
  OAI211_X1 g0991(.A(G407), .B(G213), .C1(G343), .C2(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT124), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(G409));
  INV_X1    g0994(.A(G213), .ZN(new_n1195));
  NOR2_X1   g0995(.A1(new_n1195), .A2(G343), .ZN(new_n1196));
  INV_X1    g0996(.A(new_n1196), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1109), .A2(new_n1120), .A3(new_n946), .A4(new_n1124), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1156), .A2(new_n1106), .A3(new_n1198), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1197), .B(new_n1199), .C1(new_n1188), .C2(new_n1106), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1196), .A2(G2897), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT60), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n657), .B1(new_n1159), .B2(new_n1203), .ZN(new_n1204));
  OAI211_X1 g1004(.A(new_n1204), .B(new_n1101), .C1(new_n1203), .C2(new_n1159), .ZN(new_n1205));
  AND3_X1   g1005(.A1(new_n1205), .A2(G384), .A3(new_n1178), .ZN(new_n1206));
  AOI21_X1  g1006(.A(G384), .B1(new_n1205), .B2(new_n1178), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1202), .B1(new_n1206), .B2(new_n1207), .ZN(new_n1208));
  NAND2_X1  g1008(.A1(new_n1205), .A2(new_n1178), .ZN(new_n1209));
  INV_X1    g1009(.A(G384), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1209), .A2(new_n1210), .ZN(new_n1211));
  NAND3_X1  g1011(.A1(new_n1205), .A2(G384), .A3(new_n1178), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1211), .A2(new_n1212), .A3(new_n1201), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1208), .A2(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1200), .A2(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1215), .A2(KEYINPUT63), .ZN(new_n1216));
  AOI21_X1  g1016(.A(new_n1196), .B1(G375), .B2(G378), .ZN(new_n1217));
  NOR2_X1   g1017(.A1(new_n1206), .A2(new_n1207), .ZN(new_n1218));
  NAND3_X1  g1018(.A1(new_n1217), .A2(new_n1218), .A3(new_n1199), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1216), .A2(new_n1219), .ZN(new_n1220));
  INV_X1    g1020(.A(KEYINPUT61), .ZN(new_n1221));
  AOI21_X1  g1021(.A(new_n1181), .B1(new_n935), .B2(new_n940), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1222), .A2(new_n943), .A3(new_n916), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n946), .B1(new_n1223), .B2(new_n687), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n976), .B1(new_n1224), .B2(new_n690), .ZN(new_n1225));
  OAI21_X1  g1025(.A(G390), .B1(new_n1225), .B2(new_n907), .ZN(new_n1226));
  INV_X1    g1026(.A(KEYINPUT125), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1226), .A2(new_n1185), .A3(new_n1227), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(G393), .B(new_n757), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1228), .A2(new_n1229), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1229), .B1(new_n978), .B2(KEYINPUT126), .ZN(new_n1231));
  NAND4_X1  g1031(.A1(new_n1231), .A2(new_n1227), .A3(new_n1185), .A4(new_n1226), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1226), .A2(new_n1185), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT126), .ZN(new_n1234));
  AND4_X1   g1034(.A1(new_n1221), .A2(new_n1230), .A3(new_n1232), .A4(new_n1234), .ZN(new_n1235));
  NAND4_X1  g1035(.A1(new_n1217), .A2(KEYINPUT63), .A3(new_n1218), .A4(new_n1199), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1236), .A2(KEYINPUT127), .ZN(new_n1237));
  INV_X1    g1037(.A(new_n1218), .ZN(new_n1238));
  NOR2_X1   g1038(.A1(new_n1200), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT127), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1239), .A2(new_n1240), .A3(KEYINPUT63), .ZN(new_n1241));
  NAND4_X1  g1041(.A1(new_n1220), .A2(new_n1235), .A3(new_n1237), .A4(new_n1241), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1217), .A2(new_n1243), .A3(new_n1218), .A4(new_n1199), .ZN(new_n1244));
  OAI21_X1  g1044(.A(KEYINPUT62), .B1(new_n1200), .B2(new_n1238), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n1244), .A2(new_n1245), .A3(new_n1221), .A4(new_n1215), .ZN(new_n1246));
  AOI22_X1  g1046(.A1(new_n1228), .A2(new_n1229), .B1(new_n1233), .B2(KEYINPUT126), .ZN(new_n1247));
  NAND2_X1  g1047(.A1(new_n1247), .A2(new_n1232), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1246), .A2(new_n1248), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1242), .A2(new_n1249), .ZN(G405));
  NAND2_X1  g1050(.A1(G375), .A2(G378), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1251), .A2(new_n1191), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1252), .A2(new_n1218), .ZN(new_n1253));
  NAND3_X1  g1053(.A1(new_n1251), .A2(new_n1191), .A3(new_n1238), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1253), .A2(new_n1254), .ZN(new_n1255));
  AND2_X1   g1055(.A1(new_n1255), .A2(new_n1248), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1255), .A2(new_n1248), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1256), .A2(new_n1257), .ZN(G402));
endmodule


