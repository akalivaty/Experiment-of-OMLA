//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 0 0 1 1 0 1 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:39 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n642, new_n643, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n749, new_n750, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n902, new_n903, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n937, new_n938,
    new_n939, new_n940, new_n942, new_n943, new_n944, new_n945, new_n946;
  XNOR2_X1  g000(.A(G141gat), .B(G148gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT2), .ZN(new_n203));
  AOI21_X1  g002(.A(new_n203), .B1(G155gat), .B2(G162gat), .ZN(new_n204));
  INV_X1    g003(.A(G155gat), .ZN(new_n205));
  INV_X1    g004(.A(G162gat), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  OAI22_X1  g006(.A1(new_n202), .A2(new_n204), .B1(KEYINPUT75), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G155gat), .B(G162gat), .Z(new_n209));
  OR2_X1    g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n208), .A2(new_n209), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G113gat), .ZN(new_n213));
  INV_X1    g012(.A(G120gat), .ZN(new_n214));
  AOI21_X1  g013(.A(KEYINPUT1), .B1(new_n213), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n215), .B1(new_n213), .B2(new_n214), .ZN(new_n216));
  XNOR2_X1  g015(.A(G127gat), .B(G134gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n216), .B(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n212), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT4), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT4), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n212), .A2(new_n221), .A3(new_n218), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n220), .A2(new_n222), .ZN(new_n223));
  NAND2_X1  g022(.A1(G225gat), .A2(G233gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT3), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n212), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(new_n218), .ZN(new_n227));
  NAND3_X1  g026(.A1(new_n210), .A2(KEYINPUT3), .A3(new_n211), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n226), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  XOR2_X1   g028(.A(KEYINPUT77), .B(KEYINPUT5), .Z(new_n230));
  NAND4_X1  g029(.A1(new_n223), .A2(new_n224), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT76), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n222), .A2(new_n232), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n212), .A2(KEYINPUT76), .A3(new_n221), .A4(new_n218), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n233), .A2(new_n234), .A3(new_n220), .ZN(new_n235));
  INV_X1    g034(.A(new_n224), .ZN(new_n236));
  AND2_X1   g035(.A1(new_n228), .A2(new_n227), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n236), .B1(new_n237), .B2(new_n226), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n235), .A2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n210), .A2(new_n211), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n240), .A2(new_n227), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n241), .A2(new_n219), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n230), .B1(new_n242), .B2(new_n236), .ZN(new_n243));
  AND3_X1   g042(.A1(new_n239), .A2(KEYINPUT78), .A3(new_n243), .ZN(new_n244));
  AOI21_X1  g043(.A(KEYINPUT78), .B1(new_n239), .B2(new_n243), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n231), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(G1gat), .B(G29gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(KEYINPUT0), .ZN(new_n248));
  XNOR2_X1  g047(.A(G57gat), .B(G85gat), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n248), .B(new_n249), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  AOI21_X1  g050(.A(KEYINPUT6), .B1(new_n246), .B2(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n239), .A2(new_n243), .ZN(new_n253));
  INV_X1    g052(.A(KEYINPUT78), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n239), .A2(KEYINPUT78), .A3(new_n243), .ZN(new_n256));
  NAND2_X1  g055(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT79), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n257), .A2(new_n258), .A3(new_n250), .A4(new_n231), .ZN(new_n259));
  OAI211_X1 g058(.A(new_n250), .B(new_n231), .C1(new_n244), .C2(new_n245), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT79), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n252), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n246), .A2(KEYINPUT6), .A3(new_n251), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n262), .A2(new_n263), .ZN(new_n264));
  XNOR2_X1  g063(.A(G197gat), .B(G204gat), .ZN(new_n265));
  XNOR2_X1  g064(.A(KEYINPUT71), .B(G211gat), .ZN(new_n266));
  INV_X1    g065(.A(G218gat), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n265), .B1(new_n268), .B2(KEYINPUT22), .ZN(new_n269));
  XNOR2_X1  g068(.A(G211gat), .B(G218gat), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT72), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(new_n269), .B(new_n272), .Z(new_n273));
  INV_X1    g072(.A(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(G169gat), .ZN(new_n275));
  INV_X1    g074(.A(G176gat), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(G169gat), .A2(G176gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(KEYINPUT64), .A3(KEYINPUT23), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n279), .A2(KEYINPUT23), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT23), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n282), .B1(G169gat), .B2(G176gat), .ZN(new_n283));
  NOR2_X1   g082(.A1(KEYINPUT64), .A2(KEYINPUT25), .ZN(new_n284));
  NAND3_X1  g083(.A1(new_n281), .A2(new_n283), .A3(new_n284), .ZN(new_n285));
  AOI21_X1  g084(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  INV_X1    g086(.A(G190gat), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  AOI22_X1  g089(.A1(new_n280), .A2(new_n285), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT25), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(KEYINPUT65), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n278), .B1(new_n291), .B2(new_n293), .ZN(new_n294));
  OAI22_X1  g093(.A1(KEYINPUT69), .A2(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(KEYINPUT69), .A2(KEYINPUT26), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n277), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OR2_X1    g096(.A1(new_n295), .A2(new_n296), .ZN(new_n298));
  AOI22_X1  g097(.A1(new_n297), .A2(new_n298), .B1(G183gat), .B2(G190gat), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT27), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n300), .A2(G183gat), .ZN(new_n301));
  NAND2_X1  g100(.A1(new_n287), .A2(KEYINPUT27), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT68), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  AOI21_X1  g104(.A(G190gat), .B1(new_n301), .B2(KEYINPUT68), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT28), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT28), .ZN(new_n308));
  NOR3_X1   g107(.A1(new_n303), .A2(new_n308), .A3(G190gat), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n299), .B1(new_n307), .B2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n281), .A2(new_n283), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n277), .A2(KEYINPUT65), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT66), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n290), .B(new_n313), .ZN(new_n314));
  OR3_X1    g113(.A1(KEYINPUT67), .A2(G183gat), .A3(G190gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n286), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n315), .A2(new_n316), .A3(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n311), .B(new_n312), .C1(new_n314), .C2(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(KEYINPUT25), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n294), .A2(new_n310), .A3(new_n320), .ZN(new_n321));
  AND2_X1   g120(.A1(G226gat), .A2(G233gat), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n324));
  AND2_X1   g123(.A1(new_n321), .A2(new_n324), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n274), .B(new_n323), .C1(new_n325), .C2(new_n322), .ZN(new_n326));
  INV_X1    g125(.A(new_n323), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n322), .B1(new_n321), .B2(new_n324), .ZN(new_n328));
  OAI21_X1  g127(.A(new_n273), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n326), .A2(new_n329), .ZN(new_n330));
  XOR2_X1   g129(.A(G8gat), .B(G36gat), .Z(new_n331));
  XNOR2_X1  g130(.A(new_n331), .B(KEYINPUT73), .ZN(new_n332));
  XNOR2_X1  g131(.A(G64gat), .B(G92gat), .ZN(new_n333));
  XNOR2_X1  g132(.A(new_n332), .B(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n334), .B(KEYINPUT74), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n330), .A2(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(new_n334), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n330), .A2(new_n337), .ZN(new_n338));
  OAI21_X1  g137(.A(KEYINPUT30), .B1(new_n336), .B2(new_n338), .ZN(new_n339));
  OR2_X1    g138(.A1(new_n338), .A2(KEYINPUT30), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n321), .B(new_n227), .ZN(new_n343));
  INV_X1    g142(.A(G227gat), .ZN(new_n344));
  INV_X1    g143(.A(G233gat), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(KEYINPUT33), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  XNOR2_X1  g146(.A(G15gat), .B(G43gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(G71gat), .B(G99gat), .ZN(new_n349));
  XNOR2_X1  g148(.A(new_n348), .B(new_n349), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n347), .A2(new_n350), .ZN(new_n351));
  XNOR2_X1  g150(.A(new_n321), .B(new_n218), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT34), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n352), .B(new_n353), .C1(new_n344), .C2(new_n345), .ZN(new_n354));
  OAI21_X1  g153(.A(KEYINPUT34), .B1(new_n343), .B2(new_n346), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n351), .A2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n343), .A2(new_n346), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n358), .A2(KEYINPUT32), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  OAI211_X1 g159(.A(new_n354), .B(new_n355), .C1(new_n347), .C2(new_n350), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n357), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n360), .B1(new_n357), .B2(new_n361), .ZN(new_n364));
  OAI21_X1  g163(.A(new_n225), .B1(new_n273), .B2(KEYINPUT29), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n365), .A2(new_n240), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n226), .A2(new_n324), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n273), .ZN(new_n368));
  NAND4_X1  g167(.A1(new_n366), .A2(G228gat), .A3(G233gat), .A4(new_n368), .ZN(new_n369));
  XNOR2_X1  g168(.A(G78gat), .B(G106gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(KEYINPUT31), .B(G50gat), .ZN(new_n371));
  XNOR2_X1  g170(.A(new_n370), .B(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  NOR2_X1   g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(KEYINPUT81), .A2(G22gat), .ZN(new_n375));
  AOI21_X1  g174(.A(new_n374), .B1(new_n375), .B2(new_n372), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT29), .B1(new_n269), .B2(new_n270), .ZN(new_n378));
  OAI21_X1  g177(.A(new_n378), .B1(new_n269), .B2(new_n270), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(new_n225), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(new_n240), .ZN(new_n381));
  AOI22_X1  g180(.A1(new_n381), .A2(KEYINPUT80), .B1(new_n273), .B2(new_n367), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT80), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n380), .A2(new_n383), .A3(new_n240), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n382), .A2(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(G228gat), .ZN(new_n386));
  NOR2_X1   g185(.A1(new_n386), .A2(new_n345), .ZN(new_n387));
  OAI211_X1 g186(.A(new_n369), .B(new_n377), .C1(new_n385), .C2(new_n387), .ZN(new_n388));
  AOI22_X1  g187(.A1(new_n382), .A2(new_n384), .B1(G228gat), .B2(G233gat), .ZN(new_n389));
  INV_X1    g188(.A(new_n369), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n376), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n388), .A2(new_n391), .ZN(new_n392));
  NOR3_X1   g191(.A1(new_n363), .A2(new_n364), .A3(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n264), .A2(new_n342), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT83), .B(KEYINPUT35), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  AOI21_X1  g195(.A(new_n341), .B1(new_n262), .B2(new_n263), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT83), .ZN(new_n398));
  NAND4_X1  g197(.A1(new_n397), .A2(new_n398), .A3(KEYINPUT35), .A4(new_n393), .ZN(new_n399));
  INV_X1    g198(.A(new_n364), .ZN(new_n400));
  AND2_X1   g199(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n401));
  NOR2_X1   g200(.A1(KEYINPUT70), .A2(KEYINPUT36), .ZN(new_n402));
  NOR2_X1   g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND3_X1  g203(.A1(new_n400), .A2(new_n362), .A3(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n363), .A2(new_n364), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n405), .B1(new_n406), .B2(new_n401), .ZN(new_n407));
  INV_X1    g206(.A(new_n392), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n407), .B1(new_n397), .B2(new_n408), .ZN(new_n409));
  NOR2_X1   g208(.A1(KEYINPUT82), .A2(KEYINPUT40), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n223), .A2(new_n229), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT39), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n412), .A3(new_n236), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n413), .A2(new_n250), .ZN(new_n414));
  OAI21_X1  g213(.A(KEYINPUT39), .B1(new_n242), .B2(new_n236), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n415), .B1(new_n236), .B2(new_n411), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n410), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n411), .A2(new_n236), .ZN(new_n418));
  INV_X1    g217(.A(new_n415), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(new_n410), .ZN(new_n421));
  NAND4_X1  g220(.A1(new_n420), .A2(new_n250), .A3(new_n421), .A4(new_n413), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n417), .A2(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n423), .B1(new_n251), .B2(new_n246), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n392), .B1(new_n424), .B2(new_n341), .ZN(new_n425));
  INV_X1    g224(.A(KEYINPUT37), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n326), .A2(new_n329), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT38), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(new_n428), .A3(new_n335), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n426), .B1(new_n326), .B2(new_n329), .ZN(new_n430));
  OAI22_X1  g229(.A1(new_n429), .A2(new_n430), .B1(new_n330), .B2(new_n337), .ZN(new_n431));
  INV_X1    g230(.A(new_n430), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n432), .A2(new_n337), .A3(new_n427), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n431), .B1(KEYINPUT38), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n262), .A3(new_n263), .ZN(new_n435));
  AND2_X1   g234(.A1(new_n425), .A2(new_n435), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n396), .B(new_n399), .C1(new_n409), .C2(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G113gat), .B(G141gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(G197gat), .ZN(new_n439));
  XOR2_X1   g238(.A(KEYINPUT11), .B(G169gat), .Z(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  XNOR2_X1  g240(.A(new_n441), .B(KEYINPUT12), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  XNOR2_X1  g242(.A(G15gat), .B(G22gat), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n444), .A2(G1gat), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT16), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n444), .B1(new_n448), .B2(G1gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n445), .A2(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n447), .A2(new_n450), .A3(G8gat), .ZN(new_n451));
  INV_X1    g250(.A(G8gat), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n445), .B(new_n449), .C1(new_n446), .C2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  NOR2_X1   g253(.A1(G29gat), .A2(G36gat), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT85), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT14), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n455), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  AND2_X1   g259(.A1(new_n455), .A2(new_n459), .ZN(new_n461));
  OAI21_X1  g260(.A(KEYINPUT86), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  AND2_X1   g261(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n463));
  NOR2_X1   g262(.A1(KEYINPUT85), .A2(KEYINPUT14), .ZN(new_n464));
  OAI22_X1  g263(.A1(new_n463), .A2(new_n464), .B1(G29gat), .B2(G36gat), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT86), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n455), .A2(new_n459), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n465), .A2(new_n466), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(G29gat), .A2(G36gat), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT87), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT87), .ZN(new_n471));
  NAND3_X1  g270(.A1(new_n471), .A2(G29gat), .A3(G36gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  NAND3_X1  g273(.A1(new_n462), .A2(new_n468), .A3(new_n474), .ZN(new_n475));
  AND2_X1   g274(.A1(G43gat), .A2(G50gat), .ZN(new_n476));
  NOR2_X1   g275(.A1(G43gat), .A2(G50gat), .ZN(new_n477));
  OAI21_X1  g276(.A(KEYINPUT84), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(G43gat), .ZN(new_n479));
  INV_X1    g278(.A(G50gat), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT84), .ZN(new_n482));
  NAND2_X1  g281(.A1(G43gat), .A2(G50gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n481), .A2(new_n482), .A3(new_n483), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n478), .A2(new_n484), .A3(KEYINPUT15), .ZN(new_n485));
  INV_X1    g284(.A(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n475), .A2(new_n486), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n476), .A2(new_n477), .A3(KEYINPUT15), .ZN(new_n488));
  NOR2_X1   g287(.A1(new_n488), .A2(new_n473), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n465), .A2(new_n467), .ZN(new_n490));
  NAND3_X1  g289(.A1(new_n489), .A2(new_n485), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n487), .A2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT17), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n454), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT89), .ZN(new_n495));
  AND3_X1   g294(.A1(new_n489), .A2(new_n485), .A3(new_n490), .ZN(new_n496));
  AOI21_X1  g295(.A(new_n496), .B1(new_n486), .B2(new_n475), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n495), .B1(new_n497), .B2(KEYINPUT17), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n487), .A2(new_n495), .A3(KEYINPUT17), .A4(new_n491), .ZN(new_n499));
  INV_X1    g298(.A(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n494), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(G229gat), .A2(G233gat), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n492), .A2(new_n454), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n501), .A2(KEYINPUT18), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n454), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(new_n497), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(new_n503), .ZN(new_n507));
  XOR2_X1   g306(.A(new_n502), .B(KEYINPUT13), .Z(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n503), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n487), .A2(KEYINPUT17), .A3(new_n491), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(KEYINPUT89), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(new_n499), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n511), .B1(new_n514), .B2(new_n494), .ZN(new_n515));
  AOI21_X1  g314(.A(KEYINPUT18), .B1(new_n515), .B2(new_n502), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n443), .B1(new_n510), .B2(new_n516), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n518));
  INV_X1    g317(.A(KEYINPUT18), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  NAND4_X1  g319(.A1(new_n520), .A2(new_n442), .A3(new_n504), .A4(new_n509), .ZN(new_n521));
  AND3_X1   g320(.A1(new_n517), .A2(KEYINPUT90), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g321(.A(KEYINPUT90), .B1(new_n517), .B2(new_n521), .ZN(new_n523));
  NOR2_X1   g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n437), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(G99gat), .A2(G106gat), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n527), .A2(KEYINPUT8), .ZN(new_n528));
  NAND2_X1  g327(.A1(G85gat), .A2(G92gat), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  INV_X1    g330(.A(G85gat), .ZN(new_n532));
  INV_X1    g331(.A(G92gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n535));
  NAND4_X1  g334(.A1(new_n528), .A2(new_n531), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(G99gat), .B(G106gat), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n536), .A2(new_n538), .ZN(new_n539));
  AOI22_X1  g338(.A1(KEYINPUT8), .A2(new_n527), .B1(new_n532), .B2(new_n533), .ZN(new_n540));
  NAND4_X1  g339(.A1(new_n540), .A2(new_n537), .A3(new_n531), .A4(new_n535), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n539), .A2(KEYINPUT95), .A3(new_n541), .ZN(new_n542));
  AND2_X1   g341(.A1(new_n531), .A2(new_n535), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT95), .ZN(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n537), .A4(new_n540), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(KEYINPUT96), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n542), .A2(KEYINPUT96), .A3(new_n545), .ZN(new_n549));
  AND3_X1   g348(.A1(new_n492), .A2(new_n548), .A3(new_n549), .ZN(new_n550));
  AND2_X1   g349(.A1(G232gat), .A2(G233gat), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n550), .B1(KEYINPUT41), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT97), .ZN(new_n553));
  AOI22_X1  g352(.A1(new_n493), .A2(new_n492), .B1(new_n548), .B2(new_n549), .ZN(new_n554));
  AND3_X1   g353(.A1(new_n514), .A2(new_n553), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g354(.A(new_n553), .B1(new_n514), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n552), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G190gat), .B(G218gat), .Z(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n551), .A2(KEYINPUT41), .ZN(new_n560));
  XNOR2_X1  g359(.A(new_n560), .B(KEYINPUT94), .ZN(new_n561));
  XOR2_X1   g360(.A(G134gat), .B(G162gat), .Z(new_n562));
  XNOR2_X1  g361(.A(new_n561), .B(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT98), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n558), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n552), .B(new_n566), .C1(new_n555), .C2(new_n556), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n559), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n563), .B(KEYINPUT98), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n570), .B1(new_n559), .B2(new_n567), .ZN(new_n571));
  NOR2_X1   g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(KEYINPUT21), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT91), .ZN(new_n574));
  INV_X1    g373(.A(G64gat), .ZN(new_n575));
  OAI21_X1  g374(.A(new_n574), .B1(new_n575), .B2(G57gat), .ZN(new_n576));
  INV_X1    g375(.A(G57gat), .ZN(new_n577));
  NAND3_X1  g376(.A1(new_n577), .A2(KEYINPUT91), .A3(G64gat), .ZN(new_n578));
  OAI211_X1 g377(.A(new_n576), .B(new_n578), .C1(new_n577), .C2(G64gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(G71gat), .A2(G78gat), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  INV_X1    g380(.A(KEYINPUT92), .ZN(new_n582));
  NAND2_X1  g381(.A1(G71gat), .A2(G78gat), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n583), .ZN(new_n585));
  OAI21_X1  g384(.A(KEYINPUT92), .B1(new_n585), .B2(new_n580), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g387(.A1(new_n579), .A2(new_n584), .A3(new_n586), .A4(new_n588), .ZN(new_n589));
  XNOR2_X1  g388(.A(G57gat), .B(G64gat), .ZN(new_n590));
  OAI211_X1 g389(.A(new_n583), .B(new_n581), .C1(new_n590), .C2(new_n587), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  OAI21_X1  g391(.A(new_n505), .B1(new_n573), .B2(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n592), .A2(new_n573), .ZN(new_n594));
  XNOR2_X1  g393(.A(G127gat), .B(G155gat), .ZN(new_n595));
  XNOR2_X1  g394(.A(new_n594), .B(new_n595), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n593), .B(new_n596), .ZN(new_n597));
  NAND2_X1  g396(.A1(G231gat), .A2(G233gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT93), .ZN(new_n599));
  XOR2_X1   g398(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  XNOR2_X1  g400(.A(G183gat), .B(G211gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n597), .B(new_n603), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n572), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g404(.A1(G230gat), .A2(G233gat), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT10), .ZN(new_n608));
  NOR2_X1   g407(.A1(new_n592), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n548), .A2(new_n549), .A3(new_n609), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n592), .A2(new_n545), .A3(new_n542), .ZN(new_n611));
  NAND4_X1  g410(.A1(new_n589), .A2(new_n539), .A3(new_n591), .A4(new_n541), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n611), .A2(new_n608), .A3(new_n612), .ZN(new_n613));
  AOI21_X1  g412(.A(new_n607), .B1(new_n610), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n606), .B1(new_n611), .B2(new_n612), .ZN(new_n615));
  XNOR2_X1  g414(.A(G120gat), .B(G148gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G176gat), .B(G204gat), .ZN(new_n617));
  XOR2_X1   g416(.A(new_n616), .B(new_n617), .Z(new_n618));
  INV_X1    g417(.A(new_n618), .ZN(new_n619));
  NOR3_X1   g418(.A1(new_n614), .A2(new_n615), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n614), .B2(new_n615), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n605), .A2(new_n624), .ZN(new_n625));
  INV_X1    g424(.A(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n526), .A2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n264), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XNOR2_X1  g429(.A(new_n630), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g430(.A(new_n452), .B1(new_n628), .B2(new_n341), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT16), .B(G8gat), .ZN(new_n633));
  NOR3_X1   g432(.A1(new_n627), .A2(new_n342), .A3(new_n633), .ZN(new_n634));
  OAI21_X1  g433(.A(KEYINPUT42), .B1(new_n632), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n635), .B1(KEYINPUT42), .B2(new_n634), .ZN(G1325gat));
  AOI21_X1  g435(.A(G15gat), .B1(new_n628), .B2(new_n406), .ZN(new_n637));
  INV_X1    g436(.A(new_n407), .ZN(new_n638));
  NAND2_X1  g437(.A1(new_n638), .A2(G15gat), .ZN(new_n639));
  XOR2_X1   g438(.A(new_n639), .B(KEYINPUT99), .Z(new_n640));
  AOI21_X1  g439(.A(new_n637), .B1(new_n628), .B2(new_n640), .ZN(G1326gat));
  NOR2_X1   g440(.A1(new_n627), .A2(new_n408), .ZN(new_n642));
  XOR2_X1   g441(.A(KEYINPUT43), .B(G22gat), .Z(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(G1327gat));
  NAND3_X1  g443(.A1(new_n572), .A2(new_n604), .A3(new_n624), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n645), .B(KEYINPUT100), .Z(new_n646));
  NOR2_X1   g445(.A1(new_n264), .A2(G29gat), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n526), .A2(new_n646), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(KEYINPUT45), .ZN(new_n649));
  INV_X1    g448(.A(KEYINPUT45), .ZN(new_n650));
  NAND4_X1  g449(.A1(new_n526), .A2(new_n650), .A3(new_n646), .A4(new_n647), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n437), .A2(new_n572), .ZN(new_n653));
  INV_X1    g452(.A(KEYINPUT44), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n437), .A2(KEYINPUT44), .A3(new_n572), .ZN(new_n656));
  AND2_X1   g455(.A1(new_n517), .A2(new_n521), .ZN(new_n657));
  INV_X1    g456(.A(new_n604), .ZN(new_n658));
  NOR3_X1   g457(.A1(new_n657), .A2(new_n658), .A3(new_n623), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n655), .A2(new_n629), .A3(new_n656), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n660), .A2(G29gat), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n652), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n662), .A2(KEYINPUT101), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT101), .ZN(new_n664));
  NAND3_X1  g463(.A1(new_n652), .A2(new_n664), .A3(new_n661), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(G1328gat));
  NAND2_X1  g465(.A1(new_n526), .A2(new_n646), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n342), .A2(G36gat), .ZN(new_n668));
  OAI22_X1  g467(.A1(new_n667), .A2(new_n668), .B1(KEYINPUT102), .B2(KEYINPUT46), .ZN(new_n669));
  AND2_X1   g468(.A1(KEYINPUT102), .A2(KEYINPUT46), .ZN(new_n670));
  XNOR2_X1  g469(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(new_n656), .ZN(new_n672));
  AOI21_X1  g471(.A(KEYINPUT44), .B1(new_n437), .B2(new_n572), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n674), .A2(new_n341), .A3(new_n659), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(G36gat), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n671), .A2(new_n676), .ZN(G1329gat));
  INV_X1    g476(.A(new_n406), .ZN(new_n678));
  NOR2_X1   g477(.A1(new_n678), .A2(G43gat), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n526), .A2(new_n646), .A3(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND4_X1  g481(.A1(new_n526), .A2(KEYINPUT103), .A3(new_n646), .A4(new_n679), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  NAND4_X1  g483(.A1(new_n655), .A2(new_n638), .A3(new_n656), .A4(new_n659), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G43gat), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT47), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n684), .A2(KEYINPUT47), .A3(new_n686), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(G1330gat));
  NAND4_X1  g490(.A1(new_n655), .A2(new_n392), .A3(new_n656), .A4(new_n659), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n692), .A2(G50gat), .ZN(new_n693));
  NAND4_X1  g492(.A1(new_n526), .A2(new_n480), .A3(new_n392), .A4(new_n646), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n693), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT48), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1331gat));
  INV_X1    g496(.A(new_n657), .ZN(new_n698));
  NOR4_X1   g497(.A1(new_n572), .A2(new_n698), .A3(new_n604), .A4(new_n624), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n437), .A2(new_n699), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n700), .A2(new_n264), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(new_n577), .ZN(G1332gat));
  AND2_X1   g501(.A1(new_n437), .A2(new_n699), .ZN(new_n703));
  AOI21_X1  g502(.A(new_n342), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT104), .ZN(new_n706));
  OR2_X1    g505(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n707));
  XNOR2_X1  g506(.A(new_n706), .B(new_n707), .ZN(G1333gat));
  INV_X1    g507(.A(G71gat), .ZN(new_n709));
  AOI21_X1  g508(.A(new_n709), .B1(new_n703), .B2(new_n638), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT105), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n703), .A2(new_n711), .A3(new_n406), .ZN(new_n712));
  OAI21_X1  g511(.A(KEYINPUT105), .B1(new_n700), .B2(new_n678), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n710), .B1(new_n714), .B2(new_n709), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g515(.A1(new_n703), .A2(new_n392), .ZN(new_n717));
  XNOR2_X1  g516(.A(new_n717), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g517(.A1(new_n657), .A2(new_n604), .ZN(new_n719));
  XNOR2_X1  g518(.A(new_n719), .B(KEYINPUT106), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(new_n623), .ZN(new_n721));
  XOR2_X1   g520(.A(new_n721), .B(KEYINPUT107), .Z(new_n722));
  NAND2_X1  g521(.A1(new_n674), .A2(new_n722), .ZN(new_n723));
  OAI21_X1  g522(.A(G85gat), .B1(new_n723), .B2(new_n264), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n437), .A2(new_n572), .A3(new_n720), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT51), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g526(.A1(new_n437), .A2(KEYINPUT51), .A3(new_n572), .A4(new_n720), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(new_n729), .ZN(new_n730));
  NOR3_X1   g529(.A1(new_n264), .A2(G85gat), .A3(new_n624), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(KEYINPUT108), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n724), .B1(new_n730), .B2(new_n732), .ZN(G1336gat));
  NAND4_X1  g532(.A1(new_n655), .A2(new_n722), .A3(new_n341), .A4(new_n656), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(G92gat), .ZN(new_n735));
  INV_X1    g534(.A(new_n735), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT109), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n725), .A2(new_n737), .A3(KEYINPUT51), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n725), .B2(new_n737), .ZN(new_n739));
  NOR3_X1   g538(.A1(new_n342), .A2(G92gat), .A3(new_n624), .ZN(new_n740));
  INV_X1    g539(.A(new_n740), .ZN(new_n741));
  NOR3_X1   g540(.A1(new_n738), .A2(new_n739), .A3(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT52), .B1(new_n736), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT52), .B1(new_n729), .B2(new_n740), .ZN(new_n744));
  INV_X1    g543(.A(KEYINPUT110), .ZN(new_n745));
  AND3_X1   g544(.A1(new_n744), .A2(new_n745), .A3(new_n735), .ZN(new_n746));
  AOI21_X1  g545(.A(new_n745), .B1(new_n744), .B2(new_n735), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n743), .B1(new_n746), .B2(new_n747), .ZN(G1337gat));
  OAI21_X1  g547(.A(G99gat), .B1(new_n723), .B2(new_n407), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n678), .A2(G99gat), .A3(new_n624), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n730), .B2(new_n750), .ZN(G1338gat));
  NAND3_X1  g550(.A1(new_n674), .A2(new_n392), .A3(new_n722), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G106gat), .ZN(new_n753));
  NOR3_X1   g552(.A1(new_n408), .A2(G106gat), .A3(new_n624), .ZN(new_n754));
  AOI21_X1  g553(.A(KEYINPUT53), .B1(new_n729), .B2(new_n754), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n753), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n738), .A2(new_n739), .ZN(new_n757));
  AOI22_X1  g556(.A1(G106gat), .A2(new_n752), .B1(new_n757), .B2(new_n754), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT53), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n756), .B1(new_n758), .B2(new_n759), .ZN(G1339gat));
  INV_X1    g559(.A(KEYINPUT112), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n515), .B2(new_n502), .ZN(new_n762));
  INV_X1    g561(.A(new_n502), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n473), .B1(new_n490), .B2(KEYINPUT86), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n485), .B1(new_n764), .B2(new_n468), .ZN(new_n765));
  OAI21_X1  g564(.A(new_n493), .B1(new_n765), .B2(new_n496), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(new_n505), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n767), .B1(new_n513), .B2(new_n499), .ZN(new_n768));
  OAI211_X1 g567(.A(KEYINPUT112), .B(new_n763), .C1(new_n768), .C2(new_n511), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n507), .A2(new_n508), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n762), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n771), .A2(new_n441), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n772), .A2(new_n521), .A3(new_n623), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n610), .A2(new_n613), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n774), .A2(new_n606), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n610), .A2(new_n607), .A3(new_n613), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(KEYINPUT54), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT54), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n618), .B1(new_n614), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT55), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n620), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n777), .A2(new_n779), .A3(KEYINPUT111), .A4(KEYINPUT55), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n777), .A2(KEYINPUT55), .A3(new_n779), .ZN(new_n784));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n773), .B1(new_n657), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(KEYINPUT114), .ZN(new_n789));
  INV_X1    g588(.A(new_n572), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT114), .ZN(new_n791));
  OAI211_X1 g590(.A(new_n773), .B(new_n791), .C1(new_n657), .C2(new_n787), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n789), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT113), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n772), .A2(new_n794), .A3(new_n521), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n782), .A2(new_n783), .A3(new_n786), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n559), .A2(new_n565), .A3(new_n567), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n559), .A2(new_n567), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n798), .A2(new_n569), .ZN(new_n799));
  NAND4_X1  g598(.A1(new_n795), .A2(new_n796), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  AOI21_X1  g599(.A(new_n794), .B1(new_n772), .B2(new_n521), .ZN(new_n801));
  OR2_X1    g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  AOI21_X1  g601(.A(new_n658), .B1(new_n793), .B2(new_n802), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n625), .A2(new_n698), .ZN(new_n804));
  OR2_X1    g603(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(new_n393), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n806), .A2(new_n341), .ZN(new_n807));
  NAND3_X1  g606(.A1(new_n805), .A2(new_n807), .A3(new_n629), .ZN(new_n808));
  INV_X1    g607(.A(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n213), .A3(new_n698), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n805), .A2(new_n807), .A3(new_n629), .A4(new_n525), .ZN(new_n811));
  AND3_X1   g610(.A1(new_n811), .A2(KEYINPUT115), .A3(G113gat), .ZN(new_n812));
  AOI21_X1  g611(.A(KEYINPUT115), .B1(new_n811), .B2(G113gat), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n810), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n814), .A2(KEYINPUT116), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT116), .ZN(new_n816));
  OAI211_X1 g615(.A(new_n816), .B(new_n810), .C1(new_n812), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n815), .A2(new_n817), .ZN(G1340gat));
  OAI21_X1  g617(.A(G120gat), .B1(new_n808), .B2(new_n624), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n623), .A2(new_n214), .ZN(new_n820));
  XNOR2_X1  g619(.A(new_n820), .B(KEYINPUT117), .ZN(new_n821));
  OAI21_X1  g620(.A(new_n819), .B1(new_n808), .B2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT118), .ZN(new_n823));
  XNOR2_X1  g622(.A(new_n822), .B(new_n823), .ZN(G1341gat));
  NAND2_X1  g623(.A1(new_n809), .A2(new_n658), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G127gat), .ZN(G1342gat));
  INV_X1    g625(.A(KEYINPUT119), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n808), .A2(new_n790), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT56), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n827), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n809), .A2(new_n572), .ZN(new_n832));
  AOI21_X1  g631(.A(G134gat), .B1(new_n832), .B2(KEYINPUT56), .ZN(new_n833));
  NOR4_X1   g632(.A1(new_n808), .A2(KEYINPUT119), .A3(KEYINPUT56), .A4(new_n790), .ZN(new_n834));
  INV_X1    g633(.A(new_n834), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  NOR2_X1   g635(.A1(new_n828), .A2(new_n829), .ZN(new_n837));
  OAI22_X1  g636(.A1(new_n830), .A2(new_n834), .B1(new_n837), .B2(G134gat), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n836), .A2(new_n838), .ZN(G1343gat));
  AND2_X1   g638(.A1(new_n805), .A2(new_n629), .ZN(new_n840));
  NOR3_X1   g639(.A1(new_n638), .A2(new_n408), .A3(new_n341), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  INV_X1    g641(.A(new_n842), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n524), .A2(G141gat), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT58), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT57), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n847), .B(new_n392), .C1(new_n803), .C2(new_n804), .ZN(new_n848));
  NOR3_X1   g647(.A1(new_n638), .A2(new_n264), .A3(new_n341), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n796), .B1(new_n522), .B2(new_n523), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n572), .B1(new_n850), .B2(new_n773), .ZN(new_n851));
  NOR2_X1   g650(.A1(new_n800), .A2(new_n801), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n604), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n804), .B1(new_n853), .B2(KEYINPUT120), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n855));
  OAI211_X1 g654(.A(new_n855), .B(new_n604), .C1(new_n851), .C2(new_n852), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n408), .B1(new_n854), .B2(new_n856), .ZN(new_n857));
  OAI211_X1 g656(.A(new_n848), .B(new_n849), .C1(new_n857), .C2(new_n847), .ZN(new_n858));
  OAI21_X1  g657(.A(G141gat), .B1(new_n858), .B2(new_n524), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n845), .A2(new_n846), .A3(new_n859), .ZN(new_n860));
  OR2_X1    g659(.A1(new_n857), .A2(new_n847), .ZN(new_n861));
  AND2_X1   g660(.A1(new_n848), .A2(new_n849), .ZN(new_n862));
  NAND3_X1  g661(.A1(new_n861), .A2(new_n698), .A3(new_n862), .ZN(new_n863));
  AOI22_X1  g662(.A1(new_n863), .A2(G141gat), .B1(new_n843), .B2(new_n844), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n860), .B1(new_n864), .B2(new_n846), .ZN(G1344gat));
  INV_X1    g664(.A(G148gat), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n843), .A2(new_n866), .A3(new_n623), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n408), .A2(KEYINPUT57), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n605), .A2(new_n524), .A3(new_n624), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n869), .B1(new_n853), .B2(new_n870), .ZN(new_n871));
  OAI21_X1  g670(.A(new_n392), .B1(new_n803), .B2(new_n804), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n871), .B1(new_n872), .B2(KEYINPUT57), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n849), .A2(new_n623), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n866), .B1(new_n873), .B2(new_n875), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT59), .ZN(new_n877));
  OAI21_X1  g676(.A(KEYINPUT122), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n866), .A2(KEYINPUT59), .ZN(new_n879));
  OAI211_X1 g678(.A(KEYINPUT121), .B(new_n879), .C1(new_n858), .C2(new_n624), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT122), .ZN(new_n881));
  AOI211_X1 g680(.A(new_n871), .B(new_n874), .C1(new_n872), .C2(KEYINPUT57), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n881), .B(KEYINPUT59), .C1(new_n882), .C2(new_n866), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n861), .A2(new_n623), .A3(new_n862), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT121), .B1(new_n885), .B2(new_n879), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n867), .B1(new_n884), .B2(new_n886), .ZN(G1345gat));
  OAI21_X1  g686(.A(G155gat), .B1(new_n858), .B2(new_n604), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n658), .A2(new_n205), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n888), .B1(new_n842), .B2(new_n889), .ZN(G1346gat));
  NOR3_X1   g689(.A1(new_n858), .A2(new_n206), .A3(new_n790), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n843), .A2(new_n572), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(new_n206), .ZN(G1347gat));
  AND2_X1   g692(.A1(new_n805), .A2(new_n264), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n806), .A2(new_n342), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NOR3_X1   g695(.A1(new_n896), .A2(new_n275), .A3(new_n524), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n894), .A2(new_n698), .A3(new_n895), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n897), .B1(new_n275), .B2(new_n898), .ZN(G1348gat));
  NOR2_X1   g698(.A1(new_n896), .A2(new_n624), .ZN(new_n900));
  XNOR2_X1  g699(.A(new_n900), .B(new_n276), .ZN(G1349gat));
  NAND4_X1  g700(.A1(new_n805), .A2(new_n895), .A3(new_n264), .A4(new_n658), .ZN(new_n902));
  OR3_X1    g701(.A1(new_n902), .A2(KEYINPUT123), .A3(new_n303), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n303), .ZN(new_n904));
  AOI21_X1  g703(.A(KEYINPUT123), .B1(new_n902), .B2(G183gat), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n903), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(KEYINPUT60), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n908));
  OAI211_X1 g707(.A(new_n903), .B(new_n908), .C1(new_n904), .C2(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(G1350gat));
  NOR2_X1   g709(.A1(new_n896), .A2(new_n790), .ZN(new_n911));
  NAND2_X1  g710(.A1(KEYINPUT61), .A2(G190gat), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  XOR2_X1   g712(.A(KEYINPUT61), .B(G190gat), .Z(new_n914));
  OAI21_X1  g713(.A(new_n913), .B1(new_n911), .B2(new_n914), .ZN(G1351gat));
  INV_X1    g714(.A(G197gat), .ZN(new_n916));
  NOR3_X1   g715(.A1(new_n638), .A2(new_n629), .A3(new_n342), .ZN(new_n917));
  XNOR2_X1  g716(.A(new_n917), .B(KEYINPUT124), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n873), .A2(new_n525), .A3(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n916), .B1(new_n919), .B2(KEYINPUT125), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n920), .B1(KEYINPUT125), .B2(new_n919), .ZN(new_n921));
  NOR3_X1   g720(.A1(new_n638), .A2(new_n408), .A3(new_n342), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n894), .A2(new_n922), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  NAND3_X1  g723(.A1(new_n924), .A2(new_n916), .A3(new_n698), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n921), .A2(new_n925), .ZN(G1352gat));
  NAND3_X1  g725(.A1(new_n873), .A2(new_n623), .A3(new_n918), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G204gat), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n624), .A2(G204gat), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n894), .A2(new_n922), .A3(new_n929), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n930), .A2(KEYINPUT62), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT126), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n930), .A2(KEYINPUT126), .A3(KEYINPUT62), .ZN(new_n935));
  OAI211_X1 g734(.A(new_n928), .B(new_n931), .C1(new_n934), .C2(new_n935), .ZN(G1353gat));
  NAND3_X1  g735(.A1(new_n924), .A2(new_n266), .A3(new_n658), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n873), .A2(new_n658), .A3(new_n917), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n938), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT63), .B1(new_n938), .B2(G211gat), .ZN(new_n940));
  OAI21_X1  g739(.A(new_n937), .B1(new_n939), .B2(new_n940), .ZN(G1354gat));
  OAI21_X1  g740(.A(new_n267), .B1(new_n923), .B2(new_n790), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(KEYINPUT127), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT127), .ZN(new_n944));
  OAI211_X1 g743(.A(new_n944), .B(new_n267), .C1(new_n923), .C2(new_n790), .ZN(new_n945));
  NAND4_X1  g744(.A1(new_n873), .A2(G218gat), .A3(new_n572), .A4(new_n918), .ZN(new_n946));
  AND3_X1   g745(.A1(new_n943), .A2(new_n945), .A3(new_n946), .ZN(G1355gat));
endmodule


