//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 1 1 0 0 1 0 0 0 0 0 0 1 0 0 0 1 1 0 0 0 1 0 1 1 1 1 1 1 0 1 1 1 0 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:33:34 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n494, new_n495, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n515, new_n516, new_n517, new_n518, new_n519,
    new_n520, new_n523, new_n524, new_n525, new_n526, new_n527, new_n528,
    new_n529, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n541, new_n543, new_n544, new_n546, new_n547,
    new_n548, new_n549, new_n550, new_n551, new_n552, new_n553, new_n554,
    new_n555, new_n556, new_n557, new_n558, new_n559, new_n560, new_n562,
    new_n563, new_n564, new_n565, new_n567, new_n568, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n621, new_n624, new_n626,
    new_n627, new_n628, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  XNOR2_X1  g016(.A(KEYINPUT65), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(KEYINPUT66), .ZN(new_n459));
  INV_X1    g034(.A(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(KEYINPUT3), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n461), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G125), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n459), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G113), .A2(G2104), .ZN(new_n467));
  XNOR2_X1  g042(.A(KEYINPUT3), .B(G2104), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT66), .A3(G125), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n466), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(G2105), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n460), .A2(G2105), .ZN(new_n473));
  AOI22_X1  g048(.A1(new_n472), .A2(G137), .B1(G101), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n471), .A2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(new_n475), .ZN(G160));
  NAND2_X1  g051(.A1(new_n472), .A2(G136), .ZN(new_n477));
  OAI21_X1  g052(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n478));
  INV_X1    g053(.A(G2105), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n479), .A2(G112), .ZN(new_n480));
  OAI21_X1  g055(.A(new_n477), .B1(new_n478), .B2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n464), .A2(new_n479), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G124), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT67), .ZN(G162));
  NAND3_X1  g059(.A1(new_n468), .A2(G126), .A3(G2105), .ZN(new_n485));
  OR2_X1    g060(.A1(G102), .A2(G2105), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G114), .C2(new_n479), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND4_X1  g063(.A1(new_n461), .A2(new_n463), .A3(G138), .A4(new_n479), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n468), .A2(new_n491), .A3(G138), .A4(new_n479), .ZN(new_n492));
  AOI21_X1  g067(.A(new_n488), .B1(new_n490), .B2(new_n492), .ZN(G164));
  INV_X1    g068(.A(KEYINPUT5), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n494), .A2(G543), .ZN(new_n495));
  INV_X1    g070(.A(G543), .ZN(new_n496));
  OAI21_X1  g071(.A(KEYINPUT68), .B1(new_n496), .B2(KEYINPUT5), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT68), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n498), .A2(new_n494), .A3(G543), .ZN(new_n499));
  AOI21_X1  g074(.A(new_n495), .B1(new_n497), .B2(new_n499), .ZN(new_n500));
  AOI22_X1  g075(.A1(new_n500), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  OR3_X1    g077(.A1(new_n501), .A2(KEYINPUT69), .A3(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n497), .A2(new_n499), .ZN(new_n504));
  XNOR2_X1  g079(.A(KEYINPUT6), .B(G651), .ZN(new_n505));
  INV_X1    g080(.A(new_n495), .ZN(new_n506));
  NAND3_X1  g081(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n505), .A2(G543), .ZN(new_n509));
  INV_X1    g084(.A(new_n509), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n508), .A2(G88), .B1(G50), .B2(new_n510), .ZN(new_n511));
  OAI21_X1  g086(.A(KEYINPUT69), .B1(new_n501), .B2(new_n502), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n503), .A2(new_n511), .A3(new_n512), .ZN(G303));
  INV_X1    g088(.A(G303), .ZN(G166));
  NAND2_X1  g089(.A1(new_n508), .A2(G89), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n510), .A2(G51), .ZN(new_n516));
  NAND3_X1  g091(.A1(new_n500), .A2(G63), .A3(G651), .ZN(new_n517));
  XOR2_X1   g092(.A(KEYINPUT70), .B(KEYINPUT7), .Z(new_n518));
  NAND3_X1  g093(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n519));
  XNOR2_X1  g094(.A(new_n518), .B(new_n519), .ZN(new_n520));
  NAND4_X1  g095(.A1(new_n515), .A2(new_n516), .A3(new_n517), .A4(new_n520), .ZN(G286));
  INV_X1    g096(.A(G286), .ZN(G168));
  AND2_X1   g097(.A1(new_n500), .A2(G64), .ZN(new_n523));
  AND2_X1   g098(.A1(G77), .A2(G543), .ZN(new_n524));
  OAI211_X1 g099(.A(KEYINPUT71), .B(G651), .C1(new_n523), .C2(new_n524), .ZN(new_n525));
  AOI22_X1  g100(.A1(new_n508), .A2(G90), .B1(G52), .B2(new_n510), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT71), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n524), .B1(new_n500), .B2(G64), .ZN(new_n528));
  OAI21_X1  g103(.A(new_n527), .B1(new_n528), .B2(new_n502), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n525), .A2(new_n526), .A3(new_n529), .ZN(G301));
  INV_X1    g105(.A(G301), .ZN(G171));
  NAND2_X1  g106(.A1(new_n508), .A2(G81), .ZN(new_n532));
  XOR2_X1   g107(.A(KEYINPUT73), .B(G43), .Z(new_n533));
  NAND2_X1  g108(.A1(new_n510), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n500), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  INV_X1    g111(.A(KEYINPUT72), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n536), .B(new_n537), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n538), .B2(G651), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(G860), .ZN(G153));
  AND3_X1   g115(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(G36), .ZN(G176));
  NAND2_X1  g117(.A1(G1), .A2(G3), .ZN(new_n543));
  XNOR2_X1  g118(.A(new_n543), .B(KEYINPUT8), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n541), .A2(new_n544), .ZN(G188));
  INV_X1    g120(.A(G91), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n507), .A2(KEYINPUT76), .ZN(new_n547));
  INV_X1    g122(.A(KEYINPUT76), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n500), .A2(new_n548), .A3(new_n505), .ZN(new_n549));
  AOI21_X1  g124(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  INV_X1    g125(.A(KEYINPUT74), .ZN(new_n551));
  NAND4_X1  g126(.A1(new_n551), .A2(KEYINPUT75), .A3(KEYINPUT9), .A4(G53), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n509), .A2(new_n552), .ZN(new_n553));
  NOR2_X1   g128(.A1(new_n550), .A2(new_n553), .ZN(new_n554));
  AOI22_X1  g129(.A1(new_n500), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n555), .A2(new_n502), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n551), .A2(KEYINPUT9), .ZN(new_n558));
  OAI21_X1  g133(.A(G53), .B1(KEYINPUT75), .B2(KEYINPUT9), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n509), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n554), .A2(new_n557), .A3(new_n560), .ZN(G299));
  NAND2_X1  g136(.A1(new_n547), .A2(new_n549), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G87), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n500), .B2(G74), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n510), .A2(G49), .ZN(new_n565));
  NAND3_X1  g140(.A1(new_n563), .A2(new_n564), .A3(new_n565), .ZN(G288));
  INV_X1    g141(.A(KEYINPUT80), .ZN(new_n567));
  AOI21_X1  g142(.A(KEYINPUT79), .B1(new_n562), .B2(G86), .ZN(new_n568));
  INV_X1    g143(.A(KEYINPUT79), .ZN(new_n569));
  INV_X1    g144(.A(G86), .ZN(new_n570));
  AOI211_X1 g145(.A(new_n569), .B(new_n570), .C1(new_n547), .C2(new_n549), .ZN(new_n571));
  INV_X1    g146(.A(G48), .ZN(new_n572));
  OAI22_X1  g147(.A1(new_n568), .A2(new_n571), .B1(new_n572), .B2(new_n509), .ZN(new_n573));
  INV_X1    g148(.A(KEYINPUT78), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT77), .ZN(new_n575));
  AOI21_X1  g150(.A(new_n498), .B1(new_n494), .B2(G543), .ZN(new_n576));
  NOR3_X1   g151(.A1(new_n496), .A2(KEYINPUT68), .A3(KEYINPUT5), .ZN(new_n577));
  OAI211_X1 g152(.A(G61), .B(new_n506), .C1(new_n576), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n575), .B1(new_n580), .B2(G651), .ZN(new_n581));
  AOI211_X1 g156(.A(KEYINPUT77), .B(new_n502), .C1(new_n578), .C2(new_n579), .ZN(new_n582));
  OAI21_X1  g157(.A(new_n574), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  INV_X1    g158(.A(new_n579), .ZN(new_n584));
  AOI21_X1  g159(.A(new_n584), .B1(new_n500), .B2(G61), .ZN(new_n585));
  OAI21_X1  g160(.A(KEYINPUT77), .B1(new_n585), .B2(new_n502), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n580), .A2(new_n575), .A3(G651), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT78), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n567), .B1(new_n573), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n509), .A2(new_n572), .ZN(new_n591));
  AND4_X1   g166(.A1(new_n548), .A2(new_n504), .A3(new_n505), .A4(new_n506), .ZN(new_n592));
  AOI21_X1  g167(.A(new_n548), .B1(new_n500), .B2(new_n505), .ZN(new_n593));
  OAI21_X1  g168(.A(G86), .B1(new_n592), .B2(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(new_n569), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n562), .A2(KEYINPUT79), .A3(G86), .ZN(new_n596));
  AOI21_X1  g171(.A(new_n591), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n597), .A2(KEYINPUT80), .A3(new_n583), .A4(new_n588), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n590), .A2(new_n598), .ZN(G305));
  AOI22_X1  g174(.A1(new_n500), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n600));
  NOR2_X1   g175(.A1(new_n600), .A2(new_n502), .ZN(new_n601));
  INV_X1    g176(.A(G85), .ZN(new_n602));
  INV_X1    g177(.A(G47), .ZN(new_n603));
  OAI22_X1  g178(.A1(new_n507), .A2(new_n602), .B1(new_n603), .B2(new_n509), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n601), .A2(new_n604), .ZN(G290));
  NAND2_X1  g180(.A1(G301), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(G92), .B1(new_n592), .B2(new_n593), .ZN(new_n607));
  NAND2_X1  g182(.A1(new_n607), .A2(KEYINPUT10), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n500), .A2(G66), .ZN(new_n609));
  INV_X1    g184(.A(G79), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(new_n496), .ZN(new_n611));
  AOI22_X1  g186(.A1(new_n611), .A2(G651), .B1(G54), .B2(new_n510), .ZN(new_n612));
  INV_X1    g187(.A(KEYINPUT10), .ZN(new_n613));
  NAND3_X1  g188(.A1(new_n562), .A2(new_n613), .A3(G92), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n608), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  INV_X1    g190(.A(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n606), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(new_n560), .ZN(new_n620));
  NOR4_X1   g195(.A1(new_n550), .A2(new_n556), .A3(new_n620), .A4(new_n553), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n619), .B1(new_n621), .B2(G868), .ZN(G297));
  OAI21_X1  g197(.A(new_n619), .B1(new_n621), .B2(G868), .ZN(G280));
  XNOR2_X1  g198(.A(KEYINPUT81), .B(G559), .ZN(new_n624));
  OAI21_X1  g199(.A(new_n616), .B1(G860), .B2(new_n624), .ZN(G148));
  OAI21_X1  g200(.A(KEYINPUT82), .B1(new_n539), .B2(G868), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n616), .A2(new_n624), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n627), .A2(G868), .ZN(new_n628));
  MUX2_X1   g203(.A(KEYINPUT82), .B(new_n626), .S(new_n628), .Z(G323));
  XNOR2_X1  g204(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g205(.A1(new_n468), .A2(new_n473), .ZN(new_n631));
  XOR2_X1   g206(.A(new_n631), .B(KEYINPUT12), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT13), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT83), .B(G2100), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n482), .A2(G123), .ZN(new_n636));
  NAND2_X1  g211(.A1(new_n472), .A2(G135), .ZN(new_n637));
  OR2_X1    g212(.A1(G99), .A2(G2105), .ZN(new_n638));
  OAI211_X1 g213(.A(new_n638), .B(G2104), .C1(G111), .C2(new_n479), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n636), .A2(new_n637), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2096), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n635), .A2(new_n641), .ZN(G156));
  XNOR2_X1  g217(.A(KEYINPUT15), .B(G2435), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2438), .ZN(new_n644));
  XOR2_X1   g219(.A(G2427), .B(G2430), .Z(new_n645));
  XNOR2_X1  g220(.A(new_n644), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT84), .B(KEYINPUT14), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2443), .B(G2446), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n648), .B(new_n649), .ZN(new_n650));
  XOR2_X1   g225(.A(G1341), .B(G1348), .Z(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT16), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n650), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G2451), .B(G2454), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n653), .B(new_n654), .ZN(new_n655));
  NAND2_X1  g230(.A1(new_n655), .A2(G14), .ZN(new_n656));
  INV_X1    g231(.A(new_n656), .ZN(G401));
  XOR2_X1   g232(.A(G2067), .B(G2678), .Z(new_n658));
  XNOR2_X1  g233(.A(new_n658), .B(KEYINPUT85), .ZN(new_n659));
  XOR2_X1   g234(.A(G2084), .B(G2090), .Z(new_n660));
  AND2_X1   g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2072), .B(G2078), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  XOR2_X1   g238(.A(new_n663), .B(KEYINPUT18), .Z(new_n664));
  OR2_X1    g239(.A1(new_n659), .A2(new_n660), .ZN(new_n665));
  AOI21_X1  g240(.A(new_n662), .B1(new_n665), .B2(KEYINPUT17), .ZN(new_n666));
  OR2_X1    g241(.A1(new_n666), .A2(new_n661), .ZN(new_n667));
  AND3_X1   g242(.A1(new_n665), .A2(KEYINPUT17), .A3(new_n662), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n664), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(G2096), .B(G2100), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n669), .B(new_n670), .ZN(new_n671));
  INV_X1    g246(.A(new_n671), .ZN(G227));
  XNOR2_X1  g247(.A(G1971), .B(G1976), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n673), .B(KEYINPUT19), .ZN(new_n674));
  XOR2_X1   g249(.A(G1956), .B(G2474), .Z(new_n675));
  XOR2_X1   g250(.A(G1961), .B(G1966), .Z(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT86), .ZN(new_n679));
  XOR2_X1   g254(.A(new_n679), .B(KEYINPUT20), .Z(new_n680));
  NOR2_X1   g255(.A1(new_n675), .A2(new_n676), .ZN(new_n681));
  INV_X1    g256(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n682), .A2(new_n674), .A3(new_n677), .ZN(new_n683));
  OAI211_X1 g258(.A(new_n680), .B(new_n683), .C1(new_n674), .C2(new_n682), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1991), .B(G1996), .ZN(new_n687));
  INV_X1    g262(.A(G1981), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n687), .B(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n686), .B(new_n690), .ZN(new_n691));
  INV_X1    g266(.A(new_n691), .ZN(G229));
  INV_X1    g267(.A(KEYINPUT91), .ZN(new_n693));
  NOR2_X1   g268(.A1(new_n693), .A2(KEYINPUT36), .ZN(new_n694));
  MUX2_X1   g269(.A(G6), .B(G305), .S(G16), .Z(new_n695));
  XOR2_X1   g270(.A(KEYINPUT32), .B(G1981), .Z(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(new_n697));
  OR2_X1    g272(.A1(new_n695), .A2(new_n697), .ZN(new_n698));
  INV_X1    g273(.A(G16), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n699), .A2(G22), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n700), .B1(G166), .B2(new_n699), .ZN(new_n701));
  XOR2_X1   g276(.A(new_n701), .B(G1971), .Z(new_n702));
  NAND2_X1  g277(.A1(new_n695), .A2(new_n697), .ZN(new_n703));
  AND2_X1   g278(.A1(new_n699), .A2(G23), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n704), .B1(G288), .B2(G16), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT33), .ZN(new_n706));
  INV_X1    g281(.A(G1976), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND4_X1  g283(.A1(new_n698), .A2(new_n702), .A3(new_n703), .A4(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT34), .ZN(new_n710));
  OR2_X1    g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n709), .A2(new_n710), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(G24), .ZN(new_n714));
  OAI21_X1  g289(.A(KEYINPUT88), .B1(new_n714), .B2(G16), .ZN(new_n715));
  OR3_X1    g290(.A1(new_n714), .A2(KEYINPUT88), .A3(G16), .ZN(new_n716));
  INV_X1    g291(.A(G290), .ZN(new_n717));
  OAI211_X1 g292(.A(new_n715), .B(new_n716), .C1(new_n717), .C2(new_n699), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT90), .ZN(new_n719));
  XNOR2_X1  g294(.A(KEYINPUT89), .B(G1986), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n482), .A2(G119), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n472), .A2(G131), .ZN(new_n723));
  OAI21_X1  g298(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n479), .A2(G107), .ZN(new_n725));
  OAI211_X1 g300(.A(new_n722), .B(new_n723), .C1(new_n724), .C2(new_n725), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT87), .B(G29), .ZN(new_n727));
  MUX2_X1   g302(.A(G25), .B(new_n726), .S(new_n727), .Z(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT35), .B(G1991), .ZN(new_n729));
  XOR2_X1   g304(.A(new_n728), .B(new_n729), .Z(new_n730));
  INV_X1    g305(.A(KEYINPUT36), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n730), .B1(KEYINPUT91), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(new_n721), .A2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n694), .B1(new_n713), .B2(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n734), .B1(new_n711), .B2(new_n712), .ZN(new_n736));
  INV_X1    g311(.A(new_n694), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(G171), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G1961), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  INV_X1    g317(.A(G29), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G32), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n472), .A2(G141), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n473), .A2(G105), .ZN(new_n746));
  NAND3_X1  g321(.A1(new_n468), .A2(G129), .A3(G2105), .ZN(new_n747));
  NAND3_X1  g322(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n748));
  XOR2_X1   g323(.A(new_n748), .B(KEYINPUT26), .Z(new_n749));
  NAND4_X1  g324(.A1(new_n745), .A2(new_n746), .A3(new_n747), .A4(new_n749), .ZN(new_n750));
  INV_X1    g325(.A(KEYINPUT95), .ZN(new_n751));
  XNOR2_X1  g326(.A(new_n750), .B(new_n751), .ZN(new_n752));
  OAI21_X1  g327(.A(new_n744), .B1(new_n752), .B2(new_n743), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT27), .B(G1996), .Z(new_n754));
  NOR2_X1   g329(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT96), .Z(new_n756));
  NAND2_X1  g331(.A1(G115), .A2(G2104), .ZN(new_n757));
  INV_X1    g332(.A(G127), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n757), .B1(new_n464), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n759), .A2(G2105), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n760), .A2(KEYINPUT93), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT93), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n759), .A2(new_n762), .A3(G2105), .ZN(new_n763));
  AOI22_X1  g338(.A1(new_n761), .A2(new_n763), .B1(G139), .B2(new_n472), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n473), .A2(G103), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(KEYINPUT25), .Z(new_n766));
  NAND2_X1  g341(.A1(new_n764), .A2(new_n766), .ZN(new_n767));
  MUX2_X1   g342(.A(G33), .B(new_n767), .S(G29), .Z(new_n768));
  XOR2_X1   g343(.A(new_n768), .B(G2072), .Z(new_n769));
  INV_X1    g344(.A(G2084), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT94), .B(KEYINPUT24), .Z(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G34), .ZN(new_n772));
  OAI22_X1  g347(.A1(new_n475), .A2(new_n743), .B1(new_n727), .B2(new_n772), .ZN(new_n773));
  OAI211_X1 g348(.A(new_n756), .B(new_n769), .C1(new_n770), .C2(new_n773), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(KEYINPUT97), .ZN(new_n775));
  NOR2_X1   g350(.A1(new_n740), .A2(new_n741), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(KEYINPUT100), .ZN(new_n777));
  NAND3_X1  g352(.A1(new_n699), .A2(KEYINPUT23), .A3(G20), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT23), .ZN(new_n779));
  INV_X1    g354(.A(G20), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n779), .B1(new_n780), .B2(G16), .ZN(new_n781));
  OAI211_X1 g356(.A(new_n778), .B(new_n781), .C1(new_n621), .C2(new_n699), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1956), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n699), .A2(G4), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(new_n616), .B2(new_n699), .ZN(new_n786));
  INV_X1    g361(.A(G1348), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n784), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n699), .A2(G19), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n539), .B2(new_n699), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n791), .B(G1341), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n699), .A2(G21), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(G168), .B2(new_n699), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(G1966), .ZN(new_n795));
  OR2_X1    g370(.A1(new_n792), .A2(new_n795), .ZN(new_n796));
  INV_X1    g371(.A(new_n727), .ZN(new_n797));
  NAND3_X1  g372(.A1(new_n797), .A2(KEYINPUT28), .A3(G26), .ZN(new_n798));
  NAND2_X1  g373(.A1(new_n482), .A2(G128), .ZN(new_n799));
  XNOR2_X1  g374(.A(new_n799), .B(KEYINPUT92), .ZN(new_n800));
  NAND2_X1  g375(.A1(new_n472), .A2(G140), .ZN(new_n801));
  OAI21_X1  g376(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n479), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n801), .B1(new_n802), .B2(new_n803), .ZN(new_n804));
  NOR2_X1   g379(.A1(new_n800), .A2(new_n804), .ZN(new_n805));
  OAI21_X1  g380(.A(new_n798), .B1(new_n805), .B2(new_n743), .ZN(new_n806));
  AOI21_X1  g381(.A(KEYINPUT28), .B1(new_n797), .B2(G26), .ZN(new_n807));
  NOR2_X1   g382(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2067), .ZN(new_n809));
  XOR2_X1   g384(.A(KEYINPUT99), .B(KEYINPUT30), .Z(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(G28), .ZN(new_n811));
  AOI22_X1  g386(.A1(new_n753), .A2(new_n754), .B1(new_n743), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g387(.A1(new_n797), .A2(G27), .ZN(new_n813));
  OAI21_X1  g388(.A(new_n813), .B1(G164), .B2(new_n797), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(G2078), .Z(new_n815));
  NOR2_X1   g390(.A1(new_n640), .A2(new_n797), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n816), .B1(new_n773), .B2(new_n770), .ZN(new_n817));
  NAND4_X1  g392(.A1(new_n809), .A2(new_n812), .A3(new_n815), .A4(new_n817), .ZN(new_n818));
  NOR4_X1   g393(.A1(new_n775), .A2(new_n789), .A3(new_n796), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g394(.A1(new_n735), .A2(new_n738), .A3(new_n742), .A4(new_n819), .ZN(new_n820));
  XNOR2_X1  g395(.A(KEYINPUT98), .B(KEYINPUT31), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(G11), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n797), .A2(G35), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n823), .B1(G162), .B2(new_n797), .ZN(new_n824));
  XNOR2_X1  g399(.A(KEYINPUT29), .B(G2090), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n824), .B(new_n825), .ZN(new_n826));
  NOR3_X1   g401(.A1(new_n820), .A2(new_n822), .A3(new_n826), .ZN(G311));
  INV_X1    g402(.A(new_n738), .ZN(new_n828));
  OAI21_X1  g403(.A(new_n819), .B1(new_n736), .B2(new_n737), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n822), .ZN(new_n831));
  INV_X1    g406(.A(new_n826), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n830), .A2(new_n831), .A3(new_n832), .A4(new_n742), .ZN(G150));
  AOI22_X1  g408(.A1(new_n508), .A2(G93), .B1(G55), .B2(new_n510), .ZN(new_n834));
  AND3_X1   g409(.A1(new_n504), .A2(G67), .A3(new_n506), .ZN(new_n835));
  AND2_X1   g410(.A1(G80), .A2(G543), .ZN(new_n836));
  OAI211_X1 g411(.A(KEYINPUT101), .B(G651), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  INV_X1    g412(.A(KEYINPUT101), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n836), .B1(new_n500), .B2(G67), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n838), .B1(new_n839), .B2(new_n502), .ZN(new_n840));
  NAND3_X1  g415(.A1(new_n834), .A2(new_n837), .A3(new_n840), .ZN(new_n841));
  INV_X1    g416(.A(KEYINPUT102), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND4_X1  g418(.A1(new_n834), .A2(new_n837), .A3(new_n840), .A4(KEYINPUT102), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(G860), .A3(new_n844), .ZN(new_n845));
  XOR2_X1   g420(.A(new_n845), .B(KEYINPUT37), .Z(new_n846));
  NAND2_X1  g421(.A1(new_n843), .A2(new_n844), .ZN(new_n847));
  INV_X1    g422(.A(new_n539), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n539), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n851), .B(KEYINPUT39), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n616), .A2(G559), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(KEYINPUT38), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n852), .B(new_n854), .ZN(new_n855));
  OAI21_X1  g430(.A(new_n846), .B1(new_n855), .B2(G860), .ZN(G145));
  NAND2_X1  g431(.A1(new_n482), .A2(G130), .ZN(new_n857));
  NAND2_X1  g432(.A1(new_n472), .A2(G142), .ZN(new_n858));
  OAI21_X1  g433(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n859));
  NOR2_X1   g434(.A1(new_n479), .A2(G118), .ZN(new_n860));
  OAI211_X1 g435(.A(new_n857), .B(new_n858), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  XOR2_X1   g436(.A(new_n805), .B(new_n861), .Z(new_n862));
  INV_X1    g437(.A(new_n862), .ZN(new_n863));
  XNOR2_X1  g438(.A(new_n750), .B(KEYINPUT95), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n767), .ZN(new_n865));
  INV_X1    g440(.A(new_n750), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n866), .B1(new_n764), .B2(new_n766), .ZN(new_n867));
  OAI21_X1  g442(.A(new_n632), .B1(new_n865), .B2(new_n867), .ZN(new_n868));
  NAND3_X1  g443(.A1(new_n752), .A2(new_n764), .A3(new_n766), .ZN(new_n869));
  INV_X1    g444(.A(new_n867), .ZN(new_n870));
  INV_X1    g445(.A(new_n632), .ZN(new_n871));
  NAND3_X1  g446(.A1(new_n869), .A2(new_n870), .A3(new_n871), .ZN(new_n872));
  XOR2_X1   g447(.A(G164), .B(new_n726), .Z(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n868), .A2(new_n872), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n875), .ZN(new_n876));
  AOI21_X1  g451(.A(new_n874), .B1(new_n868), .B2(new_n872), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n863), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n475), .B(new_n640), .ZN(new_n879));
  XNOR2_X1  g454(.A(G162), .B(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n868), .A2(new_n872), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n873), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n882), .A2(new_n862), .A3(new_n875), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n878), .A2(new_n880), .A3(new_n883), .ZN(new_n884));
  INV_X1    g459(.A(G37), .ZN(new_n885));
  AND2_X1   g460(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n880), .ZN(new_n887));
  NOR3_X1   g462(.A1(new_n876), .A2(new_n863), .A3(new_n877), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n862), .B1(new_n882), .B2(new_n875), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n890), .A2(KEYINPUT103), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT103), .ZN(new_n892));
  OAI211_X1 g467(.A(new_n892), .B(new_n887), .C1(new_n888), .C2(new_n889), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n886), .A2(new_n891), .A3(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n894), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n896));
  XNOR2_X1  g471(.A(G288), .B(G290), .ZN(new_n897));
  INV_X1    g472(.A(new_n897), .ZN(new_n898));
  AND3_X1   g473(.A1(new_n590), .A2(G303), .A3(new_n598), .ZN(new_n899));
  AOI21_X1  g474(.A(G303), .B1(new_n590), .B2(new_n598), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n898), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NOR3_X1   g476(.A1(new_n573), .A2(new_n589), .A3(new_n567), .ZN(new_n902));
  AND3_X1   g477(.A1(new_n586), .A2(new_n587), .A3(KEYINPUT78), .ZN(new_n903));
  AOI21_X1  g478(.A(KEYINPUT78), .B1(new_n586), .B2(new_n587), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(KEYINPUT80), .B1(new_n905), .B2(new_n597), .ZN(new_n906));
  OAI21_X1  g481(.A(G166), .B1(new_n902), .B2(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n590), .A2(G303), .A3(new_n598), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n897), .A3(new_n908), .ZN(new_n909));
  AND3_X1   g484(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(KEYINPUT104), .B1(new_n901), .B2(new_n909), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(KEYINPUT42), .ZN(new_n913));
  NOR2_X1   g488(.A1(new_n912), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g489(.A(KEYINPUT42), .B1(new_n901), .B2(new_n909), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  XNOR2_X1  g491(.A(new_n851), .B(new_n627), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n616), .A2(G299), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n621), .A2(new_n615), .ZN(new_n919));
  NAND2_X1  g494(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g495(.A(new_n920), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n917), .A2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT41), .ZN(new_n923));
  INV_X1    g498(.A(new_n919), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n621), .A2(new_n615), .ZN(new_n925));
  OAI21_X1  g500(.A(new_n923), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n918), .A2(KEYINPUT41), .A3(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  AOI21_X1  g503(.A(new_n922), .B1(new_n917), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n916), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n929), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n931), .B1(new_n914), .B2(new_n915), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n933), .A2(G868), .ZN(new_n934));
  NOR2_X1   g509(.A1(new_n847), .A2(G868), .ZN(new_n935));
  INV_X1    g510(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n896), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(G868), .ZN(new_n938));
  AOI21_X1  g513(.A(new_n938), .B1(new_n930), .B2(new_n932), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n939), .A2(KEYINPUT105), .A3(new_n935), .ZN(new_n940));
  NOR2_X1   g515(.A1(new_n937), .A2(new_n940), .ZN(G295));
  NAND2_X1  g516(.A1(new_n934), .A2(new_n936), .ZN(G331));
  XNOR2_X1  g517(.A(G168), .B(G301), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n539), .B1(new_n843), .B2(new_n844), .ZN(new_n944));
  AND2_X1   g519(.A1(new_n539), .A2(new_n841), .ZN(new_n945));
  OAI21_X1  g520(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(G301), .B(G286), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n849), .A2(new_n850), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n946), .A2(new_n948), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n949), .A2(new_n928), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT107), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n946), .A2(new_n948), .A3(new_n920), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n950), .A2(new_n951), .A3(new_n952), .ZN(new_n953));
  AOI22_X1  g528(.A1(new_n948), .A2(new_n946), .B1(new_n926), .B2(new_n927), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT107), .ZN(new_n955));
  OAI211_X1 g530(.A(new_n953), .B(new_n955), .C1(new_n910), .C2(new_n911), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT43), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  NAND3_X1  g533(.A1(new_n949), .A2(new_n928), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n952), .A2(KEYINPUT106), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n959), .B1(new_n960), .B2(new_n954), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT104), .ZN(new_n962));
  NOR3_X1   g537(.A1(new_n899), .A2(new_n900), .A3(new_n898), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n897), .B1(new_n907), .B2(new_n908), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n962), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND3_X1  g540(.A1(new_n901), .A2(KEYINPUT104), .A3(new_n909), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n961), .A2(new_n965), .A3(new_n966), .ZN(new_n967));
  NAND4_X1  g542(.A1(new_n956), .A2(new_n957), .A3(new_n967), .A4(new_n885), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT108), .ZN(new_n969));
  AOI21_X1  g544(.A(G37), .B1(new_n912), .B2(new_n961), .ZN(new_n970));
  INV_X1    g545(.A(KEYINPUT108), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n970), .A2(new_n971), .A3(new_n957), .A4(new_n956), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n967), .A2(new_n885), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n961), .B1(new_n966), .B2(new_n965), .ZN(new_n974));
  OAI21_X1  g549(.A(KEYINPUT43), .B1(new_n973), .B2(new_n974), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n969), .A2(new_n972), .A3(new_n975), .ZN(new_n976));
  NAND3_X1  g551(.A1(new_n970), .A2(KEYINPUT43), .A3(new_n956), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n957), .B1(new_n973), .B2(new_n974), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  MUX2_X1   g554(.A(new_n976), .B(new_n979), .S(KEYINPUT44), .Z(G397));
  INV_X1    g555(.A(G2067), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n805), .B(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n488), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n490), .A2(new_n492), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  XNOR2_X1  g560(.A(KEYINPUT109), .B(KEYINPUT45), .ZN(new_n986));
  NOR2_X1   g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  AND3_X1   g562(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n982), .A2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n990), .A2(new_n750), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  XNOR2_X1  g568(.A(new_n993), .B(KEYINPUT125), .ZN(new_n994));
  NOR2_X1   g569(.A1(new_n989), .A2(G1996), .ZN(new_n995));
  XOR2_X1   g570(.A(new_n995), .B(KEYINPUT46), .Z(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT126), .B(KEYINPUT47), .ZN(new_n998));
  XNOR2_X1  g573(.A(new_n997), .B(new_n998), .ZN(new_n999));
  NOR3_X1   g574(.A1(new_n989), .A2(new_n864), .A3(G1996), .ZN(new_n1000));
  XNOR2_X1  g575(.A(new_n1000), .B(KEYINPUT112), .ZN(new_n1001));
  INV_X1    g576(.A(G1996), .ZN(new_n1002));
  OAI211_X1 g577(.A(new_n1001), .B(new_n991), .C1(new_n1002), .C2(new_n992), .ZN(new_n1003));
  XNOR2_X1  g578(.A(new_n1003), .B(KEYINPUT113), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n726), .A2(new_n729), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n805), .A2(new_n981), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n989), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n726), .A2(new_n729), .ZN(new_n1009));
  OAI21_X1  g584(.A(new_n990), .B1(new_n1009), .B2(new_n1005), .ZN(new_n1010));
  AND2_X1   g585(.A1(new_n1004), .A2(new_n1010), .ZN(new_n1011));
  NOR2_X1   g586(.A1(G290), .A2(G1986), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n990), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT48), .ZN(new_n1014));
  AOI211_X1 g589(.A(new_n999), .B(new_n1008), .C1(new_n1011), .C2(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT124), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n905), .A2(new_n688), .A3(new_n597), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n591), .B1(new_n508), .B2(G86), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n586), .A2(new_n1018), .A3(new_n587), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1019), .A2(G1981), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1017), .A2(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT49), .ZN(new_n1022));
  AOI21_X1  g597(.A(new_n1021), .B1(KEYINPUT115), .B2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n988), .A2(new_n985), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1024), .A2(G8), .ZN(new_n1025));
  XNOR2_X1  g600(.A(KEYINPUT115), .B(KEYINPUT49), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1017), .B2(new_n1020), .ZN(new_n1027));
  OR3_X1    g602(.A1(new_n1023), .A2(new_n1025), .A3(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(G288), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1025), .B1(G1976), .B2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT52), .ZN(new_n1031));
  OR2_X1    g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1030), .B(new_n1031), .C1(G1976), .C2(new_n1029), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1028), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT55), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1036), .A2(KEYINPUT117), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT114), .ZN(new_n1038));
  INV_X1    g613(.A(new_n986), .ZN(new_n1039));
  OAI211_X1 g614(.A(new_n1038), .B(new_n1039), .C1(G164), .C2(G1384), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1041));
  AND2_X1   g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n471), .A2(G40), .A3(new_n474), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n1039), .B1(G164), .B2(G1384), .ZN(new_n1044));
  AOI21_X1  g619(.A(new_n1043), .B1(new_n1044), .B2(KEYINPUT114), .ZN(new_n1045));
  AOI21_X1  g620(.A(G1971), .B1(new_n1042), .B2(new_n1045), .ZN(new_n1046));
  OAI21_X1  g621(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT50), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n985), .A2(new_n1048), .ZN(new_n1049));
  NAND3_X1  g624(.A1(new_n988), .A2(new_n1047), .A3(new_n1049), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1050), .A2(G2090), .ZN(new_n1051));
  OAI21_X1  g626(.A(G8), .B1(new_n1046), .B2(new_n1051), .ZN(new_n1052));
  OR2_X1    g627(.A1(new_n1037), .A2(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT45), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1054), .B1(G164), .B2(G1384), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n985), .A2(new_n986), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n988), .A2(new_n1055), .A3(new_n1056), .ZN(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1059), .A2(KEYINPUT116), .ZN(new_n1060));
  OR2_X1    g635(.A1(new_n1050), .A2(G2084), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT116), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1057), .A2(new_n1062), .A3(new_n1058), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n1060), .A2(new_n1061), .A3(new_n1063), .ZN(new_n1064));
  AND2_X1   g639(.A1(G168), .A2(G8), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1037), .A2(new_n1052), .ZN(new_n1066));
  NAND4_X1  g641(.A1(new_n1053), .A2(new_n1064), .A3(new_n1065), .A4(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(KEYINPUT63), .B1(new_n1034), .B2(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1052), .A2(new_n1036), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1028), .A2(new_n1069), .A3(new_n1032), .A4(new_n1033), .ZN(new_n1070));
  OAI21_X1  g645(.A(new_n707), .B1(new_n1023), .B2(new_n1027), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1017), .B1(new_n1071), .B2(G288), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(G8), .A3(new_n1024), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1068), .A2(new_n1070), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(G8), .B1(new_n1064), .B2(G286), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT51), .ZN(new_n1077));
  AOI21_X1  g652(.A(new_n1077), .B1(new_n1064), .B2(G286), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  INV_X1    g654(.A(KEYINPUT53), .ZN(new_n1080));
  OAI21_X1  g655(.A(KEYINPUT114), .B1(new_n985), .B2(new_n986), .ZN(new_n1081));
  NAND4_X1  g656(.A1(new_n1081), .A2(new_n1040), .A3(new_n988), .A4(new_n1041), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1080), .B1(new_n1082), .B2(G2078), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1050), .A2(new_n741), .ZN(new_n1084));
  NOR2_X1   g659(.A1(new_n1080), .A2(G2078), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n988), .A2(new_n1055), .A3(new_n1056), .A4(new_n1085), .ZN(new_n1086));
  NAND3_X1  g661(.A1(new_n1083), .A2(new_n1084), .A3(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1087), .A2(G171), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT121), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1087), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1076), .A2(KEYINPUT51), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1079), .A2(new_n1092), .A3(KEYINPUT62), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(KEYINPUT63), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  AOI21_X1  g672(.A(KEYINPUT62), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1098));
  INV_X1    g673(.A(new_n1098), .ZN(new_n1099));
  XNOR2_X1  g674(.A(KEYINPUT56), .B(G2072), .ZN(new_n1100));
  XOR2_X1   g675(.A(new_n1100), .B(KEYINPUT119), .Z(new_n1101));
  NAND3_X1  g676(.A1(new_n1042), .A2(new_n1045), .A3(new_n1101), .ZN(new_n1102));
  INV_X1    g677(.A(G1956), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1050), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(KEYINPUT118), .B(KEYINPUT57), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n621), .A2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(new_n1105), .ZN(new_n1107));
  NAND2_X1  g682(.A1(G299), .A2(new_n1107), .ZN(new_n1108));
  NAND4_X1  g683(.A1(new_n1102), .A2(new_n1104), .A3(new_n1106), .A4(new_n1108), .ZN(new_n1109));
  NAND2_X1  g684(.A1(new_n1050), .A2(new_n787), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1043), .A2(G1384), .A3(G164), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(new_n981), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1110), .A2(new_n1112), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n616), .A3(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1101), .ZN(new_n1115));
  OAI21_X1  g690(.A(new_n1104), .B1(new_n1082), .B2(new_n1115), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1108), .A2(new_n1106), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  XOR2_X1   g694(.A(KEYINPUT58), .B(G1341), .Z(new_n1120));
  NAND2_X1  g695(.A1(new_n1024), .A2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1121), .B1(new_n1082), .B2(G1996), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT120), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI211_X1 g699(.A(new_n1121), .B(KEYINPUT120), .C1(new_n1082), .C2(G1996), .ZN(new_n1125));
  NAND3_X1  g700(.A1(new_n1124), .A2(new_n539), .A3(new_n1125), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT59), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND4_X1  g703(.A1(new_n1124), .A2(KEYINPUT59), .A3(new_n539), .A4(new_n1125), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT60), .ZN(new_n1132));
  OAI21_X1  g707(.A(new_n616), .B1(new_n1113), .B2(new_n1132), .ZN(new_n1133));
  AOI22_X1  g708(.A1(new_n787), .A2(new_n1050), .B1(new_n1111), .B2(new_n981), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1134), .A2(KEYINPUT60), .A3(new_n615), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1133), .A2(new_n1135), .B1(new_n1132), .B2(new_n1113), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1118), .A2(new_n1109), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1137), .A2(KEYINPUT61), .ZN(new_n1138));
  INV_X1    g713(.A(KEYINPUT61), .ZN(new_n1139));
  NAND3_X1  g714(.A1(new_n1118), .A2(new_n1109), .A3(new_n1139), .ZN(new_n1140));
  AOI21_X1  g715(.A(new_n1136), .B1(new_n1138), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1119), .B1(new_n1131), .B2(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT54), .ZN(new_n1143));
  INV_X1    g718(.A(KEYINPUT122), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1084), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1050), .A2(KEYINPUT122), .A3(new_n741), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  XOR2_X1   g722(.A(new_n474), .B(KEYINPUT123), .Z(new_n1148));
  AND3_X1   g723(.A1(new_n1148), .A2(G40), .A3(new_n471), .ZN(new_n1149));
  NAND4_X1  g724(.A1(new_n1149), .A2(new_n1044), .A3(new_n1041), .A4(new_n1085), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1147), .A2(G301), .A3(new_n1083), .A4(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1090), .A2(new_n1143), .A3(new_n1091), .A4(new_n1151), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1143), .B1(new_n1087), .B2(G301), .ZN(new_n1153));
  NAND3_X1  g728(.A1(new_n1147), .A2(new_n1083), .A3(new_n1150), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1153), .B1(G301), .B2(new_n1154), .ZN(new_n1155));
  AND2_X1   g730(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(new_n1099), .B1(new_n1142), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1079), .A2(new_n1093), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1097), .B1(new_n1157), .B2(new_n1158), .ZN(new_n1159));
  AND2_X1   g734(.A1(new_n1052), .A2(new_n1036), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1034), .A2(new_n1160), .A3(new_n1069), .ZN(new_n1161));
  INV_X1    g736(.A(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n1075), .B1(new_n1159), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n1012), .ZN(new_n1164));
  INV_X1    g739(.A(KEYINPUT110), .ZN(new_n1165));
  NAND2_X1  g740(.A1(G290), .A2(G1986), .ZN(new_n1166));
  NAND3_X1  g741(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .ZN(new_n1167));
  OAI211_X1 g742(.A(new_n1167), .B(new_n990), .C1(new_n1165), .C2(new_n1166), .ZN(new_n1168));
  XOR2_X1   g743(.A(new_n1168), .B(KEYINPUT111), .Z(new_n1169));
  NAND2_X1  g744(.A1(new_n1011), .A2(new_n1169), .ZN(new_n1170));
  INV_X1    g745(.A(new_n1170), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1016), .B1(new_n1163), .B2(new_n1171), .ZN(new_n1172));
  AND2_X1   g747(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1119), .ZN(new_n1174));
  NOR3_X1   g749(.A1(new_n1113), .A2(new_n1132), .A3(new_n616), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n615), .B1(new_n1134), .B2(KEYINPUT60), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1175), .A2(new_n1176), .B1(KEYINPUT60), .B2(new_n1134), .ZN(new_n1177));
  AND3_X1   g752(.A1(new_n1118), .A2(new_n1109), .A3(new_n1139), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1139), .B1(new_n1118), .B2(new_n1109), .ZN(new_n1179));
  OAI21_X1  g754(.A(new_n1177), .B1(new_n1178), .B2(new_n1179), .ZN(new_n1180));
  OAI21_X1  g755(.A(new_n1174), .B1(new_n1180), .B2(new_n1130), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1152), .A2(new_n1155), .ZN(new_n1182));
  AOI21_X1  g757(.A(new_n1098), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1183));
  INV_X1    g758(.A(new_n1158), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1173), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g760(.A(new_n1074), .B1(new_n1185), .B2(new_n1161), .ZN(new_n1186));
  NOR3_X1   g761(.A1(new_n1186), .A2(KEYINPUT124), .A3(new_n1170), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1015), .B1(new_n1172), .B2(new_n1187), .ZN(G329));
  assign    G231 = 1'b0;
  AND4_X1   g763(.A1(G319), .A2(new_n894), .A3(new_n656), .A4(new_n671), .ZN(new_n1190));
  NAND3_X1  g764(.A1(new_n976), .A2(new_n691), .A3(new_n1190), .ZN(new_n1191));
  NAND2_X1  g765(.A1(new_n1191), .A2(KEYINPUT127), .ZN(new_n1192));
  INV_X1    g766(.A(KEYINPUT127), .ZN(new_n1193));
  NAND4_X1  g767(.A1(new_n976), .A2(new_n1190), .A3(new_n1193), .A4(new_n691), .ZN(new_n1194));
  AND2_X1   g768(.A1(new_n1192), .A2(new_n1194), .ZN(G308));
  NAND2_X1  g769(.A1(new_n1192), .A2(new_n1194), .ZN(G225));
endmodule


