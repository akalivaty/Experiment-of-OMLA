

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817;

  XNOR2_X1 U378 ( .A(n536), .B(n535), .ZN(n539) );
  BUF_X1 U379 ( .A(G128), .Z(n356) );
  XNOR2_X2 U380 ( .A(n609), .B(n393), .ZN(n731) );
  XNOR2_X1 U381 ( .A(n789), .B(n475), .ZN(n703) );
  AND2_X1 U382 ( .A1(n385), .A2(n481), .ZN(n429) );
  INV_X2 U383 ( .A(n489), .ZN(n784) );
  AND2_X2 U384 ( .A1(n376), .A2(n483), .ZN(n482) );
  NAND2_X2 U385 ( .A1(n429), .A2(n362), .ZN(n681) );
  XNOR2_X2 U386 ( .A(n478), .B(n477), .ZN(n789) );
  INV_X1 U387 ( .A(n693), .ZN(n357) );
  INV_X2 U388 ( .A(G953), .ZN(n792) );
  NAND2_X1 U389 ( .A1(n423), .A2(n422), .ZN(n421) );
  NOR2_X1 U390 ( .A1(n812), .A2(n817), .ZN(n616) );
  AND2_X1 U391 ( .A1(n748), .A2(n618), .ZN(n551) );
  XNOR2_X1 U392 ( .A(n618), .B(n617), .ZN(n662) );
  AND2_X1 U393 ( .A1(n508), .A2(n507), .ZN(n506) );
  NAND2_X2 U394 ( .A1(n439), .A2(n443), .ZN(n618) );
  XNOR2_X1 U395 ( .A(n780), .B(KEYINPUT122), .ZN(n781) );
  INV_X2 U396 ( .A(G128), .ZN(n518) );
  XNOR2_X2 U397 ( .A(n595), .B(n519), .ZN(n536) );
  XNOR2_X2 U398 ( .A(n518), .B(G143), .ZN(n595) );
  XNOR2_X2 U399 ( .A(n539), .B(n538), .ZN(n802) );
  XNOR2_X2 U400 ( .A(n391), .B(n558), .ZN(n774) );
  XNOR2_X2 U401 ( .A(n802), .B(G146), .ZN(n391) );
  NOR2_X1 U402 ( .A1(G953), .A2(G237), .ZN(n542) );
  XNOR2_X1 U403 ( .A(n614), .B(n613), .ZN(n615) );
  XOR2_X1 U404 ( .A(G131), .B(G140), .Z(n554) );
  XNOR2_X1 U405 ( .A(n525), .B(n596), .ZN(n569) );
  XNOR2_X1 U406 ( .A(n476), .B(n598), .ZN(n475) );
  AND2_X1 U407 ( .A1(n440), .A2(n442), .ZN(n439) );
  NAND2_X1 U408 ( .A1(G902), .A2(G472), .ZN(n442) );
  INV_X1 U409 ( .A(KEYINPUT64), .ZN(n691) );
  XNOR2_X1 U410 ( .A(n396), .B(KEYINPUT39), .ZN(n644) );
  NAND2_X1 U411 ( .A1(n395), .A2(n358), .ZN(n396) );
  INV_X1 U412 ( .A(KEYINPUT22), .ZN(n455) );
  XNOR2_X1 U413 ( .A(n660), .B(KEYINPUT103), .ZN(n661) );
  XNOR2_X1 U414 ( .A(n532), .B(n460), .ZN(n628) );
  XNOR2_X1 U415 ( .A(n531), .B(G475), .ZN(n460) );
  XNOR2_X1 U416 ( .A(n524), .B(n523), .ZN(n627) );
  NAND2_X1 U417 ( .A1(n470), .A2(n467), .ZN(n631) );
  AND2_X1 U418 ( .A1(n682), .A2(n469), .ZN(n467) );
  INV_X1 U419 ( .A(KEYINPUT47), .ZN(n496) );
  NOR2_X1 U420 ( .A1(n720), .A2(n633), .ZN(n464) );
  NAND2_X1 U421 ( .A1(n463), .A2(KEYINPUT47), .ZN(n465) );
  NAND2_X1 U422 ( .A1(n447), .A2(n445), .ZN(n463) );
  AND2_X1 U423 ( .A1(n446), .A2(n635), .ZN(n445) );
  XNOR2_X1 U424 ( .A(n560), .B(G902), .ZN(n689) );
  XNOR2_X1 U425 ( .A(n639), .B(n638), .ZN(n448) );
  XOR2_X1 U426 ( .A(KEYINPUT48), .B(KEYINPUT70), .Z(n638) );
  INV_X1 U427 ( .A(KEYINPUT69), .ZN(n535) );
  XNOR2_X1 U428 ( .A(n500), .B(n499), .ZN(n589) );
  XNOR2_X1 U429 ( .A(G119), .B(G113), .ZN(n499) );
  XNOR2_X1 U430 ( .A(n547), .B(G101), .ZN(n500) );
  INV_X1 U431 ( .A(KEYINPUT3), .ZN(n547) );
  NOR2_X1 U432 ( .A1(n627), .A2(n622), .ZN(n751) );
  NAND2_X1 U433 ( .A1(n505), .A2(n504), .ZN(n503) );
  AND2_X1 U434 ( .A1(n748), .A2(KEYINPUT88), .ZN(n504) );
  XNOR2_X1 U435 ( .A(n495), .B(n493), .ZN(n530) );
  XNOR2_X1 U436 ( .A(n529), .B(n494), .ZN(n493) );
  XNOR2_X1 U437 ( .A(n528), .B(n527), .ZN(n495) );
  XOR2_X1 U438 ( .A(KEYINPUT92), .B(G140), .Z(n566) );
  XNOR2_X1 U439 ( .A(n356), .B(G110), .ZN(n565) );
  XNOR2_X1 U440 ( .A(n573), .B(n568), .ZN(n474) );
  INV_X1 U441 ( .A(KEYINPUT24), .ZN(n567) );
  INV_X1 U442 ( .A(n569), .ZN(n472) );
  XNOR2_X1 U443 ( .A(KEYINPUT100), .B(KEYINPUT98), .ZN(n513) );
  INV_X1 U444 ( .A(G134), .ZN(n519) );
  INV_X1 U445 ( .A(G107), .ZN(n514) );
  INV_X1 U446 ( .A(G475), .ZN(n487) );
  XNOR2_X1 U447 ( .A(KEYINPUT33), .B(KEYINPUT71), .ZN(n647) );
  AND2_X1 U448 ( .A1(n387), .A2(n386), .ZN(n640) );
  INV_X1 U449 ( .A(n724), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n388), .B(KEYINPUT107), .ZN(n387) );
  XNOR2_X1 U451 ( .A(n587), .B(n431), .ZN(n395) );
  INV_X1 U452 ( .A(KEYINPUT75), .ZN(n431) );
  NOR2_X1 U453 ( .A1(n679), .A2(n586), .ZN(n587) );
  INV_X1 U454 ( .A(n656), .ZN(n469) );
  BUF_X1 U455 ( .A(n618), .Z(n737) );
  XNOR2_X1 U456 ( .A(n400), .B(KEYINPUT85), .ZN(n383) );
  OR2_X1 U457 ( .A1(n456), .A2(n432), .ZN(n380) );
  NOR2_X1 U458 ( .A1(n411), .A2(n788), .ZN(n410) );
  NOR2_X1 U459 ( .A1(n357), .A2(n708), .ZN(n411) );
  NOR2_X1 U460 ( .A1(n403), .A2(n788), .ZN(n402) );
  NOR2_X1 U461 ( .A1(n357), .A2(n704), .ZN(n403) );
  NAND2_X1 U462 ( .A1(n470), .A2(n469), .ZN(n721) );
  XNOR2_X1 U463 ( .A(n497), .B(KEYINPUT102), .ZN(n727) );
  NAND2_X1 U464 ( .A1(n466), .A2(n634), .ZN(n446) );
  XOR2_X1 U465 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n541) );
  XNOR2_X1 U466 ( .A(G116), .B(G131), .ZN(n540) );
  XOR2_X1 U467 ( .A(KEYINPUT93), .B(KEYINPUT5), .Z(n544) );
  XNOR2_X1 U468 ( .A(n436), .B(KEYINPUT72), .ZN(n636) );
  AND2_X1 U469 ( .A1(n465), .A2(n464), .ZN(n438) );
  INV_X1 U470 ( .A(KEYINPUT67), .ZN(n537) );
  XNOR2_X1 U471 ( .A(G146), .B(G125), .ZN(n596) );
  AND2_X1 U472 ( .A1(n498), .A2(n727), .ZN(n745) );
  OR2_X1 U473 ( .A1(n748), .A2(KEYINPUT88), .ZN(n507) );
  XNOR2_X1 U474 ( .A(KEYINPUT12), .B(KEYINPUT11), .ZN(n494) );
  AND2_X1 U475 ( .A1(n550), .A2(n444), .ZN(n441) );
  INV_X1 U476 ( .A(KEYINPUT1), .ZN(n393) );
  AND2_X1 U477 ( .A1(n448), .A2(n687), .ZN(n688) );
  NAND2_X1 U478 ( .A1(G234), .A2(G237), .ZN(n580) );
  INV_X1 U479 ( .A(G237), .ZN(n533) );
  NAND2_X1 U480 ( .A1(n655), .A2(n657), .ZN(n481) );
  INV_X1 U481 ( .A(n589), .ZN(n477) );
  INV_X1 U482 ( .A(KEYINPUT2), .ZN(n766) );
  AND2_X1 U483 ( .A1(n618), .A2(n368), .ZN(n608) );
  XNOR2_X1 U484 ( .A(n435), .B(n434), .ZN(n768) );
  INV_X1 U485 ( .A(KEYINPUT41), .ZN(n434) );
  XNOR2_X1 U486 ( .A(n551), .B(n452), .ZN(n451) );
  INV_X1 U487 ( .A(n646), .ZN(n392) );
  XNOR2_X1 U488 ( .A(n473), .B(n471), .ZN(n786) );
  XNOR2_X1 U489 ( .A(n570), .B(n472), .ZN(n471) );
  XNOR2_X1 U490 ( .A(n572), .B(n474), .ZN(n473) );
  XNOR2_X1 U491 ( .A(n588), .B(n427), .ZN(n522) );
  XNOR2_X1 U492 ( .A(n516), .B(n367), .ZN(n427) );
  NOR2_X1 U493 ( .A1(n419), .A2(n788), .ZN(n418) );
  NOR2_X1 U494 ( .A1(n357), .A2(n696), .ZN(n419) );
  XNOR2_X1 U495 ( .A(n430), .B(n375), .ZN(n812) );
  XNOR2_X1 U496 ( .A(n389), .B(n449), .ZN(n814) );
  INV_X1 U497 ( .A(KEYINPUT110), .ZN(n449) );
  XNOR2_X1 U498 ( .A(n450), .B(n621), .ZN(n390) );
  INV_X1 U499 ( .A(n658), .ZN(n510) );
  NOR2_X1 U500 ( .A1(n664), .A2(n399), .ZN(n398) );
  XNOR2_X1 U501 ( .A(n678), .B(n461), .ZN(n726) );
  XNOR2_X1 U502 ( .A(n462), .B(KEYINPUT31), .ZN(n461) );
  INV_X1 U503 ( .A(KEYINPUT95), .ZN(n462) );
  INV_X1 U504 ( .A(n737), .ZN(n665) );
  NAND2_X1 U505 ( .A1(n379), .A2(n377), .ZN(n709) );
  NAND2_X1 U506 ( .A1(n378), .A2(KEYINPUT86), .ZN(n377) );
  AND2_X1 U507 ( .A1(n381), .A2(n371), .ZN(n379) );
  NAND2_X1 U508 ( .A1(n415), .A2(n414), .ZN(n413) );
  NAND2_X1 U509 ( .A1(n407), .A2(n406), .ZN(n405) );
  INV_X1 U510 ( .A(n721), .ZN(n468) );
  AND2_X1 U511 ( .A1(n397), .A2(n749), .ZN(n358) );
  NOR2_X1 U512 ( .A1(n667), .A2(n666), .ZN(n359) );
  OR2_X1 U513 ( .A1(n626), .A2(n374), .ZN(n360) );
  AND2_X1 U514 ( .A1(n709), .A2(n373), .ZN(n361) );
  XNOR2_X1 U515 ( .A(n604), .B(KEYINPUT38), .ZN(n749) );
  OR2_X1 U516 ( .A1(n656), .A2(n480), .ZN(n362) );
  AND2_X1 U517 ( .A1(n454), .A2(n398), .ZN(n363) );
  AND2_X1 U518 ( .A1(n357), .A2(n708), .ZN(n364) );
  AND2_X1 U519 ( .A1(n357), .A2(n696), .ZN(n365) );
  AND2_X1 U520 ( .A1(n357), .A2(n704), .ZN(n366) );
  XNOR2_X1 U521 ( .A(n578), .B(n577), .ZN(n605) );
  XNOR2_X1 U522 ( .A(KEYINPUT7), .B(KEYINPUT9), .ZN(n367) );
  AND2_X1 U523 ( .A1(n605), .A2(n607), .ZN(n368) );
  OR2_X1 U524 ( .A1(KEYINPUT79), .A2(n632), .ZN(n369) );
  AND2_X1 U525 ( .A1(n395), .A2(n397), .ZN(n370) );
  AND2_X1 U526 ( .A1(n380), .A2(n733), .ZN(n371) );
  AND2_X1 U527 ( .A1(n686), .A2(n689), .ZN(n372) );
  NAND2_X1 U528 ( .A1(n683), .A2(n682), .ZN(n373) );
  BUF_X1 U529 ( .A(n731), .Z(n456) );
  NAND2_X1 U530 ( .A1(n469), .A2(KEYINPUT79), .ZN(n374) );
  XOR2_X1 U531 ( .A(KEYINPUT40), .B(KEYINPUT108), .Z(n375) );
  INV_X1 U532 ( .A(n469), .ZN(n466) );
  INV_X1 U533 ( .A(KEYINPUT86), .ZN(n432) );
  AND2_X1 U534 ( .A1(n697), .A2(G953), .ZN(n788) );
  INV_X1 U535 ( .A(G469), .ZN(n394) );
  INV_X1 U536 ( .A(G472), .ZN(n444) );
  NAND2_X1 U537 ( .A1(n669), .A2(n668), .ZN(n376) );
  NAND2_X1 U538 ( .A1(n490), .A2(n690), .ZN(n433) );
  INV_X1 U539 ( .A(n383), .ZN(n378) );
  NAND2_X1 U540 ( .A1(n383), .A2(n382), .ZN(n381) );
  AND2_X1 U541 ( .A1(n456), .A2(n432), .ZN(n382) );
  NAND2_X1 U542 ( .A1(n384), .A2(n688), .ZN(n492) );
  NAND2_X1 U543 ( .A1(n501), .A2(n384), .ZN(n502) );
  AND2_X1 U544 ( .A1(n384), .A2(n803), .ZN(n692) );
  NAND2_X1 U545 ( .A1(n384), .A2(n792), .ZN(n793) );
  XNOR2_X2 U546 ( .A(n684), .B(KEYINPUT45), .ZN(n384) );
  NAND2_X1 U547 ( .A1(n656), .A2(n657), .ZN(n385) );
  XNOR2_X2 U548 ( .A(n625), .B(n624), .ZN(n656) );
  NAND2_X1 U549 ( .A1(n662), .A2(n368), .ZN(n388) );
  NOR2_X1 U550 ( .A1(n636), .A2(n814), .ZN(n426) );
  NAND2_X1 U551 ( .A1(n390), .A2(n666), .ZN(n389) );
  XNOR2_X1 U552 ( .A(n391), .B(n549), .ZN(n707) );
  NAND2_X1 U553 ( .A1(n609), .A2(n392), .ZN(n679) );
  XNOR2_X2 U554 ( .A(n559), .B(n394), .ZN(n609) );
  INV_X1 U555 ( .A(n451), .ZN(n397) );
  NAND2_X1 U556 ( .A1(n454), .A2(n453), .ZN(n400) );
  INV_X1 U557 ( .A(n453), .ZN(n399) );
  NAND2_X1 U558 ( .A1(n401), .A2(n700), .ZN(n671) );
  XNOR2_X2 U559 ( .A(n363), .B(n479), .ZN(n401) );
  XNOR2_X1 U560 ( .A(n401), .B(G119), .ZN(G21) );
  AND2_X1 U561 ( .A1(n404), .A2(n402), .ZN(n408) );
  NAND2_X1 U562 ( .A1(n485), .A2(n366), .ZN(n404) );
  NAND2_X1 U563 ( .A1(n408), .A2(n405), .ZN(n409) );
  INV_X1 U564 ( .A(n704), .ZN(n406) );
  INV_X1 U565 ( .A(n485), .ZN(n407) );
  XNOR2_X1 U566 ( .A(n409), .B(n705), .ZN(G51) );
  AND2_X1 U567 ( .A1(n412), .A2(n410), .ZN(n416) );
  NAND2_X1 U568 ( .A1(n486), .A2(n364), .ZN(n412) );
  NAND2_X1 U569 ( .A1(n416), .A2(n413), .ZN(n417) );
  INV_X1 U570 ( .A(n708), .ZN(n414) );
  INV_X1 U571 ( .A(n486), .ZN(n415) );
  XNOR2_X1 U572 ( .A(n417), .B(KEYINPUT63), .ZN(G57) );
  AND2_X1 U573 ( .A1(n420), .A2(n418), .ZN(n424) );
  NAND2_X1 U574 ( .A1(n484), .A2(n365), .ZN(n420) );
  NAND2_X1 U575 ( .A1(n424), .A2(n421), .ZN(n425) );
  INV_X1 U576 ( .A(n696), .ZN(n422) );
  INV_X1 U577 ( .A(n484), .ZN(n423) );
  XNOR2_X1 U578 ( .A(n425), .B(n698), .ZN(G60) );
  NAND2_X1 U579 ( .A1(n426), .A2(n637), .ZN(n639) );
  NAND2_X1 U580 ( .A1(n369), .A2(n496), .ZN(n437) );
  XNOR2_X2 U581 ( .A(n428), .B(n455), .ZN(n454) );
  NAND2_X1 U582 ( .A1(n681), .A2(n661), .ZN(n428) );
  NAND2_X1 U583 ( .A1(n644), .A2(n629), .ZN(n430) );
  NOR2_X2 U584 ( .A1(n731), .A2(n646), .ZN(n675) );
  NOR2_X2 U585 ( .A1(n767), .A2(n677), .ZN(n512) );
  XNOR2_X1 U586 ( .A(n512), .B(KEYINPUT34), .ZN(n511) );
  NOR2_X2 U587 ( .A1(n765), .A2(n766), .ZN(n693) );
  XNOR2_X2 U588 ( .A(n433), .B(n691), .ZN(n694) );
  NAND2_X1 U589 ( .A1(n746), .A2(n751), .ZN(n435) );
  NAND2_X1 U590 ( .A1(n438), .A2(n437), .ZN(n436) );
  NAND2_X1 U591 ( .A1(n707), .A2(n441), .ZN(n440) );
  OR2_X1 U592 ( .A1(n707), .A2(n444), .ZN(n443) );
  NAND2_X1 U593 ( .A1(n626), .A2(n634), .ZN(n447) );
  AND2_X1 U594 ( .A1(n448), .A2(n372), .ZN(n501) );
  AND2_X1 U595 ( .A1(n448), .A2(n686), .ZN(n803) );
  NAND2_X1 U596 ( .A1(n640), .A2(n625), .ZN(n450) );
  INV_X1 U597 ( .A(KEYINPUT30), .ZN(n452) );
  INV_X1 U598 ( .A(n662), .ZN(n453) );
  NAND2_X1 U599 ( .A1(n454), .A2(n359), .ZN(n700) );
  NAND2_X1 U600 ( .A1(n482), .A2(n361), .ZN(n684) );
  NAND2_X1 U601 ( .A1(n458), .A2(n457), .ZN(n659) );
  INV_X1 U602 ( .A(KEYINPUT44), .ZN(n457) );
  INV_X1 U603 ( .A(n813), .ZN(n458) );
  NAND2_X1 U604 ( .A1(n459), .A2(n674), .ZN(n483) );
  NAND2_X1 U605 ( .A1(n672), .A2(n673), .ZN(n459) );
  NOR2_X1 U606 ( .A1(n694), .A2(n487), .ZN(n484) );
  NAND2_X1 U607 ( .A1(n511), .A2(n510), .ZN(n509) );
  NOR2_X1 U608 ( .A1(n787), .A2(n788), .ZN(G66) );
  OR2_X2 U609 ( .A1(n703), .A2(n689), .ZN(n603) );
  INV_X1 U610 ( .A(n626), .ZN(n470) );
  NAND2_X1 U611 ( .A1(n468), .A2(n717), .ZN(n718) );
  XNOR2_X1 U612 ( .A(n595), .B(n594), .ZN(n476) );
  XNOR2_X1 U613 ( .A(n591), .B(n588), .ZN(n478) );
  INV_X1 U614 ( .A(KEYINPUT32), .ZN(n479) );
  OR2_X1 U615 ( .A1(n655), .A2(n657), .ZN(n480) );
  OR2_X2 U616 ( .A1(n694), .A2(n693), .ZN(n489) );
  NOR2_X1 U617 ( .A1(n694), .A2(n488), .ZN(n485) );
  NOR2_X1 U618 ( .A1(n694), .A2(n444), .ZN(n486) );
  INV_X1 U619 ( .A(G210), .ZN(n488) );
  NOR2_X1 U620 ( .A1(n489), .A2(n394), .ZN(n778) );
  XNOR2_X1 U621 ( .A(n616), .B(n615), .ZN(n637) );
  NAND2_X1 U622 ( .A1(n491), .A2(n689), .ZN(n490) );
  NAND2_X1 U623 ( .A1(n492), .A2(n766), .ZN(n491) );
  INV_X1 U624 ( .A(n727), .ZN(n717) );
  NAND2_X1 U625 ( .A1(n628), .A2(n627), .ZN(n497) );
  INV_X1 U626 ( .A(n629), .ZN(n498) );
  XNOR2_X2 U627 ( .A(n515), .B(n514), .ZN(n588) );
  NAND2_X1 U628 ( .A1(n502), .A2(n685), .ZN(n690) );
  NAND2_X1 U629 ( .A1(n619), .A2(n620), .ZN(n508) );
  NAND2_X2 U630 ( .A1(n506), .A2(n503), .ZN(n625) );
  INV_X1 U631 ( .A(n619), .ZN(n505) );
  XNOR2_X2 U632 ( .A(n509), .B(KEYINPUT35), .ZN(n813) );
  XNOR2_X2 U633 ( .A(G110), .B(G104), .ZN(n590) );
  AND2_X1 U634 ( .A1(n734), .A2(n606), .ZN(n607) );
  XNOR2_X1 U635 ( .A(n567), .B(KEYINPUT23), .ZN(n568) );
  INV_X1 U636 ( .A(KEYINPUT60), .ZN(n698) );
  XNOR2_X1 U637 ( .A(n513), .B(KEYINPUT99), .ZN(n516) );
  XNOR2_X2 U638 ( .A(G122), .B(G116), .ZN(n515) );
  NAND2_X1 U639 ( .A1(G234), .A2(n792), .ZN(n517) );
  XOR2_X1 U640 ( .A(KEYINPUT8), .B(n517), .Z(n571) );
  NAND2_X1 U641 ( .A1(G217), .A2(n571), .ZN(n520) );
  XNOR2_X1 U642 ( .A(n536), .B(n520), .ZN(n521) );
  XNOR2_X1 U643 ( .A(n522), .B(n521), .ZN(n780) );
  NOR2_X1 U644 ( .A1(G902), .A2(n780), .ZN(n524) );
  XNOR2_X1 U645 ( .A(KEYINPUT101), .B(G478), .ZN(n523) );
  XNOR2_X1 U646 ( .A(KEYINPUT10), .B(KEYINPUT68), .ZN(n525) );
  XNOR2_X1 U647 ( .A(n569), .B(n554), .ZN(n801) );
  XNOR2_X1 U648 ( .A(G113), .B(G122), .ZN(n526) );
  XNOR2_X1 U649 ( .A(n526), .B(KEYINPUT96), .ZN(n528) );
  XNOR2_X1 U650 ( .A(G143), .B(G104), .ZN(n527) );
  NAND2_X1 U651 ( .A1(G214), .A2(n542), .ZN(n529) );
  XNOR2_X1 U652 ( .A(n801), .B(n530), .ZN(n695) );
  NOR2_X1 U653 ( .A1(G902), .A2(n695), .ZN(n532) );
  XNOR2_X1 U654 ( .A(KEYINPUT13), .B(KEYINPUT97), .ZN(n531) );
  NOR2_X1 U655 ( .A1(n627), .A2(n628), .ZN(n629) );
  INV_X1 U656 ( .A(G902), .ZN(n550) );
  NAND2_X1 U657 ( .A1(n550), .A2(n533), .ZN(n599) );
  NAND2_X1 U658 ( .A1(n599), .A2(G214), .ZN(n534) );
  XNOR2_X1 U659 ( .A(n534), .B(KEYINPUT90), .ZN(n748) );
  XNOR2_X1 U660 ( .A(n537), .B(KEYINPUT4), .ZN(n597) );
  XNOR2_X1 U661 ( .A(G137), .B(n597), .ZN(n538) );
  XNOR2_X1 U662 ( .A(n541), .B(n540), .ZN(n546) );
  NAND2_X1 U663 ( .A1(n542), .A2(G210), .ZN(n543) );
  XNOR2_X1 U664 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U665 ( .A(n546), .B(n545), .ZN(n548) );
  XNOR2_X1 U666 ( .A(n548), .B(n589), .ZN(n549) );
  XNOR2_X1 U667 ( .A(G101), .B(G107), .ZN(n552) );
  XNOR2_X1 U668 ( .A(n590), .B(n552), .ZN(n553) );
  XNOR2_X1 U669 ( .A(n554), .B(n553), .ZN(n555) );
  XOR2_X1 U670 ( .A(KEYINPUT91), .B(n555), .Z(n557) );
  NAND2_X1 U671 ( .A1(G227), .A2(n792), .ZN(n556) );
  XNOR2_X1 U672 ( .A(n557), .B(n556), .ZN(n558) );
  NOR2_X2 U673 ( .A1(G902), .A2(n774), .ZN(n559) );
  INV_X1 U674 ( .A(KEYINPUT15), .ZN(n560) );
  INV_X1 U675 ( .A(n689), .ZN(n561) );
  NAND2_X1 U676 ( .A1(n561), .A2(G234), .ZN(n562) );
  XNOR2_X1 U677 ( .A(n562), .B(KEYINPUT20), .ZN(n574) );
  NAND2_X1 U678 ( .A1(n574), .A2(G221), .ZN(n563) );
  XOR2_X1 U679 ( .A(KEYINPUT21), .B(n563), .Z(n734) );
  XNOR2_X1 U680 ( .A(G119), .B(G137), .ZN(n564) );
  XNOR2_X1 U681 ( .A(n564), .B(KEYINPUT77), .ZN(n573) );
  XNOR2_X1 U682 ( .A(n566), .B(n565), .ZN(n570) );
  NAND2_X1 U683 ( .A1(G221), .A2(n571), .ZN(n572) );
  NOR2_X1 U684 ( .A1(n786), .A2(G902), .ZN(n578) );
  NAND2_X1 U685 ( .A1(n574), .A2(G217), .ZN(n576) );
  XOR2_X1 U686 ( .A(KEYINPUT76), .B(KEYINPUT25), .Z(n575) );
  XNOR2_X1 U687 ( .A(n576), .B(n575), .ZN(n577) );
  INV_X1 U688 ( .A(n605), .ZN(n579) );
  NAND2_X1 U689 ( .A1(n734), .A2(n579), .ZN(n646) );
  XNOR2_X1 U690 ( .A(n580), .B(KEYINPUT14), .ZN(n654) );
  NAND2_X1 U691 ( .A1(G953), .A2(G902), .ZN(n649) );
  NOR2_X1 U692 ( .A1(G900), .A2(n649), .ZN(n581) );
  NAND2_X1 U693 ( .A1(n654), .A2(n581), .ZN(n582) );
  XOR2_X1 U694 ( .A(KEYINPUT106), .B(n582), .Z(n584) );
  INV_X1 U695 ( .A(n654), .ZN(n761) );
  NAND2_X1 U696 ( .A1(G952), .A2(n792), .ZN(n650) );
  NOR2_X1 U697 ( .A1(n761), .A2(n650), .ZN(n583) );
  NOR2_X1 U698 ( .A1(n584), .A2(n583), .ZN(n585) );
  XOR2_X1 U699 ( .A(KEYINPUT78), .B(n585), .Z(n606) );
  INV_X1 U700 ( .A(n606), .ZN(n586) );
  XNOR2_X1 U701 ( .A(n590), .B(KEYINPUT16), .ZN(n591) );
  XNOR2_X1 U702 ( .A(KEYINPUT17), .B(KEYINPUT18), .ZN(n593) );
  NAND2_X1 U703 ( .A1(n792), .A2(G224), .ZN(n592) );
  XNOR2_X1 U704 ( .A(n593), .B(n592), .ZN(n594) );
  XNOR2_X1 U705 ( .A(n597), .B(n596), .ZN(n598) );
  NAND2_X1 U706 ( .A1(n599), .A2(G210), .ZN(n601) );
  INV_X1 U707 ( .A(KEYINPUT89), .ZN(n600) );
  XNOR2_X1 U708 ( .A(n601), .B(n600), .ZN(n602) );
  XNOR2_X2 U709 ( .A(n603), .B(n602), .ZN(n619) );
  BUF_X1 U710 ( .A(n619), .Z(n604) );
  XNOR2_X1 U711 ( .A(KEYINPUT28), .B(n608), .ZN(n610) );
  NAND2_X1 U712 ( .A1(n610), .A2(n609), .ZN(n626) );
  INV_X1 U713 ( .A(n628), .ZN(n622) );
  NAND2_X1 U714 ( .A1(n749), .A2(n748), .ZN(n611) );
  XNOR2_X1 U715 ( .A(n611), .B(KEYINPUT109), .ZN(n746) );
  NOR2_X1 U716 ( .A1(n626), .A2(n768), .ZN(n612) );
  XNOR2_X1 U717 ( .A(n612), .B(KEYINPUT42), .ZN(n817) );
  INV_X1 U718 ( .A(KEYINPUT46), .ZN(n614) );
  INV_X1 U719 ( .A(KEYINPUT84), .ZN(n613) );
  XNOR2_X1 U720 ( .A(KEYINPUT36), .B(KEYINPUT87), .ZN(n621) );
  XNOR2_X1 U721 ( .A(KEYINPUT105), .B(n629), .ZN(n724) );
  INV_X1 U722 ( .A(KEYINPUT6), .ZN(n617) );
  INV_X1 U723 ( .A(KEYINPUT88), .ZN(n620) );
  NAND2_X1 U724 ( .A1(n627), .A2(n622), .ZN(n658) );
  NOR2_X1 U725 ( .A1(n658), .A2(n604), .ZN(n623) );
  AND2_X1 U726 ( .A1(n370), .A2(n623), .ZN(n720) );
  XNOR2_X1 U727 ( .A(KEYINPUT66), .B(KEYINPUT19), .ZN(n624) );
  OR2_X1 U728 ( .A1(KEYINPUT80), .A2(n745), .ZN(n630) );
  NAND2_X1 U729 ( .A1(n360), .A2(n630), .ZN(n633) );
  XNOR2_X1 U730 ( .A(n745), .B(KEYINPUT81), .ZN(n682) );
  NAND2_X1 U731 ( .A1(KEYINPUT80), .A2(n631), .ZN(n632) );
  NAND2_X1 U732 ( .A1(KEYINPUT80), .A2(n745), .ZN(n635) );
  INV_X1 U733 ( .A(KEYINPUT79), .ZN(n634) );
  INV_X1 U734 ( .A(n456), .ZN(n666) );
  NAND2_X1 U735 ( .A1(n748), .A2(n640), .ZN(n641) );
  NOR2_X1 U736 ( .A1(n666), .A2(n641), .ZN(n642) );
  XNOR2_X1 U737 ( .A(n642), .B(KEYINPUT43), .ZN(n643) );
  NOR2_X1 U738 ( .A1(n643), .A2(n505), .ZN(n701) );
  NAND2_X1 U739 ( .A1(n644), .A2(n717), .ZN(n729) );
  INV_X1 U740 ( .A(n729), .ZN(n645) );
  NOR2_X1 U741 ( .A1(n701), .A2(n645), .ZN(n686) );
  NAND2_X1 U742 ( .A1(n662), .A2(n675), .ZN(n648) );
  XNOR2_X2 U743 ( .A(n648), .B(n647), .ZN(n767) );
  NOR2_X1 U744 ( .A1(G898), .A2(n649), .ZN(n652) );
  INV_X1 U745 ( .A(n650), .ZN(n651) );
  OR2_X1 U746 ( .A1(n652), .A2(n651), .ZN(n653) );
  NAND2_X1 U747 ( .A1(n654), .A2(n653), .ZN(n655) );
  INV_X1 U748 ( .A(KEYINPUT0), .ZN(n657) );
  INV_X1 U749 ( .A(n681), .ZN(n677) );
  INV_X1 U750 ( .A(KEYINPUT65), .ZN(n670) );
  NAND2_X1 U751 ( .A1(n659), .A2(n670), .ZN(n669) );
  NAND2_X1 U752 ( .A1(n751), .A2(n734), .ZN(n660) );
  INV_X1 U753 ( .A(KEYINPUT104), .ZN(n663) );
  XNOR2_X1 U754 ( .A(n605), .B(n663), .ZN(n733) );
  OR2_X1 U755 ( .A1(n733), .A2(n456), .ZN(n664) );
  NAND2_X1 U756 ( .A1(n605), .A2(n665), .ZN(n667) );
  INV_X1 U757 ( .A(n671), .ZN(n668) );
  NOR2_X1 U758 ( .A1(n813), .A2(n457), .ZN(n673) );
  NAND2_X1 U759 ( .A1(n671), .A2(n670), .ZN(n672) );
  OR2_X1 U760 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n674) );
  NAND2_X1 U761 ( .A1(n675), .A2(n737), .ZN(n676) );
  XNOR2_X1 U762 ( .A(n676), .B(KEYINPUT94), .ZN(n741) );
  NOR2_X1 U763 ( .A1(n741), .A2(n677), .ZN(n678) );
  NOR2_X1 U764 ( .A1(n737), .A2(n679), .ZN(n680) );
  NAND2_X1 U765 ( .A1(n681), .A2(n680), .ZN(n712) );
  NAND2_X1 U766 ( .A1(n726), .A2(n712), .ZN(n683) );
  INV_X1 U767 ( .A(KEYINPUT82), .ZN(n685) );
  AND2_X1 U768 ( .A1(n686), .A2(KEYINPUT82), .ZN(n687) );
  INV_X1 U769 ( .A(n692), .ZN(n765) );
  XNOR2_X1 U770 ( .A(n695), .B(KEYINPUT59), .ZN(n696) );
  INV_X1 U771 ( .A(G952), .ZN(n697) );
  XNOR2_X1 U772 ( .A(G110), .B(KEYINPUT114), .ZN(n699) );
  XNOR2_X1 U773 ( .A(n700), .B(n699), .ZN(G12) );
  XOR2_X1 U774 ( .A(G140), .B(n701), .Z(G42) );
  XNOR2_X1 U775 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n702) );
  XNOR2_X1 U776 ( .A(n703), .B(n702), .ZN(n704) );
  XNOR2_X1 U777 ( .A(KEYINPUT83), .B(KEYINPUT56), .ZN(n705) );
  XOR2_X1 U778 ( .A(KEYINPUT111), .B(KEYINPUT62), .Z(n706) );
  XNOR2_X1 U779 ( .A(n707), .B(n706), .ZN(n708) );
  XNOR2_X1 U780 ( .A(G101), .B(n709), .ZN(G3) );
  NOR2_X1 U781 ( .A1(n724), .A2(n712), .ZN(n710) );
  XOR2_X1 U782 ( .A(KEYINPUT112), .B(n710), .Z(n711) );
  XNOR2_X1 U783 ( .A(G104), .B(n711), .ZN(G6) );
  NOR2_X1 U784 ( .A1(n712), .A2(n727), .ZN(n716) );
  XOR2_X1 U785 ( .A(KEYINPUT26), .B(KEYINPUT113), .Z(n714) );
  XNOR2_X1 U786 ( .A(G107), .B(KEYINPUT27), .ZN(n713) );
  XNOR2_X1 U787 ( .A(n714), .B(n713), .ZN(n715) );
  XNOR2_X1 U788 ( .A(n716), .B(n715), .ZN(G9) );
  XOR2_X1 U789 ( .A(n356), .B(KEYINPUT29), .Z(n719) );
  XNOR2_X1 U790 ( .A(n719), .B(n718), .ZN(G30) );
  XOR2_X1 U791 ( .A(G143), .B(n720), .Z(G45) );
  NOR2_X1 U792 ( .A1(n721), .A2(n724), .ZN(n723) );
  XNOR2_X1 U793 ( .A(G146), .B(KEYINPUT115), .ZN(n722) );
  XNOR2_X1 U794 ( .A(n723), .B(n722), .ZN(G48) );
  NOR2_X1 U795 ( .A1(n724), .A2(n726), .ZN(n725) );
  XOR2_X1 U796 ( .A(G113), .B(n725), .Z(G15) );
  NOR2_X1 U797 ( .A1(n727), .A2(n726), .ZN(n728) );
  XOR2_X1 U798 ( .A(G116), .B(n728), .Z(G18) );
  XNOR2_X1 U799 ( .A(G134), .B(n729), .ZN(G36) );
  XNOR2_X1 U800 ( .A(KEYINPUT52), .B(KEYINPUT119), .ZN(n730) );
  XNOR2_X1 U801 ( .A(n730), .B(KEYINPUT118), .ZN(n759) );
  NAND2_X1 U802 ( .A1(n456), .A2(n646), .ZN(n732) );
  XNOR2_X1 U803 ( .A(KEYINPUT50), .B(n732), .ZN(n739) );
  NOR2_X1 U804 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U805 ( .A(KEYINPUT49), .B(n735), .Z(n736) );
  NOR2_X1 U806 ( .A1(n737), .A2(n736), .ZN(n738) );
  NAND2_X1 U807 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U808 ( .A(KEYINPUT116), .B(n740), .ZN(n742) );
  NAND2_X1 U809 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U810 ( .A(KEYINPUT51), .B(n743), .ZN(n744) );
  NOR2_X1 U811 ( .A1(n768), .A2(n744), .ZN(n757) );
  INV_X1 U812 ( .A(n745), .ZN(n747) );
  NAND2_X1 U813 ( .A1(n747), .A2(n746), .ZN(n754) );
  NOR2_X1 U814 ( .A1(n749), .A2(n748), .ZN(n750) );
  XNOR2_X1 U815 ( .A(KEYINPUT117), .B(n750), .ZN(n752) );
  NAND2_X1 U816 ( .A1(n752), .A2(n751), .ZN(n753) );
  AND2_X1 U817 ( .A1(n754), .A2(n753), .ZN(n755) );
  NOR2_X1 U818 ( .A1(n755), .A2(n767), .ZN(n756) );
  NOR2_X1 U819 ( .A1(n757), .A2(n756), .ZN(n758) );
  XOR2_X1 U820 ( .A(n759), .B(n758), .Z(n760) );
  NOR2_X1 U821 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U822 ( .A1(n762), .A2(G952), .ZN(n763) );
  XOR2_X1 U823 ( .A(KEYINPUT120), .B(n763), .Z(n764) );
  NOR2_X1 U824 ( .A1(G953), .A2(n764), .ZN(n772) );
  XNOR2_X1 U825 ( .A(n692), .B(n766), .ZN(n770) );
  NOR2_X1 U826 ( .A1(n768), .A2(n767), .ZN(n769) );
  NOR2_X1 U827 ( .A1(n770), .A2(n769), .ZN(n771) );
  NAND2_X1 U828 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U829 ( .A(KEYINPUT53), .B(n773), .Z(G75) );
  XOR2_X1 U830 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n776) );
  XNOR2_X1 U831 ( .A(n774), .B(KEYINPUT121), .ZN(n775) );
  XNOR2_X1 U832 ( .A(n776), .B(n775), .ZN(n777) );
  XNOR2_X1 U833 ( .A(n778), .B(n777), .ZN(n779) );
  NOR2_X1 U834 ( .A1(n788), .A2(n779), .ZN(G54) );
  NAND2_X1 U835 ( .A1(n784), .A2(G478), .ZN(n782) );
  XNOR2_X1 U836 ( .A(n782), .B(n781), .ZN(n783) );
  NOR2_X1 U837 ( .A1(n788), .A2(n783), .ZN(G63) );
  NAND2_X1 U838 ( .A1(n784), .A2(G217), .ZN(n785) );
  XNOR2_X1 U839 ( .A(n786), .B(n785), .ZN(n787) );
  XNOR2_X1 U840 ( .A(n789), .B(KEYINPUT125), .ZN(n791) );
  NOR2_X1 U841 ( .A1(n792), .A2(G898), .ZN(n790) );
  NOR2_X1 U842 ( .A1(n791), .A2(n790), .ZN(n800) );
  XNOR2_X1 U843 ( .A(n793), .B(KEYINPUT124), .ZN(n798) );
  XOR2_X1 U844 ( .A(KEYINPUT123), .B(KEYINPUT61), .Z(n795) );
  NAND2_X1 U845 ( .A1(G224), .A2(G953), .ZN(n794) );
  XNOR2_X1 U846 ( .A(n795), .B(n794), .ZN(n796) );
  NAND2_X1 U847 ( .A1(n796), .A2(G898), .ZN(n797) );
  NAND2_X1 U848 ( .A1(n798), .A2(n797), .ZN(n799) );
  XNOR2_X1 U849 ( .A(n800), .B(n799), .ZN(G69) );
  XNOR2_X1 U850 ( .A(n802), .B(n801), .ZN(n805) );
  XNOR2_X1 U851 ( .A(n803), .B(n805), .ZN(n804) );
  NOR2_X1 U852 ( .A1(G953), .A2(n804), .ZN(n810) );
  XNOR2_X1 U853 ( .A(G227), .B(n805), .ZN(n806) );
  NAND2_X1 U854 ( .A1(n806), .A2(G900), .ZN(n807) );
  NAND2_X1 U855 ( .A1(G953), .A2(n807), .ZN(n808) );
  XOR2_X1 U856 ( .A(KEYINPUT126), .B(n808), .Z(n809) );
  NOR2_X1 U857 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U858 ( .A(KEYINPUT127), .B(n811), .ZN(G72) );
  XOR2_X1 U859 ( .A(n812), .B(G131), .Z(G33) );
  XOR2_X1 U860 ( .A(n813), .B(G122), .Z(G24) );
  INV_X1 U861 ( .A(n814), .ZN(n815) );
  XOR2_X1 U862 ( .A(G125), .B(n815), .Z(n816) );
  XNOR2_X1 U863 ( .A(KEYINPUT37), .B(n816), .ZN(G27) );
  XOR2_X1 U864 ( .A(n817), .B(G137), .Z(G39) );
endmodule

