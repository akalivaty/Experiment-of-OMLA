//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 1 1 1 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 1 0 1 0 0 0 0 1 0 0 0 0 0 1 1 1 1 0 0 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n666, new_n667, new_n668,
    new_n669, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n744, new_n745, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n794, new_n795, new_n796, new_n797, new_n799, new_n801,
    new_n802, new_n803, new_n804, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n889, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n943, new_n944;
  XNOR2_X1  g000(.A(KEYINPUT0), .B(G57gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G85gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(G1gat), .B(G29gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G127gat), .B(G134gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n207), .B(KEYINPUT69), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT1), .ZN(new_n209));
  INV_X1    g008(.A(G120gat), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n210), .A2(G113gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n210), .A2(G113gat), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n211), .B1(KEYINPUT68), .B2(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n213), .B1(KEYINPUT68), .B2(new_n212), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n208), .A2(new_n209), .A3(new_n214), .ZN(new_n215));
  XNOR2_X1  g014(.A(new_n207), .B(KEYINPUT67), .ZN(new_n216));
  INV_X1    g015(.A(new_n212), .ZN(new_n217));
  OAI21_X1  g016(.A(new_n209), .B1(new_n217), .B2(new_n211), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n215), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G141gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(G148gat), .ZN(new_n222));
  XOR2_X1   g021(.A(KEYINPUT80), .B(G148gat), .Z(new_n223));
  OAI21_X1  g022(.A(new_n222), .B1(new_n223), .B2(new_n221), .ZN(new_n224));
  XNOR2_X1  g023(.A(KEYINPUT81), .B(G162gat), .ZN(new_n225));
  INV_X1    g024(.A(G155gat), .ZN(new_n226));
  OAI21_X1  g025(.A(KEYINPUT2), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(G155gat), .A2(G162gat), .ZN(new_n228));
  INV_X1    g027(.A(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(G155gat), .A2(G162gat), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n224), .B(new_n227), .C1(new_n229), .C2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n228), .A2(KEYINPUT2), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n232), .A2(KEYINPUT79), .ZN(new_n233));
  INV_X1    g032(.A(G148gat), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n234), .A2(G141gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n222), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT79), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n228), .A2(new_n237), .A3(KEYINPUT2), .ZN(new_n238));
  NAND3_X1  g037(.A1(new_n233), .A2(new_n236), .A3(new_n238), .ZN(new_n239));
  XOR2_X1   g038(.A(new_n228), .B(KEYINPUT78), .Z(new_n240));
  OAI211_X1 g039(.A(new_n239), .B(new_n240), .C1(G155gat), .C2(G162gat), .ZN(new_n241));
  AND2_X1   g040(.A1(new_n231), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n220), .A2(new_n242), .ZN(new_n243));
  NAND2_X1  g042(.A1(new_n215), .A2(new_n219), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n231), .A2(new_n241), .ZN(new_n245));
  NAND2_X1  g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(G225gat), .A2(G233gat), .ZN(new_n248));
  INV_X1    g047(.A(new_n248), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n250), .A2(KEYINPUT5), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT4), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n243), .A2(new_n252), .ZN(new_n253));
  NAND3_X1  g052(.A1(new_n220), .A2(new_n242), .A3(KEYINPUT4), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n245), .A2(KEYINPUT3), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT3), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n256), .A3(new_n241), .ZN(new_n257));
  NAND3_X1  g056(.A1(new_n255), .A2(new_n244), .A3(new_n257), .ZN(new_n258));
  NAND4_X1  g057(.A1(new_n253), .A2(new_n248), .A3(new_n254), .A4(new_n258), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT82), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n260), .A2(KEYINPUT5), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n251), .A2(new_n259), .A3(new_n261), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n251), .B1(new_n259), .B2(new_n261), .ZN(new_n263));
  OAI21_X1  g062(.A(new_n206), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT6), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n259), .A2(new_n261), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT5), .A3(new_n250), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n251), .A2(new_n259), .A3(new_n261), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n205), .B(KEYINPUT87), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n267), .A2(new_n268), .A3(new_n269), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n264), .A2(new_n265), .A3(new_n270), .ZN(new_n271));
  NOR2_X1   g070(.A1(new_n262), .A2(new_n263), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n272), .A2(KEYINPUT83), .A3(KEYINPUT6), .A4(new_n205), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT83), .ZN(new_n274));
  NAND3_X1  g073(.A1(new_n267), .A2(new_n268), .A3(new_n205), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n274), .B1(new_n275), .B2(new_n265), .ZN(new_n276));
  AND3_X1   g075(.A1(new_n271), .A2(new_n273), .A3(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G183gat), .A2(G190gat), .ZN(new_n278));
  XNOR2_X1  g077(.A(new_n278), .B(KEYINPUT24), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n279), .B1(G183gat), .B2(G190gat), .ZN(new_n280));
  NAND2_X1  g079(.A1(G169gat), .A2(G176gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(KEYINPUT23), .ZN(new_n282));
  INV_X1    g081(.A(G169gat), .ZN(new_n283));
  INV_X1    g082(.A(G176gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n282), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g085(.A1(G169gat), .A2(G176gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(KEYINPUT23), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n280), .A2(new_n286), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n289), .A2(KEYINPUT25), .ZN(new_n290));
  XNOR2_X1  g089(.A(KEYINPUT27), .B(G183gat), .ZN(new_n291));
  INV_X1    g090(.A(G190gat), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  OR2_X1    g092(.A1(new_n293), .A2(KEYINPUT28), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n293), .A2(KEYINPUT28), .B1(G183gat), .B2(G190gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n287), .A2(KEYINPUT26), .ZN(new_n296));
  INV_X1    g095(.A(KEYINPUT26), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n285), .A2(new_n297), .A3(new_n281), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n294), .A2(new_n295), .A3(new_n296), .A4(new_n298), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT66), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT25), .ZN(new_n301));
  NAND4_X1  g100(.A1(new_n286), .A2(new_n300), .A3(new_n301), .A4(new_n288), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n302), .B1(new_n300), .B2(new_n288), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT65), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n304), .B1(G183gat), .B2(G190gat), .ZN(new_n305));
  INV_X1    g104(.A(G183gat), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n306), .A2(new_n292), .A3(KEYINPUT65), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n279), .A2(new_n305), .A3(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n303), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g108(.A1(new_n290), .A2(new_n299), .A3(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(KEYINPUT29), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(G226gat), .A2(G233gat), .ZN(new_n313));
  XNOR2_X1  g112(.A(new_n313), .B(KEYINPUT71), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  XOR2_X1   g114(.A(new_n314), .B(KEYINPUT72), .Z(new_n316));
  NAND2_X1  g115(.A1(new_n310), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G197gat), .B(G204gat), .ZN(new_n320));
  INV_X1    g119(.A(G211gat), .ZN(new_n321));
  INV_X1    g120(.A(G218gat), .ZN(new_n322));
  NOR2_X1   g121(.A1(new_n321), .A2(new_n322), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n320), .B1(KEYINPUT22), .B2(new_n323), .ZN(new_n324));
  XNOR2_X1  g123(.A(G211gat), .B(G218gat), .ZN(new_n325));
  XNOR2_X1  g124(.A(new_n324), .B(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n316), .ZN(new_n328));
  NAND4_X1  g127(.A1(new_n315), .A2(new_n319), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  OR2_X1    g128(.A1(new_n329), .A2(KEYINPUT74), .ZN(new_n330));
  INV_X1    g129(.A(new_n316), .ZN(new_n331));
  INV_X1    g130(.A(new_n314), .ZN(new_n332));
  AOI22_X1  g131(.A1(new_n312), .A2(new_n331), .B1(new_n310), .B2(new_n332), .ZN(new_n333));
  OAI211_X1 g132(.A(new_n329), .B(KEYINPUT74), .C1(new_n333), .C2(new_n327), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n330), .A2(new_n334), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT37), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G64gat), .B(G92gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(G36gat), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n339), .B(KEYINPUT75), .ZN(new_n340));
  INV_X1    g139(.A(G8gat), .ZN(new_n341));
  XNOR2_X1  g140(.A(new_n340), .B(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n337), .A2(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n335), .A2(new_n336), .ZN(new_n345));
  OAI21_X1  g144(.A(KEYINPUT38), .B1(new_n344), .B2(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n343), .B1(new_n330), .B2(new_n334), .ZN(new_n347));
  NOR2_X1   g146(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT76), .ZN(new_n349));
  AOI211_X1 g148(.A(new_n349), .B(new_n343), .C1(new_n330), .C2(new_n334), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n348), .A2(new_n350), .ZN(new_n351));
  INV_X1    g150(.A(KEYINPUT38), .ZN(new_n352));
  NAND4_X1  g151(.A1(new_n315), .A2(new_n319), .A3(new_n326), .A4(new_n328), .ZN(new_n353));
  OAI211_X1 g152(.A(new_n353), .B(KEYINPUT37), .C1(new_n326), .C2(new_n333), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n337), .A2(new_n352), .A3(new_n343), .A4(new_n354), .ZN(new_n355));
  NAND4_X1  g154(.A1(new_n277), .A2(new_n346), .A3(new_n351), .A4(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n253), .A2(new_n254), .A3(new_n258), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n357), .A2(new_n249), .ZN(new_n358));
  OR2_X1    g157(.A1(new_n358), .A2(KEYINPUT39), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n358), .B(KEYINPUT39), .C1(new_n249), .C2(new_n247), .ZN(new_n360));
  INV_X1    g159(.A(new_n269), .ZN(new_n361));
  NAND3_X1  g160(.A1(new_n359), .A2(new_n360), .A3(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT40), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n359), .A2(new_n360), .A3(KEYINPUT40), .A4(new_n361), .ZN(new_n365));
  AND3_X1   g164(.A1(new_n364), .A2(new_n365), .A3(new_n270), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT77), .B(KEYINPUT30), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  NOR3_X1   g167(.A1(new_n348), .A2(new_n350), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n347), .A2(KEYINPUT30), .ZN(new_n370));
  OAI21_X1  g169(.A(new_n370), .B1(new_n335), .B2(new_n342), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n366), .B1(new_n369), .B2(new_n371), .ZN(new_n372));
  XNOR2_X1  g171(.A(G78gat), .B(G106gat), .ZN(new_n373));
  INV_X1    g172(.A(G22gat), .ZN(new_n374));
  XNOR2_X1  g173(.A(new_n373), .B(new_n374), .ZN(new_n375));
  XNOR2_X1  g174(.A(new_n375), .B(G50gat), .ZN(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  XNOR2_X1  g176(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n378));
  XOR2_X1   g177(.A(new_n378), .B(KEYINPUT85), .Z(new_n379));
  AND2_X1   g178(.A1(G228gat), .A2(G233gat), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n257), .A2(new_n311), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT86), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n257), .A2(KEYINPUT86), .A3(new_n311), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n384), .A2(new_n326), .A3(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n256), .B1(new_n326), .B2(KEYINPUT29), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n245), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n381), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n388), .A2(new_n381), .ZN(new_n390));
  AOI21_X1  g189(.A(new_n390), .B1(new_n326), .B2(new_n382), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n379), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NOR3_X1   g192(.A1(new_n389), .A2(new_n391), .A3(new_n379), .ZN(new_n394));
  OAI21_X1  g193(.A(new_n377), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  NAND3_X1  g195(.A1(new_n396), .A2(new_n376), .A3(new_n392), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n356), .A2(new_n372), .A3(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n335), .A2(new_n342), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n401), .A2(new_n349), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n347), .A2(KEYINPUT76), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n402), .A2(new_n403), .A3(new_n367), .ZN(new_n404));
  NOR2_X1   g203(.A1(new_n335), .A2(new_n342), .ZN(new_n405));
  AOI21_X1  g204(.A(new_n405), .B1(new_n347), .B2(KEYINPUT30), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n404), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n264), .A2(new_n265), .A3(new_n275), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n408), .A2(new_n273), .A3(new_n276), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n398), .B1(new_n407), .B2(new_n409), .ZN(new_n410));
  XNOR2_X1  g209(.A(G15gat), .B(G43gat), .ZN(new_n411));
  XNOR2_X1  g210(.A(new_n411), .B(G71gat), .ZN(new_n412));
  INV_X1    g211(.A(G99gat), .ZN(new_n413));
  XNOR2_X1  g212(.A(new_n412), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(G227gat), .A2(G233gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(new_n415), .B(KEYINPUT64), .ZN(new_n416));
  INV_X1    g215(.A(new_n416), .ZN(new_n417));
  OR2_X1    g216(.A1(new_n310), .A2(new_n244), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n310), .A2(new_n244), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(KEYINPUT70), .B(KEYINPUT33), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n414), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n418), .A2(new_n417), .A3(new_n419), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT34), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT34), .ZN(new_n425));
  NAND4_X1  g224(.A1(new_n418), .A2(new_n425), .A3(new_n417), .A4(new_n419), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT32), .ZN(new_n428));
  NOR2_X1   g227(.A1(new_n420), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(new_n427), .A2(new_n429), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n427), .A2(new_n429), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n422), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  AND2_X1   g231(.A1(new_n418), .A2(new_n419), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT32), .B1(new_n433), .B2(new_n417), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n434), .A2(new_n424), .A3(new_n426), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n427), .A2(new_n429), .ZN(new_n436));
  INV_X1    g235(.A(new_n422), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n435), .A2(new_n436), .A3(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n432), .A2(new_n438), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(KEYINPUT36), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n400), .A2(new_n410), .A3(new_n441), .ZN(new_n442));
  NOR2_X1   g241(.A1(new_n407), .A2(new_n409), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n432), .A2(new_n395), .A3(new_n438), .A4(new_n397), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT35), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(new_n444), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n271), .A2(new_n273), .A3(new_n276), .ZN(new_n448));
  NAND4_X1  g247(.A1(new_n447), .A2(new_n448), .A3(new_n406), .A4(new_n404), .ZN(new_n449));
  AOI22_X1  g248(.A1(new_n443), .A2(new_n446), .B1(new_n449), .B2(new_n445), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n442), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(G230gat), .A2(G233gat), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT91), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(G57gat), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n454), .B(G64gat), .ZN(new_n455));
  INV_X1    g254(.A(G71gat), .ZN(new_n456));
  INV_X1    g255(.A(G78gat), .ZN(new_n457));
  NOR2_X1   g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(new_n458), .ZN(new_n459));
  NOR2_X1   g258(.A1(G71gat), .A2(G78gat), .ZN(new_n460));
  INV_X1    g259(.A(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT9), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n455), .A2(new_n463), .ZN(new_n464));
  NOR2_X1   g263(.A1(new_n458), .A2(new_n460), .ZN(new_n465));
  OR2_X1    g264(.A1(G57gat), .A2(G64gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(G57gat), .A2(G64gat), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n466), .A2(KEYINPUT9), .A3(new_n467), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g269(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n471));
  NOR2_X1   g270(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n472));
  NAND2_X1  g271(.A1(G85gat), .A2(G92gat), .ZN(new_n473));
  NOR3_X1   g272(.A1(new_n471), .A2(new_n472), .A3(new_n473), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n473), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  NOR2_X1   g275(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT95), .B(G92gat), .ZN(new_n478));
  INV_X1    g277(.A(G85gat), .ZN(new_n479));
  NAND2_X1  g278(.A1(G99gat), .A2(G106gat), .ZN(new_n480));
  AOI22_X1  g279(.A1(new_n478), .A2(new_n479), .B1(KEYINPUT8), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n480), .ZN(new_n482));
  NOR2_X1   g281(.A1(G99gat), .A2(G106gat), .ZN(new_n483));
  OAI21_X1  g282(.A(KEYINPUT96), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n483), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT96), .ZN(new_n486));
  NAND3_X1  g285(.A1(new_n485), .A2(new_n486), .A3(new_n480), .ZN(new_n487));
  AOI22_X1  g286(.A1(new_n477), .A2(new_n481), .B1(new_n484), .B2(new_n487), .ZN(new_n488));
  AND2_X1   g287(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n489));
  NOR2_X1   g288(.A1(KEYINPUT95), .A2(G92gat), .ZN(new_n490));
  OAI21_X1  g289(.A(new_n479), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(KEYINPUT94), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT7), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  AND2_X1   g293(.A1(G85gat), .A2(G92gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(KEYINPUT94), .A2(KEYINPUT7), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n495), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n480), .A2(KEYINPUT8), .ZN(new_n498));
  NAND4_X1  g297(.A1(new_n491), .A2(new_n497), .A3(new_n498), .A4(new_n475), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n487), .A2(new_n484), .ZN(new_n500));
  NOR2_X1   g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g300(.A(new_n470), .B1(new_n488), .B2(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT10), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n477), .A2(new_n481), .A3(new_n484), .A4(new_n487), .ZN(new_n504));
  AOI22_X1  g303(.A1(new_n455), .A2(new_n463), .B1(new_n468), .B2(new_n465), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n499), .A2(new_n500), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n504), .A2(new_n505), .A3(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n502), .A2(new_n503), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n509));
  NOR2_X1   g308(.A1(new_n488), .A2(new_n501), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n510), .A2(KEYINPUT10), .A3(new_n505), .ZN(new_n511));
  AND3_X1   g310(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n509), .B1(new_n508), .B2(new_n511), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n452), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  AOI21_X1  g313(.A(new_n452), .B1(new_n502), .B2(new_n507), .ZN(new_n515));
  INV_X1    g314(.A(new_n515), .ZN(new_n516));
  XNOR2_X1  g315(.A(G120gat), .B(G148gat), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n517), .B(new_n284), .ZN(new_n518));
  INV_X1    g317(.A(G204gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n514), .A2(new_n516), .A3(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n508), .A2(new_n511), .ZN(new_n523));
  AND2_X1   g322(.A1(new_n523), .A2(new_n452), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n520), .B1(new_n524), .B2(new_n515), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n522), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(new_n526), .ZN(new_n527));
  OR2_X1    g326(.A1(G15gat), .A2(G22gat), .ZN(new_n528));
  NAND2_X1  g327(.A1(G15gat), .A2(G22gat), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(G1gat), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n531), .A2(KEYINPUT16), .ZN(new_n532));
  AOI21_X1  g331(.A(KEYINPUT89), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n528), .A2(new_n531), .A3(new_n529), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(new_n535), .B(G8gat), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n505), .A2(KEYINPUT21), .ZN(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  OAI21_X1  g337(.A(G183gat), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  XNOR2_X1  g338(.A(G127gat), .B(G155gat), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  NOR2_X1   g340(.A1(new_n535), .A2(G8gat), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n341), .B1(new_n533), .B2(new_n534), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n544), .A2(new_n306), .A3(new_n537), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n539), .A2(new_n541), .A3(new_n545), .ZN(new_n546));
  INV_X1    g345(.A(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(KEYINPUT92), .B(KEYINPUT21), .Z(new_n548));
  NAND2_X1  g347(.A1(new_n470), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(KEYINPUT93), .B(G211gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n549), .B(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(new_n541), .B1(new_n539), .B2(new_n545), .ZN(new_n552));
  OR3_X1    g351(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n551), .B1(new_n547), .B2(new_n552), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  XNOR2_X1  g354(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n556));
  NAND2_X1  g355(.A1(G231gat), .A2(G233gat), .ZN(new_n557));
  XOR2_X1   g356(.A(new_n556), .B(new_n557), .Z(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  NOR2_X1   g358(.A1(new_n555), .A2(new_n559), .ZN(new_n560));
  INV_X1    g359(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n555), .A2(new_n559), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT88), .ZN(new_n564));
  INV_X1    g363(.A(G50gat), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(G43gat), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT15), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(G29gat), .A2(G36gat), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT14), .ZN(new_n570));
  OAI21_X1  g369(.A(new_n570), .B1(G29gat), .B2(G36gat), .ZN(new_n571));
  INV_X1    g370(.A(G29gat), .ZN(new_n572));
  INV_X1    g371(.A(G36gat), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n572), .A2(new_n573), .A3(KEYINPUT14), .ZN(new_n574));
  NAND4_X1  g373(.A1(new_n568), .A2(new_n569), .A3(new_n571), .A4(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G43gat), .B(G50gat), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n574), .A2(new_n571), .A3(new_n569), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n577), .A2(new_n567), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n575), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AND2_X1   g378(.A1(new_n574), .A2(new_n571), .ZN(new_n580));
  INV_X1    g379(.A(new_n576), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n580), .A2(new_n581), .A3(new_n568), .A4(new_n569), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G232gat), .A2(G233gat), .ZN(new_n584));
  AOI22_X1  g383(.A1(new_n510), .A2(new_n583), .B1(KEYINPUT41), .B2(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(KEYINPUT17), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n583), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n579), .A2(KEYINPUT17), .A3(new_n582), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n585), .B1(new_n589), .B2(new_n510), .ZN(new_n590));
  XOR2_X1   g389(.A(G134gat), .B(G162gat), .Z(new_n591));
  XNOR2_X1  g390(.A(new_n590), .B(new_n591), .ZN(new_n592));
  NOR2_X1   g391(.A1(new_n584), .A2(KEYINPUT41), .ZN(new_n593));
  XNOR2_X1  g392(.A(G190gat), .B(G218gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n592), .B(new_n595), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n563), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(new_n544), .A3(new_n588), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n536), .A2(new_n583), .ZN(new_n599));
  NAND2_X1  g398(.A1(G229gat), .A2(G233gat), .ZN(new_n600));
  NAND3_X1  g399(.A1(new_n598), .A2(new_n599), .A3(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT18), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n598), .A2(KEYINPUT18), .A3(new_n599), .A4(new_n600), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XNOR2_X1  g404(.A(KEYINPUT11), .B(G169gat), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(G197gat), .ZN(new_n607));
  XNOR2_X1  g406(.A(G113gat), .B(G141gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n607), .B(new_n608), .ZN(new_n609));
  XOR2_X1   g408(.A(new_n609), .B(KEYINPUT12), .Z(new_n610));
  XNOR2_X1  g409(.A(new_n536), .B(new_n583), .ZN(new_n611));
  XOR2_X1   g410(.A(new_n600), .B(KEYINPUT13), .Z(new_n612));
  NAND2_X1  g411(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NAND4_X1  g412(.A1(new_n605), .A2(KEYINPUT90), .A3(new_n610), .A4(new_n613), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(new_n603), .A3(new_n610), .A4(new_n604), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT90), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n605), .A2(new_n613), .ZN(new_n619));
  INV_X1    g418(.A(new_n610), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n618), .A2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n597), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n451), .A2(new_n527), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT98), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n409), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n627), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g427(.A1(new_n626), .A2(new_n407), .ZN(new_n629));
  NAND2_X1  g428(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n630));
  OR2_X1    g429(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n629), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(KEYINPUT42), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n629), .A2(KEYINPUT42), .A3(new_n630), .A4(new_n631), .ZN(new_n635));
  OAI211_X1 g434(.A(new_n634), .B(new_n635), .C1(new_n341), .C2(new_n629), .ZN(G1325gat));
  INV_X1    g435(.A(new_n439), .ZN(new_n637));
  AOI21_X1  g436(.A(G15gat), .B1(new_n626), .B2(new_n637), .ZN(new_n638));
  AND2_X1   g437(.A1(new_n626), .A2(G15gat), .ZN(new_n639));
  AOI21_X1  g438(.A(new_n638), .B1(new_n440), .B2(new_n639), .ZN(G1326gat));
  NAND2_X1  g439(.A1(new_n626), .A2(new_n398), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT43), .B(G22gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n596), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n451), .A2(new_n644), .ZN(new_n645));
  NOR3_X1   g444(.A1(new_n563), .A2(new_n623), .A3(new_n526), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n645), .A2(new_n647), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n572), .A3(new_n409), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(KEYINPUT45), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n443), .A2(new_n446), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n449), .A2(new_n445), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n653), .A2(KEYINPUT99), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT99), .ZN(new_n655));
  NAND3_X1  g454(.A1(new_n651), .A2(new_n652), .A3(new_n655), .ZN(new_n656));
  NAND3_X1  g455(.A1(new_n654), .A2(new_n442), .A3(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(KEYINPUT44), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n657), .A2(new_n658), .A3(new_n644), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n645), .A2(KEYINPUT44), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n647), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n409), .ZN(new_n663));
  OAI21_X1  g462(.A(G29gat), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n650), .A2(new_n664), .ZN(G1328gat));
  NAND3_X1  g464(.A1(new_n648), .A2(new_n573), .A3(new_n407), .ZN(new_n666));
  XOR2_X1   g465(.A(new_n666), .B(KEYINPUT46), .Z(new_n667));
  INV_X1    g466(.A(new_n407), .ZN(new_n668));
  OAI21_X1  g467(.A(G36gat), .B1(new_n662), .B2(new_n668), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n667), .A2(new_n669), .ZN(G1329gat));
  AOI21_X1  g469(.A(new_n596), .B1(new_n442), .B2(new_n450), .ZN(new_n671));
  INV_X1    g470(.A(G43gat), .ZN(new_n672));
  NAND4_X1  g471(.A1(new_n671), .A2(new_n672), .A3(new_n637), .A4(new_n646), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT100), .ZN(new_n674));
  OR2_X1    g473(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n441), .B(new_n647), .C1(new_n659), .C2(new_n660), .ZN(new_n678));
  OAI21_X1  g477(.A(new_n677), .B1(new_n678), .B2(new_n672), .ZN(new_n679));
  INV_X1    g478(.A(KEYINPUT47), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n679), .A2(KEYINPUT101), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(KEYINPUT101), .B1(new_n679), .B2(new_n680), .ZN(new_n682));
  INV_X1    g481(.A(KEYINPUT102), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n659), .A2(new_n660), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n684), .A2(new_n440), .A3(new_n646), .ZN(new_n685));
  AOI22_X1  g484(.A1(new_n685), .A2(G43gat), .B1(new_n676), .B2(new_n675), .ZN(new_n686));
  AOI21_X1  g485(.A(new_n683), .B1(new_n686), .B2(KEYINPUT47), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n672), .B1(new_n661), .B2(new_n440), .ZN(new_n688));
  XNOR2_X1  g487(.A(new_n673), .B(KEYINPUT100), .ZN(new_n689));
  NOR4_X1   g488(.A1(new_n688), .A2(new_n689), .A3(KEYINPUT102), .A4(new_n680), .ZN(new_n690));
  OAI22_X1  g489(.A1(new_n681), .A2(new_n682), .B1(new_n687), .B2(new_n690), .ZN(G1330gat));
  NOR2_X1   g490(.A1(new_n662), .A2(new_n399), .ZN(new_n692));
  INV_X1    g491(.A(new_n648), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n398), .A2(new_n565), .ZN(new_n694));
  XOR2_X1   g493(.A(new_n694), .B(KEYINPUT103), .Z(new_n695));
  OAI22_X1  g494(.A1(new_n692), .A2(new_n565), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT48), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  OAI221_X1 g497(.A(KEYINPUT48), .B1(new_n693), .B2(new_n695), .C1(new_n692), .C2(new_n565), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(G1331gat));
  NOR2_X1   g499(.A1(new_n597), .A2(new_n622), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n657), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n702), .A2(new_n526), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(new_n409), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(G57gat), .ZN(G1332gat));
  AOI211_X1 g505(.A(new_n668), .B(new_n703), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(G1333gat));
  XNOR2_X1  g508(.A(new_n439), .B(KEYINPUT104), .ZN(new_n710));
  OAI21_X1  g509(.A(new_n456), .B1(new_n703), .B2(new_n710), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n440), .A2(G71gat), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n711), .B1(new_n703), .B2(new_n712), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n713), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g513(.A1(new_n703), .A2(new_n399), .ZN(new_n715));
  XNOR2_X1  g514(.A(new_n715), .B(new_n457), .ZN(G1335gat));
  INV_X1    g515(.A(new_n563), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n623), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n684), .A2(new_n526), .A3(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(new_n479), .A3(new_n663), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n657), .A2(new_n644), .A3(new_n719), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT51), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n722), .A2(new_n723), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n527), .B1(new_n724), .B2(new_n725), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(new_n409), .ZN(new_n727));
  AOI21_X1  g526(.A(new_n721), .B1(new_n727), .B2(new_n479), .ZN(G1336gat));
  NAND2_X1  g527(.A1(new_n724), .A2(new_n725), .ZN(new_n729));
  NOR3_X1   g528(.A1(new_n668), .A2(G92gat), .A3(new_n527), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT106), .B1(new_n729), .B2(new_n730), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT106), .ZN(new_n732));
  INV_X1    g531(.A(new_n730), .ZN(new_n733));
  AOI211_X1 g532(.A(new_n732), .B(new_n733), .C1(new_n724), .C2(new_n725), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  NAND4_X1  g534(.A1(new_n684), .A2(new_n526), .A3(new_n407), .A4(new_n719), .ZN(new_n736));
  INV_X1    g535(.A(new_n478), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  INV_X1    g537(.A(KEYINPUT52), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n730), .B(KEYINPUT105), .Z(new_n741));
  AOI22_X1  g540(.A1(new_n729), .A2(new_n741), .B1(new_n736), .B2(new_n737), .ZN(new_n742));
  OAI22_X1  g541(.A1(new_n735), .A2(new_n740), .B1(new_n739), .B2(new_n742), .ZN(G1337gat));
  NOR3_X1   g542(.A1(new_n720), .A2(new_n413), .A3(new_n441), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n726), .A2(new_n637), .ZN(new_n745));
  AOI21_X1  g544(.A(new_n744), .B1(new_n745), .B2(new_n413), .ZN(G1338gat));
  INV_X1    g545(.A(G106gat), .ZN(new_n747));
  NAND4_X1  g546(.A1(new_n729), .A2(new_n747), .A3(new_n526), .A4(new_n398), .ZN(new_n748));
  OAI21_X1  g547(.A(G106gat), .B1(new_n720), .B2(new_n399), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT53), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1339gat));
  OR2_X1    g553(.A1(new_n523), .A2(new_n452), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n514), .A2(KEYINPUT54), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(KEYINPUT107), .B(KEYINPUT54), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n521), .B1(new_n524), .B2(new_n757), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT55), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT109), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  AOI21_X1  g562(.A(KEYINPUT55), .B1(new_n756), .B2(new_n758), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT109), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n756), .A2(KEYINPUT55), .A3(new_n758), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(KEYINPUT108), .ZN(new_n768));
  INV_X1    g567(.A(KEYINPUT108), .ZN(new_n769));
  NAND4_X1  g568(.A1(new_n756), .A2(new_n769), .A3(KEYINPUT55), .A4(new_n758), .ZN(new_n770));
  NAND3_X1  g569(.A1(new_n768), .A2(new_n522), .A3(new_n770), .ZN(new_n771));
  NOR3_X1   g570(.A1(new_n766), .A2(new_n623), .A3(new_n771), .ZN(new_n772));
  INV_X1    g571(.A(new_n609), .ZN(new_n773));
  NOR2_X1   g572(.A1(new_n611), .A2(new_n612), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n600), .B1(new_n598), .B2(new_n599), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n774), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n618), .A2(new_n526), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n596), .B1(new_n772), .B2(new_n778), .ZN(new_n779));
  INV_X1    g578(.A(new_n771), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n764), .B(new_n762), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n618), .A2(new_n776), .ZN(new_n782));
  INV_X1    g581(.A(new_n782), .ZN(new_n783));
  NAND4_X1  g582(.A1(new_n780), .A2(new_n781), .A3(new_n644), .A4(new_n783), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n563), .B1(new_n779), .B2(new_n784), .ZN(new_n785));
  NOR3_X1   g584(.A1(new_n597), .A2(new_n526), .A3(new_n622), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR4_X1   g586(.A1(new_n787), .A2(new_n663), .A3(new_n444), .A4(new_n407), .ZN(new_n788));
  INV_X1    g587(.A(new_n788), .ZN(new_n789));
  OAI21_X1  g588(.A(G113gat), .B1(new_n789), .B2(new_n623), .ZN(new_n790));
  NOR2_X1   g589(.A1(new_n623), .A2(G113gat), .ZN(new_n791));
  XNOR2_X1  g590(.A(new_n791), .B(KEYINPUT110), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n789), .B2(new_n792), .ZN(G1340gat));
  AOI21_X1  g592(.A(new_n210), .B1(new_n788), .B2(new_n526), .ZN(new_n794));
  XNOR2_X1  g593(.A(new_n794), .B(KEYINPUT111), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n526), .A2(new_n210), .ZN(new_n796));
  XOR2_X1   g595(.A(new_n796), .B(KEYINPUT112), .Z(new_n797));
  OAI21_X1  g596(.A(new_n795), .B1(new_n789), .B2(new_n797), .ZN(G1341gat));
  NAND2_X1  g597(.A1(new_n788), .A2(new_n563), .ZN(new_n799));
  XNOR2_X1  g598(.A(new_n799), .B(G127gat), .ZN(G1342gat));
  NAND2_X1  g599(.A1(new_n788), .A2(new_n644), .ZN(new_n801));
  OR3_X1    g600(.A1(new_n801), .A2(KEYINPUT56), .A3(G134gat), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(G134gat), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT56), .B1(new_n801), .B2(G134gat), .ZN(new_n804));
  NAND3_X1  g603(.A1(new_n802), .A2(new_n803), .A3(new_n804), .ZN(G1343gat));
  NAND2_X1  g604(.A1(new_n779), .A2(new_n784), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n806), .A2(new_n717), .ZN(new_n807));
  INV_X1    g606(.A(new_n786), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(KEYINPUT57), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n809), .A2(new_n810), .A3(new_n398), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n764), .B1(new_n618), .B2(new_n621), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n778), .B1(new_n780), .B2(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n784), .B1(new_n813), .B2(new_n644), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n786), .B1(new_n814), .B2(new_n717), .ZN(new_n815));
  OAI21_X1  g614(.A(KEYINPUT57), .B1(new_n815), .B2(new_n399), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n440), .A2(new_n663), .A3(new_n407), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n811), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  OAI21_X1  g617(.A(G141gat), .B1(new_n818), .B2(new_n623), .ZN(new_n819));
  INV_X1    g618(.A(KEYINPUT58), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n819), .B1(KEYINPUT113), .B2(new_n820), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n787), .A2(KEYINPUT114), .A3(new_n663), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(KEYINPUT114), .B1(new_n787), .B2(new_n663), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n407), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n441), .A2(new_n398), .ZN(new_n826));
  XOR2_X1   g625(.A(new_n826), .B(KEYINPUT115), .Z(new_n827));
  NAND4_X1  g626(.A1(new_n825), .A2(new_n221), .A3(new_n622), .A4(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT116), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n821), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  INV_X1    g629(.A(KEYINPUT114), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n831), .B1(new_n809), .B2(new_n409), .ZN(new_n832));
  OAI211_X1 g631(.A(new_n668), .B(new_n827), .C1(new_n832), .C2(new_n822), .ZN(new_n833));
  NOR3_X1   g632(.A1(new_n833), .A2(G141gat), .A3(new_n623), .ZN(new_n834));
  OAI22_X1  g633(.A1(new_n834), .A2(KEYINPUT116), .B1(KEYINPUT113), .B2(new_n819), .ZN(new_n835));
  OAI21_X1  g634(.A(KEYINPUT58), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  OR2_X1    g635(.A1(new_n821), .A2(new_n834), .ZN(new_n837));
  NAND2_X1  g636(.A1(new_n836), .A2(new_n837), .ZN(G1344gat));
  INV_X1    g637(.A(KEYINPUT119), .ZN(new_n839));
  NAND4_X1  g638(.A1(new_n811), .A2(new_n816), .A3(new_n526), .A4(new_n817), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT59), .ZN(new_n841));
  AND3_X1   g640(.A1(new_n840), .A2(new_n841), .A3(new_n223), .ZN(new_n842));
  INV_X1    g641(.A(KEYINPUT117), .ZN(new_n843));
  NAND4_X1  g642(.A1(new_n812), .A2(new_n522), .A3(new_n768), .A4(new_n770), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n644), .B1(new_n844), .B2(new_n777), .ZN(new_n845));
  NOR4_X1   g644(.A1(new_n766), .A2(new_n771), .A3(new_n596), .A4(new_n782), .ZN(new_n846));
  OAI21_X1  g645(.A(new_n717), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n399), .B1(new_n847), .B2(new_n808), .ZN(new_n848));
  OAI21_X1  g647(.A(new_n843), .B1(new_n848), .B2(KEYINPUT57), .ZN(new_n849));
  OAI211_X1 g648(.A(KEYINPUT57), .B(new_n398), .C1(new_n785), .C2(new_n786), .ZN(new_n850));
  OAI211_X1 g649(.A(KEYINPUT117), .B(new_n810), .C1(new_n815), .C2(new_n399), .ZN(new_n851));
  NAND3_X1  g650(.A1(new_n849), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n852), .A2(new_n526), .A3(new_n817), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g654(.A1(new_n852), .A2(KEYINPUT118), .A3(new_n526), .A4(new_n817), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(G148gat), .A3(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n842), .B1(new_n857), .B2(KEYINPUT59), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n833), .A2(new_n223), .A3(new_n527), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n839), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(new_n859), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n234), .B1(new_n853), .B2(new_n854), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n841), .B1(new_n862), .B2(new_n856), .ZN(new_n863));
  OAI211_X1 g662(.A(KEYINPUT119), .B(new_n861), .C1(new_n863), .C2(new_n842), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n860), .A2(new_n864), .ZN(G1345gat));
  NOR3_X1   g664(.A1(new_n818), .A2(new_n226), .A3(new_n717), .ZN(new_n866));
  INV_X1    g665(.A(new_n833), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n563), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n866), .B1(new_n868), .B2(new_n226), .ZN(G1346gat));
  NOR3_X1   g668(.A1(new_n818), .A2(new_n225), .A3(new_n596), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n867), .A2(new_n644), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n870), .B1(new_n871), .B2(new_n225), .ZN(G1347gat));
  NOR2_X1   g671(.A1(new_n668), .A2(new_n409), .ZN(new_n873));
  NOR2_X1   g672(.A1(new_n710), .A2(new_n398), .ZN(new_n874));
  NAND3_X1  g673(.A1(new_n809), .A2(new_n873), .A3(new_n874), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n875), .A2(new_n623), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT121), .ZN(new_n877));
  AND3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(G169gat), .ZN(new_n878));
  AOI21_X1  g677(.A(new_n877), .B1(new_n876), .B2(G169gat), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT120), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n809), .A2(new_n880), .A3(new_n663), .ZN(new_n881));
  OAI21_X1  g680(.A(KEYINPUT120), .B1(new_n787), .B2(new_n409), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n883), .A2(new_n447), .A3(new_n407), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n622), .A2(new_n283), .ZN(new_n885));
  OAI22_X1  g684(.A1(new_n878), .A2(new_n879), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT122), .ZN(new_n887));
  XNOR2_X1  g686(.A(new_n886), .B(new_n887), .ZN(G1348gat));
  NOR3_X1   g687(.A1(new_n875), .A2(new_n284), .A3(new_n527), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n444), .B1(new_n881), .B2(new_n882), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n890), .A2(new_n526), .A3(new_n407), .ZN(new_n891));
  AOI21_X1  g690(.A(new_n889), .B1(new_n891), .B2(new_n284), .ZN(G1349gat));
  INV_X1    g691(.A(KEYINPUT123), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n563), .A2(new_n291), .ZN(new_n894));
  OAI21_X1  g693(.A(new_n893), .B1(new_n884), .B2(new_n894), .ZN(new_n895));
  INV_X1    g694(.A(new_n894), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n890), .A2(KEYINPUT123), .A3(new_n407), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  OAI21_X1  g697(.A(G183gat), .B1(new_n875), .B2(new_n717), .ZN(new_n899));
  NAND2_X1  g698(.A1(new_n898), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n900), .A2(KEYINPUT60), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT60), .ZN(new_n902));
  NAND3_X1  g701(.A1(new_n898), .A2(new_n902), .A3(new_n899), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n901), .A2(new_n903), .ZN(G1350gat));
  NOR2_X1   g703(.A1(new_n596), .A2(G190gat), .ZN(new_n905));
  INV_X1    g704(.A(new_n905), .ZN(new_n906));
  OAI21_X1  g705(.A(KEYINPUT124), .B1(new_n884), .B2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(KEYINPUT124), .ZN(new_n908));
  NAND4_X1  g707(.A1(new_n890), .A2(new_n908), .A3(new_n407), .A4(new_n905), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n907), .A2(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(G190gat), .B1(new_n875), .B2(new_n596), .ZN(new_n911));
  XNOR2_X1  g710(.A(new_n911), .B(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n913), .A2(KEYINPUT125), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT125), .ZN(new_n915));
  NAND3_X1  g714(.A1(new_n910), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n914), .A2(new_n916), .ZN(G1351gat));
  NOR3_X1   g716(.A1(new_n440), .A2(new_n668), .A3(new_n409), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n852), .A2(new_n622), .A3(new_n918), .ZN(new_n919));
  XNOR2_X1  g718(.A(KEYINPUT126), .B(G197gat), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n826), .B1(new_n881), .B2(new_n882), .ZN(new_n922));
  AND2_X1   g721(.A1(new_n922), .A2(new_n407), .ZN(new_n923));
  INV_X1    g722(.A(new_n923), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n623), .A2(new_n920), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1352gat));
  INV_X1    g725(.A(KEYINPUT62), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n923), .A2(new_n927), .A3(new_n519), .A4(new_n526), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n852), .A2(new_n526), .A3(new_n918), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(G204gat), .ZN(new_n930));
  NAND4_X1  g729(.A1(new_n922), .A2(new_n519), .A3(new_n526), .A4(new_n407), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT62), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT127), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NAND4_X1  g734(.A1(new_n928), .A2(KEYINPUT127), .A3(new_n930), .A4(new_n932), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1353gat));
  NAND3_X1  g736(.A1(new_n923), .A2(new_n321), .A3(new_n563), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n852), .A2(new_n563), .A3(new_n918), .ZN(new_n939));
  AND3_X1   g738(.A1(new_n939), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n940));
  AOI21_X1  g739(.A(KEYINPUT63), .B1(new_n939), .B2(G211gat), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n938), .B1(new_n940), .B2(new_n941), .ZN(G1354gat));
  NAND3_X1  g741(.A1(new_n923), .A2(new_n322), .A3(new_n644), .ZN(new_n943));
  AND3_X1   g742(.A1(new_n852), .A2(new_n644), .A3(new_n918), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n943), .B1(new_n322), .B2(new_n944), .ZN(G1355gat));
endmodule


