//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 0 1 1 0 0 1 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:08 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n592, new_n593, new_n594,
    new_n595, new_n596, new_n597, new_n598, new_n599, new_n601, new_n602,
    new_n603, new_n604, new_n605, new_n606, new_n607, new_n609, new_n610,
    new_n611, new_n612, new_n613, new_n614, new_n615, new_n616, new_n617,
    new_n618, new_n619, new_n620, new_n621, new_n622, new_n623, new_n624,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n650, new_n651, new_n652, new_n653, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n664, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n922, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000;
  INV_X1    g000(.A(G146), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G143), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT64), .B(G146), .ZN(new_n190));
  INV_X1    g004(.A(G143), .ZN(new_n191));
  AOI21_X1  g005(.A(new_n189), .B1(new_n190), .B2(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT0), .B(G128), .ZN(new_n193));
  NOR2_X1   g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT64), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT64), .A2(G146), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n195), .A2(G143), .A3(new_n196), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n187), .A2(G143), .ZN(new_n198));
  INV_X1    g012(.A(new_n198), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(KEYINPUT0), .A2(G128), .ZN(new_n201));
  NOR2_X1   g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n194), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G134), .ZN(new_n204));
  OAI21_X1  g018(.A(KEYINPUT11), .B1(new_n204), .B2(G137), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT11), .ZN(new_n206));
  INV_X1    g020(.A(G137), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n206), .A2(new_n207), .A3(G134), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n205), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(KEYINPUT65), .B1(new_n207), .B2(G134), .ZN(new_n210));
  OR3_X1    g024(.A1(new_n207), .A2(KEYINPUT65), .A3(G134), .ZN(new_n211));
  NAND3_X1  g025(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G131), .ZN(new_n213));
  INV_X1    g027(.A(G131), .ZN(new_n214));
  NAND4_X1  g028(.A1(new_n209), .A2(new_n214), .A3(new_n211), .A4(new_n210), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n207), .B2(G134), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n207), .A2(G134), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NOR3_X1   g033(.A1(new_n207), .A2(KEYINPUT66), .A3(G134), .ZN(new_n220));
  OAI21_X1  g034(.A(G131), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  AND2_X1   g035(.A1(new_n215), .A2(new_n221), .ZN(new_n222));
  XNOR2_X1  g036(.A(KEYINPUT67), .B(KEYINPUT1), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n197), .A2(G128), .A3(new_n223), .A4(new_n199), .ZN(new_n224));
  XNOR2_X1  g038(.A(KEYINPUT68), .B(G128), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT1), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n226), .A2(KEYINPUT67), .ZN(new_n227));
  INV_X1    g041(.A(KEYINPUT67), .ZN(new_n228));
  NAND2_X1  g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n227), .A2(new_n229), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n225), .B1(new_n197), .B2(new_n230), .ZN(new_n231));
  OAI21_X1  g045(.A(new_n224), .B1(new_n231), .B2(new_n192), .ZN(new_n232));
  AOI22_X1  g046(.A1(new_n203), .A2(new_n216), .B1(new_n222), .B2(new_n232), .ZN(new_n233));
  XOR2_X1   g047(.A(KEYINPUT2), .B(G113), .Z(new_n234));
  XNOR2_X1  g048(.A(G116), .B(G119), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n234), .B(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n233), .A2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(new_n238), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n203), .A2(new_n216), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n222), .A2(new_n232), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT69), .A3(KEYINPUT30), .ZN(new_n243));
  OR2_X1    g057(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n244));
  NAND2_X1  g058(.A1(KEYINPUT69), .A2(KEYINPUT30), .ZN(new_n245));
  NAND3_X1  g059(.A1(new_n233), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n243), .A2(new_n246), .ZN(new_n247));
  AOI21_X1  g061(.A(new_n239), .B1(new_n247), .B2(new_n236), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT31), .ZN(new_n249));
  INV_X1    g063(.A(G237), .ZN(new_n250));
  INV_X1    g064(.A(G953), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n250), .A2(new_n251), .A3(G210), .ZN(new_n252));
  XOR2_X1   g066(.A(new_n252), .B(KEYINPUT27), .Z(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT26), .B(G101), .ZN(new_n254));
  XNOR2_X1  g068(.A(new_n253), .B(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n248), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  AOI211_X1 g071(.A(new_n239), .B(new_n255), .C1(new_n247), .C2(new_n236), .ZN(new_n258));
  NOR2_X1   g072(.A1(KEYINPUT70), .A2(KEYINPUT28), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n238), .A2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(KEYINPUT28), .ZN(new_n261));
  OAI21_X1  g075(.A(new_n236), .B1(new_n242), .B2(new_n261), .ZN(new_n262));
  OAI211_X1 g076(.A(new_n233), .B(new_n237), .C1(KEYINPUT70), .C2(KEYINPUT28), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  AOI21_X1  g078(.A(KEYINPUT31), .B1(new_n264), .B2(new_n255), .ZN(new_n265));
  OAI21_X1  g079(.A(new_n257), .B1(new_n258), .B2(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n266), .A2(KEYINPUT71), .ZN(new_n267));
  NOR2_X1   g081(.A1(G472), .A2(G902), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n269));
  OAI211_X1 g083(.A(new_n257), .B(new_n269), .C1(new_n258), .C2(new_n265), .ZN(new_n270));
  NAND3_X1  g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT32), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  OR2_X1    g087(.A1(new_n264), .A2(new_n255), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT29), .ZN(new_n275));
  NOR2_X1   g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NOR2_X1   g090(.A1(new_n276), .A2(G902), .ZN(new_n277));
  INV_X1    g091(.A(new_n248), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(new_n255), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n279), .A2(new_n275), .A3(new_n274), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n277), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G472), .ZN(new_n282));
  NAND4_X1  g096(.A1(new_n267), .A2(KEYINPUT32), .A3(new_n268), .A4(new_n270), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n273), .A2(new_n282), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT76), .ZN(new_n285));
  XNOR2_X1  g099(.A(G125), .B(G140), .ZN(new_n286));
  INV_X1    g100(.A(KEYINPUT72), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G140), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n289), .A2(KEYINPUT72), .A3(G125), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n288), .A2(KEYINPUT16), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT16), .ZN(new_n292));
  INV_X1    g106(.A(G125), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n292), .B1(new_n293), .B2(G140), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n291), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(G146), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n291), .A2(new_n187), .A3(new_n294), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n225), .A2(KEYINPUT23), .A3(G119), .ZN(new_n299));
  INV_X1    g113(.A(G128), .ZN(new_n300));
  AOI21_X1  g114(.A(KEYINPUT23), .B1(new_n300), .B2(G119), .ZN(new_n301));
  NOR2_X1   g115(.A1(new_n300), .A2(G119), .ZN(new_n302));
  NOR2_X1   g116(.A1(new_n301), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n299), .A2(new_n303), .ZN(new_n304));
  AOI21_X1  g118(.A(new_n302), .B1(new_n225), .B2(G119), .ZN(new_n305));
  XOR2_X1   g119(.A(KEYINPUT24), .B(G110), .Z(new_n306));
  AOI22_X1  g120(.A1(new_n304), .A2(G110), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n298), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g122(.A(KEYINPUT73), .B(G110), .ZN(new_n309));
  OAI22_X1  g123(.A1(new_n304), .A2(new_n309), .B1(new_n305), .B2(new_n306), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n286), .A2(new_n195), .A3(new_n196), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n296), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n308), .A2(new_n312), .ZN(new_n313));
  XNOR2_X1  g127(.A(KEYINPUT22), .B(G137), .ZN(new_n314));
  INV_X1    g128(.A(G221), .ZN(new_n315));
  INV_X1    g129(.A(G234), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(G953), .ZN(new_n317));
  XOR2_X1   g131(.A(new_n314), .B(new_n317), .Z(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(G902), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n308), .A2(new_n312), .A3(new_n318), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  AND3_X1   g137(.A1(new_n323), .A2(KEYINPUT74), .A3(KEYINPUT25), .ZN(new_n324));
  AOI21_X1  g138(.A(KEYINPUT25), .B1(new_n323), .B2(KEYINPUT74), .ZN(new_n325));
  OAI21_X1  g139(.A(G217), .B1(new_n316), .B2(G902), .ZN(new_n326));
  NOR3_X1   g140(.A1(new_n324), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n321), .ZN(new_n328));
  INV_X1    g142(.A(new_n322), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n318), .B1(new_n308), .B2(new_n312), .ZN(new_n330));
  NOR2_X1   g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT75), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(KEYINPUT75), .B1(new_n329), .B2(new_n330), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n328), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n285), .B1(new_n327), .B2(new_n335), .ZN(new_n336));
  NOR2_X1   g150(.A1(new_n325), .A2(new_n326), .ZN(new_n337));
  INV_X1    g151(.A(new_n324), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g153(.A(new_n335), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n339), .A2(new_n340), .A3(KEYINPUT76), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n336), .A2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  XNOR2_X1  g157(.A(G110), .B(G140), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n251), .A2(G227), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n344), .B(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT77), .ZN(new_n347));
  INV_X1    g161(.A(G107), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n347), .A2(new_n348), .A3(G104), .ZN(new_n349));
  INV_X1    g163(.A(G104), .ZN(new_n350));
  OAI21_X1  g164(.A(KEYINPUT77), .B1(new_n350), .B2(G107), .ZN(new_n351));
  NOR2_X1   g165(.A1(new_n348), .A2(G104), .ZN(new_n352));
  OAI211_X1 g166(.A(G101), .B(new_n349), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(KEYINPUT3), .B1(new_n350), .B2(G107), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT3), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n348), .A3(G104), .ZN(new_n356));
  INV_X1    g170(.A(G101), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n350), .A2(G107), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n354), .A2(new_n356), .A3(new_n357), .A4(new_n358), .ZN(new_n359));
  AND2_X1   g173(.A1(new_n353), .A2(new_n359), .ZN(new_n360));
  AND4_X1   g174(.A1(G128), .A2(new_n197), .A3(new_n199), .A4(new_n223), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n188), .A2(KEYINPUT1), .ZN(new_n362));
  AOI22_X1  g176(.A1(new_n197), .A2(new_n199), .B1(new_n362), .B2(G128), .ZN(new_n363));
  OAI21_X1  g177(.A(new_n360), .B1(new_n361), .B2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT10), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n353), .A2(new_n359), .ZN(new_n367));
  INV_X1    g181(.A(KEYINPUT78), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n353), .A2(new_n359), .A3(KEYINPUT78), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n232), .A2(new_n369), .A3(KEYINPUT10), .A4(new_n370), .ZN(new_n371));
  OR2_X1    g185(.A1(new_n192), .A2(new_n193), .ZN(new_n372));
  OR2_X1    g186(.A1(new_n200), .A2(new_n201), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n354), .A2(new_n356), .A3(new_n358), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n374), .A2(G101), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n375), .A2(KEYINPUT4), .A3(new_n359), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT4), .ZN(new_n377));
  NAND3_X1  g191(.A1(new_n374), .A2(new_n377), .A3(G101), .ZN(new_n378));
  NAND4_X1  g192(.A1(new_n372), .A2(new_n373), .A3(new_n376), .A4(new_n378), .ZN(new_n379));
  AND3_X1   g193(.A1(new_n366), .A2(new_n371), .A3(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n216), .ZN(new_n381));
  NOR2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND4_X1  g196(.A1(new_n366), .A2(new_n371), .A3(new_n379), .A4(new_n381), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n346), .B1(new_n382), .B2(new_n384), .ZN(new_n385));
  INV_X1    g199(.A(new_n346), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n383), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n362), .A2(G128), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n200), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g203(.A(new_n367), .B1(new_n389), .B2(new_n224), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n369), .A2(new_n370), .ZN(new_n391));
  INV_X1    g205(.A(new_n232), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n390), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT12), .ZN(new_n394));
  NOR3_X1   g208(.A1(new_n393), .A2(new_n394), .A3(new_n381), .ZN(new_n395));
  AND3_X1   g209(.A1(new_n353), .A2(new_n359), .A3(KEYINPUT78), .ZN(new_n396));
  AOI21_X1  g210(.A(KEYINPUT78), .B1(new_n353), .B2(new_n359), .ZN(new_n397));
  NOR2_X1   g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n364), .B1(new_n398), .B2(new_n232), .ZN(new_n399));
  AOI21_X1  g213(.A(KEYINPUT12), .B1(new_n399), .B2(new_n216), .ZN(new_n400));
  NOR2_X1   g214(.A1(new_n395), .A2(new_n400), .ZN(new_n401));
  OAI21_X1  g215(.A(new_n385), .B1(new_n387), .B2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(G469), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(new_n403), .A3(new_n321), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n403), .A2(new_n321), .ZN(new_n405));
  INV_X1    g219(.A(new_n405), .ZN(new_n406));
  OR2_X1    g220(.A1(new_n380), .A2(new_n381), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT80), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n387), .A2(new_n408), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n383), .A2(KEYINPUT80), .A3(new_n386), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n407), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n394), .B1(new_n393), .B2(new_n381), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n399), .A2(KEYINPUT12), .A3(new_n216), .ZN(new_n413));
  AOI22_X1  g227(.A1(new_n412), .A2(new_n413), .B1(new_n380), .B2(new_n381), .ZN(new_n414));
  INV_X1    g228(.A(KEYINPUT79), .ZN(new_n415));
  OAI21_X1  g229(.A(new_n346), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  OAI211_X1 g230(.A(new_n415), .B(new_n383), .C1(new_n395), .C2(new_n400), .ZN(new_n417));
  INV_X1    g231(.A(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n411), .B1(new_n416), .B2(new_n418), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n404), .B(new_n406), .C1(new_n419), .C2(new_n403), .ZN(new_n420));
  XNOR2_X1  g234(.A(KEYINPUT9), .B(G234), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n315), .B1(new_n422), .B2(new_n321), .ZN(new_n423));
  INV_X1    g237(.A(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n420), .A2(new_n424), .ZN(new_n425));
  NOR2_X1   g239(.A1(G475), .A2(G902), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n288), .A2(G146), .A3(new_n290), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n427), .A2(new_n311), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n250), .A2(new_n251), .A3(G214), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(new_n191), .ZN(new_n430));
  AND2_X1   g244(.A1(KEYINPUT18), .A2(G131), .ZN(new_n431));
  AND3_X1   g245(.A1(new_n430), .A2(KEYINPUT85), .A3(new_n431), .ZN(new_n432));
  AOI21_X1  g246(.A(KEYINPUT85), .B1(new_n430), .B2(new_n431), .ZN(new_n433));
  OAI221_X1 g247(.A(new_n428), .B1(new_n430), .B2(new_n431), .C1(new_n432), .C2(new_n433), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(G131), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n429), .B(G143), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n436), .A2(new_n214), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT17), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n435), .A2(new_n437), .A3(new_n438), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n430), .A2(KEYINPUT17), .A3(G131), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n439), .A2(new_n296), .A3(new_n297), .A4(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G113), .B(G122), .ZN(new_n442));
  XNOR2_X1  g256(.A(new_n442), .B(new_n350), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n434), .A2(new_n441), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n435), .A2(new_n437), .ZN(new_n445));
  NOR2_X1   g259(.A1(new_n286), .A2(KEYINPUT19), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n288), .A2(new_n290), .ZN(new_n447));
  AOI21_X1  g261(.A(new_n446), .B1(new_n447), .B2(KEYINPUT19), .ZN(new_n448));
  OAI211_X1 g262(.A(new_n296), .B(new_n445), .C1(new_n190), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g263(.A(new_n443), .B1(new_n434), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n426), .B1(new_n444), .B2(new_n450), .ZN(new_n451));
  XOR2_X1   g265(.A(KEYINPUT84), .B(KEYINPUT20), .Z(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n451), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  OAI211_X1 g269(.A(new_n455), .B(new_n426), .C1(new_n444), .C2(new_n450), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n443), .B1(new_n434), .B2(new_n441), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n321), .B1(new_n444), .B2(new_n457), .ZN(new_n458));
  AOI22_X1  g272(.A1(new_n454), .A2(new_n456), .B1(G475), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(G234), .A2(G237), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n460), .A2(G952), .A3(new_n251), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  NAND3_X1  g276(.A1(new_n460), .A2(G902), .A3(G953), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  XNOR2_X1  g278(.A(KEYINPUT21), .B(G898), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT86), .ZN(new_n468));
  XNOR2_X1  g282(.A(G116), .B(G122), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n469), .A2(new_n348), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT14), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(G122), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n473), .A2(G116), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n348), .B1(new_n474), .B2(KEYINPUT14), .ZN(new_n475));
  AOI22_X1  g289(.A1(new_n468), .A2(new_n470), .B1(new_n472), .B2(new_n475), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n469), .A2(KEYINPUT86), .A3(new_n348), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n225), .A2(G143), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n191), .A2(G128), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n478), .A2(new_n204), .A3(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n204), .B1(new_n478), .B2(new_n479), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n476), .B(new_n477), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(new_n478), .ZN(new_n484));
  INV_X1    g298(.A(KEYINPUT13), .ZN(new_n485));
  XNOR2_X1  g299(.A(new_n479), .B(new_n485), .ZN(new_n486));
  OAI21_X1  g300(.A(G134), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  XNOR2_X1  g301(.A(new_n469), .B(new_n348), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n487), .A2(new_n480), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n422), .A2(G217), .A3(new_n251), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n483), .A2(new_n489), .A3(new_n491), .ZN(new_n492));
  INV_X1    g306(.A(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n491), .B1(new_n483), .B2(new_n489), .ZN(new_n494));
  OAI21_X1  g308(.A(new_n321), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(G478), .ZN(new_n496));
  NOR2_X1   g310(.A1(new_n496), .A2(KEYINPUT15), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n495), .B(new_n497), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n459), .A2(new_n467), .A3(new_n499), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n425), .A2(new_n500), .ZN(new_n501));
  OAI21_X1  g315(.A(G214), .B1(G237), .B2(G902), .ZN(new_n502));
  INV_X1    g316(.A(new_n502), .ZN(new_n503));
  OAI21_X1  g317(.A(G210), .B1(G237), .B2(G902), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n392), .A2(new_n293), .ZN(new_n506));
  OAI21_X1  g320(.A(G125), .B1(new_n194), .B2(new_n202), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n251), .A2(G224), .ZN(new_n509));
  XNOR2_X1  g323(.A(new_n508), .B(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT81), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT6), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n234), .A2(new_n235), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n235), .A2(KEYINPUT5), .ZN(new_n515));
  INV_X1    g329(.A(G119), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n516), .A2(G116), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n515), .B(G113), .C1(KEYINPUT5), .C2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n398), .A2(new_n514), .A3(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n236), .A2(new_n376), .A3(new_n378), .ZN(new_n520));
  XNOR2_X1  g334(.A(G110), .B(G122), .ZN(new_n521));
  AND3_X1   g335(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n521), .B1(new_n519), .B2(new_n520), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n513), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  AND2_X1   g338(.A1(new_n519), .A2(new_n520), .ZN(new_n525));
  OAI22_X1  g339(.A1(new_n525), .A2(new_n521), .B1(new_n511), .B2(new_n512), .ZN(new_n526));
  AOI21_X1  g340(.A(new_n510), .B1(new_n524), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(KEYINPUT83), .A2(KEYINPUT7), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n506), .A2(new_n507), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n509), .A2(KEYINPUT7), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  NAND3_X1  g345(.A1(new_n519), .A2(new_n520), .A3(new_n521), .ZN(new_n532));
  INV_X1    g346(.A(new_n530), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n506), .A2(new_n507), .A3(new_n533), .A4(new_n528), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  XNOR2_X1  g349(.A(new_n521), .B(KEYINPUT8), .ZN(new_n536));
  INV_X1    g350(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n518), .A2(new_n514), .ZN(new_n538));
  AOI22_X1  g352(.A1(new_n519), .A2(KEYINPUT82), .B1(new_n367), .B2(new_n538), .ZN(new_n539));
  OR3_X1    g353(.A1(new_n391), .A2(KEYINPUT82), .A3(new_n538), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n537), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n321), .B1(new_n535), .B2(new_n541), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n505), .B1(new_n527), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n524), .A2(new_n526), .ZN(new_n544));
  INV_X1    g358(.A(new_n510), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n531), .A2(new_n532), .A3(new_n534), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n519), .A2(KEYINPUT82), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n367), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n548), .A2(new_n540), .A3(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n536), .ZN(new_n551));
  AOI21_X1  g365(.A(G902), .B1(new_n547), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n546), .A2(new_n552), .A3(new_n504), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n503), .B1(new_n543), .B2(new_n553), .ZN(new_n554));
  NAND4_X1  g368(.A1(new_n284), .A2(new_n343), .A3(new_n501), .A4(new_n554), .ZN(new_n555));
  XNOR2_X1  g369(.A(KEYINPUT87), .B(G101), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n555), .B(new_n556), .ZN(G3));
  NOR2_X1   g371(.A1(new_n342), .A2(new_n425), .ZN(new_n558));
  AND2_X1   g372(.A1(new_n267), .A2(new_n270), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n267), .A2(new_n321), .A3(new_n270), .ZN(new_n560));
  AOI22_X1  g374(.A1(new_n559), .A2(new_n268), .B1(new_n560), .B2(G472), .ZN(new_n561));
  NAND2_X1  g375(.A1(new_n554), .A2(new_n467), .ZN(new_n562));
  NAND2_X1  g376(.A1(KEYINPUT88), .A2(KEYINPUT33), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n563), .B1(new_n493), .B2(new_n494), .ZN(new_n564));
  INV_X1    g378(.A(new_n494), .ZN(new_n565));
  XNOR2_X1  g379(.A(KEYINPUT88), .B(KEYINPUT33), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n565), .A2(new_n492), .A3(new_n566), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n496), .A2(G902), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n569), .A2(KEYINPUT89), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n495), .A2(new_n496), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT89), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n564), .A2(new_n567), .A3(new_n572), .A4(new_n568), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n562), .A2(new_n459), .A3(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n558), .A2(new_n561), .A3(new_n575), .ZN(new_n576));
  XOR2_X1   g390(.A(KEYINPUT34), .B(G104), .Z(new_n577));
  XNOR2_X1  g391(.A(new_n576), .B(new_n577), .ZN(G6));
  NAND2_X1  g392(.A1(new_n458), .A2(G475), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(KEYINPUT91), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n451), .A2(KEYINPUT90), .A3(new_n453), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT91), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n458), .A2(new_n582), .A3(G475), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n580), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT90), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n585), .B1(new_n451), .B2(new_n453), .ZN(new_n586));
  INV_X1    g400(.A(new_n426), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n434), .A2(new_n449), .ZN(new_n588));
  INV_X1    g402(.A(new_n443), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n434), .A2(new_n441), .A3(new_n443), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n587), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n592), .A2(new_n452), .ZN(new_n593));
  NOR2_X1   g407(.A1(new_n586), .A2(new_n593), .ZN(new_n594));
  NOR2_X1   g408(.A1(new_n584), .A2(new_n594), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n498), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n596), .A2(new_n562), .ZN(new_n597));
  NAND3_X1  g411(.A1(new_n558), .A2(new_n561), .A3(new_n597), .ZN(new_n598));
  XOR2_X1   g412(.A(KEYINPUT35), .B(G107), .Z(new_n599));
  XNOR2_X1  g413(.A(new_n598), .B(new_n599), .ZN(G9));
  NOR2_X1   g414(.A1(new_n319), .A2(KEYINPUT36), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n313), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(new_n321), .A3(new_n326), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n339), .A2(new_n603), .ZN(new_n604));
  NAND4_X1  g418(.A1(new_n561), .A2(new_n501), .A3(new_n554), .A4(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT37), .B(G110), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n606), .B(KEYINPUT92), .ZN(new_n607));
  XNOR2_X1  g421(.A(new_n605), .B(new_n607), .ZN(G12));
  INV_X1    g422(.A(new_n425), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n604), .A2(new_n554), .ZN(new_n610));
  XOR2_X1   g424(.A(new_n461), .B(KEYINPUT93), .Z(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  INV_X1    g426(.A(G900), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n612), .B1(new_n613), .B2(new_n464), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n595), .A2(new_n498), .A3(new_n615), .ZN(new_n616));
  NOR2_X1   g430(.A1(new_n610), .A2(new_n616), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n284), .A2(new_n609), .A3(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT94), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  AOI22_X1  g434(.A1(new_n271), .A2(new_n272), .B1(new_n281), .B2(G472), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n425), .B1(new_n621), .B2(new_n283), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(KEYINPUT94), .A3(new_n617), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n620), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g438(.A(new_n624), .B(G128), .ZN(G30));
  NOR2_X1   g439(.A1(new_n248), .A2(new_n255), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n238), .A2(new_n255), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n233), .A2(new_n237), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n321), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g443(.A(G472), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n273), .A2(new_n283), .A3(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT95), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT96), .B(KEYINPUT39), .ZN(new_n633));
  XOR2_X1   g447(.A(new_n614), .B(new_n633), .Z(new_n634));
  NAND3_X1  g448(.A1(new_n609), .A2(KEYINPUT97), .A3(new_n634), .ZN(new_n635));
  INV_X1    g449(.A(new_n635), .ZN(new_n636));
  AOI21_X1  g450(.A(KEYINPUT97), .B1(new_n609), .B2(new_n634), .ZN(new_n637));
  OAI21_X1  g451(.A(KEYINPUT40), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n637), .ZN(new_n639));
  INV_X1    g453(.A(KEYINPUT40), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n639), .A2(new_n640), .A3(new_n635), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n543), .A2(new_n553), .ZN(new_n642));
  XOR2_X1   g456(.A(new_n642), .B(KEYINPUT38), .Z(new_n643));
  NAND2_X1  g457(.A1(new_n498), .A2(new_n502), .ZN(new_n644));
  NOR2_X1   g458(.A1(new_n459), .A2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(new_n645), .ZN(new_n646));
  NOR3_X1   g460(.A1(new_n643), .A2(new_n604), .A3(new_n646), .ZN(new_n647));
  NAND4_X1  g461(.A1(new_n632), .A2(new_n638), .A3(new_n641), .A4(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(G143), .ZN(G45));
  NOR3_X1   g463(.A1(new_n574), .A2(new_n459), .A3(new_n614), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g465(.A1(new_n610), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n622), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(G146), .ZN(G48));
  AOI21_X1  g468(.A(new_n386), .B1(new_n407), .B2(new_n383), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n401), .A2(new_n387), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n321), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(G469), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n424), .A3(new_n404), .ZN(new_n659));
  INV_X1    g473(.A(new_n659), .ZN(new_n660));
  NAND4_X1  g474(.A1(new_n284), .A2(new_n343), .A3(new_n575), .A4(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(KEYINPUT41), .B(G113), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G15));
  NAND4_X1  g477(.A1(new_n284), .A2(new_n343), .A3(new_n597), .A4(new_n660), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G116), .ZN(G18));
  INV_X1    g479(.A(new_n554), .ZN(new_n666));
  NOR3_X1   g480(.A1(new_n666), .A2(new_n500), .A3(new_n659), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n284), .A2(new_n604), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n668), .B(G119), .ZN(G21));
  NAND2_X1  g483(.A1(new_n560), .A2(G472), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(KEYINPUT98), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n339), .A2(new_n340), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(KEYINPUT98), .ZN(new_n674));
  NAND3_X1  g488(.A1(new_n560), .A2(new_n674), .A3(G472), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n266), .A2(new_n268), .ZN(new_n676));
  NAND4_X1  g490(.A1(new_n671), .A2(new_n673), .A3(new_n675), .A4(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n642), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n646), .A2(new_n678), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n679), .A2(new_n467), .A3(new_n660), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n681), .B(new_n473), .ZN(G24));
  NAND2_X1  g496(.A1(new_n675), .A2(new_n676), .ZN(new_n683));
  INV_X1    g497(.A(new_n604), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n674), .B1(new_n560), .B2(G472), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n683), .A2(new_n684), .A3(new_n685), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n666), .A2(new_n659), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n686), .A2(new_n650), .A3(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G125), .ZN(G27));
  OR2_X1    g503(.A1(new_n283), .A2(KEYINPUT100), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n283), .A2(KEYINPUT100), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n690), .A2(new_n621), .A3(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n692), .A2(new_n673), .ZN(new_n693));
  INV_X1    g507(.A(new_n693), .ZN(new_n694));
  INV_X1    g508(.A(KEYINPUT42), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n543), .A2(new_n553), .A3(new_n502), .ZN(new_n696));
  NOR4_X1   g510(.A1(new_n425), .A2(new_n651), .A3(new_n695), .A4(new_n696), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n694), .A2(new_n697), .ZN(new_n698));
  NOR2_X1   g512(.A1(new_n425), .A2(new_n696), .ZN(new_n699));
  NAND4_X1  g513(.A1(new_n284), .A2(new_n343), .A3(new_n650), .A4(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n701), .A3(new_n695), .ZN(new_n702));
  INV_X1    g516(.A(new_n702), .ZN(new_n703));
  AOI21_X1  g517(.A(new_n701), .B1(new_n700), .B2(new_n695), .ZN(new_n704));
  OAI21_X1  g518(.A(new_n698), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G131), .ZN(G33));
  INV_X1    g520(.A(new_n616), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n284), .A2(new_n343), .A3(new_n707), .A4(new_n699), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G134), .ZN(G36));
  INV_X1    g523(.A(KEYINPUT105), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n570), .A2(new_n571), .A3(new_n573), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n459), .A2(new_n711), .ZN(new_n712));
  INV_X1    g526(.A(KEYINPUT104), .ZN(new_n713));
  NOR2_X1   g527(.A1(new_n713), .A2(KEYINPUT43), .ZN(new_n714));
  NOR2_X1   g528(.A1(new_n712), .A2(new_n714), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n713), .A2(KEYINPUT43), .ZN(new_n716));
  INV_X1    g530(.A(new_n714), .ZN(new_n717));
  AOI22_X1  g531(.A1(new_n459), .A2(new_n711), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  OAI21_X1  g532(.A(new_n710), .B1(new_n715), .B2(new_n718), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n717), .A2(new_n716), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n712), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n721), .B(KEYINPUT105), .C1(new_n712), .C2(new_n714), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n684), .B1(new_n719), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n670), .A2(new_n271), .ZN(new_n724));
  AND3_X1   g538(.A1(new_n723), .A2(KEYINPUT44), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g539(.A(KEYINPUT44), .B1(new_n723), .B2(new_n724), .ZN(new_n726));
  NOR3_X1   g540(.A1(new_n725), .A2(new_n726), .A3(new_n696), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT103), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT45), .B(new_n411), .C1(new_n416), .C2(new_n418), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT101), .ZN(new_n730));
  NAND2_X1  g544(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  INV_X1    g545(.A(KEYINPUT45), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n419), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g547(.A(new_n383), .B1(new_n395), .B2(new_n400), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n734), .A2(KEYINPUT79), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n735), .A2(new_n346), .A3(new_n417), .ZN(new_n736));
  NAND4_X1  g550(.A1(new_n736), .A2(KEYINPUT101), .A3(KEYINPUT45), .A4(new_n411), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n731), .A2(new_n733), .A3(G469), .A4(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n738), .A2(new_n406), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT46), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n405), .A2(new_n740), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n738), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n743), .A2(KEYINPUT102), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT102), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n738), .A2(new_n745), .A3(new_n742), .ZN(new_n746));
  NAND4_X1  g560(.A1(new_n741), .A2(new_n744), .A3(new_n404), .A4(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(new_n424), .ZN(new_n748));
  INV_X1    g562(.A(new_n634), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n728), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  NAND4_X1  g564(.A1(new_n747), .A2(KEYINPUT103), .A3(new_n424), .A4(new_n634), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n727), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g566(.A(KEYINPUT106), .B(G137), .Z(new_n753));
  XNOR2_X1  g567(.A(new_n752), .B(new_n753), .ZN(G39));
  INV_X1    g568(.A(KEYINPUT47), .ZN(new_n755));
  INV_X1    g569(.A(KEYINPUT107), .ZN(new_n756));
  AND3_X1   g570(.A1(new_n747), .A2(new_n756), .A3(new_n424), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n756), .B1(new_n747), .B2(new_n424), .ZN(new_n758));
  OAI211_X1 g572(.A(KEYINPUT108), .B(new_n755), .C1(new_n757), .C2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n748), .A2(KEYINPUT107), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n755), .A2(KEYINPUT108), .ZN(new_n762));
  NAND3_X1  g576(.A1(new_n747), .A2(new_n756), .A3(new_n424), .ZN(new_n763));
  NAND4_X1  g577(.A1(new_n760), .A2(new_n761), .A3(new_n762), .A4(new_n763), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g579(.A(new_n696), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n342), .A2(new_n650), .A3(new_n766), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n284), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(KEYINPUT109), .B1(new_n765), .B2(new_n768), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  INV_X1    g584(.A(new_n768), .ZN(new_n771));
  AOI211_X1 g585(.A(new_n770), .B(new_n771), .C1(new_n759), .C2(new_n764), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(new_n289), .ZN(G42));
  XOR2_X1   g588(.A(new_n631), .B(KEYINPUT95), .Z(new_n775));
  NAND2_X1  g589(.A1(new_n658), .A2(new_n404), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n776), .A2(KEYINPUT49), .ZN(new_n777));
  NAND2_X1  g591(.A1(new_n776), .A2(KEYINPUT49), .ZN(new_n778));
  NOR3_X1   g592(.A1(new_n712), .A2(new_n423), .A3(new_n503), .ZN(new_n779));
  AND4_X1   g593(.A1(new_n673), .A2(new_n777), .A3(new_n778), .A4(new_n779), .ZN(new_n780));
  NAND3_X1  g594(.A1(new_n775), .A2(new_n643), .A3(new_n780), .ZN(new_n781));
  INV_X1    g595(.A(KEYINPUT51), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n683), .A2(new_n685), .ZN(new_n783));
  OAI21_X1  g597(.A(new_n612), .B1(new_n715), .B2(new_n718), .ZN(new_n784));
  INV_X1    g598(.A(new_n784), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n783), .A2(new_n673), .A3(new_n785), .ZN(new_n786));
  NOR2_X1   g600(.A1(new_n786), .A2(new_n696), .ZN(new_n787));
  INV_X1    g601(.A(new_n787), .ZN(new_n788));
  OR2_X1    g602(.A1(new_n765), .A2(KEYINPUT116), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n776), .A2(new_n424), .ZN(new_n790));
  AOI21_X1  g604(.A(new_n790), .B1(new_n765), .B2(KEYINPUT116), .ZN(new_n791));
  AOI21_X1  g605(.A(new_n788), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n660), .A2(new_n766), .ZN(new_n793));
  NOR3_X1   g607(.A1(new_n793), .A2(new_n342), .A3(new_n461), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n775), .A2(new_n459), .A3(new_n574), .A4(new_n794), .ZN(new_n795));
  NOR2_X1   g609(.A1(new_n784), .A2(new_n793), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n686), .A2(new_n796), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n795), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n643), .A2(new_n503), .A3(new_n660), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n786), .A2(new_n800), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n801), .A2(KEYINPUT50), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT50), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n786), .A2(new_n803), .A3(new_n800), .ZN(new_n804));
  OAI211_X1 g618(.A(new_n798), .B(new_n799), .C1(new_n802), .C2(new_n804), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n802), .A2(new_n804), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n795), .A2(new_n797), .ZN(new_n807));
  OAI21_X1  g621(.A(KEYINPUT117), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n805), .A2(new_n808), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n782), .B1(new_n792), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT118), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT118), .ZN(new_n812));
  OAI211_X1 g626(.A(new_n812), .B(new_n782), .C1(new_n792), .C2(new_n809), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n684), .A2(new_n615), .ZN(new_n815));
  OR3_X1    g629(.A1(new_n815), .A2(KEYINPUT113), .A3(new_n425), .ZN(new_n816));
  OAI21_X1  g630(.A(KEYINPUT113), .B1(new_n815), .B2(new_n425), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n816), .A2(new_n817), .A3(new_n631), .A4(new_n679), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n624), .A2(new_n653), .A3(new_n688), .A4(new_n818), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT114), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(KEYINPUT52), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n661), .A2(new_n664), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n681), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n456), .B1(new_n592), .B2(new_n452), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n826), .A2(new_n498), .A3(new_n579), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n642), .A2(new_n827), .A3(new_n467), .A4(new_n502), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT111), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  INV_X1    g644(.A(KEYINPUT110), .ZN(new_n831));
  OAI21_X1  g645(.A(new_n831), .B1(new_n574), .B2(new_n459), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n826), .A2(new_n579), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n833), .A2(new_n711), .A3(KEYINPUT110), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n832), .A2(new_n554), .A3(new_n467), .A4(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n554), .A2(KEYINPUT111), .A3(new_n467), .A4(new_n827), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n830), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n558), .A3(new_n561), .ZN(new_n838));
  AND4_X1   g652(.A1(new_n555), .A2(new_n838), .A3(new_n605), .A4(new_n668), .ZN(new_n839));
  NAND3_X1  g653(.A1(new_n686), .A2(new_n650), .A3(new_n699), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n580), .A2(new_n583), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n586), .A2(new_n593), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n498), .A2(new_n614), .ZN(new_n844));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n843), .A3(new_n581), .A4(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n841), .B1(new_n845), .B2(new_n696), .ZN(new_n846));
  NAND4_X1  g660(.A1(new_n766), .A2(KEYINPUT112), .A3(new_n595), .A4(new_n844), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n425), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g662(.A1(new_n848), .A2(new_n284), .A3(new_n604), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n849), .A2(new_n708), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n825), .A2(new_n839), .A3(new_n840), .A4(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n700), .A2(new_n695), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n852), .A2(KEYINPUT99), .ZN(new_n853));
  AOI22_X1  g667(.A1(new_n853), .A2(new_n702), .B1(new_n694), .B2(new_n697), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n851), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g669(.A1(new_n819), .A2(new_n820), .A3(KEYINPUT52), .ZN(new_n856));
  NAND4_X1  g670(.A1(new_n823), .A2(new_n855), .A3(KEYINPUT53), .A4(new_n856), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT54), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n555), .A2(new_n838), .A3(new_n605), .A4(new_n668), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n859), .A2(new_n824), .A3(new_n681), .ZN(new_n860));
  AND3_X1   g674(.A1(new_n840), .A2(new_n708), .A3(new_n849), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n705), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n819), .A2(new_n822), .ZN(new_n863));
  AOI22_X1  g677(.A1(new_n620), .A2(new_n623), .B1(new_n622), .B2(new_n652), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(KEYINPUT52), .A3(new_n688), .A4(new_n818), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n862), .B1(new_n863), .B2(new_n865), .ZN(new_n866));
  OAI211_X1 g680(.A(new_n857), .B(new_n858), .C1(new_n866), .C2(KEYINPUT53), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n867), .A2(KEYINPUT115), .ZN(new_n868));
  AOI21_X1  g682(.A(KEYINPUT52), .B1(new_n819), .B2(new_n820), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n862), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT53), .B1(new_n870), .B2(new_n856), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n863), .A2(new_n865), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n872), .A2(new_n855), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(KEYINPUT54), .B1(new_n871), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n873), .A2(new_n874), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT115), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n877), .A2(new_n878), .A3(new_n858), .A4(new_n857), .ZN(new_n879));
  AND3_X1   g693(.A1(new_n868), .A2(new_n876), .A3(new_n879), .ZN(new_n880));
  NOR3_X1   g694(.A1(new_n693), .A2(new_n784), .A3(new_n793), .ZN(new_n881));
  OR2_X1    g695(.A1(new_n881), .A2(KEYINPUT48), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n251), .A2(G952), .ZN(new_n883));
  INV_X1    g697(.A(new_n786), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n883), .B1(new_n884), .B2(new_n687), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n881), .A2(KEYINPUT48), .ZN(new_n886));
  NAND4_X1  g700(.A1(new_n775), .A2(new_n833), .A3(new_n711), .A4(new_n794), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n882), .A2(new_n885), .A3(new_n886), .A4(new_n887), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n806), .A2(new_n782), .A3(new_n807), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n787), .B1(new_n765), .B2(new_n790), .ZN(new_n890));
  AOI21_X1  g704(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n814), .A2(new_n880), .A3(new_n891), .ZN(new_n892));
  NOR2_X1   g706(.A1(G952), .A2(G953), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n781), .B1(new_n892), .B2(new_n893), .ZN(G75));
  AOI21_X1  g708(.A(new_n321), .B1(new_n877), .B2(new_n857), .ZN(new_n895));
  AOI21_X1  g709(.A(KEYINPUT56), .B1(new_n895), .B2(G210), .ZN(new_n896));
  INV_X1    g710(.A(KEYINPUT120), .ZN(new_n897));
  XNOR2_X1  g711(.A(new_n544), .B(KEYINPUT119), .ZN(new_n898));
  XOR2_X1   g712(.A(new_n510), .B(KEYINPUT55), .Z(new_n899));
  XNOR2_X1  g713(.A(new_n898), .B(new_n899), .ZN(new_n900));
  OR3_X1    g714(.A1(new_n896), .A2(new_n897), .A3(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n897), .B1(new_n896), .B2(new_n900), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n251), .A2(G952), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n903), .B1(new_n896), .B2(new_n900), .ZN(new_n904));
  AND3_X1   g718(.A1(new_n901), .A2(new_n902), .A3(new_n904), .ZN(G51));
  NAND2_X1  g719(.A1(new_n877), .A2(new_n857), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(KEYINPUT54), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n867), .ZN(new_n908));
  XNOR2_X1  g722(.A(new_n405), .B(KEYINPUT57), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  XNOR2_X1  g724(.A(new_n402), .B(KEYINPUT121), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n895), .ZN(new_n913));
  OR2_X1    g727(.A1(new_n913), .A2(new_n738), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n903), .B1(new_n912), .B2(new_n914), .ZN(G54));
  NAND3_X1  g729(.A1(new_n895), .A2(KEYINPUT58), .A3(G475), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n590), .A2(new_n591), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n916), .A2(new_n918), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n916), .A2(new_n918), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n919), .A2(new_n920), .A3(new_n903), .ZN(G60));
  NAND2_X1  g735(.A1(new_n564), .A2(new_n567), .ZN(new_n922));
  NAND2_X1  g736(.A1(G478), .A2(G902), .ZN(new_n923));
  XOR2_X1   g737(.A(new_n923), .B(KEYINPUT59), .Z(new_n924));
  NOR2_X1   g738(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n908), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n903), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g742(.A1(new_n880), .A2(new_n924), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n928), .B1(new_n929), .B2(new_n922), .ZN(G63));
  NAND2_X1  g744(.A1(G217), .A2(G902), .ZN(new_n931));
  XOR2_X1   g745(.A(new_n931), .B(KEYINPUT60), .Z(new_n932));
  NAND3_X1  g746(.A1(new_n906), .A2(new_n602), .A3(new_n932), .ZN(new_n933));
  AND2_X1   g747(.A1(new_n906), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n333), .A2(new_n334), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n927), .B(new_n933), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT61), .ZN(new_n937));
  XNOR2_X1  g751(.A(new_n936), .B(new_n937), .ZN(G66));
  INV_X1    g752(.A(G224), .ZN(new_n939));
  OAI21_X1  g753(.A(G953), .B1(new_n465), .B2(new_n939), .ZN(new_n940));
  OAI21_X1  g754(.A(new_n940), .B1(new_n860), .B2(G953), .ZN(new_n941));
  OAI21_X1  g755(.A(new_n898), .B1(G898), .B2(new_n251), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT122), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n941), .B(new_n943), .ZN(G69));
  AOI21_X1  g758(.A(new_n251), .B1(G227), .B2(G900), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n945), .A2(KEYINPUT125), .ZN(new_n946));
  NOR2_X1   g760(.A1(new_n251), .A2(G900), .ZN(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n693), .A2(new_n678), .A3(new_n646), .ZN(new_n949));
  OAI211_X1 g763(.A(new_n750), .B(new_n751), .C1(new_n727), .C2(new_n949), .ZN(new_n950));
  AND3_X1   g764(.A1(new_n864), .A2(new_n688), .A3(new_n708), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n950), .A2(new_n951), .A3(new_n705), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n765), .A2(new_n768), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n770), .ZN(new_n954));
  NAND3_X1  g768(.A1(new_n765), .A2(KEYINPUT109), .A3(new_n768), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n948), .B1(new_n956), .B2(G953), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n957), .A2(KEYINPUT124), .ZN(new_n958));
  INV_X1    g772(.A(new_n952), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(new_n769), .B2(new_n772), .ZN(new_n960));
  AOI21_X1  g774(.A(new_n947), .B1(new_n960), .B2(new_n251), .ZN(new_n961));
  INV_X1    g775(.A(KEYINPUT124), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XNOR2_X1  g777(.A(new_n247), .B(new_n448), .ZN(new_n964));
  INV_X1    g778(.A(new_n964), .ZN(new_n965));
  NAND3_X1  g779(.A1(new_n958), .A2(new_n963), .A3(new_n965), .ZN(new_n966));
  INV_X1    g780(.A(KEYINPUT123), .ZN(new_n967));
  NOR2_X1   g781(.A1(new_n636), .A2(new_n637), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n827), .B1(new_n832), .B2(new_n834), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n969), .A2(new_n696), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n968), .A2(new_n284), .A3(new_n343), .A4(new_n970), .ZN(new_n971));
  AND3_X1   g785(.A1(new_n752), .A2(new_n967), .A3(new_n971), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n967), .B1(new_n752), .B2(new_n971), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n648), .A2(new_n864), .A3(new_n688), .ZN(new_n974));
  INV_X1    g788(.A(KEYINPUT62), .ZN(new_n975));
  AND2_X1   g789(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n974), .A2(new_n975), .ZN(new_n977));
  OAI22_X1  g791(.A1(new_n972), .A2(new_n973), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n251), .B1(new_n773), .B2(new_n978), .ZN(new_n979));
  AOI22_X1  g793(.A1(new_n979), .A2(new_n964), .B1(KEYINPUT125), .B2(new_n945), .ZN(new_n980));
  AOI21_X1  g794(.A(new_n946), .B1(new_n966), .B2(new_n980), .ZN(new_n981));
  OAI21_X1  g795(.A(new_n965), .B1(new_n961), .B2(new_n962), .ZN(new_n982));
  AOI211_X1 g796(.A(KEYINPUT124), .B(new_n947), .C1(new_n960), .C2(new_n251), .ZN(new_n983));
  OAI211_X1 g797(.A(new_n980), .B(new_n946), .C1(new_n982), .C2(new_n983), .ZN(new_n984));
  INV_X1    g798(.A(new_n984), .ZN(new_n985));
  NOR2_X1   g799(.A1(new_n981), .A2(new_n985), .ZN(G72));
  NAND2_X1  g800(.A1(G472), .A2(G902), .ZN(new_n987));
  XOR2_X1   g801(.A(new_n987), .B(KEYINPUT63), .Z(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  INV_X1    g803(.A(new_n258), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n989), .B1(new_n279), .B2(new_n990), .ZN(new_n991));
  XOR2_X1   g805(.A(new_n991), .B(KEYINPUT127), .Z(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n871), .B2(new_n875), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n993), .A2(new_n927), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n956), .A2(new_n860), .ZN(new_n995));
  XNOR2_X1  g809(.A(new_n988), .B(KEYINPUT126), .ZN(new_n996));
  AOI211_X1 g810(.A(new_n278), .B(new_n256), .C1(new_n995), .C2(new_n996), .ZN(new_n997));
  NOR2_X1   g811(.A1(new_n773), .A2(new_n978), .ZN(new_n998));
  NAND2_X1  g812(.A1(new_n998), .A2(new_n860), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n996), .ZN(new_n1000));
  AOI211_X1 g814(.A(new_n994), .B(new_n997), .C1(new_n626), .C2(new_n1000), .ZN(G57));
endmodule


