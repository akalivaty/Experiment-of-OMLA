//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 0 1 0 0 1 1 0 0 1 0 1 1 0 0 1 1 0 0 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:41 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n780, new_n781, new_n782, new_n783, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n794,
    new_n795, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n823, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1031,
    new_n1032, new_n1033, new_n1034, new_n1035, new_n1036, new_n1037,
    new_n1038, new_n1039, new_n1040, new_n1041;
  OAI21_X1  g000(.A(G214), .B1(G237), .B2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G953), .ZN(new_n188));
  AND2_X1   g002(.A1(new_n188), .A2(G952), .ZN(new_n189));
  NAND2_X1  g003(.A1(G234), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n189), .A2(new_n190), .ZN(new_n191));
  XNOR2_X1  g005(.A(KEYINPUT21), .B(G898), .ZN(new_n192));
  INV_X1    g006(.A(new_n192), .ZN(new_n193));
  NAND3_X1  g007(.A1(new_n190), .A2(G902), .A3(G953), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n191), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT84), .ZN(new_n196));
  INV_X1    g010(.A(G107), .ZN(new_n197));
  OAI21_X1  g011(.A(KEYINPUT82), .B1(new_n197), .B2(G104), .ZN(new_n198));
  INV_X1    g012(.A(G104), .ZN(new_n199));
  OAI21_X1  g013(.A(KEYINPUT81), .B1(new_n199), .B2(G107), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT82), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n201), .A2(new_n199), .A3(G107), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT81), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n203), .A2(new_n197), .A3(G104), .ZN(new_n204));
  NAND4_X1  g018(.A1(new_n198), .A2(new_n200), .A3(new_n202), .A4(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT83), .ZN(new_n206));
  NAND3_X1  g020(.A1(new_n205), .A2(new_n206), .A3(G101), .ZN(new_n207));
  NOR2_X1   g021(.A1(new_n199), .A2(G107), .ZN(new_n208));
  NAND2_X1  g022(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n209));
  INV_X1    g023(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g024(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n208), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  INV_X1    g026(.A(new_n211), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n197), .A2(G104), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G101), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n199), .A2(G107), .ZN(new_n217));
  NAND4_X1  g031(.A1(new_n212), .A2(new_n215), .A3(new_n216), .A4(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  AOI21_X1  g033(.A(new_n206), .B1(new_n205), .B2(G101), .ZN(new_n220));
  OAI21_X1  g034(.A(new_n196), .B1(new_n219), .B2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n205), .A2(G101), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(KEYINPUT83), .ZN(new_n223));
  NAND4_X1  g037(.A1(new_n223), .A2(KEYINPUT84), .A3(new_n218), .A4(new_n207), .ZN(new_n224));
  XNOR2_X1  g038(.A(G116), .B(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT5), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  NOR3_X1   g041(.A1(new_n227), .A2(KEYINPUT5), .A3(G119), .ZN(new_n228));
  INV_X1    g042(.A(G113), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  XOR2_X1   g044(.A(KEYINPUT2), .B(G113), .Z(new_n231));
  AOI22_X1  g045(.A1(new_n226), .A2(new_n230), .B1(new_n231), .B2(new_n225), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n221), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n234));
  NOR2_X1   g048(.A1(new_n225), .A2(new_n234), .ZN(new_n235));
  XNOR2_X1  g049(.A(new_n235), .B(new_n231), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT4), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n214), .B1(new_n213), .B2(new_n209), .ZN(new_n239));
  OAI21_X1  g053(.A(new_n217), .B1(new_n208), .B2(new_n211), .ZN(new_n240));
  OAI211_X1 g054(.A(new_n238), .B(G101), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  OAI21_X1  g055(.A(G101), .B1(new_n239), .B2(new_n240), .ZN(new_n242));
  NAND3_X1  g056(.A1(new_n242), .A2(KEYINPUT4), .A3(new_n218), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n237), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n233), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g059(.A(G110), .B(G122), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n233), .A2(new_n244), .A3(new_n246), .ZN(new_n249));
  NAND3_X1  g063(.A1(new_n248), .A2(KEYINPUT6), .A3(new_n249), .ZN(new_n250));
  AND2_X1   g064(.A1(KEYINPUT0), .A2(G128), .ZN(new_n251));
  NOR2_X1   g065(.A1(KEYINPUT0), .A2(G128), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  OR2_X1    g067(.A1(KEYINPUT64), .A2(G143), .ZN(new_n254));
  NAND2_X1  g068(.A1(KEYINPUT64), .A2(G143), .ZN(new_n255));
  AOI21_X1  g069(.A(G146), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(G146), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G143), .ZN(new_n258));
  OAI211_X1 g072(.A(KEYINPUT65), .B(new_n253), .C1(new_n256), .C2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n254), .A2(G146), .A3(new_n255), .ZN(new_n260));
  INV_X1    g074(.A(G143), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G146), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n260), .A2(new_n251), .A3(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n259), .A2(new_n264), .ZN(new_n265));
  XNOR2_X1  g079(.A(KEYINPUT0), .B(G128), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT64), .A2(G143), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT64), .A2(G143), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n257), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n258), .ZN(new_n270));
  AOI21_X1  g084(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n271), .A2(KEYINPUT65), .ZN(new_n272));
  OAI21_X1  g086(.A(G125), .B1(new_n265), .B2(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT85), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  OAI21_X1  g089(.A(KEYINPUT1), .B1(new_n261), .B2(G146), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(G128), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n277), .B1(new_n256), .B2(new_n258), .ZN(new_n278));
  INV_X1    g092(.A(G125), .ZN(new_n279));
  INV_X1    g093(.A(G128), .ZN(new_n280));
  NOR2_X1   g094(.A1(new_n280), .A2(KEYINPUT1), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n260), .A2(new_n263), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n279), .A3(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(KEYINPUT86), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT86), .ZN(new_n285));
  NAND4_X1  g099(.A1(new_n278), .A2(new_n285), .A3(new_n279), .A4(new_n282), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  OAI211_X1 g101(.A(KEYINPUT85), .B(G125), .C1(new_n265), .C2(new_n272), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n275), .A2(new_n287), .A3(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n188), .A2(G224), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n290), .B(KEYINPUT87), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n289), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n291), .ZN(new_n293));
  NAND4_X1  g107(.A1(new_n275), .A2(new_n293), .A3(new_n287), .A4(new_n288), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  INV_X1    g109(.A(KEYINPUT6), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n245), .A2(new_n296), .A3(new_n247), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n250), .A2(new_n295), .A3(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n287), .A2(new_n273), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n293), .A2(KEYINPUT7), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n299), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(new_n300), .ZN(new_n302));
  NAND4_X1  g116(.A1(new_n275), .A2(new_n287), .A3(new_n288), .A4(new_n302), .ZN(new_n303));
  OR3_X1    g117(.A1(new_n219), .A2(new_n220), .A3(new_n232), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n232), .B1(new_n219), .B2(new_n220), .ZN(new_n305));
  XNOR2_X1  g119(.A(new_n246), .B(KEYINPUT8), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n304), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n249), .A2(new_n301), .A3(new_n303), .A4(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(G902), .ZN(new_n309));
  AND2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  OAI21_X1  g124(.A(G210), .B1(G237), .B2(G902), .ZN(new_n311));
  AND3_X1   g125(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n312));
  AOI21_X1  g126(.A(new_n311), .B1(new_n298), .B2(new_n310), .ZN(new_n313));
  OAI211_X1 g127(.A(new_n187), .B(new_n195), .C1(new_n312), .C2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(new_n314), .ZN(new_n315));
  XNOR2_X1  g129(.A(KEYINPUT9), .B(G234), .ZN(new_n316));
  OAI21_X1  g130(.A(G221), .B1(new_n316), .B2(G902), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  XNOR2_X1  g132(.A(G110), .B(G140), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n188), .A2(G227), .ZN(new_n320));
  XNOR2_X1  g134(.A(new_n319), .B(new_n320), .ZN(new_n321));
  AND3_X1   g135(.A1(new_n260), .A2(new_n263), .A3(new_n281), .ZN(new_n322));
  AOI22_X1  g136(.A1(new_n269), .A2(new_n270), .B1(G128), .B2(new_n276), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g138(.A(new_n324), .B1(new_n219), .B2(new_n220), .ZN(new_n325));
  AOI21_X1  g139(.A(new_n280), .B1(new_n269), .B2(KEYINPUT1), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n267), .A2(new_n268), .ZN(new_n327));
  AOI21_X1  g141(.A(new_n262), .B1(new_n327), .B2(G146), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n282), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n329), .A2(new_n223), .A3(new_n218), .A4(new_n207), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(G134), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n332), .A2(G137), .ZN(new_n333));
  NOR2_X1   g147(.A1(new_n332), .A2(G137), .ZN(new_n334));
  INV_X1    g148(.A(KEYINPUT11), .ZN(new_n335));
  NOR2_X1   g149(.A1(new_n335), .A2(KEYINPUT66), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n333), .B1(new_n334), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(G137), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G134), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT66), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n335), .A2(KEYINPUT66), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g157(.A(G131), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  NOR2_X1   g158(.A1(new_n338), .A2(G134), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n345), .B1(new_n339), .B2(new_n341), .ZN(new_n346));
  NOR2_X1   g160(.A1(new_n340), .A2(KEYINPUT11), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n334), .B1(new_n336), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G131), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n344), .A2(new_n350), .ZN(new_n351));
  AOI21_X1  g165(.A(KEYINPUT12), .B1(new_n331), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT12), .ZN(new_n353));
  INV_X1    g167(.A(new_n351), .ZN(new_n354));
  AOI211_X1 g168(.A(new_n353), .B(new_n354), .C1(new_n325), .C2(new_n330), .ZN(new_n355));
  NOR2_X1   g169(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g170(.A1(new_n243), .A2(new_n241), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n265), .A2(new_n272), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n359));
  AOI22_X1  g173(.A1(new_n357), .A2(new_n358), .B1(new_n330), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT70), .ZN(new_n361));
  NOR3_X1   g175(.A1(new_n322), .A2(new_n323), .A3(new_n361), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT70), .B1(new_n278), .B2(new_n282), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n364), .A2(new_n221), .A3(KEYINPUT10), .A4(new_n224), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n360), .A2(new_n354), .A3(new_n365), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n321), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n221), .A2(new_n224), .ZN(new_n368));
  OAI21_X1  g182(.A(new_n361), .B1(new_n322), .B2(new_n323), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n278), .A2(KEYINPUT70), .A3(new_n282), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(KEYINPUT10), .A3(new_n370), .ZN(new_n371));
  NOR2_X1   g185(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n330), .A2(new_n359), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n358), .A2(new_n241), .A3(new_n243), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  OAI21_X1  g189(.A(new_n351), .B1(new_n372), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n360), .A2(new_n365), .A3(new_n354), .ZN(new_n377));
  INV_X1    g191(.A(new_n321), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n376), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  NAND3_X1  g193(.A1(new_n367), .A2(G469), .A3(new_n379), .ZN(new_n380));
  NAND2_X1  g194(.A1(G469), .A2(G902), .ZN(new_n381));
  AND2_X1   g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G469), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n377), .A2(new_n378), .ZN(new_n384));
  NOR2_X1   g198(.A1(new_n384), .A2(new_n356), .ZN(new_n385));
  AOI21_X1  g199(.A(new_n378), .B1(new_n376), .B2(new_n377), .ZN(new_n386));
  OAI211_X1 g200(.A(new_n383), .B(new_n309), .C1(new_n385), .C2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n318), .B1(new_n382), .B2(new_n387), .ZN(new_n388));
  INV_X1    g202(.A(G475), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT88), .ZN(new_n390));
  NOR2_X1   g204(.A1(new_n279), .A2(G140), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NOR2_X1   g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n391), .B2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n392), .A2(G125), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n279), .A2(G140), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT88), .ZN(new_n397));
  AND3_X1   g211(.A1(new_n394), .A2(G146), .A3(new_n397), .ZN(new_n398));
  NOR3_X1   g212(.A1(new_n391), .A2(new_n393), .A3(G146), .ZN(new_n399));
  INV_X1    g213(.A(G237), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(new_n188), .A3(G214), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(new_n254), .A3(new_n255), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n400), .A2(new_n188), .A3(G143), .A4(G214), .ZN(new_n403));
  AND2_X1   g217(.A1(KEYINPUT18), .A2(G131), .ZN(new_n404));
  AND3_X1   g218(.A1(new_n402), .A2(new_n403), .A3(new_n404), .ZN(new_n405));
  AOI21_X1  g219(.A(new_n404), .B1(new_n402), .B2(new_n403), .ZN(new_n406));
  OAI22_X1  g220(.A1(new_n398), .A2(new_n399), .B1(new_n405), .B2(new_n406), .ZN(new_n407));
  XNOR2_X1  g221(.A(KEYINPUT64), .B(G143), .ZN(new_n408));
  INV_X1    g222(.A(G214), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n409), .A2(G237), .A3(G953), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n403), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n411), .A2(G131), .ZN(new_n412));
  INV_X1    g226(.A(KEYINPUT17), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n402), .A2(new_n349), .A3(new_n403), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n412), .A2(new_n413), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n411), .A2(KEYINPUT17), .A3(G131), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n395), .A2(new_n396), .A3(KEYINPUT16), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT16), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n391), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(new_n257), .ZN(new_n421));
  NAND3_X1  g235(.A1(new_n417), .A2(new_n419), .A3(G146), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n416), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n407), .B1(new_n415), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g238(.A(G113), .B(G122), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(new_n199), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n427), .ZN(new_n428));
  OAI211_X1 g242(.A(new_n407), .B(new_n426), .C1(new_n415), .C2(new_n423), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  AOI21_X1  g244(.A(new_n389), .B1(new_n430), .B2(new_n309), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT89), .ZN(new_n432));
  INV_X1    g246(.A(new_n429), .ZN(new_n433));
  INV_X1    g247(.A(new_n422), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n434), .B1(new_n412), .B2(new_n414), .ZN(new_n435));
  INV_X1    g249(.A(KEYINPUT19), .ZN(new_n436));
  AOI21_X1  g250(.A(new_n436), .B1(new_n394), .B2(new_n397), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT19), .B1(new_n395), .B2(new_n396), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n257), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n435), .A2(new_n439), .ZN(new_n440));
  AOI21_X1  g254(.A(new_n426), .B1(new_n440), .B2(new_n407), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n432), .B1(new_n433), .B2(new_n441), .ZN(new_n442));
  NOR2_X1   g256(.A1(G475), .A2(G902), .ZN(new_n443));
  OR2_X1    g257(.A1(new_n398), .A2(new_n399), .ZN(new_n444));
  OR2_X1    g258(.A1(new_n405), .A2(new_n406), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n444), .A2(new_n445), .B1(new_n435), .B2(new_n439), .ZN(new_n446));
  OAI211_X1 g260(.A(KEYINPUT89), .B(new_n429), .C1(new_n446), .C2(new_n426), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n442), .A2(new_n443), .A3(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(KEYINPUT20), .ZN(new_n449));
  NOR3_X1   g263(.A1(KEYINPUT20), .A2(G475), .A3(G902), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n450), .B1(new_n433), .B2(new_n441), .ZN(new_n451));
  AOI21_X1  g265(.A(new_n431), .B1(new_n449), .B2(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(G478), .ZN(new_n453));
  OR2_X1    g267(.A1(new_n453), .A2(KEYINPUT15), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(KEYINPUT93), .ZN(new_n455));
  INV_X1    g269(.A(new_n455), .ZN(new_n456));
  NOR2_X1   g270(.A1(new_n454), .A2(KEYINPUT93), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  NOR3_X1   g273(.A1(new_n316), .A2(new_n459), .A3(G953), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT13), .ZN(new_n461));
  NAND4_X1  g275(.A1(new_n254), .A2(new_n461), .A3(G128), .A4(new_n255), .ZN(new_n462));
  AND2_X1   g276(.A1(new_n462), .A2(G134), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT90), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n254), .A2(G128), .A3(new_n255), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n261), .A2(G128), .ZN(new_n466));
  INV_X1    g280(.A(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(KEYINPUT13), .A3(new_n467), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n463), .A2(new_n464), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(new_n466), .B1(new_n327), .B2(G128), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n227), .A2(G122), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  NAND2_X1  g288(.A1(new_n474), .A2(G107), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n472), .A2(new_n473), .A3(new_n197), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n470), .A2(new_n332), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n464), .B1(new_n463), .B2(new_n468), .ZN(new_n479));
  OAI21_X1  g293(.A(KEYINPUT91), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n463), .A2(new_n468), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(KEYINPUT90), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT91), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n482), .A2(new_n483), .A3(new_n469), .A4(new_n477), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n480), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n473), .A2(KEYINPUT14), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n486), .A2(new_n472), .ZN(new_n487));
  OR2_X1    g301(.A1(new_n473), .A2(KEYINPUT14), .ZN(new_n488));
  AOI21_X1  g302(.A(new_n487), .B1(KEYINPUT92), .B2(new_n488), .ZN(new_n489));
  OR2_X1    g303(.A1(new_n488), .A2(KEYINPUT92), .ZN(new_n490));
  AOI21_X1  g304(.A(new_n197), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  AND3_X1   g305(.A1(new_n465), .A2(new_n332), .A3(new_n467), .ZN(new_n492));
  AOI21_X1  g306(.A(new_n332), .B1(new_n465), .B2(new_n467), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n476), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n491), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(new_n495), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n460), .B1(new_n485), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n460), .ZN(new_n498));
  AOI211_X1 g312(.A(new_n498), .B(new_n495), .C1(new_n480), .C2(new_n484), .ZN(new_n499));
  OAI211_X1 g313(.A(new_n309), .B(new_n458), .C1(new_n497), .C2(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n485), .A2(new_n496), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n498), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n485), .A2(new_n496), .A3(new_n460), .ZN(new_n503));
  AOI21_X1  g317(.A(G902), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OAI21_X1  g318(.A(new_n500), .B1(new_n504), .B2(new_n455), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n452), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n315), .A2(KEYINPUT94), .A3(new_n388), .A4(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT94), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n387), .A2(new_n381), .A3(new_n380), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n506), .A2(new_n509), .A3(new_n317), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n508), .B1(new_n510), .B2(new_n314), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n188), .A2(G221), .A3(G234), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT77), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT22), .B(G137), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n513), .B(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g330(.A1(new_n280), .A2(G119), .ZN(new_n517));
  INV_X1    g331(.A(G119), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  XNOR2_X1  g334(.A(KEYINPUT24), .B(G110), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  AOI21_X1  g336(.A(new_n522), .B1(new_n421), .B2(new_n422), .ZN(new_n523));
  INV_X1    g337(.A(new_n523), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT74), .B1(new_n518), .B2(G128), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT23), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT23), .ZN(new_n527));
  NAND3_X1  g341(.A1(new_n517), .A2(KEYINPUT74), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(new_n528), .A3(new_n519), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(KEYINPUT75), .ZN(new_n530));
  INV_X1    g344(.A(KEYINPUT75), .ZN(new_n531));
  NAND4_X1  g345(.A1(new_n526), .A2(new_n528), .A3(new_n531), .A4(new_n519), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n530), .A2(G110), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT76), .ZN(new_n534));
  INV_X1    g348(.A(G110), .ZN(new_n535));
  AOI21_X1  g349(.A(new_n535), .B1(new_n529), .B2(KEYINPUT75), .ZN(new_n536));
  INV_X1    g350(.A(KEYINPUT76), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n536), .A2(new_n537), .A3(new_n532), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n524), .B1(new_n534), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n434), .A2(new_n399), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n520), .A2(new_n521), .ZN(new_n541));
  OAI21_X1  g355(.A(new_n541), .B1(new_n529), .B2(G110), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n540), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  OAI21_X1  g358(.A(new_n516), .B1(new_n539), .B2(new_n544), .ZN(new_n545));
  AND3_X1   g359(.A1(new_n536), .A2(new_n537), .A3(new_n532), .ZN(new_n546));
  AOI21_X1  g360(.A(new_n537), .B1(new_n536), .B2(new_n532), .ZN(new_n547));
  OAI21_X1  g361(.A(new_n523), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n548), .A2(new_n543), .A3(new_n515), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n545), .A2(new_n549), .A3(new_n309), .ZN(new_n550));
  INV_X1    g364(.A(KEYINPUT78), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(KEYINPUT25), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n552), .A2(KEYINPUT79), .A3(new_n553), .ZN(new_n554));
  INV_X1    g368(.A(G234), .ZN(new_n555));
  OAI21_X1  g369(.A(G217), .B1(new_n555), .B2(G902), .ZN(new_n556));
  XNOR2_X1  g370(.A(new_n556), .B(KEYINPUT73), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  INV_X1    g372(.A(KEYINPUT79), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n550), .A2(new_n559), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(KEYINPUT25), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n559), .B1(new_n550), .B2(new_n551), .ZN(new_n562));
  OAI211_X1 g376(.A(new_n554), .B(new_n558), .C1(new_n561), .C2(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n545), .A2(new_n549), .ZN(new_n564));
  INV_X1    g378(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g379(.A1(new_n558), .A2(G902), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n563), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n337), .A2(new_n343), .ZN(new_n569));
  OAI211_X1 g383(.A(KEYINPUT67), .B(G131), .C1(new_n334), .C2(new_n345), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT67), .ZN(new_n571));
  XNOR2_X1  g385(.A(G134), .B(G137), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n571), .B1(new_n572), .B2(new_n349), .ZN(new_n573));
  AOI22_X1  g387(.A1(new_n569), .A2(new_n349), .B1(new_n570), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n574), .A2(new_n369), .A3(new_n370), .ZN(new_n575));
  AOI22_X1  g389(.A1(new_n271), .A2(KEYINPUT65), .B1(new_n328), .B2(new_n251), .ZN(new_n576));
  OAI21_X1  g390(.A(new_n253), .B1(new_n256), .B2(new_n258), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT65), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  NAND3_X1  g393(.A1(new_n576), .A2(new_n351), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n575), .A2(new_n236), .A3(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT28), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NAND3_X1  g397(.A1(new_n400), .A2(new_n188), .A3(G210), .ZN(new_n584));
  XNOR2_X1  g398(.A(new_n584), .B(KEYINPUT27), .ZN(new_n585));
  XNOR2_X1  g399(.A(KEYINPUT26), .B(G101), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n585), .B(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n583), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NOR2_X1   g403(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT72), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n575), .A2(new_n580), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n237), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(new_n581), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n591), .B1(new_n594), .B2(KEYINPUT28), .ZN(new_n595));
  AND3_X1   g409(.A1(new_n575), .A2(new_n236), .A3(new_n580), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n236), .B1(new_n575), .B2(new_n580), .ZN(new_n597));
  OAI211_X1 g411(.A(new_n591), .B(KEYINPUT28), .C1(new_n596), .C2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n590), .B1(new_n595), .B2(new_n599), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n575), .A2(KEYINPUT30), .A3(new_n580), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT71), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT71), .ZN(new_n603));
  NAND4_X1  g417(.A1(new_n575), .A2(new_n580), .A3(new_n603), .A4(KEYINPUT30), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n573), .A2(new_n570), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n350), .ZN(new_n607));
  OAI21_X1  g421(.A(KEYINPUT68), .B1(new_n607), .B2(new_n324), .ZN(new_n608));
  INV_X1    g422(.A(KEYINPUT68), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n278), .A2(new_n282), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n574), .A2(new_n609), .A3(new_n610), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n608), .A2(new_n611), .A3(new_n580), .ZN(new_n612));
  INV_X1    g426(.A(KEYINPUT30), .ZN(new_n613));
  AOI21_X1  g427(.A(new_n236), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  AOI21_X1  g428(.A(new_n596), .B1(new_n605), .B2(new_n614), .ZN(new_n615));
  NOR2_X1   g429(.A1(new_n615), .A2(new_n587), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n612), .A2(new_n237), .ZN(new_n617));
  AOI21_X1  g431(.A(new_n582), .B1(new_n617), .B2(new_n581), .ZN(new_n618));
  OAI21_X1  g432(.A(new_n589), .B1(new_n618), .B2(new_n588), .ZN(new_n619));
  OAI211_X1 g433(.A(new_n600), .B(new_n309), .C1(new_n616), .C2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n605), .A2(new_n614), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n581), .A2(new_n587), .ZN(new_n622));
  INV_X1    g436(.A(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT31), .ZN(new_n625));
  INV_X1    g439(.A(new_n587), .ZN(new_n626));
  INV_X1    g440(.A(new_n583), .ZN(new_n627));
  OAI21_X1  g441(.A(new_n626), .B1(new_n618), .B2(new_n627), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT31), .ZN(new_n629));
  NAND3_X1  g443(.A1(new_n621), .A2(new_n629), .A3(new_n623), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n625), .A2(new_n628), .A3(new_n630), .ZN(new_n631));
  NOR2_X1   g445(.A1(G472), .A2(G902), .ZN(new_n632));
  INV_X1    g446(.A(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(KEYINPUT32), .ZN(new_n634));
  NOR2_X1   g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g449(.A1(G472), .A2(new_n620), .B1(new_n631), .B2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(new_n628), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n629), .B1(new_n621), .B2(new_n623), .ZN(new_n638));
  AOI211_X1 g452(.A(KEYINPUT31), .B(new_n622), .C1(new_n605), .C2(new_n614), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n637), .A2(new_n638), .A3(new_n639), .ZN(new_n640));
  OAI21_X1  g454(.A(new_n634), .B1(new_n640), .B2(new_n633), .ZN(new_n641));
  AOI21_X1  g455(.A(new_n568), .B1(new_n636), .B2(new_n641), .ZN(new_n642));
  NAND3_X1  g456(.A1(new_n507), .A2(new_n511), .A3(new_n642), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n643), .B(G101), .ZN(G3));
  NOR2_X1   g458(.A1(new_n638), .A2(new_n639), .ZN(new_n645));
  AOI21_X1  g459(.A(G902), .B1(new_n645), .B2(new_n628), .ZN(new_n646));
  INV_X1    g460(.A(G472), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(KEYINPUT95), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n646), .B(new_n648), .ZN(new_n649));
  NOR2_X1   g463(.A1(new_n453), .A2(G902), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  INV_X1    g465(.A(KEYINPUT33), .ZN(new_n652));
  NAND4_X1  g466(.A1(new_n502), .A2(KEYINPUT96), .A3(new_n652), .A4(new_n503), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n652), .A2(KEYINPUT96), .ZN(new_n654));
  OR2_X1    g468(.A1(new_n652), .A2(KEYINPUT96), .ZN(new_n655));
  OAI211_X1 g469(.A(new_n654), .B(new_n655), .C1(new_n497), .C2(new_n499), .ZN(new_n656));
  AOI21_X1  g470(.A(new_n651), .B1(new_n653), .B2(new_n656), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n504), .A2(G478), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR3_X1   g473(.A1(new_n314), .A2(new_n452), .A3(new_n659), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n380), .A2(new_n381), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n354), .B1(new_n360), .B2(new_n365), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n321), .B1(new_n366), .B2(new_n662), .ZN(new_n663));
  OAI211_X1 g477(.A(new_n377), .B(new_n378), .C1(new_n355), .C2(new_n352), .ZN(new_n664));
  AOI211_X1 g478(.A(G469), .B(G902), .C1(new_n663), .C2(new_n664), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n317), .B1(new_n661), .B2(new_n665), .ZN(new_n666));
  NOR2_X1   g480(.A1(new_n666), .A2(new_n568), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n649), .A2(new_n660), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g482(.A(KEYINPUT34), .B(G104), .ZN(new_n669));
  XOR2_X1   g483(.A(new_n669), .B(KEYINPUT97), .Z(new_n670));
  XNOR2_X1  g484(.A(new_n668), .B(new_n670), .ZN(G6));
  NAND2_X1  g485(.A1(new_n449), .A2(KEYINPUT98), .ZN(new_n672));
  INV_X1    g486(.A(KEYINPUT98), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n448), .A2(new_n673), .A3(KEYINPUT20), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n442), .A2(new_n447), .ZN(new_n675));
  INV_X1    g489(.A(new_n450), .ZN(new_n676));
  OAI211_X1 g490(.A(new_n672), .B(new_n674), .C1(new_n675), .C2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n431), .ZN(new_n678));
  INV_X1    g492(.A(new_n505), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n677), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  NOR2_X1   g494(.A1(new_n680), .A2(new_n314), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n649), .A2(new_n667), .A3(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT35), .B(G107), .Z(new_n683));
  XOR2_X1   g497(.A(new_n683), .B(KEYINPUT99), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n682), .B(new_n684), .ZN(G9));
  INV_X1    g499(.A(KEYINPUT100), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n548), .A2(new_n543), .ZN(new_n687));
  NOR2_X1   g501(.A1(new_n516), .A2(KEYINPUT36), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n689), .A2(new_n566), .ZN(new_n690));
  INV_X1    g504(.A(new_n690), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n552), .A2(KEYINPUT79), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n692), .A2(KEYINPUT25), .A3(new_n560), .ZN(new_n693));
  AOI21_X1  g507(.A(new_n557), .B1(new_n562), .B2(new_n553), .ZN(new_n694));
  AOI211_X1 g508(.A(new_n686), .B(new_n691), .C1(new_n693), .C2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(KEYINPUT100), .B1(new_n563), .B2(new_n690), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n507), .A2(new_n511), .A3(new_n649), .A4(new_n697), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT37), .B(G110), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n698), .B(new_n699), .ZN(G12));
  AOI21_X1  g514(.A(new_n666), .B1(new_n636), .B2(new_n641), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n191), .B1(G900), .B2(new_n194), .ZN(new_n702));
  NAND4_X1  g516(.A1(new_n677), .A2(new_n678), .A3(new_n679), .A4(new_n702), .ZN(new_n703));
  OAI21_X1  g517(.A(new_n187), .B1(new_n312), .B2(new_n313), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n701), .A2(new_n697), .A3(new_n705), .ZN(new_n706));
  XNOR2_X1  g520(.A(new_n706), .B(G128), .ZN(G30));
  XNOR2_X1  g521(.A(new_n702), .B(KEYINPUT39), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n388), .A2(new_n708), .ZN(new_n709));
  XOR2_X1   g523(.A(new_n709), .B(KEYINPUT40), .Z(new_n710));
  INV_X1    g524(.A(KEYINPUT101), .ZN(new_n711));
  NAND2_X1  g525(.A1(new_n298), .A2(new_n310), .ZN(new_n712));
  INV_X1    g526(.A(new_n311), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND3_X1  g528(.A1(new_n298), .A2(new_n310), .A3(new_n311), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(KEYINPUT38), .ZN(new_n717));
  AOI21_X1  g531(.A(new_n691), .B1(new_n693), .B2(new_n694), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n452), .A2(new_n505), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n631), .A2(new_n635), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n615), .A2(new_n626), .ZN(new_n722));
  OAI21_X1  g536(.A(new_n309), .B1(new_n594), .B2(new_n587), .ZN(new_n723));
  OAI21_X1  g537(.A(G472), .B1(new_n722), .B2(new_n723), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n641), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n717), .A2(new_n187), .A3(new_n720), .A4(new_n725), .ZN(new_n726));
  OAI21_X1  g540(.A(new_n710), .B1(new_n711), .B2(new_n726), .ZN(new_n727));
  AND2_X1   g541(.A1(new_n726), .A2(new_n711), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(new_n327), .ZN(G45));
  INV_X1    g544(.A(new_n452), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n731), .B(new_n702), .C1(new_n658), .C2(new_n657), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n704), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n701), .A2(new_n697), .A3(new_n733), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G146), .ZN(G48));
  NAND2_X1  g549(.A1(new_n663), .A2(new_n664), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n383), .B1(new_n736), .B2(new_n309), .ZN(new_n737));
  NOR3_X1   g551(.A1(new_n737), .A2(new_n665), .A3(new_n318), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n642), .A2(new_n660), .A3(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(KEYINPUT41), .B(G113), .ZN(new_n740));
  XNOR2_X1  g554(.A(new_n739), .B(new_n740), .ZN(G15));
  NAND3_X1  g555(.A1(new_n642), .A2(new_n681), .A3(new_n738), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G116), .ZN(G18));
  NAND2_X1  g557(.A1(new_n620), .A2(G472), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n633), .B1(new_n645), .B2(new_n628), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n744), .B(new_n721), .C1(new_n745), .C2(KEYINPUT32), .ZN(new_n746));
  OAI21_X1  g560(.A(new_n309), .B1(new_n385), .B2(new_n386), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(G469), .ZN(new_n748));
  NAND3_X1  g562(.A1(new_n748), .A2(new_n317), .A3(new_n387), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n452), .A2(new_n505), .ZN(new_n750));
  NOR2_X1   g564(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  NAND4_X1  g565(.A1(new_n697), .A2(new_n315), .A3(new_n746), .A4(new_n751), .ZN(new_n752));
  XNOR2_X1  g566(.A(new_n752), .B(G119), .ZN(G21));
  INV_X1    g567(.A(new_n187), .ZN(new_n754));
  AOI21_X1  g568(.A(new_n754), .B1(new_n714), .B2(new_n715), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n738), .A2(new_n755), .A3(new_n195), .A4(new_n719), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n693), .A2(new_n694), .B1(new_n565), .B2(new_n566), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n632), .B(KEYINPUT102), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n625), .A2(new_n630), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT28), .B1(new_n596), .B2(new_n597), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n760), .A2(KEYINPUT72), .ZN(new_n761));
  NAND2_X1  g575(.A1(new_n761), .A2(new_n598), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n587), .B1(new_n762), .B2(new_n583), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n758), .B1(new_n759), .B2(new_n763), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n757), .B(new_n764), .C1(new_n646), .C2(new_n647), .ZN(new_n765));
  OAI21_X1  g579(.A(KEYINPUT103), .B1(new_n756), .B2(new_n765), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n647), .B1(new_n631), .B2(new_n309), .ZN(new_n767));
  INV_X1    g581(.A(new_n758), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n762), .A2(new_n583), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(new_n626), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n768), .B1(new_n770), .B2(new_n645), .ZN(new_n771));
  NOR3_X1   g585(.A1(new_n767), .A2(new_n568), .A3(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n719), .A2(new_n317), .A3(new_n387), .A4(new_n748), .ZN(new_n773));
  NOR2_X1   g587(.A1(new_n773), .A2(new_n314), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT103), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n772), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n766), .A2(new_n776), .ZN(new_n777));
  XOR2_X1   g591(.A(KEYINPUT104), .B(G122), .Z(new_n778));
  XNOR2_X1  g592(.A(new_n777), .B(new_n778), .ZN(G24));
  NOR3_X1   g593(.A1(new_n767), .A2(new_n718), .A3(new_n771), .ZN(new_n780));
  INV_X1    g594(.A(new_n732), .ZN(new_n781));
  NOR2_X1   g595(.A1(new_n749), .A2(new_n704), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G125), .ZN(G27));
  NAND3_X1  g598(.A1(new_n714), .A2(new_n187), .A3(new_n715), .ZN(new_n785));
  AOI211_X1 g599(.A(new_n785), .B(new_n568), .C1(new_n636), .C2(new_n641), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n786), .A2(KEYINPUT42), .A3(new_n388), .A4(new_n781), .ZN(new_n787));
  INV_X1    g601(.A(KEYINPUT42), .ZN(new_n788));
  INV_X1    g602(.A(new_n785), .ZN(new_n789));
  NAND4_X1  g603(.A1(new_n746), .A2(new_n388), .A3(new_n757), .A4(new_n789), .ZN(new_n790));
  OAI21_X1  g604(.A(new_n788), .B1(new_n790), .B2(new_n732), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G131), .ZN(G33));
  INV_X1    g607(.A(new_n703), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n642), .A2(new_n388), .A3(new_n794), .A4(new_n789), .ZN(new_n795));
  XNOR2_X1  g609(.A(new_n795), .B(G134), .ZN(G36));
  NAND2_X1  g610(.A1(new_n367), .A2(new_n379), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n383), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n798), .B2(new_n797), .ZN(new_n800));
  NAND2_X1  g614(.A1(new_n800), .A2(new_n381), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n665), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(KEYINPUT46), .A3(new_n381), .ZN(new_n804));
  AOI21_X1  g618(.A(new_n318), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n708), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(KEYINPUT105), .ZN(new_n807));
  NOR2_X1   g621(.A1(new_n659), .A2(new_n731), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT43), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT106), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n809), .A2(new_n810), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n810), .ZN(new_n812));
  NOR2_X1   g626(.A1(new_n649), .A2(new_n718), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT44), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n785), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n807), .B(new_n816), .C1(new_n815), .C2(new_n814), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(G137), .ZN(G39));
  NAND2_X1  g632(.A1(KEYINPUT107), .A2(KEYINPUT47), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n805), .A2(new_n819), .ZN(new_n820));
  NOR4_X1   g634(.A1(new_n746), .A2(new_n757), .A3(new_n732), .A4(new_n785), .ZN(new_n821));
  XOR2_X1   g635(.A(KEYINPUT107), .B(KEYINPUT47), .Z(new_n822));
  OAI211_X1 g636(.A(new_n820), .B(new_n821), .C1(new_n805), .C2(new_n822), .ZN(new_n823));
  XNOR2_X1  g637(.A(new_n823), .B(G140), .ZN(G42));
  NOR2_X1   g638(.A1(new_n725), .A2(new_n568), .ZN(new_n825));
  NOR3_X1   g639(.A1(new_n749), .A2(new_n785), .A3(new_n191), .ZN(new_n826));
  AND2_X1   g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI211_X1 g641(.A(new_n827), .B(new_n731), .C1(new_n658), .C2(new_n657), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(new_n189), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n809), .A2(new_n642), .A3(new_n826), .ZN(new_n830));
  XOR2_X1   g644(.A(new_n830), .B(KEYINPUT48), .Z(new_n831));
  AND4_X1   g645(.A1(new_n190), .A2(new_n809), .A3(new_n189), .A4(new_n772), .ZN(new_n832));
  AOI211_X1 g646(.A(new_n829), .B(new_n831), .C1(new_n782), .C2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n827), .A2(new_n452), .A3(new_n659), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n809), .A2(new_n780), .A3(new_n826), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n820), .B1(new_n805), .B2(new_n822), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n737), .A2(new_n665), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  OAI21_X1  g654(.A(new_n838), .B1(new_n317), .B2(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n832), .A2(new_n789), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n837), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  NOR3_X1   g657(.A1(new_n717), .A2(new_n187), .A3(new_n749), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n832), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g659(.A(KEYINPUT50), .B1(new_n845), .B2(KEYINPUT113), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n846), .B1(KEYINPUT113), .B2(new_n845), .ZN(new_n847));
  INV_X1    g661(.A(KEYINPUT50), .ZN(new_n848));
  OAI22_X1  g662(.A1(new_n847), .A2(KEYINPUT114), .B1(new_n848), .B2(new_n845), .ZN(new_n849));
  AND2_X1   g663(.A1(new_n847), .A2(KEYINPUT114), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n834), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT115), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(KEYINPUT115), .B1(new_n851), .B2(new_n834), .ZN(new_n855));
  OAI221_X1 g669(.A(new_n833), .B1(new_n834), .B2(new_n851), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT110), .ZN(new_n857));
  OAI211_X1 g671(.A(new_n701), .B(new_n697), .C1(new_n705), .C2(new_n733), .ZN(new_n858));
  INV_X1    g672(.A(new_n702), .ZN(new_n859));
  NOR3_X1   g673(.A1(new_n666), .A2(new_n704), .A3(new_n859), .ZN(new_n860));
  NAND3_X1  g674(.A1(new_n860), .A2(new_n720), .A3(new_n725), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n858), .A2(new_n783), .A3(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT109), .ZN(new_n863));
  XNOR2_X1  g677(.A(KEYINPUT108), .B(KEYINPUT52), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n858), .A2(KEYINPUT52), .A3(new_n783), .A4(new_n861), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(new_n866), .ZN(new_n867));
  AOI21_X1  g681(.A(new_n863), .B1(new_n862), .B2(new_n864), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n857), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n862), .A2(new_n864), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(KEYINPUT109), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n871), .A2(KEYINPUT110), .A3(new_n866), .A4(new_n865), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT112), .ZN(new_n874));
  AND2_X1   g688(.A1(new_n766), .A2(new_n776), .ZN(new_n875));
  OAI211_X1 g689(.A(new_n642), .B(new_n738), .C1(new_n660), .C2(new_n681), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n876), .A2(new_n752), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n874), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n777), .A2(KEYINPUT112), .A3(new_n752), .A4(new_n876), .ZN(new_n879));
  INV_X1    g693(.A(KEYINPUT53), .ZN(new_n880));
  AOI21_X1  g694(.A(new_n880), .B1(new_n787), .B2(new_n791), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n878), .A2(new_n879), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT111), .ZN(new_n883));
  OAI21_X1  g697(.A(new_n309), .B1(new_n497), .B2(new_n499), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(new_n456), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n859), .B1(new_n885), .B2(new_n500), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n677), .A2(new_n678), .A3(new_n886), .ZN(new_n887));
  AOI21_X1  g701(.A(new_n887), .B1(new_n636), .B2(new_n641), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n697), .A2(new_n888), .B1(new_n780), .B2(new_n781), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n789), .A2(new_n388), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n795), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n659), .A2(new_n731), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n892), .A2(new_n750), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n893), .A2(new_n314), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n894), .A2(new_n649), .A3(new_n667), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n698), .A2(new_n643), .A3(new_n895), .ZN(new_n896));
  OAI21_X1  g710(.A(new_n883), .B1(new_n891), .B2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n891), .A2(new_n896), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT111), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n882), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND2_X1  g714(.A1(new_n873), .A2(new_n900), .ZN(new_n901));
  INV_X1    g715(.A(KEYINPUT52), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n862), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(new_n866), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n875), .A2(new_n877), .ZN(new_n905));
  NAND4_X1  g719(.A1(new_n904), .A2(new_n898), .A3(new_n792), .A4(new_n905), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n906), .A2(new_n880), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n901), .A2(new_n907), .ZN(new_n908));
  OR2_X1    g722(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n909));
  AND3_X1   g723(.A1(new_n898), .A2(new_n792), .A3(new_n905), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n873), .A2(new_n880), .A3(new_n910), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n906), .A2(KEYINPUT53), .ZN(new_n912));
  NAND3_X1  g726(.A1(new_n911), .A2(KEYINPUT54), .A3(new_n912), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  OAI22_X1  g728(.A1(new_n856), .A2(new_n914), .B1(G952), .B2(G953), .ZN(new_n915));
  XNOR2_X1  g729(.A(new_n839), .B(KEYINPUT49), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n916), .A2(new_n187), .A3(new_n317), .A4(new_n808), .ZN(new_n917));
  NOR2_X1   g731(.A1(new_n917), .A2(new_n717), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n825), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n915), .A2(new_n919), .ZN(G75));
  NOR2_X1   g734(.A1(new_n188), .A2(G952), .ZN(new_n921));
  INV_X1    g735(.A(new_n921), .ZN(new_n922));
  AOI22_X1  g736(.A1(new_n873), .A2(new_n900), .B1(new_n880), .B2(new_n906), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n923), .A2(new_n309), .ZN(new_n924));
  AOI21_X1  g738(.A(KEYINPUT56), .B1(new_n924), .B2(G210), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n250), .A2(new_n297), .ZN(new_n926));
  XNOR2_X1  g740(.A(new_n926), .B(new_n295), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n927), .B(KEYINPUT55), .ZN(new_n928));
  OAI21_X1  g742(.A(new_n922), .B1(new_n925), .B2(new_n928), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n925), .B2(new_n928), .ZN(G51));
  AND2_X1   g744(.A1(new_n908), .A2(KEYINPUT54), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT116), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n931), .B1(new_n909), .B2(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(new_n932), .B2(new_n909), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n381), .B(KEYINPUT57), .Z(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(new_n736), .ZN(new_n937));
  OR3_X1    g751(.A1(new_n923), .A2(new_n309), .A3(new_n800), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n921), .B1(new_n937), .B2(new_n938), .ZN(G54));
  NAND3_X1  g753(.A1(new_n924), .A2(KEYINPUT58), .A3(G475), .ZN(new_n940));
  AND2_X1   g754(.A1(new_n940), .A2(new_n675), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n675), .ZN(new_n942));
  NOR3_X1   g756(.A1(new_n941), .A2(new_n942), .A3(new_n921), .ZN(G60));
  NAND2_X1  g757(.A1(new_n653), .A2(new_n656), .ZN(new_n944));
  XNOR2_X1  g758(.A(KEYINPUT117), .B(KEYINPUT59), .ZN(new_n945));
  NOR2_X1   g759(.A1(new_n453), .A2(new_n309), .ZN(new_n946));
  XOR2_X1   g760(.A(new_n945), .B(new_n946), .Z(new_n947));
  INV_X1    g761(.A(new_n947), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n944), .B1(new_n914), .B2(new_n948), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n947), .B1(new_n653), .B2(new_n656), .ZN(new_n950));
  AOI211_X1 g764(.A(new_n921), .B(new_n949), .C1(new_n934), .C2(new_n950), .ZN(G63));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g766(.A1(G217), .A2(G902), .ZN(new_n953));
  XNOR2_X1  g767(.A(new_n953), .B(KEYINPUT60), .ZN(new_n954));
  OAI21_X1  g768(.A(KEYINPUT119), .B1(new_n923), .B2(new_n954), .ZN(new_n955));
  INV_X1    g769(.A(KEYINPUT119), .ZN(new_n956));
  INV_X1    g770(.A(new_n954), .ZN(new_n957));
  AND2_X1   g771(.A1(new_n881), .A2(new_n879), .ZN(new_n958));
  INV_X1    g772(.A(new_n896), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n780), .A2(new_n781), .ZN(new_n960));
  INV_X1    g774(.A(new_n696), .ZN(new_n961));
  INV_X1    g775(.A(new_n887), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n718), .A2(KEYINPUT100), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n746), .A2(new_n961), .A3(new_n962), .A4(new_n963), .ZN(new_n964));
  AOI21_X1  g778(.A(new_n890), .B1(new_n960), .B2(new_n964), .ZN(new_n965));
  INV_X1    g779(.A(new_n795), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n965), .A2(new_n966), .ZN(new_n967));
  AOI21_X1  g781(.A(KEYINPUT111), .B1(new_n959), .B2(new_n967), .ZN(new_n968));
  NOR3_X1   g782(.A1(new_n891), .A2(new_n896), .A3(new_n883), .ZN(new_n969));
  OAI211_X1 g783(.A(new_n958), .B(new_n878), .C1(new_n968), .C2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n970), .B1(new_n869), .B2(new_n872), .ZN(new_n971));
  INV_X1    g785(.A(new_n907), .ZN(new_n972));
  OAI211_X1 g786(.A(new_n956), .B(new_n957), .C1(new_n971), .C2(new_n972), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n955), .A2(new_n973), .A3(new_n564), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n974), .A2(KEYINPUT121), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT121), .ZN(new_n976));
  NAND4_X1  g790(.A1(new_n955), .A2(new_n973), .A3(new_n976), .A4(new_n564), .ZN(new_n977));
  AND2_X1   g791(.A1(new_n975), .A2(new_n977), .ZN(new_n978));
  AOI21_X1  g792(.A(new_n956), .B1(new_n908), .B2(new_n957), .ZN(new_n979));
  NOR3_X1   g793(.A1(new_n923), .A2(KEYINPUT119), .A3(new_n954), .ZN(new_n980));
  OAI21_X1  g794(.A(new_n689), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n922), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n952), .B1(new_n978), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n975), .A2(new_n977), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n981), .A2(KEYINPUT61), .A3(new_n922), .ZN(new_n985));
  NOR3_X1   g799(.A1(new_n984), .A2(new_n985), .A3(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n955), .A2(new_n973), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n921), .B1(new_n987), .B2(new_n689), .ZN(new_n988));
  NAND2_X1  g802(.A1(new_n988), .A2(new_n974), .ZN(new_n989));
  XNOR2_X1  g803(.A(KEYINPUT118), .B(KEYINPUT61), .ZN(new_n990));
  INV_X1    g804(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g805(.A(KEYINPUT120), .B1(new_n989), .B2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(KEYINPUT120), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n993), .B(new_n990), .C1(new_n988), .C2(new_n974), .ZN(new_n994));
  OAI22_X1  g808(.A1(new_n983), .A2(new_n986), .B1(new_n992), .B2(new_n994), .ZN(G66));
  AOI21_X1  g809(.A(new_n188), .B1(new_n193), .B2(G224), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n905), .A2(new_n959), .ZN(new_n997));
  AOI21_X1  g811(.A(new_n996), .B1(new_n997), .B2(new_n188), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n926), .B1(G898), .B2(new_n188), .ZN(new_n999));
  XOR2_X1   g813(.A(new_n999), .B(KEYINPUT123), .Z(new_n1000));
  XNOR2_X1  g814(.A(new_n998), .B(new_n1000), .ZN(G69));
  INV_X1    g815(.A(KEYINPUT125), .ZN(new_n1002));
  NAND2_X1  g816(.A1(new_n858), .A2(new_n783), .ZN(new_n1003));
  OR3_X1    g817(.A1(new_n729), .A2(KEYINPUT62), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g818(.A(new_n823), .ZN(new_n1005));
  NOR2_X1   g819(.A1(new_n709), .A2(new_n893), .ZN(new_n1006));
  AOI21_X1  g820(.A(new_n1005), .B1(new_n786), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g821(.A(KEYINPUT62), .B1(new_n729), .B2(new_n1003), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1004), .A2(new_n817), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1009), .A2(new_n188), .ZN(new_n1010));
  NAND2_X1  g824(.A1(new_n612), .A2(new_n613), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n605), .A2(new_n1011), .ZN(new_n1012));
  XNOR2_X1  g826(.A(new_n1012), .B(KEYINPUT124), .ZN(new_n1013));
  NOR2_X1   g827(.A1(new_n437), .A2(new_n438), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n1002), .B1(new_n1010), .B2(new_n1015), .ZN(new_n1016));
  AOI21_X1  g830(.A(new_n1015), .B1(G900), .B2(G953), .ZN(new_n1017));
  NAND4_X1  g831(.A1(new_n807), .A2(new_n755), .A3(new_n642), .A4(new_n719), .ZN(new_n1018));
  AOI211_X1 g832(.A(new_n966), .B(new_n1003), .C1(new_n791), .C2(new_n787), .ZN(new_n1019));
  NAND4_X1  g833(.A1(new_n817), .A2(new_n1018), .A3(new_n823), .A4(new_n1019), .ZN(new_n1020));
  OAI21_X1  g834(.A(new_n1017), .B1(new_n1020), .B2(G953), .ZN(new_n1021));
  NAND2_X1  g835(.A1(new_n1016), .A2(new_n1021), .ZN(new_n1022));
  OR2_X1    g836(.A1(new_n1022), .A2(KEYINPUT126), .ZN(new_n1023));
  NAND2_X1  g837(.A1(new_n1022), .A2(KEYINPUT126), .ZN(new_n1024));
  NAND2_X1  g838(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n188), .B1(G227), .B2(G900), .ZN(new_n1026));
  INV_X1    g840(.A(new_n1026), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1023), .A2(new_n1026), .A3(new_n1024), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n1028), .A2(new_n1029), .ZN(G72));
  NAND2_X1  g844(.A1(G472), .A2(G902), .ZN(new_n1031));
  XOR2_X1   g845(.A(new_n1031), .B(KEYINPUT63), .Z(new_n1032));
  OAI21_X1  g846(.A(new_n1032), .B1(new_n1009), .B2(new_n997), .ZN(new_n1033));
  AOI21_X1  g847(.A(new_n921), .B1(new_n1033), .B2(new_n722), .ZN(new_n1034));
  AND2_X1   g848(.A1(new_n615), .A2(new_n626), .ZN(new_n1035));
  INV_X1    g849(.A(new_n1032), .ZN(new_n1036));
  NOR3_X1   g850(.A1(new_n1035), .A2(new_n722), .A3(new_n1036), .ZN(new_n1037));
  XOR2_X1   g851(.A(new_n1037), .B(KEYINPUT127), .Z(new_n1038));
  NAND3_X1  g852(.A1(new_n911), .A2(new_n912), .A3(new_n1038), .ZN(new_n1039));
  OAI21_X1  g853(.A(new_n1032), .B1(new_n1020), .B2(new_n997), .ZN(new_n1040));
  NAND2_X1  g854(.A1(new_n1040), .A2(new_n1035), .ZN(new_n1041));
  AND3_X1   g855(.A1(new_n1034), .A2(new_n1039), .A3(new_n1041), .ZN(G57));
endmodule


