//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 1 0 1 0 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 1 1 0 0 0 1 1 1 0 1 0 1 0 1 1 1 1 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:27 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1101, new_n1102, new_n1103, new_n1104, new_n1105,
    new_n1106, new_n1107, new_n1108, new_n1109, new_n1110, new_n1111,
    new_n1112, new_n1113, new_n1114, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1141, new_n1142,
    new_n1143, new_n1144, new_n1145, new_n1146, new_n1147, new_n1148,
    new_n1149, new_n1150, new_n1151, new_n1152, new_n1153, new_n1154,
    new_n1155, new_n1156, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1296, new_n1297, new_n1298, new_n1299, new_n1300, new_n1301,
    new_n1302, new_n1303, new_n1304, new_n1305, new_n1306, new_n1307,
    new_n1308, new_n1309, new_n1310, new_n1311, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1320,
    new_n1321, new_n1322, new_n1323, new_n1324, new_n1325, new_n1326,
    new_n1328, new_n1329, new_n1330, new_n1331, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1374, new_n1375, new_n1376, new_n1377,
    new_n1378, new_n1379, new_n1380, new_n1381, new_n1382, new_n1383,
    new_n1384, new_n1385, new_n1386, new_n1387, new_n1388, new_n1389,
    new_n1390, new_n1391;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  OAI21_X1  g0012(.A(G50), .B1(G58), .B2(G68), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n215), .A2(new_n207), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n218));
  INV_X1    g0018(.A(G68), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n218), .B1(new_n219), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  INV_X1    g0024(.A(G77), .ZN(new_n225));
  INV_X1    g0025(.A(G244), .ZN(new_n226));
  INV_X1    g0026(.A(G107), .ZN(new_n227));
  INV_X1    g0027(.A(G264), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n224), .B1(new_n225), .B2(new_n226), .C1(new_n227), .C2(new_n228), .ZN(new_n229));
  OAI21_X1  g0029(.A(new_n209), .B1(new_n223), .B2(new_n229), .ZN(new_n230));
  OAI211_X1 g0030(.A(new_n212), .B(new_n217), .C1(KEYINPUT1), .C2(new_n230), .ZN(new_n231));
  AOI21_X1  g0031(.A(new_n231), .B1(KEYINPUT1), .B2(new_n230), .ZN(G361));
  XOR2_X1   g0032(.A(G250), .B(G257), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n233), .B(KEYINPUT64), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G264), .B(G270), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n236), .B(new_n241), .ZN(G358));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n243), .B(KEYINPUT65), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XOR2_X1   g0046(.A(G87), .B(G97), .Z(new_n247));
  XNOR2_X1  g0047(.A(G107), .B(G116), .ZN(new_n248));
  XOR2_X1   g0048(.A(new_n247), .B(new_n248), .Z(new_n249));
  XNOR2_X1  g0049(.A(new_n246), .B(new_n249), .ZN(G351));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n215), .ZN(new_n252));
  XNOR2_X1  g0052(.A(KEYINPUT8), .B(G58), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n207), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(G150), .ZN(new_n255));
  INV_X1    g0055(.A(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n207), .A2(new_n256), .ZN(new_n257));
  OAI22_X1  g0057(.A1(new_n253), .A2(new_n254), .B1(new_n255), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n203), .A2(G20), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g0060(.A(new_n252), .B1(new_n258), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g0061(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n262));
  INV_X1    g0062(.A(new_n262), .ZN(new_n263));
  NOR2_X1   g0063(.A1(new_n263), .A2(new_n252), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n207), .A2(G1), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(new_n202), .ZN(new_n266));
  AOI22_X1  g0066(.A1(new_n264), .A2(new_n266), .B1(new_n202), .B2(new_n263), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n261), .A2(KEYINPUT70), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  AOI21_X1  g0069(.A(KEYINPUT70), .B1(new_n261), .B2(new_n267), .ZN(new_n270));
  NOR2_X1   g0070(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AND2_X1   g0071(.A1(G33), .A2(G41), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n272), .A2(new_n215), .ZN(new_n273));
  XNOR2_X1  g0073(.A(KEYINPUT3), .B(G33), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT66), .ZN(new_n275));
  INV_X1    g0075(.A(G1698), .ZN(new_n276));
  NAND4_X1  g0076(.A1(new_n274), .A2(new_n275), .A3(G222), .A4(new_n276), .ZN(new_n277));
  NAND3_X1  g0077(.A1(new_n274), .A2(G222), .A3(new_n276), .ZN(new_n278));
  INV_X1    g0078(.A(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(KEYINPUT66), .B1(new_n282), .B2(G77), .ZN(new_n283));
  OAI21_X1  g0083(.A(new_n277), .B1(new_n279), .B2(new_n283), .ZN(new_n284));
  INV_X1    g0084(.A(G223), .ZN(new_n285));
  OAI21_X1  g0085(.A(KEYINPUT67), .B1(new_n282), .B2(new_n276), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT67), .ZN(new_n287));
  OAI211_X1 g0087(.A(new_n287), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n288));
  AOI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g0089(.A(new_n273), .B1(new_n284), .B2(new_n289), .ZN(new_n290));
  INV_X1    g0090(.A(G41), .ZN(new_n291));
  INV_X1    g0091(.A(G45), .ZN(new_n292));
  AOI21_X1  g0092(.A(G1), .B1(new_n291), .B2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(G33), .A2(G41), .ZN(new_n294));
  NAND3_X1  g0094(.A1(new_n294), .A2(G1), .A3(G13), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n293), .A2(new_n295), .A3(G274), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(new_n299), .ZN(new_n300));
  AOI21_X1  g0100(.A(new_n297), .B1(G226), .B2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n290), .A2(new_n301), .ZN(new_n302));
  AOI22_X1  g0102(.A1(new_n271), .A2(KEYINPUT9), .B1(new_n302), .B2(G200), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n290), .A2(G190), .A3(new_n301), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT9), .ZN(new_n306));
  OAI21_X1  g0106(.A(new_n306), .B1(new_n269), .B2(new_n270), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n303), .A2(new_n304), .A3(new_n305), .A4(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(new_n301), .ZN(new_n309));
  AOI21_X1  g0109(.A(new_n287), .B1(new_n274), .B2(G1698), .ZN(new_n310));
  INV_X1    g0110(.A(new_n288), .ZN(new_n311));
  OAI21_X1  g0111(.A(G223), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  OAI211_X1 g0112(.A(new_n312), .B(new_n277), .C1(new_n283), .C2(new_n279), .ZN(new_n313));
  AOI21_X1  g0113(.A(new_n309), .B1(new_n313), .B2(new_n273), .ZN(new_n314));
  INV_X1    g0114(.A(G200), .ZN(new_n315));
  INV_X1    g0115(.A(KEYINPUT70), .ZN(new_n316));
  INV_X1    g0116(.A(new_n252), .ZN(new_n317));
  NOR2_X1   g0117(.A1(new_n257), .A2(new_n255), .ZN(new_n318));
  XOR2_X1   g0118(.A(KEYINPUT8), .B(G58), .Z(new_n319));
  INV_X1    g0119(.A(new_n254), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n318), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n317), .B1(new_n321), .B2(new_n259), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n317), .A2(new_n262), .ZN(new_n323));
  INV_X1    g0123(.A(new_n266), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n323), .A2(new_n324), .B1(G50), .B2(new_n262), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n316), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n326), .A2(new_n268), .ZN(new_n327));
  OAI22_X1  g0127(.A1(new_n314), .A2(new_n315), .B1(new_n327), .B2(new_n306), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n307), .A2(new_n305), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT10), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n308), .A2(new_n330), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n302), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n261), .A2(new_n267), .ZN(new_n334));
  OAI211_X1 g0134(.A(new_n333), .B(new_n334), .C1(G179), .C2(new_n302), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n331), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G13), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n337), .A2(G1), .ZN(new_n338));
  NAND3_X1  g0138(.A1(new_n338), .A2(KEYINPUT68), .A3(G20), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT68), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n262), .A2(new_n340), .ZN(new_n341));
  AOI21_X1  g0141(.A(new_n252), .B1(new_n339), .B2(new_n341), .ZN(new_n342));
  INV_X1    g0142(.A(new_n265), .ZN(new_n343));
  AND3_X1   g0143(.A1(new_n342), .A2(G77), .A3(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n257), .ZN(new_n345));
  AOI22_X1  g0145(.A1(new_n319), .A2(new_n345), .B1(G20), .B2(G77), .ZN(new_n346));
  XNOR2_X1  g0146(.A(KEYINPUT15), .B(G87), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n320), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n317), .B1(new_n346), .B2(new_n349), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n339), .A2(new_n341), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n351), .A2(G77), .ZN(new_n352));
  OR3_X1    g0152(.A1(new_n344), .A2(new_n350), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT69), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n297), .B1(G244), .B2(new_n300), .ZN(new_n355));
  INV_X1    g0155(.A(new_n355), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n274), .A2(new_n276), .ZN(new_n357));
  OAI22_X1  g0157(.A1(new_n357), .A2(new_n238), .B1(new_n227), .B2(new_n274), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(G238), .B1(new_n310), .B2(new_n311), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n356), .B1(new_n361), .B2(new_n273), .ZN(new_n362));
  OAI211_X1 g0162(.A(new_n353), .B(new_n354), .C1(new_n362), .C2(G169), .ZN(new_n363));
  INV_X1    g0163(.A(G179), .ZN(new_n364));
  NAND2_X1  g0164(.A1(new_n362), .A2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n220), .B1(new_n286), .B2(new_n288), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n273), .B1(new_n366), .B2(new_n358), .ZN(new_n367));
  AOI21_X1  g0167(.A(G169), .B1(new_n367), .B2(new_n355), .ZN(new_n368));
  NOR3_X1   g0168(.A1(new_n344), .A2(new_n350), .A3(new_n352), .ZN(new_n369));
  OAI21_X1  g0169(.A(KEYINPUT69), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n365), .A3(new_n370), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n362), .A2(G190), .ZN(new_n372));
  OAI211_X1 g0172(.A(new_n372), .B(new_n369), .C1(new_n315), .C2(new_n362), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n371), .A2(new_n373), .ZN(new_n374));
  NOR2_X1   g0174(.A1(new_n336), .A2(new_n374), .ZN(new_n375));
  OR3_X1    g0175(.A1(new_n253), .A2(KEYINPUT77), .A3(new_n265), .ZN(new_n376));
  OAI21_X1  g0176(.A(KEYINPUT77), .B1(new_n253), .B2(new_n265), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n376), .A2(new_n264), .A3(new_n377), .ZN(new_n378));
  NAND2_X1  g0178(.A1(new_n253), .A2(new_n263), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  INV_X1    g0180(.A(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT76), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT7), .B1(new_n282), .B2(new_n207), .ZN(new_n383));
  INV_X1    g0183(.A(KEYINPUT3), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(new_n256), .ZN(new_n385));
  NAND2_X1  g0185(.A1(KEYINPUT3), .A2(G33), .ZN(new_n386));
  NAND4_X1  g0186(.A1(new_n385), .A2(KEYINPUT7), .A3(new_n207), .A4(new_n386), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  OAI21_X1  g0188(.A(G68), .B1(new_n383), .B2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(G58), .ZN(new_n390));
  NOR2_X1   g0190(.A1(new_n390), .A2(new_n219), .ZN(new_n391));
  OAI21_X1  g0191(.A(G20), .B1(new_n391), .B2(new_n201), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n345), .A2(G159), .ZN(new_n393));
  AND3_X1   g0193(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n394));
  AOI21_X1  g0194(.A(new_n382), .B1(new_n389), .B2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n385), .A2(new_n207), .A3(new_n386), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n219), .B1(new_n398), .B2(new_n387), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT16), .ZN(new_n400));
  NOR3_X1   g0200(.A1(new_n399), .A2(KEYINPUT76), .A3(new_n400), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n395), .A2(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(KEYINPUT16), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n392), .A2(new_n393), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n403), .B1(new_n399), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n405), .A2(new_n252), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n381), .B1(new_n402), .B2(new_n406), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n407), .A2(KEYINPUT78), .ZN(new_n408));
  INV_X1    g0208(.A(new_n404), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n389), .A2(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n317), .B1(new_n410), .B2(new_n403), .ZN(new_n411));
  OAI21_X1  g0211(.A(KEYINPUT76), .B1(new_n399), .B2(new_n400), .ZN(new_n412));
  NAND3_X1  g0212(.A1(new_n389), .A2(new_n382), .A3(new_n394), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n380), .B1(new_n411), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT78), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  INV_X1    g0217(.A(G226), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(G1698), .ZN(new_n419));
  OAI221_X1 g0219(.A(new_n419), .B1(G223), .B2(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n420));
  NAND2_X1  g0220(.A1(G33), .A2(G87), .ZN(new_n421));
  AOI21_X1  g0221(.A(new_n295), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(new_n296), .B1(new_n299), .B2(new_n238), .ZN(new_n423));
  NOR3_X1   g0223(.A1(new_n422), .A2(new_n423), .A3(new_n364), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n420), .A2(new_n421), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n425), .A2(new_n273), .ZN(new_n426));
  INV_X1    g0226(.A(new_n423), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n424), .B1(G169), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(new_n429), .ZN(new_n430));
  NAND3_X1  g0230(.A1(new_n408), .A2(new_n417), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT18), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT18), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n408), .A2(new_n433), .A3(new_n417), .A4(new_n430), .ZN(new_n434));
  AOI21_X1  g0234(.A(new_n315), .B1(new_n426), .B2(new_n427), .ZN(new_n435));
  INV_X1    g0235(.A(G190), .ZN(new_n436));
  NOR3_X1   g0236(.A1(new_n422), .A2(new_n423), .A3(new_n436), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n435), .A2(new_n437), .ZN(new_n438));
  OAI211_X1 g0238(.A(new_n438), .B(new_n381), .C1(new_n402), .C2(new_n406), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT17), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n415), .A2(KEYINPUT17), .A3(new_n438), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n432), .A2(new_n434), .A3(new_n444), .ZN(new_n445));
  INV_X1    g0245(.A(new_n445), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n219), .A2(G20), .ZN(new_n447));
  OAI221_X1 g0247(.A(new_n447), .B1(new_n254), .B2(new_n225), .C1(new_n202), .C2(new_n257), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(new_n252), .ZN(new_n449));
  XNOR2_X1  g0249(.A(new_n449), .B(KEYINPUT11), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n342), .A2(G68), .A3(new_n343), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  AND2_X1   g0252(.A1(new_n339), .A2(new_n341), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n453), .A2(new_n219), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n447), .A2(KEYINPUT12), .ZN(new_n455));
  AOI22_X1  g0255(.A1(new_n454), .A2(KEYINPUT12), .B1(new_n338), .B2(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n452), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT72), .ZN(new_n458));
  OAI21_X1  g0258(.A(G274), .B1(new_n272), .B2(new_n215), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n459), .B2(new_n298), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n293), .A2(new_n295), .A3(KEYINPUT72), .A4(G274), .ZN(new_n461));
  AOI22_X1  g0261(.A1(new_n460), .A2(new_n461), .B1(new_n300), .B2(G238), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT71), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n418), .A2(new_n276), .ZN(new_n464));
  NAND2_X1  g0264(.A1(new_n238), .A2(G1698), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n464), .B(new_n465), .C1(new_n280), .C2(new_n281), .ZN(new_n466));
  NAND2_X1  g0266(.A1(G33), .A2(G97), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n463), .B1(new_n468), .B2(new_n273), .ZN(new_n469));
  AOI211_X1 g0269(.A(KEYINPUT71), .B(new_n295), .C1(new_n466), .C2(new_n467), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n462), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n364), .B1(new_n471), .B2(KEYINPUT13), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n295), .B1(new_n466), .B2(new_n467), .ZN(new_n473));
  XNOR2_X1  g0273(.A(new_n473), .B(new_n463), .ZN(new_n474));
  INV_X1    g0274(.A(KEYINPUT13), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n474), .A2(KEYINPUT74), .A3(new_n475), .A4(new_n462), .ZN(new_n476));
  OAI211_X1 g0276(.A(new_n462), .B(new_n475), .C1(new_n469), .C2(new_n470), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT74), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g0279(.A1(new_n472), .A2(new_n476), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(KEYINPUT75), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT75), .ZN(new_n482));
  NAND4_X1  g0282(.A1(new_n472), .A2(new_n476), .A3(new_n479), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n481), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(KEYINPUT14), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n471), .A2(KEYINPUT13), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n486), .A2(new_n477), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n485), .B1(new_n487), .B2(G169), .ZN(new_n488));
  AOI211_X1 g0288(.A(KEYINPUT14), .B(new_n332), .C1(new_n486), .C2(new_n477), .ZN(new_n489));
  NOR2_X1   g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n457), .B1(new_n484), .B2(new_n490), .ZN(new_n491));
  NAND4_X1  g0291(.A1(new_n476), .A2(new_n479), .A3(G190), .A4(new_n486), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n492), .A2(new_n457), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n315), .B1(new_n486), .B2(new_n477), .ZN(new_n494));
  OR2_X1    g0294(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n495));
  NAND2_X1  g0295(.A1(new_n494), .A2(KEYINPUT73), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  AND3_X1   g0298(.A1(new_n375), .A2(new_n446), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(G33), .A2(G283), .ZN(new_n501));
  INV_X1    g0301(.A(G97), .ZN(new_n502));
  OAI211_X1 g0302(.A(new_n501), .B(new_n207), .C1(G33), .C2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT87), .ZN(new_n504));
  INV_X1    g0304(.A(G116), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(G20), .ZN(new_n506));
  AND3_X1   g0306(.A1(new_n252), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n504), .B1(new_n252), .B2(new_n506), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n503), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT20), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n509), .A2(new_n510), .ZN(new_n511));
  OAI211_X1 g0311(.A(KEYINPUT20), .B(new_n503), .C1(new_n507), .C2(new_n508), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT86), .ZN(new_n514));
  OAI21_X1  g0314(.A(new_n514), .B1(new_n351), .B2(G116), .ZN(new_n515));
  NAND4_X1  g0315(.A1(new_n339), .A2(new_n341), .A3(KEYINPUT86), .A4(new_n505), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n505), .B1(new_n206), .B2(G33), .ZN(new_n517));
  AOI22_X1  g0317(.A1(new_n515), .A2(new_n516), .B1(new_n342), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  NOR2_X1   g0319(.A1(new_n292), .A2(G1), .ZN(new_n520));
  AND2_X1   g0320(.A1(KEYINPUT5), .A2(G41), .ZN(new_n521));
  NOR2_X1   g0321(.A1(KEYINPUT5), .A2(G41), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n523), .A2(G270), .A3(new_n295), .ZN(new_n524));
  OR2_X1    g0324(.A1(KEYINPUT5), .A2(G41), .ZN(new_n525));
  NAND2_X1  g0325(.A1(KEYINPUT5), .A2(G41), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n527), .A2(G274), .A3(new_n295), .A4(new_n520), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n524), .A2(new_n528), .ZN(new_n529));
  OAI211_X1 g0329(.A(G264), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT85), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT85), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n274), .A2(new_n532), .A3(G264), .A4(G1698), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n282), .A2(G303), .ZN(new_n534));
  NAND3_X1  g0334(.A1(new_n274), .A2(G257), .A3(new_n276), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n531), .A2(new_n533), .A3(new_n534), .A4(new_n535), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n529), .B1(new_n536), .B2(new_n273), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n537), .A2(new_n332), .ZN(new_n538));
  AOI21_X1  g0338(.A(KEYINPUT21), .B1(new_n519), .B2(new_n538), .ZN(new_n539));
  INV_X1    g0339(.A(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n519), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n537), .A2(G190), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n536), .A2(new_n273), .ZN(new_n543));
  INV_X1    g0343(.A(new_n529), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(G200), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n541), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  AOI211_X1 g0347(.A(new_n364), .B(new_n529), .C1(new_n536), .C2(new_n273), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n519), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n519), .A2(new_n538), .A3(KEYINPUT21), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n540), .A2(new_n547), .A3(new_n549), .A4(new_n550), .ZN(new_n551));
  OAI211_X1 g0351(.A(G244), .B(G1698), .C1(new_n280), .C2(new_n281), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT84), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND4_X1  g0354(.A1(new_n274), .A2(KEYINPUT84), .A3(G244), .A4(G1698), .ZN(new_n555));
  NAND2_X1  g0355(.A1(G33), .A2(G116), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n274), .A2(G238), .A3(new_n276), .ZN(new_n557));
  NAND4_X1  g0357(.A1(new_n554), .A2(new_n555), .A3(new_n556), .A4(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n558), .A2(new_n273), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n206), .A2(G45), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n459), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(KEYINPUT82), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n563), .A2(new_n206), .A3(G45), .ZN(new_n564));
  NAND2_X1  g0364(.A1(new_n562), .A2(new_n564), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n295), .A2(G250), .ZN(new_n566));
  OAI21_X1  g0366(.A(KEYINPUT83), .B1(new_n565), .B2(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(new_n215), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n222), .B1(new_n568), .B2(new_n294), .ZN(new_n569));
  INV_X1    g0369(.A(KEYINPUT83), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n569), .A2(new_n570), .A3(new_n564), .A4(new_n562), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n561), .B1(new_n567), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n559), .A2(new_n572), .A3(G190), .ZN(new_n573));
  INV_X1    g0373(.A(KEYINPUT19), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n207), .B1(new_n467), .B2(new_n574), .ZN(new_n575));
  NOR2_X1   g0375(.A1(G97), .A2(G107), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n576), .A2(new_n221), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n207), .B(G68), .C1(new_n280), .C2(new_n281), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n574), .B1(new_n254), .B2(new_n502), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(new_n252), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n453), .A2(new_n347), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n264), .B1(G1), .B2(new_n256), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n585), .A2(new_n221), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n584), .A2(new_n586), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n573), .A2(new_n587), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n559), .A2(new_n572), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G200), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n264), .B(new_n348), .C1(G1), .C2(new_n256), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n582), .A2(new_n583), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(new_n592), .B1(new_n589), .B2(new_n332), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n559), .A2(new_n572), .A3(new_n364), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n588), .A2(new_n590), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  OAI21_X1  g0395(.A(G107), .B1(new_n383), .B2(new_n388), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT6), .ZN(new_n597));
  AND2_X1   g0397(.A1(G97), .A2(G107), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n597), .B1(new_n598), .B2(new_n576), .ZN(new_n599));
  NAND3_X1  g0399(.A1(new_n227), .A2(KEYINPUT6), .A3(G97), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  AOI22_X1  g0401(.A1(new_n601), .A2(G20), .B1(G77), .B2(new_n345), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  NAND2_X1  g0403(.A1(new_n603), .A2(new_n252), .ZN(new_n604));
  NOR2_X1   g0404(.A1(new_n262), .A2(G97), .ZN(new_n605));
  INV_X1    g0405(.A(new_n605), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n606), .B1(new_n585), .B2(new_n502), .ZN(new_n607));
  INV_X1    g0407(.A(new_n607), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n604), .A2(KEYINPUT81), .A3(new_n608), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT81), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n317), .B1(new_n596), .B2(new_n602), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n610), .B1(new_n611), .B2(new_n607), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(new_n501), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n276), .A2(G244), .ZN(new_n615));
  INV_X1    g0415(.A(KEYINPUT4), .ZN(new_n616));
  OAI22_X1  g0416(.A1(new_n615), .A2(new_n616), .B1(new_n222), .B2(new_n276), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n614), .B1(new_n617), .B2(new_n274), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n616), .A2(KEYINPUT79), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT79), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n620), .A2(KEYINPUT4), .ZN(new_n621));
  OAI211_X1 g0421(.A(new_n619), .B(new_n621), .C1(new_n282), .C2(new_n615), .ZN(new_n622));
  AOI21_X1  g0422(.A(new_n295), .B1(new_n618), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n523), .A2(new_n295), .ZN(new_n624));
  INV_X1    g0424(.A(G257), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n528), .B1(new_n624), .B2(new_n625), .ZN(new_n626));
  NOR2_X1   g0426(.A1(new_n623), .A2(new_n626), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(G179), .ZN(new_n628));
  OAI21_X1  g0428(.A(G169), .B1(new_n623), .B2(new_n626), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n613), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g0431(.A1(new_n585), .A2(new_n227), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n262), .A2(G107), .ZN(new_n633));
  XNOR2_X1  g0433(.A(new_n633), .B(KEYINPUT25), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  OAI211_X1 g0435(.A(new_n207), .B(G87), .C1(new_n280), .C2(new_n281), .ZN(new_n636));
  AND2_X1   g0436(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n637));
  NOR2_X1   g0437(.A1(KEYINPUT88), .A2(KEYINPUT22), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n636), .A2(new_n639), .ZN(new_n640));
  NAND4_X1  g0440(.A1(new_n274), .A2(new_n207), .A3(G87), .A4(new_n637), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n556), .A2(G20), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT23), .ZN(new_n643));
  OAI21_X1  g0443(.A(new_n643), .B1(new_n207), .B2(G107), .ZN(new_n644));
  NAND3_X1  g0444(.A1(new_n227), .A2(KEYINPUT23), .A3(G20), .ZN(new_n645));
  AOI21_X1  g0445(.A(new_n642), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n640), .A2(new_n641), .A3(new_n646), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(KEYINPUT24), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT24), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n640), .A2(new_n641), .A3(new_n646), .A4(new_n649), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n635), .B1(new_n252), .B2(new_n651), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT89), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n560), .B1(new_n525), .B2(new_n526), .ZN(new_n654));
  NOR3_X1   g0454(.A1(new_n654), .A2(new_n228), .A3(new_n273), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n222), .A2(new_n276), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n625), .A2(G1698), .ZN(new_n657));
  OAI211_X1 g0457(.A(new_n656), .B(new_n657), .C1(new_n280), .C2(new_n281), .ZN(new_n658));
  NAND2_X1  g0458(.A1(G33), .A2(G294), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n295), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n653), .B1(new_n655), .B2(new_n660), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n523), .A2(G264), .A3(new_n295), .ZN(new_n662));
  NOR2_X1   g0462(.A1(G250), .A2(G1698), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n663), .B1(new_n625), .B2(G1698), .ZN(new_n664));
  AOI22_X1  g0464(.A1(new_n664), .A2(new_n274), .B1(G33), .B2(G294), .ZN(new_n665));
  OAI211_X1 g0465(.A(KEYINPUT89), .B(new_n662), .C1(new_n665), .C2(new_n295), .ZN(new_n666));
  NAND3_X1  g0466(.A1(new_n661), .A2(new_n666), .A3(new_n528), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(new_n315), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n523), .A2(new_n459), .ZN(new_n669));
  NOR3_X1   g0469(.A1(new_n655), .A2(new_n660), .A3(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n670), .A2(KEYINPUT90), .A3(new_n436), .ZN(new_n671));
  INV_X1    g0471(.A(KEYINPUT90), .ZN(new_n672));
  OAI211_X1 g0472(.A(new_n528), .B(new_n662), .C1(new_n665), .C2(new_n295), .ZN(new_n673));
  OAI21_X1  g0473(.A(new_n672), .B1(new_n673), .B2(G190), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n652), .B1(new_n668), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(G200), .B1(new_n623), .B2(new_n626), .ZN(new_n677));
  OR2_X1    g0477(.A1(new_n677), .A2(KEYINPUT80), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n677), .A2(KEYINPUT80), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n611), .A2(new_n607), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n627), .A2(G190), .ZN(new_n681));
  NAND4_X1  g0481(.A1(new_n678), .A2(new_n679), .A3(new_n680), .A4(new_n681), .ZN(new_n682));
  NAND4_X1  g0482(.A1(new_n595), .A2(new_n631), .A3(new_n676), .A4(new_n682), .ZN(new_n683));
  NAND2_X1  g0483(.A1(new_n651), .A2(new_n252), .ZN(new_n684));
  AND2_X1   g0484(.A1(new_n632), .A2(new_n634), .ZN(new_n685));
  NAND4_X1  g0485(.A1(new_n661), .A2(new_n666), .A3(G179), .A4(new_n528), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n673), .A2(G169), .ZN(new_n687));
  AOI22_X1  g0487(.A1(new_n684), .A2(new_n685), .B1(new_n686), .B2(new_n687), .ZN(new_n688));
  NOR4_X1   g0488(.A1(new_n500), .A2(new_n551), .A3(new_n683), .A4(new_n688), .ZN(G372));
  INV_X1    g0489(.A(new_n335), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n497), .A2(new_n371), .ZN(new_n691));
  OAI21_X1  g0491(.A(new_n444), .B1(new_n691), .B2(new_n491), .ZN(new_n692));
  XNOR2_X1  g0492(.A(KEYINPUT91), .B(KEYINPUT18), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n407), .B2(new_n430), .ZN(new_n694));
  INV_X1    g0494(.A(new_n693), .ZN(new_n695));
  NOR3_X1   g0495(.A1(new_n415), .A2(new_n429), .A3(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n694), .A2(new_n696), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n692), .A2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(new_n690), .B1(new_n699), .B2(new_n331), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n684), .A2(new_n685), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n686), .A2(new_n687), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND4_X1  g0503(.A1(new_n540), .A2(new_n703), .A3(new_n549), .A4(new_n550), .ZN(new_n704));
  AND3_X1   g0504(.A1(new_n679), .A2(new_n680), .A3(new_n681), .ZN(new_n705));
  AOI22_X1  g0505(.A1(new_n705), .A2(new_n678), .B1(new_n613), .B2(new_n630), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n704), .A2(new_n706), .A3(new_n595), .A4(new_n676), .ZN(new_n707));
  INV_X1    g0507(.A(new_n592), .ZN(new_n708));
  AND2_X1   g0508(.A1(new_n559), .A2(new_n572), .ZN(new_n709));
  OAI211_X1 g0509(.A(new_n594), .B(new_n708), .C1(new_n709), .C2(G169), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n590), .A2(new_n587), .A3(new_n573), .ZN(new_n711));
  AOI22_X1  g0511(.A1(new_n628), .A2(new_n629), .B1(new_n604), .B2(new_n608), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT26), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n713), .A2(new_n714), .ZN(new_n715));
  AOI22_X1  g0515(.A1(new_n609), .A2(new_n612), .B1(new_n628), .B2(new_n629), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(KEYINPUT26), .A3(new_n710), .A4(new_n711), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n707), .A2(new_n710), .A3(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(new_n719), .ZN(new_n720));
  OAI21_X1  g0520(.A(new_n700), .B1(new_n500), .B2(new_n720), .ZN(G369));
  NAND2_X1  g0521(.A1(new_n338), .A2(new_n207), .ZN(new_n722));
  XNOR2_X1  g0522(.A(new_n722), .B(KEYINPUT92), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n723), .A2(KEYINPUT27), .ZN(new_n724));
  OAI21_X1  g0524(.A(G213), .B1(new_n723), .B2(KEYINPUT27), .ZN(new_n725));
  INV_X1    g0525(.A(G343), .ZN(new_n726));
  NOR3_X1   g0526(.A1(new_n724), .A2(new_n725), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n701), .A2(new_n727), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n676), .A2(new_n703), .A3(new_n728), .ZN(new_n729));
  INV_X1    g0529(.A(KEYINPUT93), .ZN(new_n730));
  OR2_X1    g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n729), .A2(new_n730), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n688), .A2(new_n727), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n724), .A2(new_n725), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G343), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n541), .A2(new_n738), .ZN(new_n739));
  OR2_X1    g0539(.A1(new_n551), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g0540(.A1(new_n540), .A2(new_n549), .A3(new_n550), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n739), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n740), .A2(new_n742), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G330), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n736), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n741), .A2(new_n738), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  NAND3_X1  g0547(.A1(new_n731), .A2(new_n747), .A3(new_n732), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n688), .A2(new_n738), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  OR2_X1    g0550(.A1(new_n745), .A2(new_n750), .ZN(G399));
  NAND2_X1  g0551(.A1(new_n210), .A2(new_n291), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n577), .A2(G116), .ZN(new_n753));
  NAND3_X1  g0553(.A1(new_n752), .A2(G1), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g0554(.A(new_n754), .B1(new_n213), .B2(new_n752), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT28), .ZN(new_n756));
  INV_X1    g0556(.A(KEYINPUT29), .ZN(new_n757));
  AND3_X1   g0557(.A1(new_n719), .A2(new_n757), .A3(new_n738), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n713), .A2(KEYINPUT26), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n595), .A2(new_n714), .A3(new_n716), .ZN(new_n761));
  NAND4_X1  g0561(.A1(new_n707), .A2(new_n710), .A3(new_n760), .A4(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n757), .B1(new_n762), .B2(new_n738), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  AND2_X1   g0564(.A1(new_n661), .A2(new_n666), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n548), .A2(new_n709), .A3(new_n627), .A4(new_n765), .ZN(new_n766));
  INV_X1    g0566(.A(KEYINPUT30), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AND3_X1   g0568(.A1(new_n559), .A2(new_n572), .A3(KEYINPUT94), .ZN(new_n769));
  AOI21_X1  g0569(.A(KEYINPUT94), .B1(new_n559), .B2(new_n572), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n226), .A2(G1698), .ZN(new_n772));
  AOI22_X1  g0572(.A1(new_n772), .A2(KEYINPUT4), .B1(G250), .B2(G1698), .ZN(new_n773));
  OAI21_X1  g0573(.A(new_n501), .B1(new_n773), .B2(new_n282), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n619), .A2(new_n621), .ZN(new_n775));
  AOI21_X1  g0575(.A(new_n775), .B1(new_n274), .B2(new_n772), .ZN(new_n776));
  OAI21_X1  g0576(.A(new_n273), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NOR2_X1   g0577(.A1(new_n654), .A2(new_n273), .ZN(new_n778));
  AOI21_X1  g0578(.A(new_n669), .B1(new_n778), .B2(G257), .ZN(new_n779));
  AOI21_X1  g0579(.A(G179), .B1(new_n777), .B2(new_n779), .ZN(new_n780));
  AND3_X1   g0580(.A1(new_n780), .A2(new_n667), .A3(new_n545), .ZN(new_n781));
  NAND2_X1  g0581(.A1(new_n771), .A2(new_n781), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n627), .A2(new_n661), .A3(new_n666), .ZN(new_n783));
  NAND4_X1  g0583(.A1(new_n783), .A2(KEYINPUT30), .A3(new_n548), .A4(new_n709), .ZN(new_n784));
  NAND3_X1  g0584(.A1(new_n768), .A2(new_n782), .A3(new_n784), .ZN(new_n785));
  AND3_X1   g0585(.A1(new_n785), .A2(KEYINPUT31), .A3(new_n727), .ZN(new_n786));
  AOI21_X1  g0586(.A(KEYINPUT31), .B1(new_n785), .B2(new_n727), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n786), .A2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n683), .ZN(new_n789));
  INV_X1    g0589(.A(new_n551), .ZN(new_n790));
  NAND4_X1  g0590(.A1(new_n789), .A2(new_n790), .A3(new_n703), .A4(new_n738), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n788), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n792), .A2(G330), .ZN(new_n793));
  NAND3_X1  g0593(.A1(new_n759), .A2(new_n764), .A3(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g0595(.A(new_n756), .B1(new_n795), .B2(G1), .ZN(G364));
  AOI21_X1  g0596(.A(new_n215), .B1(G20), .B2(new_n332), .ZN(new_n797));
  INV_X1    g0597(.A(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n207), .A2(G190), .ZN(new_n799));
  NOR2_X1   g0599(.A1(G179), .A2(G200), .ZN(new_n800));
  NAND2_X1  g0600(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g0602(.A1(new_n802), .A2(G159), .ZN(new_n803));
  XNOR2_X1  g0603(.A(new_n803), .B(KEYINPUT32), .ZN(new_n804));
  NOR2_X1   g0604(.A1(new_n207), .A2(new_n436), .ZN(new_n805));
  NOR2_X1   g0605(.A1(new_n315), .A2(G179), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OAI21_X1  g0607(.A(new_n274), .B1(new_n807), .B2(new_n221), .ZN(new_n808));
  NOR2_X1   g0608(.A1(new_n364), .A2(G200), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n799), .A2(new_n809), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n806), .A2(new_n799), .ZN(new_n811));
  OAI22_X1  g0611(.A1(new_n225), .A2(new_n810), .B1(new_n811), .B2(new_n227), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n804), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n207), .B1(new_n800), .B2(G190), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n814), .A2(new_n502), .ZN(new_n815));
  NAND3_X1  g0615(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n816));
  NOR2_X1   g0616(.A1(new_n816), .A2(new_n436), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n818), .A2(new_n202), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n816), .A2(G190), .ZN(new_n820));
  AOI211_X1 g0620(.A(new_n815), .B(new_n819), .C1(G68), .C2(new_n820), .ZN(new_n821));
  AND3_X1   g0621(.A1(new_n805), .A2(KEYINPUT95), .A3(new_n809), .ZN(new_n822));
  AOI21_X1  g0622(.A(KEYINPUT95), .B1(new_n805), .B2(new_n809), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XOR2_X1   g0624(.A(new_n824), .B(KEYINPUT96), .Z(new_n825));
  OAI211_X1 g0625(.A(new_n813), .B(new_n821), .C1(new_n390), .C2(new_n825), .ZN(new_n826));
  INV_X1    g0626(.A(new_n824), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n827), .A2(G322), .ZN(new_n828));
  INV_X1    g0628(.A(G303), .ZN(new_n829));
  INV_X1    g0629(.A(G311), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n807), .A2(new_n829), .B1(new_n810), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g0631(.A(new_n831), .B1(G329), .B2(new_n802), .ZN(new_n832));
  INV_X1    g0632(.A(G283), .ZN(new_n833));
  OAI21_X1  g0633(.A(new_n282), .B1(new_n811), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g0634(.A(KEYINPUT33), .B(G317), .ZN(new_n835));
  AOI21_X1  g0635(.A(new_n834), .B1(new_n820), .B2(new_n835), .ZN(new_n836));
  INV_X1    g0636(.A(new_n814), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n837), .A2(G294), .B1(G326), .B2(new_n817), .ZN(new_n838));
  NAND4_X1  g0638(.A1(new_n828), .A2(new_n832), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n798), .B1(new_n826), .B2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(new_n752), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n337), .A2(G20), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n206), .B1(new_n842), .B2(G45), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n210), .A2(new_n274), .ZN(new_n846));
  INV_X1    g0646(.A(G355), .ZN(new_n847));
  OAI22_X1  g0647(.A1(new_n846), .A2(new_n847), .B1(G116), .B2(new_n210), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n246), .A2(G45), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n210), .A2(new_n282), .ZN(new_n850));
  AOI21_X1  g0650(.A(new_n850), .B1(new_n292), .B2(new_n214), .ZN(new_n851));
  AOI21_X1  g0651(.A(new_n848), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  NOR2_X1   g0652(.A1(G13), .A2(G33), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n854), .A2(G20), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n855), .A2(new_n797), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n845), .B1(new_n852), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g0658(.A1(new_n840), .A2(new_n858), .ZN(new_n859));
  INV_X1    g0659(.A(new_n855), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n859), .B1(new_n743), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n845), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n744), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n743), .A2(G330), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n861), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  XNOR2_X1  g0665(.A(new_n865), .B(KEYINPUT97), .ZN(G396));
  NOR2_X1   g0666(.A1(new_n738), .A2(new_n369), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n867), .A2(KEYINPUT102), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT102), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n738), .B2(new_n369), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n371), .A2(new_n868), .A3(new_n373), .A4(new_n870), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n867), .A2(new_n363), .A3(new_n365), .A4(new_n370), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n873), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n874), .B1(new_n720), .B2(new_n727), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n550), .A2(new_n549), .ZN(new_n876));
  NOR3_X1   g0676(.A1(new_n876), .A2(new_n539), .A3(new_n688), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n710), .B1(new_n683), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g0678(.A1(new_n715), .A2(new_n717), .ZN(new_n879));
  OAI211_X1 g0679(.A(new_n738), .B(new_n873), .C1(new_n878), .C2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n875), .A2(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n845), .B1(new_n881), .B2(new_n793), .ZN(new_n882));
  OAI21_X1  g0682(.A(new_n882), .B1(new_n793), .B2(new_n881), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n797), .A2(new_n853), .ZN(new_n884));
  INV_X1    g0684(.A(new_n884), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n845), .B1(new_n885), .B2(G77), .ZN(new_n886));
  INV_X1    g0686(.A(new_n807), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n274), .B(new_n815), .C1(G107), .C2(new_n887), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n888), .B1(new_n829), .B2(new_n818), .ZN(new_n889));
  OAI22_X1  g0689(.A1(new_n811), .A2(new_n221), .B1(new_n801), .B2(new_n830), .ZN(new_n890));
  XOR2_X1   g0690(.A(new_n890), .B(KEYINPUT99), .Z(new_n891));
  INV_X1    g0691(.A(new_n810), .ZN(new_n892));
  AOI22_X1  g0692(.A1(new_n892), .A2(G116), .B1(G283), .B2(new_n820), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n891), .B1(KEYINPUT98), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g0694(.A(new_n894), .B1(KEYINPUT98), .B2(new_n893), .ZN(new_n895));
  AOI211_X1 g0695(.A(new_n889), .B(new_n895), .C1(G294), .C2(new_n827), .ZN(new_n896));
  XNOR2_X1  g0696(.A(new_n896), .B(KEYINPUT100), .ZN(new_n897));
  AOI22_X1  g0697(.A1(new_n892), .A2(G159), .B1(G137), .B2(new_n817), .ZN(new_n898));
  INV_X1    g0698(.A(new_n820), .ZN(new_n899));
  INV_X1    g0699(.A(G143), .ZN(new_n900));
  OAI221_X1 g0700(.A(new_n898), .B1(new_n255), .B2(new_n899), .C1(new_n825), .C2(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT34), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n282), .B1(new_n887), .B2(G50), .ZN(new_n904));
  INV_X1    g0704(.A(new_n811), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n905), .A2(G68), .ZN(new_n906));
  INV_X1    g0706(.A(G132), .ZN(new_n907));
  OAI211_X1 g0707(.A(new_n904), .B(new_n906), .C1(new_n907), .C2(new_n801), .ZN(new_n908));
  AOI21_X1  g0708(.A(new_n908), .B1(G58), .B2(new_n837), .ZN(new_n909));
  XOR2_X1   g0709(.A(new_n909), .B(KEYINPUT101), .Z(new_n910));
  INV_X1    g0710(.A(new_n901), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(KEYINPUT34), .B2(new_n911), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n897), .B1(new_n903), .B2(new_n912), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n886), .B1(new_n913), .B2(new_n797), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n854), .B2(new_n873), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n883), .A2(new_n915), .ZN(G384));
  OR2_X1    g0716(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n601), .A2(KEYINPUT35), .ZN(new_n918));
  NAND4_X1  g0718(.A1(new_n917), .A2(G116), .A3(new_n216), .A4(new_n918), .ZN(new_n919));
  XOR2_X1   g0719(.A(new_n919), .B(KEYINPUT36), .Z(new_n920));
  OAI211_X1 g0720(.A(new_n214), .B(G77), .C1(new_n390), .C2(new_n219), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n202), .A2(G68), .ZN(new_n922));
  AOI211_X1 g0722(.A(new_n206), .B(G13), .C1(new_n921), .C2(new_n922), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NOR2_X1   g0724(.A1(new_n371), .A2(new_n727), .ZN(new_n925));
  INV_X1    g0725(.A(new_n925), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n880), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n484), .A2(new_n490), .ZN(new_n928));
  INV_X1    g0728(.A(new_n457), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g0730(.A(new_n497), .ZN(new_n931));
  NOR2_X1   g0731(.A1(new_n457), .A2(new_n738), .ZN(new_n932));
  INV_X1    g0732(.A(new_n932), .ZN(new_n933));
  NAND3_X1  g0733(.A1(new_n930), .A2(new_n931), .A3(new_n933), .ZN(new_n934));
  OAI21_X1  g0734(.A(new_n932), .B1(new_n491), .B2(new_n497), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n927), .A2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT38), .ZN(new_n939));
  AOI21_X1  g0739(.A(KEYINPUT16), .B1(new_n389), .B2(new_n409), .ZN(new_n940));
  OAI21_X1  g0740(.A(KEYINPUT103), .B1(new_n940), .B2(new_n317), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT103), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n405), .A2(new_n942), .A3(new_n252), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n941), .A2(new_n414), .A3(new_n943), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n944), .A2(new_n381), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n737), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n443), .B1(KEYINPUT18), .B2(new_n431), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n946), .B1(new_n947), .B2(new_n434), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n408), .A2(new_n417), .A3(new_n737), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT37), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n439), .A2(new_n950), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n411), .A2(new_n414), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n416), .B1(new_n952), .B2(new_n381), .ZN(new_n953));
  AOI211_X1 g0753(.A(KEYINPUT78), .B(new_n380), .C1(new_n411), .C2(new_n414), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n951), .B1(new_n955), .B2(new_n430), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n945), .A2(new_n430), .ZN(new_n957));
  NAND3_X1  g0757(.A1(new_n946), .A2(new_n957), .A3(new_n439), .ZN(new_n958));
  AOI22_X1  g0758(.A1(new_n949), .A2(new_n956), .B1(new_n958), .B2(KEYINPUT37), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n939), .B1(new_n948), .B2(new_n959), .ZN(new_n960));
  INV_X1    g0760(.A(new_n946), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n445), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n958), .A2(KEYINPUT37), .ZN(new_n963));
  INV_X1    g0763(.A(new_n951), .ZN(new_n964));
  NAND3_X1  g0764(.A1(new_n431), .A2(new_n949), .A3(new_n964), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n963), .A2(new_n965), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n962), .A2(KEYINPUT38), .A3(new_n966), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n960), .A2(new_n967), .ZN(new_n968));
  INV_X1    g0768(.A(new_n737), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n938), .A2(new_n968), .B1(new_n697), .B2(new_n969), .ZN(new_n970));
  NOR3_X1   g0770(.A1(new_n953), .A2(new_n954), .A3(new_n969), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n971), .B1(new_n697), .B2(new_n443), .ZN(new_n972));
  AND3_X1   g0772(.A1(new_n431), .A2(new_n949), .A3(new_n964), .ZN(new_n973));
  AND3_X1   g0773(.A1(new_n952), .A2(new_n381), .A3(new_n438), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n429), .B1(new_n952), .B2(new_n381), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  AOI21_X1  g0776(.A(new_n950), .B1(new_n949), .B2(new_n976), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n972), .B1(new_n973), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n978), .A2(new_n939), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n967), .A2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT39), .ZN(new_n981));
  NAND2_X1  g0781(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n930), .A2(new_n727), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n960), .A2(KEYINPUT39), .A3(new_n967), .ZN(new_n984));
  NAND3_X1  g0784(.A1(new_n982), .A2(new_n983), .A3(new_n984), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n970), .A2(new_n985), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n499), .B1(new_n758), .B2(new_n763), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n987), .A2(new_n700), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n986), .B(new_n988), .ZN(new_n989));
  INV_X1    g0789(.A(new_n989), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n439), .B1(new_n415), .B2(new_n429), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n991), .B1(new_n955), .B2(new_n737), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n965), .B1(new_n992), .B2(new_n950), .ZN(new_n993));
  AOI21_X1  g0793(.A(KEYINPUT38), .B1(new_n993), .B2(new_n972), .ZN(new_n994));
  AOI22_X1  g0794(.A1(new_n445), .A2(new_n961), .B1(new_n963), .B2(new_n965), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n994), .B1(KEYINPUT38), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n874), .B1(new_n788), .B2(new_n791), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n997), .A2(new_n936), .ZN(new_n998));
  OAI21_X1  g0798(.A(KEYINPUT40), .B1(new_n996), .B2(new_n998), .ZN(new_n999));
  AOI21_X1  g0799(.A(KEYINPUT40), .B1(new_n960), .B2(new_n967), .ZN(new_n1000));
  AND2_X1   g0800(.A1(new_n997), .A2(new_n936), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  AND2_X1   g0803(.A1(new_n499), .A2(new_n792), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1007));
  INV_X1    g0807(.A(G330), .ZN(new_n1008));
  NOR3_X1   g0808(.A1(new_n1006), .A2(new_n1007), .A3(new_n1008), .ZN(new_n1009));
  OAI22_X1  g0809(.A1(new_n990), .A2(new_n1009), .B1(new_n206), .B2(new_n842), .ZN(new_n1010));
  AND2_X1   g0810(.A1(new_n990), .A2(new_n1009), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n924), .B1(new_n1010), .B2(new_n1011), .ZN(G367));
  NOR2_X1   g0812(.A1(new_n236), .A2(new_n850), .ZN(new_n1013));
  OAI21_X1  g0813(.A(new_n856), .B1(new_n210), .B2(new_n347), .ZN(new_n1014));
  OAI21_X1  g0814(.A(new_n845), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n827), .A2(G150), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n274), .B1(new_n810), .B2(new_n202), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n1017), .B1(G159), .B2(new_n820), .ZN(new_n1018));
  INV_X1    g0818(.A(G137), .ZN(new_n1019));
  OAI22_X1  g0819(.A1(new_n811), .A2(new_n225), .B1(new_n801), .B2(new_n1019), .ZN(new_n1020));
  AOI21_X1  g0820(.A(new_n1020), .B1(G58), .B2(new_n887), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n814), .A2(new_n219), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n1022), .B1(new_n817), .B2(G143), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1016), .A2(new_n1018), .A3(new_n1021), .A4(new_n1023), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n825), .A2(new_n829), .ZN(new_n1025));
  NAND2_X1  g0825(.A1(new_n887), .A2(G116), .ZN(new_n1026));
  XNOR2_X1  g0826(.A(new_n1026), .B(KEYINPUT46), .ZN(new_n1027));
  INV_X1    g0827(.A(G294), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n899), .A2(new_n1028), .B1(new_n814), .B2(new_n227), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(G311), .B2(new_n817), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n274), .B1(new_n905), .B2(G97), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G283), .A2(new_n892), .B1(new_n802), .B2(G317), .ZN(new_n1032));
  NAND4_X1  g0832(.A1(new_n1027), .A2(new_n1030), .A3(new_n1031), .A4(new_n1032), .ZN(new_n1033));
  OAI21_X1  g0833(.A(new_n1024), .B1(new_n1025), .B2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT47), .ZN(new_n1035));
  AOI21_X1  g0835(.A(new_n1015), .B1(new_n1035), .B2(new_n797), .ZN(new_n1036));
  OAI21_X1  g0836(.A(new_n727), .B1(new_n584), .B2(new_n586), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1037), .A2(new_n710), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT104), .Z(new_n1039));
  AND2_X1   g0839(.A1(new_n595), .A2(new_n1037), .ZN(new_n1040));
  OR2_X1    g0840(.A1(new_n1040), .A2(KEYINPUT105), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n1040), .A2(KEYINPUT105), .ZN(new_n1042));
  NAND3_X1  g0842(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1036), .B1(new_n1043), .B2(new_n860), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n706), .B1(new_n680), .B2(new_n738), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n712), .A2(new_n727), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n750), .A2(new_n1048), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1049), .A2(KEYINPUT45), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT45), .ZN(new_n1051));
  NOR3_X1   g0851(.A1(new_n750), .A2(new_n1051), .A3(new_n1048), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n750), .A2(new_n1048), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT44), .ZN(new_n1054));
  NOR2_X1   g0854(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(KEYINPUT44), .B1(new_n750), .B2(new_n1048), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n1050), .A2(new_n1052), .B1(new_n1055), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n745), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n745), .ZN(new_n1059));
  OAI221_X1 g0859(.A(new_n1059), .B1(new_n1055), .B2(new_n1056), .C1(new_n1052), .C2(new_n1050), .ZN(new_n1060));
  INV_X1    g0860(.A(new_n748), .ZN(new_n1061));
  NAND3_X1  g0861(.A1(new_n733), .A2(new_n734), .A3(new_n746), .ZN(new_n1062));
  INV_X1    g0862(.A(KEYINPUT108), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1061), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n748), .A2(KEYINPUT108), .ZN(new_n1065));
  OAI211_X1 g0865(.A(G330), .B(new_n743), .C1(new_n1064), .C2(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n1065), .ZN(new_n1067));
  AND2_X1   g0867(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1068));
  OAI211_X1 g0868(.A(new_n744), .B(new_n1067), .C1(new_n1068), .C2(new_n1061), .ZN(new_n1069));
  AOI21_X1  g0869(.A(new_n794), .B1(new_n1066), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT109), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n1058), .B(new_n1060), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  INV_X1    g0873(.A(new_n1073), .ZN(new_n1074));
  OAI21_X1  g0874(.A(new_n795), .B1(new_n1072), .B2(new_n1074), .ZN(new_n1075));
  XNOR2_X1  g0875(.A(new_n752), .B(KEYINPUT41), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n844), .B1(new_n1075), .B2(new_n1077), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1047), .A2(new_n688), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n727), .B1(new_n1079), .B2(new_n631), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n1061), .A2(KEYINPUT106), .A3(new_n1047), .ZN(new_n1081));
  INV_X1    g0881(.A(KEYINPUT106), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n748), .B2(new_n1048), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1081), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT42), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1081), .A2(KEYINPUT42), .A3(new_n1083), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1080), .B1(new_n1086), .B2(new_n1087), .ZN(new_n1088));
  XNOR2_X1  g0888(.A(new_n1043), .B(KEYINPUT43), .ZN(new_n1089));
  OR2_X1    g0889(.A1(new_n1088), .A2(new_n1089), .ZN(new_n1090));
  NOR2_X1   g0890(.A1(new_n1043), .A2(KEYINPUT43), .ZN(new_n1091));
  AND3_X1   g0891(.A1(new_n1088), .A2(KEYINPUT107), .A3(new_n1091), .ZN(new_n1092));
  AOI21_X1  g0892(.A(KEYINPUT107), .B1(new_n1088), .B2(new_n1091), .ZN(new_n1093));
  OAI21_X1  g0893(.A(new_n1090), .B1(new_n1092), .B2(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n1059), .A2(new_n1048), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1094), .A2(new_n1096), .ZN(new_n1097));
  OAI211_X1 g0897(.A(new_n1095), .B(new_n1090), .C1(new_n1092), .C2(new_n1093), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1044), .B1(new_n1078), .B2(new_n1099), .ZN(G387));
  NAND2_X1  g0900(.A1(new_n1066), .A2(new_n1069), .ZN(new_n1101));
  NAND2_X1  g0901(.A1(new_n736), .A2(new_n855), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n846), .A2(new_n753), .B1(G107), .B2(new_n210), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n241), .A2(new_n292), .ZN(new_n1104));
  INV_X1    g0904(.A(new_n753), .ZN(new_n1105));
  AOI211_X1 g0905(.A(G45), .B(new_n1105), .C1(G68), .C2(G77), .ZN(new_n1106));
  NOR2_X1   g0906(.A1(new_n253), .A2(G50), .ZN(new_n1107));
  XNOR2_X1  g0907(.A(new_n1107), .B(KEYINPUT50), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n850), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1103), .B1(new_n1104), .B2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n845), .B1(new_n1110), .B2(new_n857), .ZN(new_n1111));
  NOR2_X1   g0911(.A1(new_n814), .A2(new_n347), .ZN(new_n1112));
  AOI22_X1  g0912(.A1(G77), .A2(new_n887), .B1(new_n802), .B2(G150), .ZN(new_n1113));
  OAI211_X1 g0913(.A(new_n1113), .B(new_n274), .C1(new_n502), .C2(new_n811), .ZN(new_n1114));
  AOI211_X1 g0914(.A(new_n1112), .B(new_n1114), .C1(G159), .C2(new_n817), .ZN(new_n1115));
  AOI22_X1  g0915(.A1(new_n892), .A2(G68), .B1(new_n319), .B2(new_n820), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(new_n1116), .B(KEYINPUT110), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1115), .B(new_n1117), .C1(new_n202), .C2(new_n824), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n817), .A2(G322), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n892), .A2(G303), .B1(G311), .B2(new_n820), .ZN(new_n1120));
  INV_X1    g0920(.A(G317), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1119), .B(new_n1120), .C1(new_n825), .C2(new_n1121), .ZN(new_n1122));
  INV_X1    g0922(.A(KEYINPUT48), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1124));
  OAI22_X1  g0924(.A1(new_n807), .A2(new_n1028), .B1(new_n814), .B2(new_n833), .ZN(new_n1125));
  AOI21_X1  g0925(.A(new_n1125), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1124), .A2(KEYINPUT49), .A3(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n274), .B1(new_n802), .B2(G326), .ZN(new_n1128));
  OAI211_X1 g0928(.A(new_n1127), .B(new_n1128), .C1(new_n505), .C2(new_n811), .ZN(new_n1129));
  AOI21_X1  g0929(.A(KEYINPUT49), .B1(new_n1124), .B2(new_n1126), .ZN(new_n1130));
  OAI21_X1  g0930(.A(new_n1118), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(KEYINPUT111), .ZN(new_n1132));
  OR2_X1    g0932(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n798), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1134));
  AOI21_X1  g0934(.A(new_n1111), .B1(new_n1133), .B2(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n1101), .A2(new_n844), .B1(new_n1102), .B2(new_n1135), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1101), .A2(new_n795), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1137), .A2(new_n841), .ZN(new_n1138));
  NOR2_X1   g0938(.A1(new_n1101), .A2(new_n795), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1136), .B1(new_n1138), .B2(new_n1139), .ZN(G393));
  NAND2_X1  g0940(.A1(new_n1137), .A2(KEYINPUT109), .ZN(new_n1141));
  NAND4_X1  g0941(.A1(new_n1141), .A2(new_n1073), .A3(new_n1060), .A4(new_n1058), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n752), .B1(new_n1143), .B2(new_n1137), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1142), .A2(new_n1144), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1058), .A2(new_n1060), .A3(new_n844), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n249), .ZN(new_n1147));
  OAI221_X1 g0947(.A(new_n856), .B1(new_n502), .B2(new_n210), .C1(new_n1147), .C2(new_n850), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n1148), .A2(new_n845), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n282), .B1(new_n811), .B2(new_n227), .C1(new_n899), .C2(new_n829), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1150), .B1(G116), .B2(new_n837), .ZN(new_n1151));
  NAND2_X1  g0951(.A1(new_n802), .A2(G322), .ZN(new_n1152));
  AOI22_X1  g0952(.A1(G283), .A2(new_n887), .B1(new_n892), .B2(G294), .ZN(new_n1153));
  AND3_X1   g0953(.A1(new_n1151), .A2(new_n1152), .A3(new_n1153), .ZN(new_n1154));
  OAI22_X1  g0954(.A1(new_n824), .A2(new_n830), .B1(new_n1121), .B2(new_n818), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1155), .B(KEYINPUT52), .ZN(new_n1156));
  INV_X1    g0956(.A(G159), .ZN(new_n1157));
  OAI22_X1  g0957(.A1(new_n824), .A2(new_n1157), .B1(new_n255), .B2(new_n818), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1158), .B(KEYINPUT51), .ZN(new_n1159));
  OAI22_X1  g0959(.A1(new_n807), .A2(new_n219), .B1(new_n810), .B2(new_n253), .ZN(new_n1160));
  AOI21_X1  g0960(.A(new_n282), .B1(new_n905), .B2(G87), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n225), .B2(new_n814), .C1(new_n899), .C2(new_n202), .ZN(new_n1162));
  AOI211_X1 g0962(.A(new_n1160), .B(new_n1162), .C1(G143), .C2(new_n802), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1154), .A2(new_n1156), .B1(new_n1159), .B2(new_n1163), .ZN(new_n1164));
  OAI221_X1 g0964(.A(new_n1149), .B1(new_n798), .B2(new_n1164), .C1(new_n1047), .C2(new_n860), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1145), .A2(new_n1146), .A3(new_n1165), .ZN(G390));
  AND2_X1   g0966(.A1(new_n934), .A2(new_n935), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n785), .A2(new_n727), .ZN(new_n1168));
  INV_X1    g0968(.A(KEYINPUT31), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1168), .A2(new_n1169), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n785), .A2(KEYINPUT31), .A3(new_n727), .ZN(new_n1171));
  NAND2_X1  g0971(.A1(new_n1170), .A2(new_n1171), .ZN(new_n1172));
  NOR4_X1   g0972(.A1(new_n683), .A2(new_n551), .A3(new_n688), .A4(new_n727), .ZN(new_n1173));
  OAI211_X1 g0973(.A(G330), .B(new_n873), .C1(new_n1172), .C2(new_n1173), .ZN(new_n1174));
  NOR2_X1   g0974(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n983), .B1(new_n927), .B2(new_n936), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n982), .B2(new_n984), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n761), .A2(new_n760), .ZN(new_n1178));
  OAI211_X1 g0978(.A(new_n738), .B(new_n873), .C1(new_n878), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n926), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1180), .A2(new_n936), .ZN(new_n1181));
  INV_X1    g0981(.A(new_n983), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1181), .A2(new_n1182), .A3(new_n980), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1183), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1175), .B1(new_n1177), .B2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n937), .A2(new_n1182), .ZN(new_n1186));
  AND3_X1   g0986(.A1(new_n960), .A2(KEYINPUT39), .A3(new_n967), .ZN(new_n1187));
  AOI21_X1  g0987(.A(KEYINPUT39), .B1(new_n967), .B2(new_n979), .ZN(new_n1188));
  OAI21_X1  g0988(.A(new_n1186), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1189));
  NAND3_X1  g0989(.A1(new_n997), .A2(G330), .A3(new_n936), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1189), .A2(new_n1190), .A3(new_n1183), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1008), .B1(new_n788), .B2(new_n791), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n499), .A2(new_n1192), .ZN(new_n1193));
  NAND3_X1  g0993(.A1(new_n987), .A2(new_n700), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n936), .B1(new_n997), .B2(G330), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n927), .B1(new_n1175), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1167), .A2(new_n1174), .ZN(new_n1197));
  NAND4_X1  g0997(.A1(new_n1197), .A2(new_n1190), .A3(new_n926), .A4(new_n1179), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1194), .B1(new_n1196), .B2(new_n1198), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1185), .A2(new_n1191), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(new_n841), .ZN(new_n1201));
  INV_X1    g1001(.A(KEYINPUT112), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1201), .A2(new_n1202), .ZN(new_n1203));
  NAND2_X1  g1003(.A1(new_n1185), .A2(new_n1191), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1199), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1204), .A2(new_n1205), .ZN(new_n1206));
  NAND3_X1  g1006(.A1(new_n1200), .A2(KEYINPUT112), .A3(new_n841), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1203), .A2(new_n1206), .A3(new_n1207), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1204), .A2(new_n843), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n853), .B1(new_n1187), .B2(new_n1188), .ZN(new_n1210));
  OR3_X1    g1010(.A1(new_n807), .A2(KEYINPUT53), .A3(new_n255), .ZN(new_n1211));
  OAI21_X1  g1011(.A(KEYINPUT53), .B1(new_n807), .B2(new_n255), .ZN(new_n1212));
  OAI211_X1 g1012(.A(new_n1211), .B(new_n1212), .C1(new_n1157), .C2(new_n814), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(KEYINPUT54), .B(G143), .ZN(new_n1214));
  INV_X1    g1014(.A(G125), .ZN(new_n1215));
  OAI22_X1  g1015(.A1(new_n810), .A2(new_n1214), .B1(new_n801), .B2(new_n1215), .ZN(new_n1216));
  AOI211_X1 g1016(.A(new_n282), .B(new_n1216), .C1(G50), .C2(new_n905), .ZN(new_n1217));
  INV_X1    g1017(.A(G128), .ZN(new_n1218));
  OAI221_X1 g1018(.A(new_n1217), .B1(new_n1218), .B2(new_n818), .C1(new_n1019), .C2(new_n899), .ZN(new_n1219));
  AOI211_X1 g1019(.A(new_n1213), .B(new_n1219), .C1(G132), .C2(new_n827), .ZN(new_n1220));
  OAI22_X1  g1020(.A1(new_n824), .A2(new_n505), .B1(new_n225), .B2(new_n814), .ZN(new_n1221));
  XOR2_X1   g1021(.A(new_n1221), .B(KEYINPUT114), .Z(new_n1222));
  OAI221_X1 g1022(.A(new_n906), .B1(new_n502), .B2(new_n810), .C1(new_n1028), .C2(new_n801), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n274), .B1(new_n887), .B2(G87), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n899), .B2(new_n227), .C1(new_n833), .C2(new_n818), .ZN(new_n1225));
  NOR3_X1   g1025(.A1(new_n1222), .A2(new_n1223), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n797), .B1(new_n1220), .B2(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n845), .B1(new_n885), .B2(new_n319), .ZN(new_n1228));
  XOR2_X1   g1028(.A(new_n1228), .B(KEYINPUT113), .Z(new_n1229));
  NAND2_X1  g1029(.A1(new_n1227), .A2(new_n1229), .ZN(new_n1230));
  XOR2_X1   g1030(.A(new_n1230), .B(KEYINPUT115), .Z(new_n1231));
  AOI21_X1  g1031(.A(new_n1209), .B1(new_n1210), .B2(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1208), .A2(new_n1232), .ZN(G378));
  INV_X1    g1033(.A(new_n1194), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1200), .A2(new_n1234), .ZN(new_n1235));
  XOR2_X1   g1035(.A(KEYINPUT119), .B(KEYINPUT56), .Z(new_n1236));
  INV_X1    g1036(.A(new_n1236), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n327), .A2(new_n737), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT55), .Z(new_n1239));
  NAND2_X1  g1039(.A1(new_n336), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1240), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n336), .A2(new_n1239), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1237), .B1(new_n1241), .B2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(new_n1242), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1244), .A2(new_n1236), .A3(new_n1240), .ZN(new_n1245));
  AND2_X1   g1045(.A1(new_n1243), .A2(new_n1245), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1246), .ZN(new_n1247));
  AOI21_X1  g1047(.A(new_n1247), .B1(new_n1003), .B2(G330), .ZN(new_n1248));
  AOI211_X1 g1048(.A(new_n1008), .B(new_n1246), .C1(new_n999), .C2(new_n1002), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n986), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1001), .A2(new_n980), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n1251), .A2(KEYINPUT40), .B1(new_n1001), .B2(new_n1000), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1246), .B1(new_n1252), .B2(new_n1008), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n986), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1003), .A2(G330), .A3(new_n1247), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1253), .A2(new_n1254), .A3(new_n1255), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1235), .A2(new_n1250), .A3(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT57), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1257), .A2(new_n1258), .ZN(new_n1259));
  NAND4_X1  g1059(.A1(new_n1235), .A2(new_n1250), .A3(new_n1256), .A4(KEYINPUT57), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n841), .A3(new_n1260), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1250), .A2(new_n1256), .A3(new_n844), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n862), .B1(new_n202), .B2(new_n884), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n905), .A2(G58), .ZN(new_n1264));
  XNOR2_X1  g1064(.A(new_n1264), .B(KEYINPUT116), .ZN(new_n1265));
  OAI22_X1  g1065(.A1(new_n807), .A2(new_n225), .B1(new_n810), .B2(new_n347), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n801), .A2(new_n833), .ZN(new_n1267));
  NAND2_X1  g1067(.A1(new_n282), .A2(new_n291), .ZN(new_n1268));
  NOR4_X1   g1068(.A1(new_n1265), .A2(new_n1266), .A3(new_n1267), .A4(new_n1268), .ZN(new_n1269));
  NOR2_X1   g1069(.A1(new_n818), .A2(new_n505), .ZN(new_n1270));
  AOI211_X1 g1070(.A(new_n1022), .B(new_n1270), .C1(G97), .C2(new_n820), .ZN(new_n1271));
  OAI211_X1 g1071(.A(new_n1269), .B(new_n1271), .C1(new_n227), .C2(new_n824), .ZN(new_n1272));
  XNOR2_X1  g1072(.A(new_n1272), .B(KEYINPUT58), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1268), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1274));
  OAI211_X1 g1074(.A(new_n256), .B(new_n291), .C1(new_n811), .C2(new_n1157), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1275), .B1(G124), .B2(new_n802), .ZN(new_n1276));
  OAI22_X1  g1076(.A1(new_n818), .A2(new_n1215), .B1(new_n807), .B2(new_n1214), .ZN(new_n1277));
  AOI21_X1  g1077(.A(new_n1277), .B1(G150), .B2(new_n837), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1218), .B2(new_n824), .ZN(new_n1279));
  OAI22_X1  g1079(.A1(new_n899), .A2(new_n907), .B1(new_n810), .B2(new_n1019), .ZN(new_n1280));
  XNOR2_X1  g1080(.A(new_n1280), .B(KEYINPUT117), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT59), .ZN(new_n1283));
  OAI21_X1  g1083(.A(new_n1276), .B1(new_n1282), .B2(new_n1283), .ZN(new_n1284));
  INV_X1    g1084(.A(new_n1282), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1285), .A2(KEYINPUT59), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1273), .B(new_n1274), .C1(new_n1284), .C2(new_n1286), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT118), .ZN(new_n1288));
  NOR2_X1   g1088(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1288), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1290), .A2(new_n797), .ZN(new_n1291));
  OAI221_X1 g1091(.A(new_n1263), .B1(new_n1289), .B2(new_n1291), .C1(new_n1246), .C2(new_n854), .ZN(new_n1292));
  XNOR2_X1  g1092(.A(new_n1292), .B(KEYINPUT120), .ZN(new_n1293));
  AND2_X1   g1093(.A1(new_n1262), .A2(new_n1293), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1261), .A2(new_n1294), .ZN(G375));
  NAND2_X1  g1095(.A1(new_n1196), .A2(new_n1198), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1296), .A2(new_n844), .ZN(new_n1297));
  OAI22_X1  g1097(.A1(new_n810), .A2(new_n255), .B1(new_n814), .B2(new_n202), .ZN(new_n1298));
  XNOR2_X1  g1098(.A(new_n1298), .B(KEYINPUT121), .ZN(new_n1299));
  OAI221_X1 g1099(.A(new_n274), .B1(new_n801), .B2(new_n1218), .C1(new_n1157), .C2(new_n807), .ZN(new_n1300));
  NOR3_X1   g1100(.A1(new_n1265), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  XNOR2_X1  g1101(.A(new_n1301), .B(KEYINPUT122), .ZN(new_n1302));
  INV_X1    g1102(.A(new_n1214), .ZN(new_n1303));
  AOI22_X1  g1103(.A1(new_n1303), .A2(new_n820), .B1(G132), .B2(new_n817), .ZN(new_n1304));
  OAI211_X1 g1104(.A(new_n1302), .B(new_n1304), .C1(new_n1019), .C2(new_n825), .ZN(new_n1305));
  AOI211_X1 g1105(.A(new_n274), .B(new_n1112), .C1(G77), .C2(new_n905), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n827), .A2(G283), .ZN(new_n1307));
  AOI22_X1  g1107(.A1(new_n820), .A2(G116), .B1(new_n817), .B2(G294), .ZN(new_n1308));
  OAI22_X1  g1108(.A1(new_n807), .A2(new_n502), .B1(new_n810), .B2(new_n227), .ZN(new_n1309));
  AOI21_X1  g1109(.A(new_n1309), .B1(G303), .B2(new_n802), .ZN(new_n1310));
  NAND4_X1  g1110(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .A4(new_n1310), .ZN(new_n1311));
  AOI21_X1  g1111(.A(new_n798), .B1(new_n1305), .B2(new_n1311), .ZN(new_n1312));
  AOI211_X1 g1112(.A(new_n862), .B(new_n1312), .C1(new_n219), .C2(new_n884), .ZN(new_n1313));
  OAI21_X1  g1113(.A(new_n1313), .B1(new_n854), .B2(new_n936), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1297), .A2(new_n1314), .ZN(new_n1315));
  INV_X1    g1115(.A(new_n1315), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1196), .A2(new_n1194), .A3(new_n1198), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1205), .A2(new_n1077), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1316), .A2(new_n1318), .ZN(G381));
  INV_X1    g1119(.A(G390), .ZN(new_n1320));
  INV_X1    g1120(.A(G384), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(G393), .A2(G396), .ZN(new_n1322));
  NAND3_X1  g1122(.A1(new_n1320), .A2(new_n1321), .A3(new_n1322), .ZN(new_n1323));
  NOR3_X1   g1123(.A1(new_n1323), .A2(G387), .A3(G381), .ZN(new_n1324));
  INV_X1    g1124(.A(G378), .ZN(new_n1325));
  INV_X1    g1125(.A(G375), .ZN(new_n1326));
  NAND3_X1  g1126(.A1(new_n1324), .A2(new_n1325), .A3(new_n1326), .ZN(G407));
  NAND2_X1  g1127(.A1(new_n726), .A2(G213), .ZN(new_n1328));
  INV_X1    g1128(.A(new_n1328), .ZN(new_n1329));
  NAND3_X1  g1129(.A1(new_n1326), .A2(new_n1325), .A3(new_n1329), .ZN(new_n1330));
  XNOR2_X1  g1130(.A(new_n1330), .B(KEYINPUT123), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1331), .A2(G213), .A3(G407), .ZN(G409));
  NAND2_X1  g1132(.A1(G387), .A2(new_n1320), .ZN(new_n1333));
  AND2_X1   g1133(.A1(G393), .A2(G396), .ZN(new_n1334));
  NOR2_X1   g1134(.A1(new_n1334), .A2(new_n1322), .ZN(new_n1335));
  OAI211_X1 g1135(.A(new_n1044), .B(G390), .C1(new_n1078), .C2(new_n1099), .ZN(new_n1336));
  AND3_X1   g1136(.A1(new_n1333), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1337));
  AOI21_X1  g1137(.A(new_n1335), .B1(new_n1333), .B2(new_n1336), .ZN(new_n1338));
  NOR3_X1   g1138(.A1(new_n1337), .A2(new_n1338), .A3(KEYINPUT61), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(new_n1261), .A2(G378), .A3(new_n1294), .ZN(new_n1340));
  OAI211_X1 g1140(.A(new_n1262), .B(new_n1292), .C1(new_n1257), .C2(new_n1076), .ZN(new_n1341));
  NAND3_X1  g1141(.A1(new_n1341), .A2(new_n1208), .A3(new_n1232), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1329), .B1(new_n1340), .B2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(new_n1317), .A2(KEYINPUT124), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT60), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND3_X1  g1146(.A1(new_n1317), .A2(KEYINPUT124), .A3(KEYINPUT60), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1346), .A2(new_n1347), .ZN(new_n1348));
  NAND3_X1  g1148(.A1(new_n1348), .A2(new_n841), .A3(new_n1205), .ZN(new_n1349));
  NAND3_X1  g1149(.A1(new_n1349), .A2(G384), .A3(new_n1316), .ZN(new_n1350));
  INV_X1    g1150(.A(new_n1350), .ZN(new_n1351));
  AOI21_X1  g1151(.A(G384), .B1(new_n1349), .B2(new_n1316), .ZN(new_n1352));
  NOR2_X1   g1152(.A1(new_n1351), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1343), .A2(new_n1353), .ZN(new_n1354));
  XNOR2_X1  g1154(.A(KEYINPUT125), .B(KEYINPUT63), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1329), .A2(G2897), .ZN(new_n1357));
  INV_X1    g1157(.A(new_n1357), .ZN(new_n1358));
  OAI21_X1  g1158(.A(new_n1358), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1359));
  INV_X1    g1159(.A(new_n1352), .ZN(new_n1360));
  NAND3_X1  g1160(.A1(new_n1360), .A2(new_n1350), .A3(new_n1357), .ZN(new_n1361));
  NAND2_X1  g1161(.A1(new_n1359), .A2(new_n1361), .ZN(new_n1362));
  OR2_X1    g1162(.A1(new_n1343), .A2(new_n1362), .ZN(new_n1363));
  NAND3_X1  g1163(.A1(new_n1343), .A2(KEYINPUT63), .A3(new_n1353), .ZN(new_n1364));
  NAND4_X1  g1164(.A1(new_n1339), .A2(new_n1356), .A3(new_n1363), .A4(new_n1364), .ZN(new_n1365));
  INV_X1    g1165(.A(KEYINPUT62), .ZN(new_n1366));
  AND3_X1   g1166(.A1(new_n1343), .A2(new_n1366), .A3(new_n1353), .ZN(new_n1367));
  XOR2_X1   g1167(.A(KEYINPUT126), .B(KEYINPUT61), .Z(new_n1368));
  OAI21_X1  g1168(.A(new_n1368), .B1(new_n1343), .B2(new_n1362), .ZN(new_n1369));
  AOI21_X1  g1169(.A(new_n1366), .B1(new_n1343), .B2(new_n1353), .ZN(new_n1370));
  NOR3_X1   g1170(.A1(new_n1367), .A2(new_n1369), .A3(new_n1370), .ZN(new_n1371));
  NOR2_X1   g1171(.A1(new_n1337), .A2(new_n1338), .ZN(new_n1372));
  OAI21_X1  g1172(.A(new_n1365), .B1(new_n1371), .B2(new_n1372), .ZN(G405));
  OAI21_X1  g1173(.A(KEYINPUT127), .B1(new_n1351), .B2(new_n1352), .ZN(new_n1374));
  INV_X1    g1174(.A(new_n1374), .ZN(new_n1375));
  NOR3_X1   g1175(.A1(new_n1337), .A2(new_n1338), .A3(new_n1375), .ZN(new_n1376));
  AOI21_X1  g1176(.A(new_n1076), .B1(new_n1142), .B2(new_n795), .ZN(new_n1377));
  OAI211_X1 g1177(.A(new_n1097), .B(new_n1098), .C1(new_n1377), .C2(new_n844), .ZN(new_n1378));
  AOI21_X1  g1178(.A(G390), .B1(new_n1378), .B2(new_n1044), .ZN(new_n1379));
  INV_X1    g1179(.A(new_n1336), .ZN(new_n1380));
  OAI22_X1  g1180(.A1(new_n1379), .A2(new_n1380), .B1(new_n1322), .B2(new_n1334), .ZN(new_n1381));
  NAND3_X1  g1181(.A1(new_n1333), .A2(new_n1335), .A3(new_n1336), .ZN(new_n1382));
  AOI21_X1  g1182(.A(new_n1374), .B1(new_n1381), .B2(new_n1382), .ZN(new_n1383));
  INV_X1    g1183(.A(KEYINPUT127), .ZN(new_n1384));
  AOI22_X1  g1184(.A1(new_n1326), .A2(G378), .B1(new_n1353), .B2(new_n1384), .ZN(new_n1385));
  NAND2_X1  g1185(.A1(G375), .A2(new_n1325), .ZN(new_n1386));
  NAND2_X1  g1186(.A1(new_n1385), .A2(new_n1386), .ZN(new_n1387));
  NOR3_X1   g1187(.A1(new_n1376), .A2(new_n1383), .A3(new_n1387), .ZN(new_n1388));
  OAI21_X1  g1188(.A(new_n1375), .B1(new_n1337), .B2(new_n1338), .ZN(new_n1389));
  NAND3_X1  g1189(.A1(new_n1381), .A2(new_n1382), .A3(new_n1374), .ZN(new_n1390));
  AOI22_X1  g1190(.A1(new_n1389), .A2(new_n1390), .B1(new_n1386), .B2(new_n1385), .ZN(new_n1391));
  NOR2_X1   g1191(.A1(new_n1388), .A2(new_n1391), .ZN(G402));
endmodule


