//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 0 0 1 0 1 0 1 1 1 0 1 0 0 0 1 0 0 0 1 1 1 0 0 1 0 1 1 0 1 1 1 0 0 0 1 1 1 0 0 1 1 1 0 1 1 0 0 0 0 0 0 1 0 0 1 0 1 1 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:18 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n785,
    new_n786, new_n787, new_n788, new_n789, new_n790, new_n791, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n801, new_n802, new_n803, new_n804, new_n805, new_n806,
    new_n807, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n874, new_n875, new_n876, new_n877,
    new_n878, new_n879, new_n880, new_n881, new_n882, new_n883, new_n884,
    new_n885, new_n886, new_n887, new_n888, new_n889, new_n890, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n896, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n963, new_n964, new_n965, new_n966, new_n967, new_n968, new_n969,
    new_n970, new_n971, new_n972, new_n973, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1010,
    new_n1011, new_n1012, new_n1013, new_n1014, new_n1015, new_n1016,
    new_n1017, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1037, new_n1038, new_n1039, new_n1040, new_n1041,
    new_n1042, new_n1043, new_n1044, new_n1045, new_n1046, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1095, new_n1096,
    new_n1097, new_n1098, new_n1099, new_n1100, new_n1101, new_n1102,
    new_n1103, new_n1104, new_n1105, new_n1106, new_n1107, new_n1108,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1149, new_n1150, new_n1151,
    new_n1152, new_n1153, new_n1154, new_n1155, new_n1156, new_n1157,
    new_n1158, new_n1159, new_n1160, new_n1161, new_n1162, new_n1163,
    new_n1164, new_n1165, new_n1166, new_n1167, new_n1169, new_n1170,
    new_n1171, new_n1173, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195, new_n1196,
    new_n1197, new_n1198, new_n1199, new_n1200, new_n1201, new_n1202,
    new_n1203, new_n1204, new_n1205, new_n1206, new_n1207, new_n1208,
    new_n1209, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1249, new_n1250, new_n1251,
    new_n1252;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0004(.A1(G1), .A2(G20), .ZN(new_n205));
  XNOR2_X1  g0005(.A(new_n205), .B(KEYINPUT64), .ZN(new_n206));
  AOI22_X1  g0006(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n207));
  XNOR2_X1  g0007(.A(new_n207), .B(KEYINPUT65), .ZN(new_n208));
  AOI22_X1  g0008(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n211));
  NAND3_X1  g0011(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g0012(.A(new_n206), .B1(new_n208), .B2(new_n212), .ZN(new_n213));
  XNOR2_X1  g0013(.A(new_n213), .B(KEYINPUT1), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n206), .A2(G13), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G257), .ZN(new_n218));
  INV_X1    g0018(.A(G264), .ZN(new_n219));
  AOI211_X1 g0019(.A(new_n215), .B(new_n217), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G1), .A2(G13), .ZN(new_n221));
  INV_X1    g0021(.A(G20), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  INV_X1    g0023(.A(new_n223), .ZN(new_n224));
  NAND2_X1  g0024(.A1(new_n202), .A2(G50), .ZN(new_n225));
  OAI22_X1  g0025(.A1(new_n220), .A2(KEYINPUT0), .B1(new_n224), .B2(new_n225), .ZN(new_n226));
  AOI211_X1 g0026(.A(new_n214), .B(new_n226), .C1(KEYINPUT0), .C2(new_n220), .ZN(G361));
  XNOR2_X1  g0027(.A(G238), .B(G244), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(KEYINPUT2), .B(G226), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n229), .B(new_n230), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n232), .B(KEYINPUT66), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n231), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G116), .Z(new_n237));
  XNOR2_X1  g0037(.A(G97), .B(G107), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(G13), .ZN(new_n248));
  NOR3_X1   g0048(.A1(new_n248), .A2(new_n222), .A3(G1), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G50), .ZN(new_n250));
  NAND3_X1  g0050(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(new_n221), .ZN(new_n252));
  INV_X1    g0052(.A(new_n252), .ZN(new_n253));
  OAI21_X1  g0053(.A(new_n253), .B1(G1), .B2(new_n222), .ZN(new_n254));
  AOI21_X1  g0054(.A(new_n250), .B1(new_n254), .B2(G50), .ZN(new_n255));
  XOR2_X1   g0055(.A(new_n255), .B(KEYINPUT69), .Z(new_n256));
  XOR2_X1   g0056(.A(KEYINPUT8), .B(G58), .Z(new_n257));
  INV_X1    g0057(.A(G33), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n258), .A2(G20), .ZN(new_n259));
  NOR2_X1   g0059(.A1(G20), .A2(G33), .ZN(new_n260));
  AOI22_X1  g0060(.A1(new_n257), .A2(new_n259), .B1(G150), .B2(new_n260), .ZN(new_n261));
  AND2_X1   g0061(.A1(new_n261), .A2(KEYINPUT68), .ZN(new_n262));
  OAI21_X1  g0062(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n263), .B1(new_n261), .B2(KEYINPUT68), .ZN(new_n264));
  OAI21_X1  g0064(.A(new_n252), .B1(new_n262), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n256), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(KEYINPUT72), .ZN(new_n267));
  XNOR2_X1  g0067(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(KEYINPUT9), .ZN(new_n269));
  XNOR2_X1  g0069(.A(new_n266), .B(KEYINPUT72), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT9), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT10), .ZN(new_n273));
  NOR2_X1   g0073(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n274));
  INV_X1    g0074(.A(G1), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n275), .B1(G41), .B2(G45), .ZN(new_n276));
  INV_X1    g0076(.A(G274), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT67), .ZN(new_n279));
  AND2_X1   g0079(.A1(new_n276), .A2(new_n279), .ZN(new_n280));
  NOR2_X1   g0080(.A1(new_n276), .A2(new_n279), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n221), .B1(G33), .B2(G41), .ZN(new_n282));
  NOR3_X1   g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n278), .B1(new_n283), .B2(G226), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT3), .B(G33), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(G1698), .ZN(new_n286));
  INV_X1    g0086(.A(G223), .ZN(new_n287));
  INV_X1    g0087(.A(G77), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n286), .A2(new_n287), .B1(new_n288), .B2(new_n285), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n258), .A2(KEYINPUT3), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT3), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n291), .A2(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NOR2_X1   g0093(.A1(new_n293), .A2(G1698), .ZN(new_n294));
  AOI21_X1  g0094(.A(new_n289), .B1(G222), .B2(new_n294), .ZN(new_n295));
  INV_X1    g0095(.A(new_n282), .ZN(new_n296));
  OAI21_X1  g0096(.A(new_n284), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G190), .ZN(new_n298));
  NOR2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  AOI211_X1 g0099(.A(new_n274), .B(new_n299), .C1(G200), .C2(new_n297), .ZN(new_n300));
  NAND3_X1  g0100(.A1(new_n269), .A2(new_n272), .A3(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n273), .A2(KEYINPUT73), .ZN(new_n302));
  INV_X1    g0102(.A(new_n302), .ZN(new_n303));
  OR2_X1    g0103(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(new_n301), .A2(new_n303), .ZN(new_n305));
  INV_X1    g0105(.A(G169), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n266), .B(new_n307), .C1(G179), .C2(new_n297), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n304), .A2(new_n305), .A3(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(G33), .A2(G97), .ZN(new_n310));
  INV_X1    g0110(.A(G232), .ZN(new_n311));
  INV_X1    g0111(.A(G226), .ZN(new_n312));
  INV_X1    g0112(.A(G1698), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n285), .A2(new_n313), .ZN(new_n314));
  OAI221_X1 g0114(.A(new_n310), .B1(new_n286), .B2(new_n311), .C1(new_n312), .C2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(new_n282), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT13), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n278), .B1(new_n283), .B2(G238), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n317), .B1(new_n316), .B2(new_n318), .ZN(new_n321));
  OAI21_X1  g0121(.A(G200), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(new_n321), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n323), .A2(G190), .A3(new_n319), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n249), .A2(new_n242), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n325), .B(KEYINPUT12), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT11), .ZN(new_n327));
  INV_X1    g0127(.A(new_n259), .ZN(new_n328));
  OAI22_X1  g0128(.A1(new_n328), .A2(new_n288), .B1(new_n222), .B2(G68), .ZN(new_n329));
  INV_X1    g0129(.A(new_n260), .ZN(new_n330));
  NOR2_X1   g0130(.A1(new_n330), .A2(new_n240), .ZN(new_n331));
  OAI21_X1  g0131(.A(new_n252), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  OAI221_X1 g0132(.A(new_n326), .B1(new_n242), .B2(new_n254), .C1(new_n327), .C2(new_n332), .ZN(new_n333));
  AND2_X1   g0133(.A1(new_n332), .A2(new_n327), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n322), .A2(new_n324), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT74), .ZN(new_n337));
  XNOR2_X1  g0137(.A(new_n336), .B(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n306), .B1(new_n323), .B2(new_n319), .ZN(new_n339));
  INV_X1    g0139(.A(KEYINPUT14), .ZN(new_n340));
  AND2_X1   g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n323), .A2(G179), .A3(new_n319), .ZN(new_n342));
  OAI21_X1  g0142(.A(new_n342), .B1(new_n339), .B2(new_n340), .ZN(new_n343));
  OAI22_X1  g0143(.A1(new_n341), .A2(new_n343), .B1(new_n334), .B2(new_n333), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n338), .A2(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n293), .A2(G107), .ZN(new_n346));
  INV_X1    g0146(.A(G238), .ZN(new_n347));
  OAI221_X1 g0147(.A(new_n346), .B1(new_n286), .B2(new_n347), .C1(new_n311), .C2(new_n314), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(new_n282), .ZN(new_n349));
  AOI21_X1  g0149(.A(new_n278), .B1(new_n283), .B2(G244), .ZN(new_n350));
  AND2_X1   g0150(.A1(new_n349), .A2(new_n350), .ZN(new_n351));
  INV_X1    g0151(.A(G200), .ZN(new_n352));
  NOR2_X1   g0152(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n353), .B1(G190), .B2(new_n351), .ZN(new_n354));
  INV_X1    g0154(.A(new_n257), .ZN(new_n355));
  OAI22_X1  g0155(.A1(new_n355), .A2(new_n330), .B1(new_n222), .B2(new_n288), .ZN(new_n356));
  XNOR2_X1  g0156(.A(KEYINPUT15), .B(G87), .ZN(new_n357));
  INV_X1    g0157(.A(KEYINPUT70), .ZN(new_n358));
  OR2_X1    g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(new_n358), .ZN(new_n360));
  AND2_X1   g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(new_n259), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT71), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n356), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n364), .B1(new_n363), .B2(new_n362), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n252), .ZN(new_n366));
  INV_X1    g0166(.A(new_n249), .ZN(new_n367));
  MUX2_X1   g0167(.A(new_n367), .B(new_n254), .S(G77), .Z(new_n368));
  NAND3_X1  g0168(.A1(new_n354), .A2(new_n366), .A3(new_n368), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n366), .A2(new_n368), .ZN(new_n370));
  OR2_X1    g0170(.A1(new_n351), .A2(G169), .ZN(new_n371));
  INV_X1    g0171(.A(G179), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n351), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g0173(.A1(new_n370), .A2(new_n371), .A3(new_n373), .ZN(new_n374));
  AND2_X1   g0174(.A1(new_n369), .A2(new_n374), .ZN(new_n375));
  INV_X1    g0175(.A(new_n375), .ZN(new_n376));
  NOR3_X1   g0176(.A1(new_n309), .A2(new_n345), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g0177(.A1(G33), .A2(G87), .ZN(new_n378));
  OAI221_X1 g0178(.A(new_n378), .B1(new_n286), .B2(new_n312), .C1(new_n287), .C2(new_n314), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(new_n282), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n278), .B1(new_n283), .B2(G232), .ZN(new_n381));
  AND2_X1   g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(G179), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n383), .B1(new_n306), .B2(new_n382), .ZN(new_n384));
  NAND2_X1  g0184(.A1(G58), .A2(G68), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n202), .A2(new_n385), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n386), .A2(G20), .B1(G159), .B2(new_n260), .ZN(new_n387));
  AOI21_X1  g0187(.A(KEYINPUT7), .B1(new_n293), .B2(new_n222), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT75), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n242), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT7), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n285), .B2(G20), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n293), .A2(KEYINPUT7), .A3(new_n222), .ZN(new_n393));
  NAND3_X1  g0193(.A1(new_n392), .A2(new_n393), .A3(KEYINPUT75), .ZN(new_n394));
  AND3_X1   g0194(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g0195(.A(KEYINPUT76), .B1(new_n390), .B2(new_n394), .ZN(new_n396));
  OAI211_X1 g0196(.A(KEYINPUT16), .B(new_n387), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT16), .ZN(new_n398));
  AOI21_X1  g0198(.A(new_n242), .B1(new_n392), .B2(new_n393), .ZN(new_n399));
  INV_X1    g0199(.A(new_n387), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n398), .B1(new_n399), .B2(new_n400), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n397), .A2(new_n401), .A3(new_n252), .ZN(new_n402));
  NOR2_X1   g0202(.A1(new_n257), .A2(new_n249), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n403), .B1(new_n254), .B2(new_n257), .ZN(new_n404));
  INV_X1    g0204(.A(new_n404), .ZN(new_n405));
  AND3_X1   g0205(.A1(new_n402), .A2(KEYINPUT77), .A3(new_n405), .ZN(new_n406));
  AOI21_X1  g0206(.A(KEYINPUT77), .B1(new_n402), .B2(new_n405), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n384), .B1(new_n406), .B2(new_n407), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n408), .A2(KEYINPUT18), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT18), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n410), .B(new_n384), .C1(new_n406), .C2(new_n407), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n352), .B1(new_n380), .B2(new_n381), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n412), .B1(G190), .B2(new_n382), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n413), .A2(new_n402), .A3(new_n405), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(KEYINPUT17), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT17), .ZN(new_n416));
  NAND4_X1  g0216(.A1(new_n413), .A2(new_n402), .A3(new_n416), .A4(new_n405), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n415), .A2(new_n417), .ZN(new_n418));
  NAND3_X1  g0218(.A1(new_n409), .A2(new_n411), .A3(new_n418), .ZN(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n377), .A2(new_n420), .ZN(new_n421));
  INV_X1    g0221(.A(KEYINPUT21), .ZN(new_n422));
  XOR2_X1   g0222(.A(KEYINPUT5), .B(G41), .Z(new_n423));
  INV_X1    g0223(.A(G45), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n424), .A2(G1), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(new_n296), .B1(new_n423), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n428), .A2(G270), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n425), .A2(G274), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n423), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(KEYINPUT78), .ZN(new_n432));
  INV_X1    g0232(.A(KEYINPUT78), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n433), .B1(new_n423), .B2(new_n430), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n429), .A2(new_n435), .ZN(new_n436));
  OR3_X1    g0236(.A1(new_n286), .A2(KEYINPUT82), .A3(new_n219), .ZN(new_n437));
  OAI21_X1  g0237(.A(KEYINPUT82), .B1(new_n286), .B2(new_n219), .ZN(new_n438));
  AOI22_X1  g0238(.A1(new_n294), .A2(G257), .B1(G303), .B2(new_n293), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(new_n436), .B1(new_n282), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(G33), .A2(G283), .ZN(new_n442));
  INV_X1    g0242(.A(G97), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n442), .B(new_n222), .C1(G33), .C2(new_n443), .ZN(new_n444));
  OAI211_X1 g0244(.A(new_n444), .B(new_n252), .C1(new_n222), .C2(G116), .ZN(new_n445));
  XNOR2_X1  g0245(.A(new_n445), .B(KEYINPUT20), .ZN(new_n446));
  INV_X1    g0246(.A(G116), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n249), .A2(new_n447), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n367), .B(new_n253), .C1(G1), .C2(new_n258), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n448), .B1(new_n449), .B2(new_n447), .ZN(new_n450));
  OAI21_X1  g0250(.A(G169), .B1(new_n446), .B2(new_n450), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n422), .B1(new_n441), .B2(new_n451), .ZN(new_n452));
  OR2_X1    g0252(.A1(new_n446), .A2(new_n450), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n441), .A2(G179), .A3(new_n453), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n440), .A2(new_n282), .ZN(new_n455));
  AOI22_X1  g0255(.A1(G270), .A2(new_n428), .B1(new_n432), .B2(new_n434), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND4_X1  g0257(.A1(new_n457), .A2(new_n453), .A3(KEYINPUT21), .A4(G169), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n452), .A2(new_n454), .A3(new_n458), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n441), .A2(G190), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n453), .B1(new_n457), .B2(G200), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n459), .B1(new_n460), .B2(new_n461), .ZN(new_n462));
  INV_X1    g0262(.A(new_n434), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n423), .A2(new_n430), .A3(new_n433), .ZN(new_n464));
  OAI22_X1  g0264(.A1(new_n463), .A2(new_n464), .B1(new_n218), .B2(new_n427), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n294), .A2(KEYINPUT4), .A3(G244), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT4), .ZN(new_n467));
  INV_X1    g0267(.A(G244), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n467), .B1(new_n314), .B2(new_n468), .ZN(new_n469));
  NOR2_X1   g0269(.A1(new_n293), .A2(new_n313), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(G250), .ZN(new_n471));
  NAND4_X1  g0271(.A1(new_n466), .A2(new_n469), .A3(new_n442), .A4(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n465), .B1(new_n282), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n473), .A2(new_n372), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(KEYINPUT6), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n238), .A2(new_n476), .ZN(new_n477));
  INV_X1    g0277(.A(G107), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G97), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n477), .B1(new_n476), .B2(new_n479), .ZN(new_n480));
  AOI22_X1  g0280(.A1(new_n480), .A2(G20), .B1(G77), .B2(new_n260), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n392), .A2(new_n393), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n482), .A2(G107), .ZN(new_n483));
  AOI21_X1  g0283(.A(new_n253), .B1(new_n481), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n249), .A2(new_n443), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n485), .B1(new_n449), .B2(new_n443), .ZN(new_n486));
  OAI22_X1  g0286(.A1(new_n473), .A2(G169), .B1(new_n484), .B2(new_n486), .ZN(new_n487));
  OAI21_X1  g0287(.A(KEYINPUT79), .B1(new_n475), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n472), .A2(new_n282), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n428), .A2(G257), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n489), .A2(new_n435), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n491), .A2(new_n306), .ZN(new_n492));
  OR2_X1    g0292(.A1(new_n484), .A2(new_n486), .ZN(new_n493));
  INV_X1    g0293(.A(KEYINPUT79), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n492), .A2(new_n493), .A3(new_n474), .A4(new_n494), .ZN(new_n495));
  AOI21_X1  g0295(.A(new_n493), .B1(G200), .B2(new_n491), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n473), .A2(G190), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n488), .A2(new_n495), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AND2_X1   g0298(.A1(new_n462), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g0299(.A1(G33), .A2(G294), .ZN(new_n500));
  OAI221_X1 g0300(.A(new_n500), .B1(new_n286), .B2(new_n218), .C1(new_n215), .C2(new_n314), .ZN(new_n501));
  NAND3_X1  g0301(.A1(new_n501), .A2(KEYINPUT84), .A3(new_n282), .ZN(new_n502));
  INV_X1    g0302(.A(new_n502), .ZN(new_n503));
  AOI21_X1  g0303(.A(KEYINPUT84), .B1(new_n501), .B2(new_n282), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n428), .A2(G264), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n505), .A2(new_n435), .ZN(new_n506));
  NOR3_X1   g0306(.A1(new_n503), .A2(new_n504), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n501), .A2(new_n282), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n508), .A2(new_n435), .A3(new_n505), .ZN(new_n509));
  OAI22_X1  g0309(.A1(new_n507), .A2(new_n306), .B1(new_n372), .B2(new_n509), .ZN(new_n510));
  INV_X1    g0310(.A(KEYINPUT24), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n285), .A2(new_n222), .A3(G87), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT83), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT83), .ZN(new_n514));
  NAND4_X1  g0314(.A1(new_n285), .A2(new_n514), .A3(new_n222), .A4(G87), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n513), .A2(KEYINPUT22), .A3(new_n515), .ZN(new_n516));
  NOR3_X1   g0316(.A1(new_n222), .A2(KEYINPUT23), .A3(G107), .ZN(new_n517));
  INV_X1    g0317(.A(KEYINPUT23), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n518), .B1(G20), .B2(new_n478), .ZN(new_n519));
  AOI211_X1 g0319(.A(new_n517), .B(new_n519), .C1(G116), .C2(new_n259), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g0321(.A(KEYINPUT22), .B1(new_n513), .B2(new_n515), .ZN(new_n522));
  OAI21_X1  g0322(.A(new_n511), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(new_n522), .ZN(new_n524));
  NAND4_X1  g0324(.A1(new_n524), .A2(KEYINPUT24), .A3(new_n516), .A4(new_n520), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n523), .A2(new_n525), .A3(new_n252), .ZN(new_n526));
  INV_X1    g0326(.A(new_n449), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT25), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n367), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n249), .A2(KEYINPUT25), .A3(new_n478), .ZN(new_n530));
  AOI22_X1  g0330(.A1(new_n527), .A2(G107), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n526), .A2(new_n531), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n510), .A2(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(new_n532), .ZN(new_n535));
  NAND2_X1  g0335(.A1(new_n509), .A2(new_n352), .ZN(new_n536));
  NOR2_X1   g0336(.A1(new_n504), .A2(new_n506), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n537), .A2(new_n502), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n536), .B1(new_n538), .B2(G190), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n534), .B1(new_n535), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n294), .A2(G238), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n285), .A2(G244), .A3(G1698), .ZN(new_n542));
  NAND2_X1  g0342(.A1(G33), .A2(G116), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT80), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n541), .A2(KEYINPUT80), .A3(new_n542), .A4(new_n543), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n282), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n296), .A2(G250), .A3(new_n426), .ZN(new_n550));
  NAND2_X1  g0350(.A1(new_n550), .A2(new_n430), .ZN(new_n551));
  INV_X1    g0351(.A(new_n551), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n549), .A2(new_n372), .A3(new_n552), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(KEYINPUT81), .ZN(new_n554));
  AOI21_X1  g0354(.A(new_n296), .B1(new_n546), .B2(new_n547), .ZN(new_n555));
  NOR2_X1   g0355(.A1(new_n555), .A2(new_n551), .ZN(new_n556));
  INV_X1    g0356(.A(KEYINPUT81), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n556), .A2(new_n557), .A3(new_n372), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n306), .B1(new_n555), .B2(new_n551), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n359), .A2(new_n360), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(new_n249), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT19), .ZN(new_n562));
  OAI21_X1  g0362(.A(new_n562), .B1(new_n328), .B2(new_n443), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n285), .A2(new_n222), .A3(G68), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n222), .B1(new_n310), .B2(new_n562), .ZN(new_n565));
  INV_X1    g0365(.A(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n566), .A2(new_n443), .A3(new_n478), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n563), .A2(new_n564), .A3(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n252), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n561), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n560), .B2(new_n449), .ZN(new_n573));
  NAND4_X1  g0373(.A1(new_n554), .A2(new_n558), .A3(new_n559), .A4(new_n573), .ZN(new_n574));
  NAND3_X1  g0374(.A1(new_n549), .A2(G190), .A3(new_n552), .ZN(new_n575));
  OAI21_X1  g0375(.A(new_n572), .B1(new_n566), .B2(new_n449), .ZN(new_n576));
  INV_X1    g0376(.A(new_n576), .ZN(new_n577));
  OAI211_X1 g0377(.A(new_n575), .B(new_n577), .C1(new_n352), .C2(new_n556), .ZN(new_n578));
  AND2_X1   g0378(.A1(new_n574), .A2(new_n578), .ZN(new_n579));
  AND4_X1   g0379(.A1(new_n421), .A2(new_n499), .A3(new_n540), .A4(new_n579), .ZN(G372));
  NAND4_X1  g0380(.A1(new_n574), .A2(new_n488), .A3(new_n495), .A4(new_n578), .ZN(new_n581));
  NAND2_X1  g0381(.A1(new_n581), .A2(KEYINPUT26), .ZN(new_n582));
  XNOR2_X1  g0382(.A(new_n551), .B(KEYINPUT85), .ZN(new_n583));
  NOR2_X1   g0383(.A1(new_n555), .A2(new_n583), .ZN(new_n584));
  OAI211_X1 g0384(.A(new_n553), .B(new_n573), .C1(new_n584), .C2(G169), .ZN(new_n585));
  OAI211_X1 g0385(.A(new_n575), .B(new_n577), .C1(new_n584), .C2(new_n352), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n475), .A2(new_n487), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OR2_X1    g0388(.A1(new_n588), .A2(KEYINPUT26), .ZN(new_n589));
  AND3_X1   g0389(.A1(new_n452), .A2(new_n458), .A3(new_n454), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n533), .A2(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n584), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(G200), .ZN(new_n593));
  AOI21_X1  g0393(.A(new_n576), .B1(new_n556), .B2(G190), .ZN(new_n594));
  AOI22_X1  g0394(.A1(new_n535), .A2(new_n539), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n591), .A2(new_n498), .A3(new_n595), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n582), .A2(new_n589), .A3(new_n596), .A4(new_n585), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n421), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n374), .A2(KEYINPUT86), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT86), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n370), .A2(new_n600), .A3(new_n371), .A4(new_n373), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n338), .ZN(new_n603));
  AOI22_X1  g0403(.A1(new_n603), .A2(new_n344), .B1(new_n415), .B2(new_n417), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n402), .A2(new_n405), .ZN(new_n605));
  AND2_X1   g0405(.A1(new_n605), .A2(new_n384), .ZN(new_n606));
  AND2_X1   g0406(.A1(new_n606), .A2(KEYINPUT18), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n606), .A2(KEYINPUT18), .ZN(new_n608));
  NOR2_X1   g0408(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  OAI211_X1 g0409(.A(new_n305), .B(new_n304), .C1(new_n604), .C2(new_n609), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n598), .A2(new_n308), .A3(new_n610), .ZN(G369));
  NOR2_X1   g0411(.A1(new_n248), .A2(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n612), .A2(new_n275), .ZN(new_n613));
  OR2_X1    g0413(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n613), .A2(KEYINPUT27), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n614), .A2(G213), .A3(new_n615), .ZN(new_n616));
  XOR2_X1   g0416(.A(KEYINPUT87), .B(G343), .Z(new_n617));
  INV_X1    g0417(.A(new_n617), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n616), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n534), .A2(new_n619), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT88), .ZN(new_n621));
  INV_X1    g0421(.A(new_n619), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n540), .B1(new_n535), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g0423(.A1(new_n621), .A2(new_n623), .ZN(new_n624));
  NOR2_X1   g0424(.A1(new_n590), .A2(new_n619), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n624), .A2(new_n625), .B1(new_n534), .B2(new_n622), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n453), .A2(new_n619), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n462), .A2(new_n627), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n628), .B1(new_n590), .B2(new_n627), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(G330), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n624), .A2(new_n631), .ZN(new_n632));
  NAND2_X1  g0432(.A1(new_n626), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g0433(.A(new_n633), .B(KEYINPUT89), .Z(G399));
  NOR2_X1   g0434(.A1(new_n217), .A2(G41), .ZN(new_n635));
  NOR2_X1   g0435(.A1(new_n567), .A2(G116), .ZN(new_n636));
  INV_X1    g0436(.A(new_n636), .ZN(new_n637));
  NOR3_X1   g0437(.A1(new_n635), .A2(new_n275), .A3(new_n637), .ZN(new_n638));
  INV_X1    g0438(.A(new_n225), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n638), .B1(new_n639), .B2(new_n635), .ZN(new_n640));
  XOR2_X1   g0440(.A(new_n640), .B(KEYINPUT28), .Z(new_n641));
  NAND2_X1  g0441(.A1(new_n597), .A2(new_n622), .ZN(new_n642));
  INV_X1    g0442(.A(new_n642), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n643), .A2(KEYINPUT29), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n596), .A2(new_n585), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n588), .A2(KEYINPUT26), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n646), .B1(new_n581), .B2(KEYINPUT26), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n622), .B1(new_n645), .B2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(KEYINPUT90), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  OAI211_X1 g0450(.A(KEYINPUT90), .B(new_n622), .C1(new_n645), .C2(new_n647), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  AOI21_X1  g0452(.A(new_n644), .B1(KEYINPUT29), .B2(new_n652), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n508), .A2(new_n505), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n491), .A2(new_n654), .ZN(new_n655));
  NAND4_X1  g0455(.A1(new_n655), .A2(G179), .A3(new_n441), .A4(new_n556), .ZN(new_n656));
  INV_X1    g0456(.A(KEYINPUT30), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n473), .A2(G179), .ZN(new_n659));
  NAND4_X1  g0459(.A1(new_n592), .A2(new_n659), .A3(new_n457), .A4(new_n509), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n658), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n656), .A2(new_n657), .ZN(new_n662));
  OAI21_X1  g0462(.A(new_n619), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  NOR2_X1   g0463(.A1(new_n663), .A2(KEYINPUT31), .ZN(new_n664));
  NAND4_X1  g0464(.A1(new_n499), .A2(new_n540), .A3(new_n579), .A4(new_n622), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n663), .A2(KEYINPUT31), .ZN(new_n666));
  AOI21_X1  g0466(.A(new_n664), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  AND2_X1   g0467(.A1(new_n667), .A2(G330), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n653), .A2(new_n668), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n641), .B1(new_n669), .B2(G1), .ZN(G364));
  XNOR2_X1  g0470(.A(new_n612), .B(KEYINPUT91), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n671), .A2(G45), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n672), .A2(G1), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n635), .A2(new_n673), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n631), .A2(new_n674), .ZN(new_n675));
  OAI21_X1  g0475(.A(new_n675), .B1(G330), .B2(new_n629), .ZN(new_n676));
  NOR2_X1   g0476(.A1(new_n217), .A2(new_n293), .ZN(new_n677));
  XOR2_X1   g0477(.A(G355), .B(KEYINPUT92), .Z(new_n678));
  AOI22_X1  g0478(.A1(new_n677), .A2(new_n678), .B1(new_n447), .B2(new_n217), .ZN(new_n679));
  NOR2_X1   g0479(.A1(new_n217), .A2(new_n285), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(G45), .B2(new_n225), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n246), .A2(new_n424), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n679), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g0483(.A(KEYINPUT93), .ZN(new_n684));
  OR2_X1    g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n683), .A2(new_n684), .ZN(new_n686));
  NOR2_X1   g0486(.A1(G13), .A2(G33), .ZN(new_n687));
  INV_X1    g0487(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G20), .ZN(new_n689));
  AOI21_X1  g0489(.A(new_n221), .B1(G20), .B2(new_n306), .ZN(new_n690));
  NOR2_X1   g0490(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n685), .A2(new_n686), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n674), .ZN(new_n693));
  INV_X1    g0493(.A(G58), .ZN(new_n694));
  NAND2_X1  g0494(.A1(G20), .A2(G179), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT94), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n298), .A2(G200), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n697), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(G190), .A2(G200), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  OAI22_X1  g0501(.A1(new_n694), .A2(new_n699), .B1(new_n701), .B2(new_n288), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n298), .A2(new_n352), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n697), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n702), .B1(G50), .B2(new_n705), .ZN(new_n706));
  NOR2_X1   g0506(.A1(new_n222), .A2(G179), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n352), .A2(G190), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n707), .A2(new_n708), .ZN(new_n709));
  OAI21_X1  g0509(.A(new_n285), .B1(new_n709), .B2(new_n478), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n698), .A2(new_n372), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n711), .A2(G20), .ZN(new_n712));
  INV_X1    g0512(.A(new_n712), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n713), .A2(new_n443), .ZN(new_n714));
  NAND2_X1  g0514(.A1(new_n703), .A2(new_n707), .ZN(new_n715));
  INV_X1    g0515(.A(new_n715), .ZN(new_n716));
  AOI211_X1 g0516(.A(new_n710), .B(new_n714), .C1(G87), .C2(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n697), .A2(new_n708), .ZN(new_n718));
  INV_X1    g0518(.A(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT32), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n707), .A2(new_n700), .ZN(new_n721));
  INV_X1    g0521(.A(G159), .ZN(new_n722));
  OAI21_X1  g0522(.A(new_n720), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(new_n721), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n724), .A2(KEYINPUT32), .A3(G159), .ZN(new_n725));
  AOI22_X1  g0525(.A1(new_n719), .A2(G68), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  NAND3_X1  g0526(.A1(new_n706), .A2(new_n717), .A3(new_n726), .ZN(new_n727));
  INV_X1    g0527(.A(G326), .ZN(new_n728));
  INV_X1    g0528(.A(G294), .ZN(new_n729));
  OAI22_X1  g0529(.A1(new_n704), .A2(new_n728), .B1(new_n713), .B2(new_n729), .ZN(new_n730));
  XNOR2_X1  g0530(.A(new_n730), .B(KEYINPUT95), .ZN(new_n731));
  INV_X1    g0531(.A(new_n699), .ZN(new_n732));
  XNOR2_X1  g0532(.A(KEYINPUT33), .B(G317), .ZN(new_n733));
  AOI22_X1  g0533(.A1(G322), .A2(new_n732), .B1(new_n719), .B2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n701), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G311), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n285), .B1(new_n716), .B2(G303), .ZN(new_n737));
  INV_X1    g0537(.A(new_n709), .ZN(new_n738));
  AOI22_X1  g0538(.A1(G283), .A2(new_n738), .B1(new_n724), .B2(G329), .ZN(new_n739));
  NAND4_X1  g0539(.A1(new_n734), .A2(new_n736), .A3(new_n737), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n727), .B1(new_n731), .B2(new_n740), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n693), .B1(new_n741), .B2(new_n690), .ZN(new_n742));
  INV_X1    g0542(.A(new_n689), .ZN(new_n743));
  OAI211_X1 g0543(.A(new_n692), .B(new_n742), .C1(new_n629), .C2(new_n743), .ZN(new_n744));
  AND2_X1   g0544(.A1(new_n676), .A2(new_n744), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(G396));
  NOR2_X1   g0546(.A1(new_n690), .A2(new_n687), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n693), .B1(new_n288), .B2(new_n747), .ZN(new_n748));
  INV_X1    g0548(.A(new_n690), .ZN(new_n749));
  AOI22_X1  g0549(.A1(G116), .A2(new_n735), .B1(new_n719), .B2(G283), .ZN(new_n750));
  INV_X1    g0550(.A(G303), .ZN(new_n751));
  OAI221_X1 g0551(.A(new_n750), .B1(new_n729), .B2(new_n699), .C1(new_n751), .C2(new_n704), .ZN(new_n752));
  OAI21_X1  g0552(.A(new_n293), .B1(new_n715), .B2(new_n478), .ZN(new_n753));
  INV_X1    g0553(.A(G311), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n709), .A2(new_n566), .B1(new_n721), .B2(new_n754), .ZN(new_n755));
  NOR4_X1   g0555(.A1(new_n752), .A2(new_n714), .A3(new_n753), .A4(new_n755), .ZN(new_n756));
  AOI22_X1  g0556(.A1(G137), .A2(new_n705), .B1(new_n732), .B2(G143), .ZN(new_n757));
  INV_X1    g0557(.A(G150), .ZN(new_n758));
  OAI221_X1 g0558(.A(new_n757), .B1(new_n758), .B2(new_n718), .C1(new_n722), .C2(new_n701), .ZN(new_n759));
  INV_X1    g0559(.A(KEYINPUT34), .ZN(new_n760));
  OR2_X1    g0560(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  AOI21_X1  g0561(.A(new_n293), .B1(new_n716), .B2(G50), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n712), .A2(G58), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n724), .A2(G132), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n738), .A2(G68), .ZN(new_n765));
  NAND4_X1  g0565(.A1(new_n762), .A2(new_n763), .A3(new_n764), .A4(new_n765), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n766), .B1(new_n759), .B2(new_n760), .ZN(new_n767));
  AOI21_X1  g0567(.A(new_n756), .B1(new_n761), .B2(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n370), .A2(new_n619), .ZN(new_n769));
  AOI21_X1  g0569(.A(new_n769), .B1(new_n599), .B2(new_n601), .ZN(new_n770));
  AND3_X1   g0570(.A1(new_n369), .A2(new_n374), .A3(new_n769), .ZN(new_n771));
  OR2_X1    g0571(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  OAI221_X1 g0572(.A(new_n748), .B1(new_n749), .B2(new_n768), .C1(new_n772), .C2(new_n688), .ZN(new_n773));
  XNOR2_X1  g0573(.A(new_n642), .B(new_n772), .ZN(new_n774));
  OR3_X1    g0574(.A1(new_n774), .A2(KEYINPUT97), .A3(new_n668), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n774), .A2(new_n668), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n776), .A2(KEYINPUT96), .ZN(new_n777));
  OAI21_X1  g0577(.A(KEYINPUT97), .B1(new_n774), .B2(new_n668), .ZN(new_n778));
  NAND3_X1  g0578(.A1(new_n775), .A2(new_n777), .A3(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n693), .B1(new_n776), .B2(KEYINPUT96), .ZN(new_n780));
  OAI21_X1  g0580(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(G384));
  NOR2_X1   g0581(.A1(new_n671), .A2(new_n275), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n770), .A2(new_n771), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n335), .A2(new_n622), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n345), .A2(new_n784), .ZN(new_n785));
  OAI211_X1 g0585(.A(new_n338), .B(new_n344), .C1(new_n335), .C2(new_n622), .ZN(new_n786));
  AOI21_X1  g0586(.A(new_n783), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n787), .A2(new_n667), .A3(KEYINPUT40), .ZN(new_n788));
  AND2_X1   g0588(.A1(new_n397), .A2(new_n252), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n387), .B1(new_n395), .B2(new_n396), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(new_n398), .ZN(new_n791));
  AOI21_X1  g0591(.A(new_n404), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n792), .A2(new_n616), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n794), .A2(new_n414), .ZN(new_n795));
  INV_X1    g0595(.A(new_n792), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n796), .A2(new_n384), .ZN(new_n797));
  OAI21_X1  g0597(.A(KEYINPUT37), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  INV_X1    g0598(.A(new_n414), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n799), .A2(KEYINPUT37), .ZN(new_n800));
  INV_X1    g0600(.A(new_n616), .ZN(new_n801));
  OAI21_X1  g0601(.A(new_n801), .B1(new_n406), .B2(new_n407), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n800), .A2(new_n408), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g0603(.A1(new_n798), .A2(new_n803), .ZN(new_n804));
  AOI22_X1  g0604(.A1(new_n408), .A2(KEYINPUT18), .B1(new_n415), .B2(new_n417), .ZN(new_n805));
  AOI211_X1 g0605(.A(KEYINPUT99), .B(new_n794), .C1(new_n805), .C2(new_n411), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT99), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n807), .B1(new_n419), .B2(new_n793), .ZN(new_n808));
  OAI211_X1 g0608(.A(KEYINPUT38), .B(new_n804), .C1(new_n806), .C2(new_n808), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n418), .B1(new_n607), .B2(new_n608), .ZN(new_n810));
  INV_X1    g0610(.A(new_n802), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g0612(.A(new_n803), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT37), .ZN(new_n814));
  NOR2_X1   g0614(.A1(new_n606), .A2(new_n799), .ZN(new_n815));
  AOI21_X1  g0615(.A(new_n814), .B1(new_n815), .B2(new_n802), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n812), .B1(new_n813), .B2(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT38), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  AOI21_X1  g0619(.A(new_n788), .B1(new_n809), .B2(new_n819), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n787), .A2(new_n667), .ZN(new_n821));
  INV_X1    g0621(.A(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n419), .A2(new_n793), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(KEYINPUT99), .ZN(new_n824));
  NAND3_X1  g0624(.A1(new_n419), .A2(new_n807), .A3(new_n793), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(KEYINPUT38), .B1(new_n826), .B2(new_n804), .ZN(new_n827));
  INV_X1    g0627(.A(new_n809), .ZN(new_n828));
  OAI21_X1  g0628(.A(new_n822), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(KEYINPUT40), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n820), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g0631(.A1(new_n831), .A2(new_n421), .A3(new_n667), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n809), .A2(new_n819), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n833), .A2(new_n822), .A3(KEYINPUT40), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n804), .B1(new_n806), .B2(new_n808), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n835), .A2(new_n818), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n821), .B1(new_n836), .B2(new_n809), .ZN(new_n837));
  OAI211_X1 g0637(.A(new_n834), .B(G330), .C1(new_n837), .C2(KEYINPUT40), .ZN(new_n838));
  NAND2_X1  g0638(.A1(new_n421), .A2(new_n668), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n832), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n610), .A2(new_n308), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(new_n653), .B2(new_n421), .ZN(new_n843));
  XNOR2_X1  g0643(.A(new_n841), .B(new_n843), .ZN(new_n844));
  NOR2_X1   g0644(.A1(new_n344), .A2(new_n619), .ZN(new_n845));
  INV_X1    g0645(.A(KEYINPUT39), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n846), .B1(new_n836), .B2(new_n809), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n809), .A2(new_n819), .A3(new_n846), .ZN(new_n848));
  INV_X1    g0648(.A(new_n848), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n845), .B1(new_n847), .B2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n772), .A2(new_n597), .A3(new_n622), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n374), .A2(new_n619), .ZN(new_n852));
  INV_X1    g0652(.A(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n851), .A2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n785), .A2(new_n786), .ZN(new_n856));
  INV_X1    g0656(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g0658(.A1(new_n836), .A2(new_n809), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n858), .A2(new_n859), .B1(new_n609), .B2(new_n616), .ZN(new_n860));
  AND2_X1   g0660(.A1(new_n850), .A2(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n782), .B1(new_n844), .B2(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n862), .B1(new_n861), .B2(new_n844), .ZN(new_n863));
  INV_X1    g0663(.A(new_n480), .ZN(new_n864));
  INV_X1    g0664(.A(KEYINPUT35), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n447), .B(new_n224), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  OAI22_X1  g0666(.A1(new_n866), .A2(KEYINPUT98), .B1(new_n865), .B2(new_n864), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n867), .B1(KEYINPUT98), .B2(new_n866), .ZN(new_n868));
  XOR2_X1   g0668(.A(new_n868), .B(KEYINPUT36), .Z(new_n869));
  NAND3_X1  g0669(.A1(new_n639), .A2(G77), .A3(new_n385), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n241), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(G1), .A3(new_n248), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n863), .A2(new_n869), .A3(new_n872), .ZN(G367));
  INV_X1    g0673(.A(new_n680), .ZN(new_n874));
  NOR2_X1   g0674(.A1(new_n235), .A2(new_n874), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n691), .B1(new_n560), .B2(new_n216), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n674), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n751), .A2(new_n699), .B1(new_n704), .B2(new_n754), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n878), .B1(G283), .B2(new_n735), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n716), .A2(KEYINPUT46), .A3(G116), .ZN(new_n880));
  INV_X1    g0680(.A(G317), .ZN(new_n881));
  OAI221_X1 g0681(.A(new_n293), .B1(new_n721), .B2(new_n881), .C1(new_n443), .C2(new_n709), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n882), .B1(new_n719), .B2(G294), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT46), .B1(new_n716), .B2(G116), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n884), .B1(G107), .B2(new_n712), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n879), .A2(new_n880), .A3(new_n883), .A4(new_n885), .ZN(new_n886));
  NOR2_X1   g0686(.A1(new_n713), .A2(new_n242), .ZN(new_n887));
  AOI211_X1 g0687(.A(new_n293), .B(new_n887), .C1(G77), .C2(new_n738), .ZN(new_n888));
  AOI22_X1  g0688(.A1(G58), .A2(new_n716), .B1(new_n724), .B2(G137), .ZN(new_n889));
  AOI22_X1  g0689(.A1(new_n705), .A2(G143), .B1(new_n889), .B2(KEYINPUT107), .ZN(new_n890));
  OAI211_X1 g0690(.A(new_n888), .B(new_n890), .C1(new_n758), .C2(new_n699), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n719), .A2(G159), .ZN(new_n892));
  OAI221_X1 g0692(.A(new_n892), .B1(KEYINPUT107), .B2(new_n889), .C1(new_n240), .C2(new_n701), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n886), .B1(new_n891), .B2(new_n893), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT47), .ZN(new_n895));
  OR2_X1    g0695(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n749), .B1(new_n894), .B2(new_n895), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n877), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g0698(.A1(new_n576), .A2(new_n619), .ZN(new_n899));
  NAND3_X1  g0699(.A1(new_n585), .A2(new_n586), .A3(new_n899), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n585), .B2(new_n899), .ZN(new_n901));
  OAI21_X1  g0701(.A(new_n898), .B1(new_n901), .B2(new_n743), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n624), .A2(new_n625), .ZN(new_n903));
  INV_X1    g0703(.A(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n493), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n498), .B1(new_n905), .B2(new_n622), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n587), .A2(new_n619), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n904), .A2(new_n908), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT100), .ZN(new_n910));
  OR3_X1    g0710(.A1(new_n909), .A2(new_n910), .A3(KEYINPUT42), .ZN(new_n911));
  OAI21_X1  g0711(.A(new_n910), .B1(new_n909), .B2(KEYINPUT42), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n908), .A2(new_n534), .B1(new_n488), .B2(new_n495), .ZN(new_n913));
  OR2_X1    g0713(.A1(new_n913), .A2(new_n619), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n909), .A2(KEYINPUT42), .ZN(new_n915));
  NAND4_X1  g0715(.A1(new_n911), .A2(new_n912), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  NAND2_X1  g0716(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g0718(.A1(new_n901), .A2(KEYINPUT43), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n920), .ZN(new_n921));
  NOR3_X1   g0721(.A1(new_n916), .A2(KEYINPUT43), .A3(new_n901), .ZN(new_n922));
  INV_X1    g0722(.A(new_n922), .ZN(new_n923));
  INV_X1    g0723(.A(new_n632), .ZN(new_n924));
  AOI22_X1  g0724(.A1(new_n921), .A2(new_n923), .B1(new_n924), .B2(new_n908), .ZN(new_n925));
  INV_X1    g0725(.A(new_n908), .ZN(new_n926));
  NOR4_X1   g0726(.A1(new_n920), .A2(new_n922), .A3(new_n632), .A4(new_n926), .ZN(new_n927));
  OR2_X1    g0727(.A1(new_n925), .A2(new_n927), .ZN(new_n928));
  OR2_X1    g0728(.A1(new_n624), .A2(new_n625), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n929), .A2(KEYINPUT106), .A3(new_n630), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n630), .B1(new_n929), .B2(KEYINPUT106), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n903), .B1(new_n931), .B2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n932), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n934), .A2(new_n904), .A3(new_n930), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n933), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n936), .A2(new_n669), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT103), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n926), .B1(new_n939), .B2(KEYINPUT44), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(KEYINPUT44), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n941), .B(KEYINPUT104), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  OR3_X1    g0743(.A1(new_n626), .A2(new_n940), .A3(new_n943), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n943), .B1(new_n626), .B2(new_n940), .ZN(new_n945));
  XNOR2_X1  g0745(.A(KEYINPUT102), .B(KEYINPUT45), .ZN(new_n946));
  INV_X1    g0746(.A(new_n946), .ZN(new_n947));
  AND3_X1   g0747(.A1(new_n626), .A2(new_n908), .A3(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n947), .B1(new_n626), .B2(new_n908), .ZN(new_n949));
  OAI211_X1 g0749(.A(new_n944), .B(new_n945), .C1(new_n948), .C2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n950), .A2(new_n924), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n938), .B1(KEYINPUT105), .B2(new_n952), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT105), .ZN(new_n954));
  NOR2_X1   g0754(.A1(new_n950), .A2(new_n924), .ZN(new_n955));
  INV_X1    g0755(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g0756(.A(new_n954), .B1(new_n956), .B2(new_n951), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n669), .B1(new_n953), .B2(new_n957), .ZN(new_n958));
  XNOR2_X1  g0758(.A(KEYINPUT101), .B(KEYINPUT41), .ZN(new_n959));
  XNOR2_X1  g0759(.A(new_n635), .B(new_n959), .ZN(new_n960));
  AOI21_X1  g0760(.A(new_n673), .B1(new_n958), .B2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n902), .B1(new_n928), .B2(new_n961), .ZN(G387));
  NAND2_X1  g0762(.A1(new_n936), .A2(new_n673), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G303), .A2(new_n735), .B1(new_n719), .B2(G311), .ZN(new_n964));
  INV_X1    g0764(.A(G322), .ZN(new_n965));
  OAI221_X1 g0765(.A(new_n964), .B1(new_n881), .B2(new_n699), .C1(new_n965), .C2(new_n704), .ZN(new_n966));
  XNOR2_X1  g0766(.A(new_n966), .B(KEYINPUT48), .ZN(new_n967));
  INV_X1    g0767(.A(G283), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n967), .B1(new_n968), .B2(new_n713), .C1(new_n729), .C2(new_n715), .ZN(new_n969));
  XOR2_X1   g0769(.A(new_n969), .B(KEYINPUT49), .Z(new_n970));
  OAI221_X1 g0770(.A(new_n293), .B1(new_n721), .B2(new_n728), .C1(new_n447), .C2(new_n709), .ZN(new_n971));
  XNOR2_X1  g0771(.A(new_n971), .B(KEYINPUT109), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  AOI22_X1  g0773(.A1(G77), .A2(new_n716), .B1(new_n724), .B2(G150), .ZN(new_n974));
  OAI211_X1 g0774(.A(new_n974), .B(new_n285), .C1(new_n443), .C2(new_n709), .ZN(new_n975));
  AOI22_X1  g0775(.A1(G159), .A2(new_n705), .B1(new_n719), .B2(new_n257), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n361), .A2(new_n712), .ZN(new_n977));
  OAI211_X1 g0777(.A(new_n976), .B(new_n977), .C1(new_n240), .C2(new_n699), .ZN(new_n978));
  AOI211_X1 g0778(.A(new_n975), .B(new_n978), .C1(G68), .C2(new_n735), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n690), .B1(new_n973), .B2(new_n979), .ZN(new_n980));
  AOI211_X1 g0780(.A(G45), .B(new_n637), .C1(G68), .C2(G77), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n982), .A2(KEYINPUT108), .ZN(new_n983));
  OAI21_X1  g0783(.A(KEYINPUT50), .B1(new_n355), .B2(G50), .ZN(new_n984));
  OR3_X1    g0784(.A1(new_n355), .A2(KEYINPUT50), .A3(G50), .ZN(new_n985));
  INV_X1    g0785(.A(KEYINPUT108), .ZN(new_n986));
  OAI211_X1 g0786(.A(new_n984), .B(new_n985), .C1(new_n981), .C2(new_n986), .ZN(new_n987));
  OAI221_X1 g0787(.A(new_n680), .B1(new_n424), .B2(new_n231), .C1(new_n983), .C2(new_n987), .ZN(new_n988));
  AOI22_X1  g0788(.A1(new_n677), .A2(new_n637), .B1(new_n478), .B2(new_n217), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n988), .A2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n693), .B1(new_n990), .B2(new_n691), .ZN(new_n991));
  OAI211_X1 g0791(.A(new_n980), .B(new_n991), .C1(new_n624), .C2(new_n743), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n937), .A2(new_n635), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n936), .A2(new_n669), .ZN(new_n994));
  OAI211_X1 g0794(.A(new_n963), .B(new_n992), .C1(new_n993), .C2(new_n994), .ZN(G393));
  INV_X1    g0795(.A(KEYINPUT113), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n937), .B1(new_n954), .B2(new_n951), .ZN(new_n997));
  NOR2_X1   g0797(.A1(new_n952), .A2(new_n955), .ZN(new_n998));
  OAI21_X1  g0798(.A(new_n997), .B1(new_n998), .B2(new_n954), .ZN(new_n999));
  INV_X1    g0799(.A(new_n635), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n956), .A2(new_n951), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n1000), .B1(new_n1001), .B2(new_n937), .ZN(new_n1002));
  AND2_X1   g0802(.A1(new_n999), .A2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT110), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n1001), .A2(new_n1004), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n998), .A2(KEYINPUT110), .ZN(new_n1006));
  NAND3_X1  g0806(.A1(new_n1005), .A2(new_n1006), .A3(new_n673), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n691), .B1(new_n216), .B2(new_n443), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n239), .ZN(new_n1009));
  AOI21_X1  g0809(.A(new_n1008), .B1(new_n680), .B2(new_n1009), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n693), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n712), .A2(G77), .ZN(new_n1012));
  OAI221_X1 g0812(.A(new_n1012), .B1(new_n701), .B2(new_n355), .C1(new_n240), .C2(new_n718), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT112), .Z(new_n1014));
  AOI22_X1  g0814(.A1(G68), .A2(new_n716), .B1(new_n724), .B2(G143), .ZN(new_n1015));
  OAI211_X1 g0815(.A(new_n1015), .B(new_n285), .C1(new_n566), .C2(new_n709), .ZN(new_n1016));
  XNOR2_X1  g0816(.A(new_n1016), .B(KEYINPUT111), .ZN(new_n1017));
  OAI22_X1  g0817(.A1(new_n758), .A2(new_n704), .B1(new_n699), .B2(new_n722), .ZN(new_n1018));
  XNOR2_X1  g0818(.A(new_n1018), .B(KEYINPUT51), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n1017), .A2(new_n1019), .ZN(new_n1020));
  AOI22_X1  g0820(.A1(G311), .A2(new_n732), .B1(new_n705), .B2(G317), .ZN(new_n1021));
  NOR2_X1   g0821(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n1021), .A2(KEYINPUT52), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n293), .B1(new_n709), .B2(new_n478), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n715), .A2(new_n968), .B1(new_n721), .B2(new_n965), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n1024), .B(new_n1025), .C1(G116), .C2(new_n712), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(G294), .A2(new_n735), .B1(new_n719), .B2(G303), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1023), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  OAI22_X1  g0828(.A1(new_n1014), .A2(new_n1020), .B1(new_n1022), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g0829(.A(new_n1029), .ZN(new_n1030));
  OAI221_X1 g0830(.A(new_n1011), .B1(new_n749), .B2(new_n1030), .C1(new_n908), .C2(new_n743), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1007), .A2(new_n1031), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n996), .B1(new_n1003), .B2(new_n1032), .ZN(new_n1033));
  OAI221_X1 g0833(.A(new_n635), .B1(new_n998), .B2(new_n938), .C1(new_n953), .C2(new_n957), .ZN(new_n1034));
  NAND4_X1  g0834(.A1(new_n1034), .A2(KEYINPUT113), .A3(new_n1031), .A4(new_n1007), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1033), .A2(new_n1035), .ZN(G390));
  NAND4_X1  g0836(.A1(new_n667), .A2(G330), .A3(new_n772), .A4(new_n856), .ZN(new_n1037));
  INV_X1    g0837(.A(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(KEYINPUT114), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1037), .A2(KEYINPUT114), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n845), .B1(new_n854), .B2(new_n856), .ZN(new_n1042));
  NOR3_X1   g0842(.A1(new_n847), .A2(new_n849), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n783), .B1(new_n650), .B2(new_n651), .ZN(new_n1044));
  OAI21_X1  g0844(.A(new_n856), .B1(new_n1044), .B2(new_n852), .ZN(new_n1045));
  INV_X1    g0845(.A(new_n845), .ZN(new_n1046));
  AND3_X1   g0846(.A1(new_n1045), .A2(new_n1046), .A3(new_n833), .ZN(new_n1047));
  OAI211_X1 g0847(.A(new_n1040), .B(new_n1041), .C1(new_n1043), .C2(new_n1047), .ZN(new_n1048));
  INV_X1    g0848(.A(new_n1042), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n859), .ZN(new_n1050));
  OAI211_X1 g0850(.A(new_n848), .B(new_n1049), .C1(new_n1050), .C2(new_n846), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1045), .A2(new_n1046), .A3(new_n833), .ZN(new_n1052));
  NAND4_X1  g0852(.A1(new_n1051), .A2(new_n1039), .A3(new_n1038), .A4(new_n1052), .ZN(new_n1053));
  NAND2_X1  g0853(.A1(new_n1048), .A2(new_n1053), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n667), .A2(G330), .A3(new_n772), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1055), .A2(new_n857), .ZN(new_n1056));
  NAND2_X1  g0856(.A1(new_n1056), .A2(new_n1037), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n854), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1044), .A2(new_n852), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n1058), .B1(new_n1059), .B2(new_n1057), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n1060), .A2(new_n843), .A3(new_n839), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NAND2_X1  g0862(.A1(new_n1054), .A2(new_n1062), .ZN(new_n1063));
  NAND3_X1  g0863(.A1(new_n1048), .A2(new_n1061), .A3(new_n1053), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n1063), .A2(new_n635), .A3(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n747), .ZN(new_n1066));
  OAI21_X1  g0866(.A(new_n674), .B1(new_n257), .B2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n765), .B1(new_n729), .B2(new_n721), .ZN(new_n1068));
  AOI211_X1 g0868(.A(new_n285), .B(new_n1068), .C1(G87), .C2(new_n716), .ZN(new_n1069));
  AOI22_X1  g0869(.A1(G97), .A2(new_n735), .B1(new_n732), .B2(G116), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(G107), .A2(new_n719), .B1(new_n705), .B2(G283), .ZN(new_n1071));
  NAND4_X1  g0871(.A1(new_n1069), .A2(new_n1012), .A3(new_n1070), .A4(new_n1071), .ZN(new_n1072));
  NOR2_X1   g0872(.A1(new_n715), .A2(new_n758), .ZN(new_n1073));
  XNOR2_X1  g0873(.A(new_n1073), .B(KEYINPUT117), .ZN(new_n1074));
  AND2_X1   g0874(.A1(new_n1074), .A2(KEYINPUT53), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(KEYINPUT53), .ZN(new_n1076));
  AOI21_X1  g0876(.A(new_n293), .B1(new_n724), .B2(G125), .ZN(new_n1077));
  OAI221_X1 g0877(.A(new_n1077), .B1(new_n240), .B2(new_n709), .C1(new_n722), .C2(new_n713), .ZN(new_n1078));
  OR3_X1    g0878(.A1(new_n1075), .A2(new_n1076), .A3(new_n1078), .ZN(new_n1079));
  AOI22_X1  g0879(.A1(G128), .A2(new_n705), .B1(new_n732), .B2(G132), .ZN(new_n1080));
  INV_X1    g0880(.A(G137), .ZN(new_n1081));
  XNOR2_X1  g0881(.A(KEYINPUT54), .B(G143), .ZN(new_n1082));
  XOR2_X1   g0882(.A(new_n1082), .B(KEYINPUT116), .Z(new_n1083));
  INV_X1    g0883(.A(new_n1083), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n1080), .B1(new_n1081), .B2(new_n718), .C1(new_n701), .C2(new_n1084), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n1072), .B1(new_n1079), .B2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1067), .B1(new_n1086), .B2(new_n690), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n848), .B1(new_n1050), .B2(new_n846), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n1087), .B1(new_n1088), .B2(new_n688), .ZN(new_n1089));
  AOI21_X1  g0889(.A(KEYINPUT115), .B1(new_n1054), .B2(new_n673), .ZN(new_n1090));
  INV_X1    g0890(.A(KEYINPUT115), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n673), .ZN(new_n1092));
  AOI211_X1 g0892(.A(new_n1091), .B(new_n1092), .C1(new_n1048), .C2(new_n1053), .ZN(new_n1093));
  OAI211_X1 g0893(.A(new_n1065), .B(new_n1089), .C1(new_n1090), .C2(new_n1093), .ZN(G378));
  AOI21_X1  g0894(.A(new_n1061), .B1(new_n1048), .B2(new_n1053), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n843), .A2(new_n839), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n268), .A2(new_n616), .ZN(new_n1097));
  OR2_X1    g0897(.A1(new_n309), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n309), .A2(new_n1097), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n1101), .ZN(new_n1102));
  NAND2_X1  g0902(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1103));
  NAND3_X1  g0903(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n1105), .B1(new_n831), .B2(G330), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n838), .A2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n850), .A2(new_n860), .ZN(new_n1109));
  NOR3_X1   g0909(.A1(new_n1106), .A2(new_n1108), .A3(new_n1109), .ZN(new_n1110));
  NAND3_X1  g0910(.A1(new_n831), .A2(G330), .A3(new_n1105), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n838), .A2(new_n1107), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n861), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI22_X1  g0913(.A1(new_n1095), .A2(new_n1096), .B1(new_n1110), .B2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(KEYINPUT57), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n635), .B1(new_n1114), .B2(new_n1115), .ZN(new_n1116));
  INV_X1    g0916(.A(new_n1096), .ZN(new_n1117));
  NAND2_X1  g0917(.A1(new_n1063), .A2(new_n1117), .ZN(new_n1118));
  OAI21_X1  g0918(.A(new_n1109), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n861), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1119), .A2(new_n1120), .ZN(new_n1121));
  AOI21_X1  g0921(.A(KEYINPUT57), .B1(new_n1118), .B2(new_n1121), .ZN(new_n1122));
  OR2_X1    g0922(.A1(new_n1116), .A2(new_n1122), .ZN(new_n1123));
  AOI22_X1  g0923(.A1(G97), .A2(new_n719), .B1(new_n705), .B2(G116), .ZN(new_n1124));
  OAI221_X1 g0924(.A(new_n1124), .B1(new_n478), .B2(new_n699), .C1(new_n560), .C2(new_n701), .ZN(new_n1125));
  INV_X1    g0925(.A(G41), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1126), .B(new_n293), .C1(new_n715), .C2(new_n288), .ZN(new_n1127));
  OAI22_X1  g0927(.A1(new_n709), .A2(new_n694), .B1(new_n721), .B2(new_n968), .ZN(new_n1128));
  NOR4_X1   g0928(.A1(new_n1125), .A2(new_n887), .A3(new_n1127), .A4(new_n1128), .ZN(new_n1129));
  OR2_X1    g0929(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n1129), .A2(KEYINPUT58), .ZN(new_n1131));
  AOI21_X1  g0931(.A(G50), .B1(new_n258), .B2(new_n1126), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1132), .B1(new_n285), .B2(G41), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1130), .A2(new_n1131), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(G128), .A2(new_n732), .B1(new_n735), .B2(G137), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n719), .A2(G132), .B1(G150), .B2(new_n712), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1083), .A2(new_n716), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n705), .A2(G125), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1135), .A2(new_n1136), .A3(new_n1137), .A4(new_n1138), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(new_n1139), .B(KEYINPUT59), .ZN(new_n1140));
  AOI211_X1 g0940(.A(G33), .B(G41), .C1(new_n724), .C2(G124), .ZN(new_n1141));
  OAI21_X1  g0941(.A(new_n1141), .B1(new_n722), .B2(new_n709), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1140), .A2(new_n1142), .ZN(new_n1143));
  OAI21_X1  g0943(.A(new_n690), .B1(new_n1134), .B2(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(new_n1144), .B(new_n674), .C1(G50), .C2(new_n1066), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n1107), .B2(new_n687), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1146), .B1(new_n1121), .B2(new_n673), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n1123), .A2(new_n1147), .ZN(G375));
  NAND2_X1  g0948(.A1(new_n857), .A2(new_n687), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n674), .B1(G68), .B2(new_n1066), .ZN(new_n1150));
  XNOR2_X1  g0950(.A(new_n1150), .B(KEYINPUT119), .ZN(new_n1151));
  AOI22_X1  g0951(.A1(G159), .A2(new_n716), .B1(new_n724), .B2(G128), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n293), .B1(new_n738), .B2(G58), .ZN(new_n1153));
  OAI211_X1 g0953(.A(new_n1152), .B(new_n1153), .C1(new_n240), .C2(new_n713), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(G132), .A2(new_n705), .B1(new_n735), .B2(G150), .ZN(new_n1155));
  OAI221_X1 g0955(.A(new_n1155), .B1(new_n1081), .B2(new_n699), .C1(new_n718), .C2(new_n1084), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(G107), .A2(new_n735), .B1(new_n719), .B2(G116), .ZN(new_n1157));
  OAI221_X1 g0957(.A(new_n1157), .B1(new_n968), .B2(new_n699), .C1(new_n729), .C2(new_n704), .ZN(new_n1158));
  AOI21_X1  g0958(.A(new_n285), .B1(new_n738), .B2(G77), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(G97), .A2(new_n716), .B1(new_n724), .B2(G303), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n977), .A2(new_n1159), .A3(new_n1160), .ZN(new_n1161));
  OAI22_X1  g0961(.A1(new_n1154), .A2(new_n1156), .B1(new_n1158), .B2(new_n1161), .ZN(new_n1162));
  AOI21_X1  g0962(.A(new_n1151), .B1(new_n1162), .B2(new_n690), .ZN(new_n1163));
  AOI22_X1  g0963(.A1(new_n1060), .A2(new_n673), .B1(new_n1149), .B2(new_n1163), .ZN(new_n1164));
  XOR2_X1   g0964(.A(new_n960), .B(KEYINPUT118), .Z(new_n1165));
  NAND2_X1  g0965(.A1(new_n1061), .A2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n1117), .A2(new_n1060), .ZN(new_n1167));
  OAI21_X1  g0967(.A(new_n1164), .B1(new_n1166), .B2(new_n1167), .ZN(G381));
  NOR2_X1   g0968(.A1(G375), .A2(G378), .ZN(new_n1169));
  NOR2_X1   g0969(.A1(G390), .A2(G387), .ZN(new_n1170));
  NOR4_X1   g0970(.A1(G393), .A2(G381), .A3(G396), .A4(G384), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1169), .A2(new_n1170), .A3(new_n1171), .ZN(G407));
  NAND2_X1  g0972(.A1(new_n1169), .A2(new_n618), .ZN(new_n1173));
  NAND3_X1  g0973(.A1(G407), .A2(G213), .A3(new_n1173), .ZN(G409));
  OAI211_X1 g0974(.A(new_n1121), .B(new_n1165), .C1(new_n1096), .C2(new_n1095), .ZN(new_n1175));
  AND2_X1   g0975(.A1(new_n1175), .A2(new_n1147), .ZN(new_n1176));
  OAI21_X1  g0976(.A(KEYINPUT120), .B1(new_n1176), .B2(G378), .ZN(new_n1177));
  OAI211_X1 g0977(.A(G378), .B(new_n1147), .C1(new_n1116), .C2(new_n1122), .ZN(new_n1178));
  AND2_X1   g0978(.A1(new_n1065), .A2(new_n1089), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1175), .A2(new_n1147), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT120), .ZN(new_n1181));
  OR2_X1    g0981(.A1(new_n1090), .A2(new_n1093), .ZN(new_n1182));
  NAND4_X1  g0982(.A1(new_n1179), .A2(new_n1180), .A3(new_n1181), .A4(new_n1182), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1177), .A2(new_n1178), .A3(new_n1183), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1167), .A2(KEYINPUT60), .ZN(new_n1185));
  INV_X1    g0985(.A(KEYINPUT60), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n1117), .B2(new_n1060), .ZN(new_n1187));
  NAND4_X1  g0987(.A1(new_n1185), .A2(new_n635), .A3(new_n1061), .A4(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT121), .ZN(new_n1189));
  OR2_X1    g0989(.A1(G384), .A2(new_n1189), .ZN(new_n1190));
  INV_X1    g0990(.A(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1188), .A2(new_n1164), .A3(new_n1191), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(G384), .B(new_n1189), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(new_n1188), .B2(new_n1164), .ZN(new_n1195));
  OAI21_X1  g0995(.A(KEYINPUT122), .B1(new_n1193), .B2(new_n1195), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT122), .ZN(new_n1197));
  AND2_X1   g0997(.A1(new_n1188), .A2(new_n1164), .ZN(new_n1198));
  OAI211_X1 g0998(.A(new_n1197), .B(new_n1192), .C1(new_n1198), .C2(new_n1194), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1196), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n618), .A2(G213), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1184), .A2(new_n1200), .A3(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1202), .A2(KEYINPUT124), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT125), .ZN(new_n1204));
  INV_X1    g1004(.A(KEYINPUT62), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1203), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  INV_X1    g1006(.A(KEYINPUT61), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1193), .A2(new_n1195), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n618), .A2(G213), .A3(G2897), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1207), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1184), .A2(new_n1201), .ZN(new_n1211));
  AND3_X1   g1011(.A1(new_n1196), .A2(new_n1199), .A3(new_n1209), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1210), .B1(new_n1211), .B2(new_n1212), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n1202), .A2(KEYINPUT125), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1214), .A2(KEYINPUT62), .ZN(new_n1215));
  AOI21_X1  g1015(.A(KEYINPUT125), .B1(new_n1202), .B2(KEYINPUT124), .ZN(new_n1216));
  OAI211_X1 g1016(.A(new_n1206), .B(new_n1213), .C1(new_n1215), .C2(new_n1216), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(G393), .B(new_n745), .ZN(new_n1218));
  NOR2_X1   g1018(.A1(new_n925), .A2(new_n927), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n960), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n1220), .B1(new_n999), .B2(new_n669), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1219), .B1(new_n1221), .B2(new_n673), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(new_n1033), .A2(new_n1035), .B1(new_n1222), .B2(new_n902), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n1218), .B1(new_n1170), .B2(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(G390), .A2(G387), .ZN(new_n1225));
  NAND4_X1  g1025(.A1(new_n1033), .A2(new_n1222), .A3(new_n902), .A4(new_n1035), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n1218), .ZN(new_n1227));
  NAND3_X1  g1027(.A1(new_n1225), .A2(new_n1226), .A3(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1224), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1217), .A2(new_n1229), .ZN(new_n1230));
  AND3_X1   g1030(.A1(new_n1213), .A2(new_n1224), .A3(new_n1228), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT63), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1202), .A2(KEYINPUT123), .A3(new_n1232), .ZN(new_n1233));
  OR2_X1    g1033(.A1(new_n1202), .A2(new_n1232), .ZN(new_n1234));
  NAND2_X1  g1034(.A1(new_n1202), .A2(new_n1232), .ZN(new_n1235));
  INV_X1    g1035(.A(KEYINPUT123), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1235), .A2(new_n1236), .ZN(new_n1237));
  NAND4_X1  g1037(.A1(new_n1231), .A2(new_n1233), .A3(new_n1234), .A4(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1230), .A2(new_n1238), .ZN(G405));
  OR2_X1    g1039(.A1(new_n1229), .A2(KEYINPUT127), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1229), .A2(KEYINPUT127), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1208), .ZN(new_n1242));
  AOI21_X1  g1042(.A(G378), .B1(new_n1123), .B2(new_n1147), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1178), .A2(KEYINPUT126), .ZN(new_n1244));
  OR2_X1    g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1242), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1247), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1245), .A2(new_n1200), .A3(new_n1246), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1240), .A2(new_n1241), .A3(new_n1248), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(new_n1249), .ZN(new_n1251));
  OAI211_X1 g1051(.A(KEYINPUT127), .B(new_n1229), .C1(new_n1251), .C2(new_n1247), .ZN(new_n1252));
  NAND2_X1  g1052(.A1(new_n1250), .A2(new_n1252), .ZN(G402));
endmodule


