//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 1 1 1 1 1 0 1 1 0 1 0 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 1 0 0 1 1 0 0 0 1 0 1 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:18:09 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n692, new_n693,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n723, new_n724,
    new_n725, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n763, new_n764,
    new_n765, new_n767, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n862,
    new_n864, new_n866, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n908, new_n909,
    new_n910, new_n911, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n952, new_n953, new_n954, new_n955, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n978,
    new_n979, new_n980, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n999, new_n1000;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  OAI21_X1  g002(.A(new_n202), .B1(new_n203), .B2(G1gat), .ZN(new_n204));
  OAI21_X1  g003(.A(new_n204), .B1(G1gat), .B2(new_n202), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n205), .B(G8gat), .ZN(new_n206));
  INV_X1    g005(.A(new_n206), .ZN(new_n207));
  INV_X1    g006(.A(KEYINPUT15), .ZN(new_n208));
  OR2_X1    g007(.A1(G43gat), .A2(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(G43gat), .A2(G50gat), .ZN(new_n210));
  AOI21_X1  g009(.A(new_n208), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n211), .B1(G29gat), .B2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(G29gat), .ZN(new_n213));
  INV_X1    g012(.A(G36gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT14), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT14), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT92), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n215), .A2(new_n217), .A3(KEYINPUT92), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT91), .B(G43gat), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n208), .B(new_n210), .C1(new_n222), .C2(G50gat), .ZN(new_n223));
  NAND4_X1  g022(.A1(new_n212), .A2(new_n220), .A3(new_n221), .A4(new_n223), .ZN(new_n224));
  OAI22_X1  g023(.A1(new_n218), .A2(KEYINPUT90), .B1(new_n213), .B2(new_n214), .ZN(new_n225));
  AND2_X1   g024(.A1(new_n218), .A2(KEYINPUT90), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n211), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT17), .ZN(new_n228));
  AND3_X1   g027(.A1(new_n224), .A2(new_n227), .A3(new_n228), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n228), .B1(new_n224), .B2(new_n227), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n207), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n224), .A2(new_n227), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n206), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G229gat), .A2(G233gat), .ZN(new_n234));
  NAND4_X1  g033(.A1(new_n231), .A2(KEYINPUT18), .A3(new_n233), .A4(new_n234), .ZN(new_n235));
  XOR2_X1   g034(.A(new_n234), .B(KEYINPUT13), .Z(new_n236));
  INV_X1    g035(.A(new_n233), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n206), .A2(new_n232), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n236), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  AND2_X1   g038(.A1(new_n235), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT93), .ZN(new_n244));
  XNOR2_X1  g043(.A(G113gat), .B(G141gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(G169gat), .B(G197gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT89), .B(KEYINPUT11), .ZN(new_n248));
  XNOR2_X1  g047(.A(new_n247), .B(new_n248), .ZN(new_n249));
  XOR2_X1   g048(.A(new_n249), .B(KEYINPUT12), .Z(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n240), .B(new_n243), .C1(new_n244), .C2(new_n251), .ZN(new_n252));
  NAND3_X1  g051(.A1(new_n235), .A2(new_n244), .A3(new_n239), .ZN(new_n253));
  AND2_X1   g052(.A1(new_n241), .A2(new_n242), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n235), .A2(new_n239), .ZN(new_n255));
  OAI211_X1 g054(.A(new_n253), .B(new_n250), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  AND2_X1   g055(.A1(new_n252), .A2(new_n256), .ZN(new_n257));
  AND2_X1   g056(.A1(G197gat), .A2(G204gat), .ZN(new_n258));
  NOR2_X1   g057(.A1(G197gat), .A2(G204gat), .ZN(new_n259));
  NOR2_X1   g058(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  AND2_X1   g059(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n261));
  NOR2_X1   g060(.A1(KEYINPUT71), .A2(G211gat), .ZN(new_n262));
  OAI21_X1  g061(.A(G218gat), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT22), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n260), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT72), .ZN(new_n266));
  XNOR2_X1  g065(.A(G211gat), .B(G218gat), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n265), .A2(new_n266), .A3(new_n268), .ZN(new_n269));
  OAI21_X1  g068(.A(new_n267), .B1(new_n265), .B2(new_n266), .ZN(new_n270));
  AOI211_X1 g069(.A(KEYINPUT72), .B(new_n260), .C1(new_n264), .C2(new_n263), .ZN(new_n271));
  OAI21_X1  g070(.A(new_n269), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n272), .A2(KEYINPUT73), .ZN(new_n273));
  AND2_X1   g072(.A1(G155gat), .A2(G162gat), .ZN(new_n274));
  NOR2_X1   g073(.A1(G155gat), .A2(G162gat), .ZN(new_n275));
  NOR2_X1   g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  XNOR2_X1  g075(.A(G141gat), .B(G148gat), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT2), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n278), .B1(G155gat), .B2(G162gat), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n276), .B1(new_n277), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(G141gat), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n281), .A2(G148gat), .ZN(new_n282));
  INV_X1    g081(.A(G148gat), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(G141gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  XNOR2_X1  g084(.A(G155gat), .B(G162gat), .ZN(new_n286));
  INV_X1    g085(.A(G155gat), .ZN(new_n287));
  INV_X1    g086(.A(G162gat), .ZN(new_n288));
  OAI21_X1  g087(.A(KEYINPUT2), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n285), .A2(new_n286), .A3(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(KEYINPUT3), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n280), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT29), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  INV_X1    g093(.A(KEYINPUT73), .ZN(new_n295));
  OAI211_X1 g094(.A(new_n295), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n273), .A2(new_n294), .A3(new_n296), .ZN(new_n297));
  OAI211_X1 g096(.A(new_n293), .B(new_n269), .C1(new_n270), .C2(new_n271), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n298), .A2(new_n291), .ZN(new_n299));
  AND3_X1   g098(.A1(new_n280), .A2(new_n290), .A3(KEYINPUT79), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT79), .B1(new_n280), .B2(new_n290), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n299), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g102(.A1(G228gat), .A2(G233gat), .ZN(new_n304));
  INV_X1    g103(.A(new_n304), .ZN(new_n305));
  AND3_X1   g104(.A1(new_n297), .A2(new_n303), .A3(new_n305), .ZN(new_n306));
  NAND2_X1  g105(.A1(new_n280), .A2(new_n290), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n299), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT82), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n280), .A2(new_n290), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n298), .B2(new_n291), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(KEYINPUT82), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n313), .A3(new_n297), .ZN(new_n314));
  AOI21_X1  g113(.A(new_n306), .B1(new_n314), .B2(new_n304), .ZN(new_n315));
  INV_X1    g114(.A(G22gat), .ZN(new_n316));
  AOI21_X1  g115(.A(KEYINPUT83), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g116(.A(G78gat), .B(G106gat), .ZN(new_n318));
  XNOR2_X1  g117(.A(KEYINPUT31), .B(G50gat), .ZN(new_n319));
  XNOR2_X1  g118(.A(new_n318), .B(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(new_n320), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n297), .B1(KEYINPUT82), .B2(new_n312), .ZN(new_n322));
  INV_X1    g121(.A(new_n313), .ZN(new_n323));
  OAI21_X1  g122(.A(new_n304), .B1(new_n322), .B2(new_n323), .ZN(new_n324));
  INV_X1    g123(.A(new_n306), .ZN(new_n325));
  AND3_X1   g124(.A1(new_n324), .A2(new_n316), .A3(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n316), .B1(new_n324), .B2(new_n325), .ZN(new_n327));
  OAI22_X1  g126(.A1(new_n317), .A2(new_n321), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  INV_X1    g127(.A(new_n327), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n315), .A2(new_n316), .ZN(new_n330));
  NAND4_X1  g129(.A1(new_n329), .A2(new_n330), .A3(KEYINPUT83), .A4(new_n320), .ZN(new_n331));
  AND2_X1   g130(.A1(new_n328), .A2(new_n331), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT36), .ZN(new_n333));
  XOR2_X1   g132(.A(G15gat), .B(G43gat), .Z(new_n334));
  XNOR2_X1  g133(.A(G71gat), .B(G99gat), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  INV_X1    g135(.A(G190gat), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT27), .ZN(new_n338));
  OAI211_X1 g137(.A(KEYINPUT65), .B(new_n337), .C1(new_n338), .C2(G183gat), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT28), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT66), .B1(new_n339), .B2(new_n340), .ZN(new_n342));
  AND2_X1   g141(.A1(new_n338), .A2(G183gat), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n337), .B1(new_n338), .B2(G183gat), .ZN(new_n344));
  OAI22_X1  g143(.A1(new_n341), .A2(new_n342), .B1(new_n343), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n339), .A2(new_n340), .ZN(new_n346));
  INV_X1    g145(.A(KEYINPUT66), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n343), .A2(new_n344), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n339), .A2(KEYINPUT66), .A3(new_n340), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n348), .A2(new_n349), .A3(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(G183gat), .A2(G190gat), .ZN(new_n352));
  AOI21_X1  g151(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G169gat), .A2(G176gat), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT67), .ZN(new_n355));
  OR3_X1    g154(.A1(new_n353), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  OR2_X1    g155(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(KEYINPUT68), .A2(KEYINPUT26), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n357), .A2(new_n354), .A3(new_n358), .ZN(new_n359));
  OAI21_X1  g158(.A(new_n355), .B1(new_n353), .B2(new_n354), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n356), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND4_X1  g160(.A1(new_n345), .A2(new_n351), .A3(new_n352), .A4(new_n361), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n354), .A2(KEYINPUT23), .ZN(new_n363));
  NAND2_X1  g162(.A1(G169gat), .A2(G176gat), .ZN(new_n364));
  INV_X1    g163(.A(KEYINPUT23), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n365), .B1(G169gat), .B2(G176gat), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n364), .A3(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n368), .B1(G183gat), .B2(G190gat), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT64), .ZN(new_n370));
  INV_X1    g169(.A(KEYINPUT24), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n352), .B2(new_n371), .ZN(new_n372));
  NOR2_X1   g171(.A1(new_n369), .A2(new_n372), .ZN(new_n373));
  NAND3_X1  g172(.A1(new_n352), .A2(new_n370), .A3(new_n371), .ZN(new_n374));
  AOI21_X1  g173(.A(new_n367), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n363), .A2(KEYINPUT25), .A3(new_n366), .A4(new_n364), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n369), .B1(new_n371), .B2(new_n352), .ZN(new_n377));
  OAI22_X1  g176(.A1(new_n375), .A2(KEYINPUT25), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  XOR2_X1   g177(.A(G127gat), .B(G134gat), .Z(new_n379));
  INV_X1    g178(.A(G120gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G113gat), .ZN(new_n381));
  INV_X1    g180(.A(G113gat), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n382), .A2(G120gat), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n381), .A2(new_n383), .A3(KEYINPUT69), .ZN(new_n384));
  INV_X1    g183(.A(KEYINPUT1), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT69), .B1(new_n381), .B2(new_n383), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n379), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n379), .A2(KEYINPUT1), .ZN(new_n389));
  OR3_X1    g188(.A1(new_n380), .A2(KEYINPUT70), .A3(G113gat), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n383), .A2(KEYINPUT70), .ZN(new_n391));
  NAND3_X1  g190(.A1(new_n390), .A2(new_n391), .A3(new_n381), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n389), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  AND3_X1   g193(.A1(new_n362), .A2(new_n378), .A3(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n394), .B1(new_n362), .B2(new_n378), .ZN(new_n396));
  NAND2_X1  g195(.A1(G227gat), .A2(G233gat), .ZN(new_n397));
  NOR3_X1   g196(.A1(new_n395), .A2(new_n396), .A3(new_n397), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n336), .B1(new_n398), .B2(KEYINPUT33), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n362), .A2(new_n378), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n381), .A2(new_n383), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT69), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n403), .A2(new_n385), .A3(new_n384), .ZN(new_n404));
  AOI22_X1  g203(.A1(new_n404), .A2(new_n379), .B1(new_n389), .B2(new_n392), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n362), .A2(new_n378), .A3(new_n394), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n408), .A2(new_n397), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(KEYINPUT34), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT34), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n411), .B(new_n397), .C1(new_n395), .C2(new_n396), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n399), .A2(new_n410), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n336), .ZN(new_n414));
  NAND4_X1  g213(.A1(new_n406), .A2(G227gat), .A3(G233gat), .A4(new_n407), .ZN(new_n415));
  INV_X1    g214(.A(KEYINPUT33), .ZN(new_n416));
  AOI21_X1  g215(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n411), .B1(new_n408), .B2(new_n397), .ZN(new_n418));
  INV_X1    g217(.A(new_n412), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n415), .A2(KEYINPUT32), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  AND3_X1   g221(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n422), .B1(new_n413), .B2(new_n420), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n333), .B1(new_n423), .B2(new_n424), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n413), .A2(new_n420), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n426), .A2(new_n421), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n413), .A2(new_n420), .A3(new_n422), .ZN(new_n428));
  NAND3_X1  g227(.A1(new_n427), .A2(KEYINPUT36), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n425), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n332), .A2(new_n430), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n328), .A2(new_n331), .ZN(new_n432));
  NAND2_X1  g231(.A1(new_n427), .A2(new_n428), .ZN(new_n433));
  INV_X1    g232(.A(new_n433), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n432), .A2(new_n434), .A3(KEYINPUT35), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n431), .A2(new_n435), .ZN(new_n436));
  XNOR2_X1  g235(.A(G8gat), .B(G36gat), .ZN(new_n437));
  XNOR2_X1  g236(.A(G64gat), .B(G92gat), .ZN(new_n438));
  XOR2_X1   g237(.A(new_n437), .B(new_n438), .Z(new_n439));
  INV_X1    g238(.A(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n296), .ZN(new_n441));
  XNOR2_X1  g240(.A(KEYINPUT71), .B(G211gat), .ZN(new_n442));
  AOI21_X1  g241(.A(KEYINPUT22), .B1(new_n442), .B2(G218gat), .ZN(new_n443));
  OAI21_X1  g242(.A(KEYINPUT72), .B1(new_n443), .B2(new_n260), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n265), .A2(new_n266), .ZN(new_n445));
  NAND3_X1  g244(.A1(new_n444), .A2(new_n445), .A3(new_n267), .ZN(new_n446));
  AOI21_X1  g245(.A(new_n295), .B1(new_n446), .B2(new_n269), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n441), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g247(.A1(G226gat), .A2(G233gat), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  AOI21_X1  g249(.A(new_n450), .B1(new_n400), .B2(new_n293), .ZN(new_n451));
  AOI21_X1  g250(.A(new_n449), .B1(new_n362), .B2(new_n378), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n273), .A2(new_n296), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n400), .A2(new_n450), .ZN(new_n455));
  AOI21_X1  g254(.A(KEYINPUT29), .B1(new_n362), .B2(new_n378), .ZN(new_n456));
  OAI211_X1 g255(.A(new_n454), .B(new_n455), .C1(new_n450), .C2(new_n456), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT74), .ZN(new_n458));
  AOI21_X1  g257(.A(KEYINPUT74), .B1(new_n453), .B2(new_n457), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n440), .B1(new_n458), .B2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT75), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n453), .A2(new_n457), .A3(new_n439), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT30), .ZN(new_n463));
  OAI21_X1  g262(.A(new_n461), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  AND2_X1   g263(.A1(new_n453), .A2(new_n457), .ZN(new_n465));
  NAND4_X1  g264(.A1(new_n465), .A2(KEYINPUT75), .A3(KEYINPUT30), .A4(new_n439), .ZN(new_n466));
  NAND3_X1  g265(.A1(new_n460), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT76), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT76), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n460), .A2(new_n466), .A3(new_n469), .A4(new_n464), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n311), .A2(new_n388), .A3(new_n393), .ZN(new_n471));
  INV_X1    g270(.A(KEYINPUT4), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n405), .A2(KEYINPUT4), .A3(new_n311), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n300), .A2(new_n301), .A3(new_n291), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n394), .A2(new_n292), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(G225gat), .A2(G233gat), .ZN(new_n478));
  INV_X1    g277(.A(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(new_n301), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n280), .A2(new_n290), .A3(KEYINPUT79), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n394), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n478), .B1(new_n482), .B2(new_n471), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT5), .ZN(new_n484));
  OAI22_X1  g283(.A1(new_n477), .A2(new_n479), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  AND2_X1   g284(.A1(new_n473), .A2(new_n474), .ZN(new_n486));
  OR2_X1    g285(.A1(new_n475), .A2(new_n476), .ZN(new_n487));
  NAND4_X1  g286(.A1(new_n486), .A2(new_n487), .A3(KEYINPUT5), .A4(new_n478), .ZN(new_n488));
  XOR2_X1   g287(.A(G1gat), .B(G29gat), .Z(new_n489));
  XNOR2_X1  g288(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n489), .B(new_n490), .ZN(new_n491));
  XNOR2_X1  g290(.A(G57gat), .B(G85gat), .ZN(new_n492));
  XNOR2_X1  g291(.A(new_n491), .B(new_n492), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n485), .A2(new_n488), .A3(new_n493), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT6), .ZN(new_n495));
  OR2_X1    g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n485), .A2(new_n488), .ZN(new_n497));
  INV_X1    g296(.A(new_n493), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT6), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n499), .A2(new_n494), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT77), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n462), .A2(new_n501), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT77), .A4(new_n439), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(KEYINPUT78), .B(KEYINPUT30), .Z(new_n505));
  INV_X1    g304(.A(new_n505), .ZN(new_n506));
  AOI22_X1  g305(.A1(new_n496), .A2(new_n500), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n468), .A2(new_n470), .A3(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT81), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND4_X1  g309(.A1(new_n468), .A2(new_n507), .A3(KEYINPUT81), .A4(new_n470), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n436), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n453), .A2(new_n457), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT88), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT88), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  AOI211_X1 g315(.A(new_n515), .B(new_n516), .C1(new_n453), .C2(new_n457), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n514), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g317(.A(new_n440), .B1(new_n513), .B2(KEYINPUT37), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT38), .ZN(new_n520));
  AOI22_X1  g319(.A1(new_n518), .A2(new_n520), .B1(new_n502), .B2(new_n503), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT84), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n493), .B(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(new_n523), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n524), .A2(new_n485), .A3(new_n488), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n499), .A2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT87), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n497), .A2(new_n498), .ZN(new_n529));
  NAND4_X1  g328(.A1(new_n529), .A2(KEYINPUT87), .A3(new_n495), .A4(new_n525), .ZN(new_n530));
  AND2_X1   g329(.A1(new_n530), .A2(new_n496), .ZN(new_n531));
  INV_X1    g330(.A(KEYINPUT74), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n513), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n453), .A2(new_n457), .A3(KEYINPUT74), .ZN(new_n534));
  AOI21_X1  g333(.A(new_n516), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT38), .B1(new_n535), .B2(new_n519), .ZN(new_n536));
  NAND4_X1  g335(.A1(new_n521), .A2(new_n528), .A3(new_n531), .A4(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n477), .A2(new_n479), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n482), .A2(new_n478), .A3(new_n471), .ZN(new_n539));
  AND3_X1   g338(.A1(new_n538), .A2(KEYINPUT39), .A3(new_n539), .ZN(new_n540));
  INV_X1    g339(.A(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(KEYINPUT39), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n477), .A2(new_n542), .A3(new_n479), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(new_n523), .ZN(new_n544));
  INV_X1    g343(.A(new_n544), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n541), .A2(KEYINPUT40), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT86), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT86), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n541), .A2(new_n548), .A3(new_n545), .A4(KEYINPUT40), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n547), .A2(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(new_n525), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT40), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n540), .B2(new_n544), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n553), .A2(KEYINPUT85), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT85), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n555), .B(new_n552), .C1(new_n540), .C2(new_n544), .ZN(new_n556));
  AOI21_X1  g355(.A(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n505), .B1(new_n502), .B2(new_n503), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n550), .B(new_n557), .C1(new_n467), .C2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n537), .A2(new_n559), .ZN(new_n560));
  AOI22_X1  g359(.A1(new_n425), .A2(new_n429), .B1(new_n328), .B2(new_n331), .ZN(new_n561));
  NAND2_X1  g360(.A1(new_n531), .A2(new_n528), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n467), .A2(new_n558), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n432), .A2(new_n434), .A3(new_n562), .A4(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT35), .ZN(new_n565));
  AOI22_X1  g364(.A1(new_n560), .A2(new_n561), .B1(new_n564), .B2(new_n565), .ZN(new_n566));
  AOI21_X1  g365(.A(new_n257), .B1(new_n512), .B2(new_n566), .ZN(new_n567));
  XOR2_X1   g366(.A(G57gat), .B(G64gat), .Z(new_n568));
  INV_X1    g367(.A(KEYINPUT9), .ZN(new_n569));
  INV_X1    g368(.A(G71gat), .ZN(new_n570));
  INV_X1    g369(.A(G78gat), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n569), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G71gat), .B(G78gat), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n573), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g375(.A1(new_n568), .A2(new_n574), .A3(new_n572), .ZN(new_n577));
  AND3_X1   g376(.A1(new_n576), .A2(KEYINPUT94), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(KEYINPUT94), .B1(new_n576), .B2(new_n577), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g379(.A1(new_n580), .A2(KEYINPUT21), .ZN(new_n581));
  AND2_X1   g380(.A1(G231gat), .A2(G233gat), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n581), .B(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(G127gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n206), .B1(new_n580), .B2(KEYINPUT21), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(new_n583), .B(G127gat), .ZN(new_n588));
  INV_X1    g387(.A(new_n586), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(new_n287), .ZN(new_n593));
  XNOR2_X1  g392(.A(G183gat), .B(G211gat), .ZN(new_n594));
  XOR2_X1   g393(.A(new_n593), .B(new_n594), .Z(new_n595));
  INV_X1    g394(.A(new_n595), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n591), .A2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n587), .A2(new_n590), .A3(new_n595), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  XNOR2_X1  g398(.A(G99gat), .B(G106gat), .ZN(new_n600));
  XNOR2_X1  g399(.A(new_n600), .B(KEYINPUT98), .ZN(new_n601));
  INV_X1    g400(.A(new_n601), .ZN(new_n602));
  NAND2_X1  g401(.A1(G85gat), .A2(G92gat), .ZN(new_n603));
  OAI21_X1  g402(.A(KEYINPUT96), .B1(new_n603), .B2(KEYINPUT7), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT96), .ZN(new_n605));
  INV_X1    g404(.A(KEYINPUT7), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n605), .A2(new_n606), .A3(G85gat), .A4(G92gat), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n604), .A2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT95), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n609), .B1(new_n603), .B2(KEYINPUT7), .ZN(new_n610));
  NAND3_X1  g409(.A1(new_n603), .A2(new_n609), .A3(KEYINPUT7), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n608), .B1(new_n610), .B2(new_n612), .ZN(new_n613));
  INV_X1    g412(.A(KEYINPUT97), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(new_n610), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n611), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n617), .A2(KEYINPUT97), .A3(new_n608), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n615), .A2(new_n618), .ZN(new_n619));
  NAND2_X1  g418(.A1(G99gat), .A2(G106gat), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n620), .A2(KEYINPUT8), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n621), .B1(G85gat), .B2(G92gat), .ZN(new_n622));
  INV_X1    g421(.A(new_n622), .ZN(new_n623));
  AOI21_X1  g422(.A(new_n602), .B1(new_n619), .B2(new_n623), .ZN(new_n624));
  AOI211_X1 g423(.A(new_n622), .B(new_n601), .C1(new_n615), .C2(new_n618), .ZN(new_n625));
  NOR2_X1   g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n232), .ZN(new_n627));
  NAND3_X1  g426(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  OR2_X1    g428(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n629), .A2(KEYINPUT99), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n229), .A2(new_n230), .ZN(new_n632));
  OAI211_X1 g431(.A(new_n630), .B(new_n631), .C1(new_n632), .C2(new_n626), .ZN(new_n633));
  XNOR2_X1  g432(.A(G190gat), .B(G218gat), .ZN(new_n634));
  INV_X1    g433(.A(KEYINPUT100), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n634), .A2(new_n635), .ZN(new_n637));
  AOI21_X1  g436(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G134gat), .B(G162gat), .Z(new_n640));
  XNOR2_X1  g439(.A(new_n639), .B(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n633), .A2(new_n636), .A3(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n641), .B1(new_n633), .B2(new_n636), .ZN(new_n643));
  OR2_X1    g442(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n599), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n580), .B1(new_n624), .B2(new_n625), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n613), .A2(new_n614), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT97), .B1(new_n617), .B2(new_n608), .ZN(new_n649));
  OAI21_X1  g448(.A(new_n623), .B1(new_n648), .B2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n601), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n576), .A2(new_n577), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n619), .A2(new_n602), .A3(new_n623), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n651), .A2(new_n652), .A3(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n647), .A2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT10), .ZN(new_n656));
  NOR3_X1   g455(.A1(new_n578), .A2(new_n579), .A3(new_n656), .ZN(new_n657));
  AOI22_X1  g456(.A1(new_n655), .A2(new_n656), .B1(new_n626), .B2(new_n657), .ZN(new_n658));
  INV_X1    g457(.A(G230gat), .ZN(new_n659));
  INV_X1    g458(.A(G233gat), .ZN(new_n660));
  NOR2_X1   g459(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  OAI21_X1  g460(.A(new_n646), .B1(new_n658), .B2(new_n661), .ZN(new_n662));
  AOI21_X1  g461(.A(KEYINPUT10), .B1(new_n647), .B2(new_n654), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n626), .A2(new_n657), .ZN(new_n664));
  INV_X1    g463(.A(new_n664), .ZN(new_n665));
  OAI221_X1 g464(.A(KEYINPUT101), .B1(new_n659), .B2(new_n660), .C1(new_n663), .C2(new_n665), .ZN(new_n666));
  NOR3_X1   g465(.A1(new_n655), .A2(new_n659), .A3(new_n660), .ZN(new_n667));
  XNOR2_X1  g466(.A(G120gat), .B(G148gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(G176gat), .B(G204gat), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n668), .B(new_n669), .Z(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n667), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n662), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n663), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n661), .B1(new_n674), .B2(new_n664), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n671), .B1(new_n675), .B2(new_n667), .ZN(new_n676));
  NAND2_X1  g475(.A1(new_n673), .A2(new_n676), .ZN(new_n677));
  NOR2_X1   g476(.A1(new_n645), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n567), .A2(new_n678), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n500), .A2(new_n496), .ZN(new_n681));
  XOR2_X1   g480(.A(new_n681), .B(KEYINPUT102), .Z(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  NAND2_X1  g482(.A1(new_n680), .A2(new_n683), .ZN(new_n684));
  XNOR2_X1  g483(.A(new_n684), .B(G1gat), .ZN(G1324gat));
  INV_X1    g484(.A(new_n563), .ZN(new_n686));
  XOR2_X1   g485(.A(KEYINPUT16), .B(G8gat), .Z(new_n687));
  NAND3_X1  g486(.A1(new_n680), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  OAI21_X1  g487(.A(G8gat), .B1(new_n679), .B2(new_n563), .ZN(new_n689));
  NAND2_X1  g488(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  MUX2_X1   g489(.A(new_n688), .B(new_n690), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g490(.A(G15gat), .B1(new_n679), .B2(new_n430), .ZN(new_n692));
  OR2_X1    g491(.A1(new_n433), .A2(G15gat), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n692), .B1(new_n679), .B2(new_n693), .ZN(G1326gat));
  NAND2_X1  g493(.A1(new_n680), .A2(new_n332), .ZN(new_n695));
  XNOR2_X1  g494(.A(new_n695), .B(KEYINPUT103), .ZN(new_n696));
  XNOR2_X1  g495(.A(KEYINPUT43), .B(G22gat), .ZN(new_n697));
  XNOR2_X1  g496(.A(new_n696), .B(new_n697), .ZN(G1327gat));
  AOI21_X1  g497(.A(new_n644), .B1(new_n512), .B2(new_n566), .ZN(new_n699));
  NOR3_X1   g498(.A1(new_n599), .A2(new_n257), .A3(new_n677), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n701), .A2(new_n213), .A3(new_n683), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT45), .ZN(new_n703));
  INV_X1    g502(.A(new_n644), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n433), .B1(new_n331), .B2(new_n328), .ZN(new_n705));
  AOI22_X1  g504(.A1(KEYINPUT35), .A2(new_n705), .B1(new_n332), .B2(new_n430), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n510), .A2(new_n511), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n560), .A2(new_n561), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n564), .A2(new_n565), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(new_n704), .B1(new_n708), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT44), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n512), .A2(new_n566), .ZN(new_n715));
  NAND3_X1  g514(.A1(new_n715), .A2(KEYINPUT44), .A3(new_n704), .ZN(new_n716));
  AND2_X1   g515(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n700), .ZN(new_n718));
  OAI21_X1  g517(.A(KEYINPUT104), .B1(new_n718), .B2(new_n682), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n719), .A2(G29gat), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(KEYINPUT104), .A3(new_n682), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n703), .B1(new_n720), .B2(new_n721), .ZN(G1328gat));
  OAI21_X1  g521(.A(G36gat), .B1(new_n718), .B2(new_n563), .ZN(new_n723));
  NOR4_X1   g522(.A1(new_n599), .A2(new_n644), .A3(G36gat), .A4(new_n677), .ZN(new_n724));
  NAND3_X1  g523(.A1(new_n567), .A2(new_n686), .A3(new_n724), .ZN(new_n725));
  XOR2_X1   g524(.A(new_n725), .B(KEYINPUT46), .Z(new_n726));
  NAND2_X1  g525(.A1(new_n723), .A2(new_n726), .ZN(G1329gat));
  INV_X1    g526(.A(new_n430), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n714), .A2(new_n728), .A3(new_n716), .A4(new_n700), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n222), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n433), .A2(new_n222), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n701), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g531(.A1(new_n730), .A2(KEYINPUT47), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g532(.A1(new_n729), .A2(KEYINPUT106), .A3(new_n222), .ZN(new_n734));
  AOI21_X1  g533(.A(KEYINPUT106), .B1(new_n729), .B2(new_n222), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n732), .A2(KEYINPUT107), .ZN(new_n736));
  INV_X1    g535(.A(KEYINPUT107), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n737), .B1(new_n701), .B2(new_n731), .ZN(new_n738));
  NOR4_X1   g537(.A1(new_n734), .A2(new_n735), .A3(new_n736), .A4(new_n738), .ZN(new_n739));
  XNOR2_X1  g538(.A(KEYINPUT105), .B(KEYINPUT47), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n733), .B1(new_n739), .B2(new_n740), .ZN(G1330gat));
  NAND4_X1  g540(.A1(new_n714), .A2(new_n332), .A3(new_n716), .A4(new_n700), .ZN(new_n742));
  NAND2_X1  g541(.A1(new_n742), .A2(G50gat), .ZN(new_n743));
  AOI21_X1  g542(.A(KEYINPUT48), .B1(new_n743), .B2(KEYINPUT108), .ZN(new_n744));
  INV_X1    g543(.A(G50gat), .ZN(new_n745));
  NAND3_X1  g544(.A1(new_n701), .A2(new_n745), .A3(new_n332), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n744), .B(new_n747), .ZN(G1331gat));
  INV_X1    g547(.A(new_n257), .ZN(new_n749));
  INV_X1    g548(.A(new_n677), .ZN(new_n750));
  NOR3_X1   g549(.A1(new_n645), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n715), .A2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(new_n683), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(G57gat), .ZN(G1332gat));
  XNOR2_X1  g554(.A(new_n563), .B(KEYINPUT109), .ZN(new_n756));
  INV_X1    g555(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g556(.A1(new_n752), .A2(new_n757), .ZN(new_n758));
  NOR2_X1   g557(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n759));
  AND2_X1   g558(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n758), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(new_n761), .B1(new_n758), .B2(new_n759), .ZN(G1333gat));
  OAI21_X1  g561(.A(G71gat), .B1(new_n752), .B2(new_n430), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n434), .A2(new_n570), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n763), .B1(new_n752), .B2(new_n764), .ZN(new_n765));
  XOR2_X1   g564(.A(new_n765), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g565(.A1(new_n752), .A2(new_n432), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(new_n571), .ZN(G1335gat));
  INV_X1    g567(.A(new_n599), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(new_n257), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n770), .A2(new_n750), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n717), .A2(new_n771), .ZN(new_n772));
  OAI21_X1  g571(.A(G85gat), .B1(new_n772), .B2(new_n682), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n770), .B1(new_n699), .B2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT110), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n712), .A2(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(KEYINPUT51), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT51), .B1(new_n774), .B2(new_n776), .ZN(new_n779));
  OAI21_X1  g578(.A(new_n677), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  OR2_X1    g579(.A1(new_n682), .A2(G85gat), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n773), .B1(new_n780), .B2(new_n781), .ZN(G1336gat));
  INV_X1    g581(.A(KEYINPUT112), .ZN(new_n783));
  OAI211_X1 g582(.A(KEYINPUT110), .B(new_n704), .C1(new_n708), .C2(new_n711), .ZN(new_n784));
  INV_X1    g583(.A(new_n770), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n699), .A2(KEYINPUT110), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n783), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT51), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n774), .A2(new_n776), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n791), .A2(new_n783), .A3(KEYINPUT51), .ZN(new_n792));
  NOR3_X1   g591(.A1(new_n757), .A2(G92gat), .A3(new_n750), .ZN(new_n793));
  AND3_X1   g592(.A1(new_n790), .A2(new_n792), .A3(new_n793), .ZN(new_n794));
  NAND4_X1  g593(.A1(new_n714), .A2(new_n686), .A3(new_n716), .A4(new_n771), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n795), .A2(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT111), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n795), .A2(KEYINPUT111), .A3(G92gat), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT52), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g600(.A(G92gat), .B1(new_n772), .B2(new_n757), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT52), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n778), .A2(new_n779), .ZN(new_n804));
  INV_X1    g603(.A(new_n793), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n802), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n801), .A2(new_n806), .ZN(G1337gat));
  INV_X1    g606(.A(KEYINPUT113), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n717), .A2(new_n728), .A3(new_n771), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(G99gat), .ZN(new_n810));
  INV_X1    g609(.A(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n433), .A2(G99gat), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n789), .B1(new_n786), .B2(new_n787), .ZN(new_n814));
  AOI211_X1 g613(.A(new_n750), .B(new_n813), .C1(new_n814), .C2(new_n777), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n808), .B1(new_n811), .B2(new_n815), .ZN(new_n816));
  OAI211_X1 g615(.A(KEYINPUT113), .B(new_n810), .C1(new_n780), .C2(new_n813), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n816), .A2(new_n817), .ZN(G1338gat));
  NAND4_X1  g617(.A1(new_n714), .A2(new_n332), .A3(new_n716), .A4(new_n771), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n819), .A2(G106gat), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(KEYINPUT53), .ZN(new_n821));
  NOR3_X1   g620(.A1(new_n432), .A2(G106gat), .A3(new_n750), .ZN(new_n822));
  INV_X1    g621(.A(new_n822), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n821), .B1(new_n804), .B2(new_n823), .ZN(new_n824));
  AOI21_X1  g623(.A(KEYINPUT51), .B1(new_n791), .B2(new_n783), .ZN(new_n825));
  AOI211_X1 g624(.A(KEYINPUT112), .B(new_n789), .C1(new_n774), .C2(new_n776), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n820), .B1(new_n827), .B2(new_n822), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT53), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n824), .B1(new_n828), .B2(new_n829), .ZN(G1339gat));
  NAND3_X1  g629(.A1(new_n240), .A2(new_n243), .A3(new_n251), .ZN(new_n831));
  AOI21_X1  g630(.A(new_n234), .B1(new_n231), .B2(new_n233), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n237), .A2(new_n238), .A3(new_n236), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n249), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n831), .A2(new_n834), .ZN(new_n835));
  NOR3_X1   g634(.A1(new_n642), .A2(new_n643), .A3(new_n835), .ZN(new_n836));
  INV_X1    g635(.A(KEYINPUT54), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n837), .B1(new_n658), .B2(new_n661), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n662), .A2(new_n838), .A3(new_n666), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n670), .B1(new_n675), .B2(new_n837), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n839), .A2(KEYINPUT55), .A3(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n841), .A2(new_n673), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n839), .A2(new_n840), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT55), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n843), .A2(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n836), .A2(new_n842), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g645(.A(new_n835), .B1(new_n673), .B2(new_n676), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n257), .B1(new_n843), .B2(new_n844), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n847), .B1(new_n842), .B2(new_n848), .ZN(new_n849));
  OAI21_X1  g648(.A(new_n846), .B1(new_n849), .B2(new_n704), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n769), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n678), .A2(new_n257), .ZN(new_n852));
  AOI21_X1  g651(.A(new_n682), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n705), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(new_n757), .ZN(new_n855));
  INV_X1    g654(.A(new_n855), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n856), .A2(new_n749), .ZN(new_n857));
  AND2_X1   g656(.A1(KEYINPUT114), .A2(G113gat), .ZN(new_n858));
  NOR2_X1   g657(.A1(KEYINPUT114), .A2(G113gat), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n857), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n860), .B1(new_n857), .B2(new_n858), .ZN(G1340gat));
  NOR2_X1   g660(.A1(new_n855), .A2(new_n750), .ZN(new_n862));
  XNOR2_X1  g661(.A(new_n862), .B(new_n380), .ZN(G1341gat));
  NOR2_X1   g662(.A1(new_n855), .A2(new_n769), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n864), .B(new_n584), .ZN(G1342gat));
  NAND2_X1  g664(.A1(new_n856), .A2(new_n704), .ZN(new_n866));
  INV_X1    g665(.A(G134gat), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n644), .A2(new_n686), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n854), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI22_X1  g668(.A1(new_n866), .A2(G134gat), .B1(KEYINPUT56), .B2(new_n869), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(KEYINPUT56), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT115), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  NOR3_X1   g672(.A1(new_n869), .A2(KEYINPUT115), .A3(KEYINPUT56), .ZN(new_n874));
  OAI21_X1  g673(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(G1343gat));
  INV_X1    g674(.A(new_n431), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n853), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n257), .A2(G141gat), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n877), .A2(new_n757), .A3(new_n878), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(KEYINPUT116), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(KEYINPUT58), .ZN(new_n881));
  NAND3_X1  g680(.A1(new_n757), .A2(new_n430), .A3(new_n683), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n851), .A2(new_n852), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n332), .ZN(new_n884));
  INV_X1    g683(.A(KEYINPUT57), .ZN(new_n885));
  NAND2_X1  g684(.A1(new_n884), .A2(new_n885), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n883), .A2(KEYINPUT57), .A3(new_n332), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n888), .A2(new_n749), .ZN(new_n889));
  OAI211_X1 g688(.A(new_n881), .B(new_n879), .C1(new_n889), .C2(new_n281), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n281), .B1(new_n888), .B2(new_n749), .ZN(new_n891));
  INV_X1    g690(.A(new_n879), .ZN(new_n892));
  OAI211_X1 g691(.A(KEYINPUT58), .B(new_n880), .C1(new_n891), .C2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n890), .A2(new_n893), .ZN(G1344gat));
  AOI211_X1 g693(.A(KEYINPUT59), .B(new_n283), .C1(new_n888), .C2(new_n677), .ZN(new_n895));
  INV_X1    g694(.A(KEYINPUT59), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n850), .A2(KEYINPUT117), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT117), .ZN(new_n898));
  OAI211_X1 g697(.A(new_n898), .B(new_n846), .C1(new_n849), .C2(new_n704), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n897), .A2(new_n769), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n432), .B1(new_n900), .B2(new_n852), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n887), .B1(new_n901), .B2(KEYINPUT57), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n882), .A2(new_n750), .ZN(new_n903));
  NAND2_X1  g702(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  AOI21_X1  g703(.A(new_n896), .B1(new_n904), .B2(G148gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n903), .A2(new_n283), .ZN(new_n906));
  OAI22_X1  g705(.A1(new_n895), .A2(new_n905), .B1(new_n884), .B2(new_n906), .ZN(G1345gat));
  NAND2_X1  g706(.A1(new_n853), .A2(new_n876), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n908), .A2(new_n756), .ZN(new_n909));
  AOI21_X1  g708(.A(G155gat), .B1(new_n909), .B2(new_n599), .ZN(new_n910));
  NOR2_X1   g709(.A1(new_n769), .A2(new_n287), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n910), .B1(new_n888), .B2(new_n911), .ZN(G1346gat));
  NAND3_X1  g711(.A1(new_n877), .A2(new_n288), .A3(new_n868), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n888), .A2(new_n704), .ZN(new_n914));
  OAI211_X1 g713(.A(KEYINPUT118), .B(new_n913), .C1(new_n914), .C2(new_n288), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT118), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n288), .B1(new_n888), .B2(new_n704), .ZN(new_n917));
  INV_X1    g716(.A(new_n913), .ZN(new_n918));
  OAI21_X1  g717(.A(new_n916), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n915), .A2(new_n919), .ZN(G1347gat));
  NOR2_X1   g719(.A1(new_n683), .A2(new_n563), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n921), .A2(new_n434), .ZN(new_n922));
  INV_X1    g721(.A(KEYINPUT120), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n432), .B1(new_n922), .B2(new_n923), .ZN(new_n924));
  AOI21_X1  g723(.A(new_n924), .B1(new_n923), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n925), .A2(new_n883), .ZN(new_n926));
  INV_X1    g725(.A(G169gat), .ZN(new_n927));
  NOR3_X1   g726(.A1(new_n926), .A2(new_n927), .A3(new_n257), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n756), .A2(new_n705), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n929), .B(KEYINPUT119), .Z(new_n930));
  AOI21_X1  g729(.A(new_n683), .B1(new_n851), .B2(new_n852), .ZN(new_n931));
  AND2_X1   g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  AOI21_X1  g731(.A(G169gat), .B1(new_n932), .B2(new_n749), .ZN(new_n933));
  NOR2_X1   g732(.A1(new_n928), .A2(new_n933), .ZN(G1348gat));
  NAND4_X1  g733(.A1(new_n925), .A2(G176gat), .A3(new_n677), .A4(new_n883), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n935), .B(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n932), .A2(new_n677), .ZN(new_n937));
  INV_X1    g736(.A(G176gat), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n937), .A2(KEYINPUT121), .A3(new_n938), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n937), .B2(new_n938), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n936), .A2(new_n939), .A3(new_n940), .ZN(G1349gat));
  NOR2_X1   g740(.A1(new_n338), .A2(G183gat), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n769), .A2(new_n343), .A3(new_n942), .ZN(new_n943));
  NAND3_X1  g742(.A1(new_n930), .A2(new_n931), .A3(new_n943), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT123), .ZN(new_n945));
  OAI21_X1  g744(.A(G183gat), .B1(new_n926), .B2(new_n769), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n947), .A2(KEYINPUT60), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT60), .ZN(new_n949));
  NAND3_X1  g748(.A1(new_n945), .A2(new_n946), .A3(new_n949), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1350gat));
  NAND3_X1  g750(.A1(new_n932), .A2(new_n337), .A3(new_n704), .ZN(new_n952));
  OAI21_X1  g751(.A(G190gat), .B1(new_n926), .B2(new_n644), .ZN(new_n953));
  AND2_X1   g752(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n954));
  NOR2_X1   g753(.A1(new_n953), .A2(KEYINPUT61), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1351gat));
  INV_X1    g755(.A(G197gat), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n921), .A2(new_n430), .ZN(new_n958));
  XNOR2_X1  g757(.A(new_n958), .B(KEYINPUT125), .ZN(new_n959));
  INV_X1    g758(.A(new_n959), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n645), .A2(new_n749), .A3(new_n677), .ZN(new_n961));
  AOI21_X1  g760(.A(new_n599), .B1(new_n850), .B2(KEYINPUT117), .ZN(new_n962));
  AOI21_X1  g761(.A(new_n961), .B1(new_n962), .B2(new_n899), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n885), .B1(new_n963), .B2(new_n432), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n960), .B1(new_n964), .B2(new_n887), .ZN(new_n965));
  AOI21_X1  g764(.A(new_n957), .B1(new_n965), .B2(new_n749), .ZN(new_n966));
  NOR2_X1   g765(.A1(new_n757), .A2(new_n431), .ZN(new_n967));
  AND2_X1   g766(.A1(new_n931), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g767(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n969));
  AND3_X1   g768(.A1(new_n931), .A2(KEYINPUT124), .A3(new_n967), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n749), .A2(new_n957), .ZN(new_n971));
  NOR3_X1   g770(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  OAI21_X1  g771(.A(KEYINPUT126), .B1(new_n966), .B2(new_n972), .ZN(new_n973));
  NAND3_X1  g772(.A1(new_n902), .A2(new_n749), .A3(new_n959), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(G197gat), .ZN(new_n975));
  OR2_X1    g774(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n976));
  INV_X1    g775(.A(new_n970), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n976), .A2(new_n957), .A3(new_n749), .A4(new_n977), .ZN(new_n978));
  INV_X1    g777(.A(KEYINPUT126), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n975), .A2(new_n978), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n973), .A2(new_n980), .ZN(G1352gat));
  INV_X1    g780(.A(G204gat), .ZN(new_n982));
  NAND3_X1  g781(.A1(new_n968), .A2(new_n982), .A3(new_n677), .ZN(new_n983));
  XNOR2_X1  g782(.A(new_n983), .B(KEYINPUT62), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n965), .B2(new_n677), .ZN(new_n985));
  OR2_X1    g784(.A1(new_n984), .A2(new_n985), .ZN(G1353gat));
  NOR2_X1   g785(.A1(new_n969), .A2(new_n970), .ZN(new_n987));
  INV_X1    g786(.A(new_n442), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n987), .A2(new_n988), .A3(new_n599), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT127), .ZN(new_n990));
  OAI21_X1  g789(.A(G211gat), .B1(new_n990), .B2(KEYINPUT63), .ZN(new_n991));
  NOR2_X1   g790(.A1(new_n958), .A2(new_n769), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n902), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n990), .A2(KEYINPUT63), .ZN(new_n994));
  INV_X1    g793(.A(new_n994), .ZN(new_n995));
  NOR2_X1   g794(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI211_X1 g795(.A(new_n994), .B(new_n991), .C1(new_n902), .C2(new_n992), .ZN(new_n997));
  OAI21_X1  g796(.A(new_n989), .B1(new_n996), .B2(new_n997), .ZN(G1354gat));
  AOI21_X1  g797(.A(G218gat), .B1(new_n987), .B2(new_n704), .ZN(new_n999));
  AND2_X1   g798(.A1(new_n704), .A2(G218gat), .ZN(new_n1000));
  AOI21_X1  g799(.A(new_n999), .B1(new_n965), .B2(new_n1000), .ZN(G1355gat));
endmodule


