//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 0 0 0 1 1 1 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 0 1 0 1 0 0 1 1 0 1 0 1 0 0 1 0 1 0 1 0 1 1 1 0 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:33 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n551, new_n552, new_n553, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n610, new_n613, new_n615, new_n616, new_n617, new_n618, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n835, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  XNOR2_X1  g009(.A(KEYINPUT65), .B(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G218), .A2(G219), .A3(G220), .A4(G221), .ZN(new_n450));
  XOR2_X1   g025(.A(KEYINPUT66), .B(KEYINPUT2), .Z(new_n451));
  XNOR2_X1  g026(.A(new_n450), .B(new_n451), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  XOR2_X1   g028(.A(new_n453), .B(KEYINPUT67), .Z(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  NAND2_X1  g031(.A1(new_n452), .A2(G2106), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n454), .A2(G567), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2105), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT68), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT68), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n466), .A2(new_n468), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n464), .A2(new_n469), .ZN(new_n470));
  AND2_X1   g045(.A1(new_n465), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G101), .ZN(new_n472));
  AND2_X1   g047(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n473));
  NOR2_X1   g048(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n474));
  OAI211_X1 g049(.A(new_n466), .B(new_n468), .C1(new_n473), .C2(new_n474), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n472), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(G160));
  XNOR2_X1  g055(.A(KEYINPUT68), .B(G2105), .ZN(new_n481));
  OAI221_X1 g056(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n481), .C2(G112), .ZN(new_n482));
  XOR2_X1   g057(.A(new_n482), .B(KEYINPUT69), .Z(new_n483));
  NAND2_X1  g058(.A1(new_n469), .A2(new_n461), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(new_n485));
  NOR2_X1   g060(.A1(new_n473), .A2(new_n474), .ZN(new_n486));
  NOR2_X1   g061(.A1(new_n486), .A2(G2105), .ZN(new_n487));
  AOI22_X1  g062(.A1(new_n485), .A2(G124), .B1(new_n487), .B2(G136), .ZN(new_n488));
  AND2_X1   g063(.A1(new_n483), .A2(new_n488), .ZN(G162));
  OAI21_X1  g064(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n490));
  INV_X1    g065(.A(G114), .ZN(new_n491));
  AOI21_X1  g066(.A(new_n490), .B1(new_n491), .B2(G2105), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n461), .A2(new_n481), .A3(G138), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT70), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n494), .A2(KEYINPUT4), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n492), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(G126), .A2(G2105), .ZN(new_n497));
  NAND3_X1  g072(.A1(new_n494), .A2(KEYINPUT4), .A3(G138), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n497), .B1(new_n469), .B2(new_n498), .ZN(new_n499));
  NAND2_X1  g074(.A1(new_n499), .A2(new_n461), .ZN(new_n500));
  AND3_X1   g075(.A1(new_n496), .A2(KEYINPUT71), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g076(.A(KEYINPUT71), .B1(new_n496), .B2(new_n500), .ZN(new_n502));
  NOR2_X1   g077(.A1(new_n501), .A2(new_n502), .ZN(G164));
  INV_X1    g078(.A(G543), .ZN(new_n504));
  INV_X1    g079(.A(KEYINPUT6), .ZN(new_n505));
  INV_X1    g080(.A(G651), .ZN(new_n506));
  OAI21_X1  g081(.A(new_n505), .B1(new_n506), .B2(KEYINPUT72), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT72), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT6), .A3(G651), .ZN(new_n509));
  AOI21_X1  g084(.A(new_n504), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G50), .ZN(new_n511));
  INV_X1    g086(.A(G88), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(new_n504), .ZN(new_n514));
  NAND2_X1  g089(.A1(KEYINPUT5), .A2(G543), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(new_n509), .ZN(new_n517));
  AOI21_X1  g092(.A(KEYINPUT6), .B1(new_n508), .B2(G651), .ZN(new_n518));
  OAI21_X1  g093(.A(new_n516), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n511), .B1(new_n512), .B2(new_n519), .ZN(new_n520));
  AOI22_X1  g095(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n521));
  NOR2_X1   g096(.A1(new_n521), .A2(new_n506), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n520), .A2(new_n522), .ZN(G166));
  NAND3_X1  g098(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT7), .ZN(new_n525));
  INV_X1    g100(.A(G89), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n519), .B2(new_n526), .ZN(new_n527));
  XOR2_X1   g102(.A(new_n527), .B(KEYINPUT74), .Z(new_n528));
  XOR2_X1   g103(.A(KEYINPUT73), .B(G51), .Z(new_n529));
  AND2_X1   g104(.A1(G63), .A2(G651), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n510), .A2(new_n529), .B1(new_n516), .B2(new_n530), .ZN(new_n531));
  AND2_X1   g106(.A1(new_n528), .A2(new_n531), .ZN(G168));
  AOI22_X1  g107(.A1(new_n507), .A2(new_n509), .B1(new_n514), .B2(new_n515), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G90), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  AOI21_X1  g110(.A(new_n535), .B1(new_n514), .B2(new_n515), .ZN(new_n536));
  AND2_X1   g111(.A1(G77), .A2(G543), .ZN(new_n537));
  OAI21_X1  g112(.A(G651), .B1(new_n536), .B2(new_n537), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n510), .A2(G52), .ZN(new_n539));
  AND3_X1   g114(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(G171));
  XNOR2_X1  g115(.A(KEYINPUT75), .B(G81), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n533), .A2(new_n541), .ZN(new_n542));
  INV_X1    g117(.A(G56), .ZN(new_n543));
  AOI21_X1  g118(.A(new_n543), .B1(new_n514), .B2(new_n515), .ZN(new_n544));
  AND2_X1   g119(.A1(G68), .A2(G543), .ZN(new_n545));
  OAI21_X1  g120(.A(G651), .B1(new_n544), .B2(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n510), .A2(G43), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  NAND4_X1  g124(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g125(.A1(G1), .A2(G3), .ZN(new_n551));
  XNOR2_X1  g126(.A(new_n551), .B(KEYINPUT76), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND4_X1  g128(.A1(G319), .A2(G483), .A3(G661), .A4(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n533), .A2(G91), .ZN(new_n555));
  AOI22_X1  g130(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT78), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n506), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n516), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(KEYINPUT78), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n555), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND3_X1  g139(.A1(new_n510), .A2(new_n564), .A3(G53), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(KEYINPUT77), .ZN(new_n567));
  AOI21_X1  g142(.A(new_n564), .B1(new_n510), .B2(G53), .ZN(new_n568));
  NOR3_X1   g143(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  OAI211_X1 g144(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(KEYINPUT9), .ZN(new_n571));
  AOI21_X1  g146(.A(KEYINPUT77), .B1(new_n571), .B2(new_n565), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n563), .B1(new_n569), .B2(new_n572), .ZN(G299));
  NAND3_X1  g148(.A1(new_n534), .A2(new_n538), .A3(new_n539), .ZN(G301));
  NAND2_X1  g149(.A1(new_n528), .A2(new_n531), .ZN(G286));
  INV_X1    g150(.A(G166), .ZN(G303));
  INV_X1    g151(.A(G74), .ZN(new_n577));
  NAND3_X1  g152(.A1(new_n514), .A2(new_n577), .A3(new_n515), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n533), .A2(G87), .B1(G651), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n510), .A2(G49), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n579), .A2(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(new_n510), .A2(G48), .ZN(new_n582));
  INV_X1    g157(.A(G86), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n583), .B2(new_n519), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n516), .A2(G61), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT79), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT79), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n516), .A2(new_n587), .A3(G61), .ZN(new_n588));
  NAND2_X1  g163(.A1(G73), .A2(G543), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  AOI21_X1  g165(.A(new_n584), .B1(G651), .B2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OR2_X1    g168(.A1(new_n593), .A2(new_n506), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n510), .A2(G47), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n533), .A2(G85), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(G290));
  NAND2_X1  g172(.A1(G301), .A2(G868), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n510), .A2(G54), .ZN(new_n599));
  AOI22_X1  g174(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n600), .B2(new_n506), .ZN(new_n601));
  INV_X1    g176(.A(KEYINPUT10), .ZN(new_n602));
  INV_X1    g177(.A(G92), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n519), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g179(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n601), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n598), .B1(new_n606), .B2(G868), .ZN(G321));
  INV_X1    g183(.A(G868), .ZN(new_n609));
  NAND2_X1  g184(.A1(G299), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G168), .B2(new_n609), .ZN(G297));
  OAI21_X1  g186(.A(new_n610), .B1(G168), .B2(new_n609), .ZN(G280));
  XNOR2_X1  g187(.A(KEYINPUT80), .B(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n606), .B1(G860), .B2(new_n613), .ZN(G148));
  NAND3_X1  g189(.A1(new_n542), .A2(new_n546), .A3(new_n547), .ZN(new_n615));
  NAND2_X1  g190(.A1(new_n615), .A2(new_n609), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n606), .A2(new_n613), .ZN(new_n617));
  INV_X1    g192(.A(new_n617), .ZN(new_n618));
  OAI21_X1  g193(.A(new_n616), .B1(new_n618), .B2(new_n609), .ZN(G323));
  XNOR2_X1  g194(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g195(.A1(new_n461), .A2(new_n471), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(KEYINPUT12), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT81), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  INV_X1    g199(.A(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT82), .ZN(new_n627));
  AOI22_X1  g202(.A1(new_n485), .A2(G123), .B1(new_n487), .B2(G135), .ZN(new_n628));
  OAI221_X1 g203(.A(G2104), .B1(G99), .B2(G2105), .C1(new_n481), .C2(G111), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  XOR2_X1   g205(.A(new_n630), .B(G2096), .Z(new_n631));
  OAI211_X1 g206(.A(new_n627), .B(new_n631), .C1(new_n625), .C2(new_n624), .ZN(G156));
  INV_X1    g207(.A(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(G2427), .B(G2438), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2430), .ZN(new_n635));
  XNOR2_X1  g210(.A(KEYINPUT15), .B(G2435), .ZN(new_n636));
  AOI21_X1  g211(.A(new_n633), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g212(.A(new_n637), .B1(new_n636), .B2(new_n635), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2451), .B(G2454), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT16), .ZN(new_n640));
  XNOR2_X1  g215(.A(G1341), .B(G1348), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n640), .B(new_n641), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n638), .B(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2443), .B(G2446), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  AND3_X1   g221(.A1(new_n645), .A2(G14), .A3(new_n646), .ZN(G401));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT17), .Z(new_n649));
  XNOR2_X1  g224(.A(G2067), .B(G2678), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n649), .A2(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(G2084), .B(G2090), .ZN(new_n653));
  OAI21_X1  g228(.A(new_n653), .B1(new_n650), .B2(new_n648), .ZN(new_n654));
  NOR2_X1   g229(.A1(new_n652), .A2(new_n654), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT83), .ZN(new_n656));
  NAND2_X1  g231(.A1(new_n650), .A2(new_n648), .ZN(new_n657));
  NOR2_X1   g232(.A1(new_n657), .A2(new_n653), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT18), .Z(new_n659));
  NOR2_X1   g234(.A1(new_n650), .A2(new_n653), .ZN(new_n660));
  AOI21_X1  g235(.A(new_n659), .B1(new_n649), .B2(new_n660), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n656), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2096), .B(G2100), .Z(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(G227));
  XOR2_X1   g239(.A(G1991), .B(G1996), .Z(new_n665));
  XNOR2_X1  g240(.A(G1956), .B(G2474), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT85), .ZN(new_n667));
  XNOR2_X1  g242(.A(G1961), .B(G1966), .ZN(new_n668));
  OR2_X1    g243(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(KEYINPUT84), .B(KEYINPUT19), .Z(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  NOR2_X1   g247(.A1(new_n669), .A2(new_n672), .ZN(new_n673));
  INV_X1    g248(.A(KEYINPUT20), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n669), .A2(new_n672), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n667), .A2(new_n668), .ZN(new_n677));
  MUX2_X1   g252(.A(new_n672), .B(new_n676), .S(new_n677), .Z(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n679));
  NAND3_X1  g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  INV_X1    g255(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n682));
  OAI21_X1  g257(.A(new_n665), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  INV_X1    g258(.A(new_n682), .ZN(new_n684));
  INV_X1    g259(.A(new_n665), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n684), .A2(new_n685), .A3(new_n680), .ZN(new_n686));
  XNOR2_X1  g261(.A(G1981), .B(G1986), .ZN(new_n687));
  AND3_X1   g262(.A1(new_n683), .A2(new_n686), .A3(new_n687), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n687), .B1(new_n683), .B2(new_n686), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(new_n689), .ZN(G229));
  AOI22_X1  g265(.A1(new_n487), .A2(G141), .B1(G105), .B2(new_n471), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n485), .A2(G129), .ZN(new_n692));
  NAND3_X1  g267(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT26), .Z(new_n694));
  NAND3_X1  g269(.A1(new_n691), .A2(new_n692), .A3(new_n694), .ZN(new_n695));
  INV_X1    g270(.A(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(G29), .ZN(new_n697));
  NOR2_X1   g272(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  AOI21_X1  g273(.A(new_n698), .B1(new_n697), .B2(G32), .ZN(new_n699));
  XNOR2_X1  g274(.A(KEYINPUT27), .B(G1996), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  OR2_X1    g276(.A1(G29), .A2(G33), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n481), .A2(G103), .A3(G2104), .ZN(new_n703));
  XOR2_X1   g278(.A(KEYINPUT96), .B(KEYINPUT25), .Z(new_n704));
  XNOR2_X1  g279(.A(new_n703), .B(new_n704), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n487), .A2(G139), .ZN(new_n706));
  AOI22_X1  g281(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n707));
  OAI211_X1 g282(.A(new_n705), .B(new_n706), .C1(new_n481), .C2(new_n707), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n702), .B1(new_n708), .B2(new_n697), .ZN(new_n709));
  INV_X1    g284(.A(G2072), .ZN(new_n710));
  OAI21_X1  g285(.A(new_n701), .B1(new_n709), .B2(new_n710), .ZN(new_n711));
  INV_X1    g286(.A(KEYINPUT24), .ZN(new_n712));
  INV_X1    g287(.A(G34), .ZN(new_n713));
  AOI21_X1  g288(.A(G29), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n712), .B2(new_n713), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G160), .B2(new_n697), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT98), .ZN(new_n717));
  INV_X1    g292(.A(G2084), .ZN(new_n718));
  NOR2_X1   g293(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n711), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n709), .A2(new_n710), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(KEYINPUT97), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(KEYINPUT99), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  NAND3_X1  g300(.A1(new_n720), .A2(KEYINPUT99), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  INV_X1    g302(.A(G16), .ZN(new_n728));
  NAND2_X1  g303(.A1(new_n728), .A2(G21), .ZN(new_n729));
  OAI21_X1  g304(.A(new_n729), .B1(G168), .B2(new_n728), .ZN(new_n730));
  NOR2_X1   g305(.A1(new_n730), .A2(G1966), .ZN(new_n731));
  XOR2_X1   g306(.A(new_n731), .B(KEYINPUT101), .Z(new_n732));
  NOR2_X1   g307(.A1(G27), .A2(G29), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G164), .B2(G29), .ZN(new_n734));
  INV_X1    g309(.A(G2078), .ZN(new_n735));
  XNOR2_X1  g310(.A(new_n734), .B(new_n735), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT31), .B(G11), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n737), .B(KEYINPUT100), .ZN(new_n738));
  INV_X1    g313(.A(G28), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n739), .A2(KEYINPUT30), .ZN(new_n740));
  AOI21_X1  g315(.A(G29), .B1(new_n739), .B2(KEYINPUT30), .ZN(new_n741));
  AOI21_X1  g316(.A(new_n738), .B1(new_n740), .B2(new_n741), .ZN(new_n742));
  OAI221_X1 g317(.A(new_n742), .B1(new_n697), .B2(new_n630), .C1(new_n699), .C2(new_n700), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(new_n717), .B2(new_n718), .ZN(new_n744));
  NOR2_X1   g319(.A1(G5), .A2(G16), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(KEYINPUT102), .ZN(new_n746));
  OAI21_X1  g321(.A(new_n746), .B1(G301), .B2(new_n728), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(KEYINPUT103), .ZN(new_n748));
  INV_X1    g323(.A(G1961), .ZN(new_n749));
  XNOR2_X1  g324(.A(new_n748), .B(new_n749), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n730), .A2(G1966), .ZN(new_n751));
  AND4_X1   g326(.A1(new_n736), .A2(new_n744), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NAND3_X1  g327(.A1(new_n727), .A2(new_n732), .A3(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT104), .ZN(new_n754));
  INV_X1    g329(.A(KEYINPUT104), .ZN(new_n755));
  NAND4_X1  g330(.A1(new_n727), .A2(new_n752), .A3(new_n755), .A4(new_n732), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n697), .A2(G35), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT105), .ZN(new_n758));
  OAI21_X1  g333(.A(new_n758), .B1(G162), .B2(new_n697), .ZN(new_n759));
  XOR2_X1   g334(.A(KEYINPUT29), .B(G2090), .Z(new_n760));
  XNOR2_X1  g335(.A(new_n759), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n697), .A2(G26), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT28), .Z(new_n763));
  AOI22_X1  g338(.A1(new_n485), .A2(G128), .B1(new_n487), .B2(G140), .ZN(new_n764));
  OAI221_X1 g339(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n481), .C2(G116), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AOI21_X1  g341(.A(new_n763), .B1(new_n766), .B2(G29), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G2067), .ZN(new_n768));
  NOR2_X1   g343(.A1(G4), .A2(G16), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(new_n606), .B2(G16), .ZN(new_n770));
  INV_X1    g345(.A(G1348), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n770), .B(new_n771), .ZN(new_n772));
  NAND3_X1  g347(.A1(new_n761), .A2(new_n768), .A3(new_n772), .ZN(new_n773));
  XOR2_X1   g348(.A(KEYINPUT89), .B(G16), .Z(new_n774));
  NAND2_X1  g349(.A1(new_n774), .A2(G20), .ZN(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(KEYINPUT23), .Z(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G299), .B2(G16), .ZN(new_n777));
  INV_X1    g352(.A(G1956), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n777), .B(new_n778), .ZN(new_n779));
  INV_X1    g354(.A(new_n774), .ZN(new_n780));
  NOR2_X1   g355(.A1(new_n780), .A2(G19), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n781), .B1(new_n548), .B2(new_n780), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(KEYINPUT95), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1341), .ZN(new_n784));
  NOR3_X1   g359(.A1(new_n773), .A2(new_n779), .A3(new_n784), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n754), .A2(new_n756), .A3(new_n785), .ZN(new_n786));
  INV_X1    g361(.A(KEYINPUT92), .ZN(new_n787));
  NAND2_X1  g362(.A1(G288), .A2(new_n787), .ZN(new_n788));
  NAND3_X1  g363(.A1(new_n579), .A2(KEYINPUT92), .A3(new_n580), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n728), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(new_n728), .B2(G23), .ZN(new_n791));
  XOR2_X1   g366(.A(KEYINPUT33), .B(G1976), .Z(new_n792));
  XNOR2_X1  g367(.A(new_n791), .B(new_n792), .ZN(new_n793));
  INV_X1    g368(.A(KEYINPUT93), .ZN(new_n794));
  XNOR2_X1  g369(.A(new_n793), .B(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n780), .A2(G22), .ZN(new_n796));
  AOI21_X1  g371(.A(new_n796), .B1(G166), .B2(new_n780), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT94), .B(G1971), .ZN(new_n798));
  XOR2_X1   g373(.A(new_n797), .B(new_n798), .Z(new_n799));
  XOR2_X1   g374(.A(KEYINPUT32), .B(G1981), .Z(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT91), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n728), .A2(G6), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(new_n591), .B2(new_n728), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT90), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n799), .B1(new_n801), .B2(new_n804), .ZN(new_n805));
  OR2_X1    g380(.A1(new_n804), .A2(new_n801), .ZN(new_n806));
  AND2_X1   g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n795), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n808), .A2(KEYINPUT34), .ZN(new_n809));
  INV_X1    g384(.A(KEYINPUT34), .ZN(new_n810));
  NAND3_X1  g385(.A1(new_n795), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  INV_X1    g386(.A(G25), .ZN(new_n812));
  OR3_X1    g387(.A1(new_n812), .A2(KEYINPUT86), .A3(G29), .ZN(new_n813));
  OAI21_X1  g388(.A(KEYINPUT86), .B1(new_n812), .B2(G29), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n487), .A2(G131), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT87), .ZN(new_n816));
  NOR2_X1   g391(.A1(G95), .A2(G2105), .ZN(new_n817));
  XOR2_X1   g392(.A(new_n817), .B(KEYINPUT88), .Z(new_n818));
  OAI211_X1 g393(.A(new_n818), .B(G2104), .C1(G107), .C2(new_n481), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n485), .A2(G119), .ZN(new_n820));
  AND3_X1   g395(.A1(new_n816), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  OAI211_X1 g396(.A(new_n813), .B(new_n814), .C1(new_n821), .C2(new_n697), .ZN(new_n822));
  XOR2_X1   g397(.A(KEYINPUT35), .B(G1991), .Z(new_n823));
  XOR2_X1   g398(.A(new_n822), .B(new_n823), .Z(new_n824));
  NOR2_X1   g399(.A1(new_n780), .A2(G24), .ZN(new_n825));
  AND3_X1   g400(.A1(new_n594), .A2(new_n595), .A3(new_n596), .ZN(new_n826));
  AOI21_X1  g401(.A(new_n825), .B1(new_n826), .B2(new_n780), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(G1986), .ZN(new_n828));
  NOR2_X1   g403(.A1(new_n824), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n809), .A2(new_n811), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n830), .A2(KEYINPUT36), .ZN(new_n831));
  INV_X1    g406(.A(KEYINPUT36), .ZN(new_n832));
  NAND4_X1  g407(.A1(new_n809), .A2(new_n811), .A3(new_n832), .A4(new_n829), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n786), .B1(new_n831), .B2(new_n833), .ZN(G311));
  NAND2_X1  g409(.A1(new_n831), .A2(new_n833), .ZN(new_n835));
  NAND4_X1  g410(.A1(new_n835), .A2(new_n754), .A3(new_n756), .A4(new_n785), .ZN(G150));
  NAND2_X1  g411(.A1(new_n606), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  XOR2_X1   g413(.A(KEYINPUT106), .B(G93), .Z(new_n839));
  NAND2_X1  g414(.A1(new_n533), .A2(new_n839), .ZN(new_n840));
  INV_X1    g415(.A(G67), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(new_n514), .B2(new_n515), .ZN(new_n842));
  AND2_X1   g417(.A1(G80), .A2(G543), .ZN(new_n843));
  OAI21_X1  g418(.A(G651), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n510), .A2(G55), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n840), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  OR2_X1    g421(.A1(new_n615), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n615), .A2(new_n846), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  XOR2_X1   g424(.A(new_n838), .B(new_n849), .Z(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  NOR2_X1   g426(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n852));
  NOR3_X1   g427(.A1(new_n851), .A2(new_n852), .A3(G860), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n846), .A2(G860), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n854), .B(KEYINPUT37), .ZN(new_n855));
  OR2_X1    g430(.A1(new_n853), .A2(new_n855), .ZN(G145));
  XOR2_X1   g431(.A(new_n821), .B(new_n622), .Z(new_n857));
  NAND2_X1  g432(.A1(new_n496), .A2(new_n500), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n766), .B(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(KEYINPUT107), .ZN(new_n861));
  OR3_X1    g436(.A1(new_n708), .A2(new_n696), .A3(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n485), .A2(G130), .ZN(new_n863));
  OAI221_X1 g438(.A(G2104), .B1(G106), .B2(G2105), .C1(new_n481), .C2(G118), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n487), .A2(G142), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n696), .B1(new_n708), .B2(new_n861), .ZN(new_n867));
  NAND3_X1  g442(.A1(new_n862), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n866), .B1(new_n862), .B2(new_n867), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n860), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g446(.A(new_n870), .ZN(new_n872));
  NAND3_X1  g447(.A1(new_n872), .A2(new_n859), .A3(new_n868), .ZN(new_n873));
  AOI21_X1  g448(.A(new_n857), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  INV_X1    g449(.A(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(KEYINPUT108), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n871), .A2(new_n873), .A3(new_n857), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n875), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(G162), .B(G160), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n879), .B(new_n630), .ZN(new_n880));
  AOI21_X1  g455(.A(G37), .B1(new_n878), .B2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n877), .A2(new_n876), .ZN(new_n882));
  OR3_X1    g457(.A1(new_n882), .A2(new_n880), .A3(new_n874), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n884), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g460(.A1(new_n846), .A2(new_n609), .ZN(new_n886));
  AOI22_X1  g461(.A1(new_n585), .A2(KEYINPUT79), .B1(G73), .B2(G543), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n506), .B1(new_n887), .B2(new_n588), .ZN(new_n888));
  OAI211_X1 g463(.A(new_n788), .B(new_n789), .C1(new_n888), .C2(new_n584), .ZN(new_n889));
  INV_X1    g464(.A(new_n789), .ZN(new_n890));
  AOI21_X1  g465(.A(KEYINPUT92), .B1(new_n579), .B2(new_n580), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n591), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n889), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(G303), .A2(new_n826), .ZN(new_n894));
  NAND2_X1  g469(.A1(G290), .A2(G166), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NAND4_X1  g472(.A1(new_n894), .A2(new_n889), .A3(new_n892), .A4(new_n895), .ZN(new_n898));
  AOI21_X1  g473(.A(KEYINPUT42), .B1(new_n897), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n897), .A2(KEYINPUT109), .A3(new_n898), .ZN(new_n900));
  AOI21_X1  g475(.A(KEYINPUT109), .B1(new_n897), .B2(new_n898), .ZN(new_n901));
  NOR2_X1   g476(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n899), .B1(new_n903), .B2(KEYINPUT42), .ZN(new_n904));
  INV_X1    g479(.A(new_n606), .ZN(new_n905));
  NOR2_X1   g480(.A1(G299), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n567), .B1(new_n566), .B2(new_n568), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n571), .A2(KEYINPUT77), .A3(new_n565), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n606), .B1(new_n909), .B2(new_n563), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n906), .A2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(KEYINPUT41), .B1(new_n906), .B2(new_n910), .ZN(new_n912));
  NAND2_X1  g487(.A1(G299), .A2(new_n905), .ZN(new_n913));
  INV_X1    g488(.A(KEYINPUT41), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n909), .A2(new_n606), .A3(new_n563), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n618), .B(new_n849), .ZN(new_n918));
  MUX2_X1   g493(.A(new_n911), .B(new_n917), .S(new_n918), .Z(new_n919));
  XNOR2_X1  g494(.A(new_n904), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n886), .B1(new_n920), .B2(new_n609), .ZN(G295));
  OAI21_X1  g496(.A(new_n886), .B1(new_n920), .B2(new_n609), .ZN(G331));
  INV_X1    g497(.A(KEYINPUT111), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT110), .ZN(new_n924));
  NAND2_X1  g499(.A1(G301), .A2(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(new_n925), .ZN(new_n926));
  NOR2_X1   g501(.A1(G301), .A2(new_n924), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n847), .B(new_n848), .C1(new_n926), .C2(new_n927), .ZN(new_n928));
  NAND2_X1  g503(.A1(G171), .A2(KEYINPUT110), .ZN(new_n929));
  AND2_X1   g504(.A1(new_n615), .A2(new_n846), .ZN(new_n930));
  NOR2_X1   g505(.A1(new_n615), .A2(new_n846), .ZN(new_n931));
  OAI211_X1 g506(.A(new_n925), .B(new_n929), .C1(new_n930), .C2(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(G168), .A2(new_n928), .A3(new_n932), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n928), .A2(new_n932), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(G286), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n917), .A2(new_n923), .A3(new_n933), .A4(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n933), .ZN(new_n937));
  AOI21_X1  g512(.A(G168), .B1(new_n928), .B2(new_n932), .ZN(new_n938));
  OAI21_X1  g513(.A(new_n911), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  AND2_X1   g514(.A1(new_n936), .A2(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n906), .A2(new_n910), .A3(KEYINPUT41), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n914), .B1(new_n913), .B2(new_n915), .ZN(new_n942));
  OAI211_X1 g517(.A(new_n935), .B(new_n933), .C1(new_n941), .C2(new_n942), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n940), .A2(KEYINPUT112), .A3(new_n902), .A4(new_n944), .ZN(new_n945));
  NAND4_X1  g520(.A1(new_n944), .A2(new_n902), .A3(new_n939), .A4(new_n936), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT112), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AND2_X1   g523(.A1(new_n943), .A2(KEYINPUT111), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n936), .A2(new_n939), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n903), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(G37), .ZN(new_n952));
  NAND4_X1  g527(.A1(new_n945), .A2(new_n948), .A3(new_n951), .A4(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT43), .ZN(new_n954));
  AND2_X1   g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(G37), .B1(new_n946), .B2(new_n947), .ZN(new_n956));
  NOR2_X1   g531(.A1(new_n917), .A2(KEYINPUT113), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT113), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n935), .B(new_n933), .C1(new_n912), .C2(new_n958), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n939), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n903), .ZN(new_n961));
  AND4_X1   g536(.A1(KEYINPUT43), .A2(new_n956), .A3(new_n945), .A4(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(KEYINPUT44), .B1(new_n955), .B2(new_n962), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n953), .A2(KEYINPUT43), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n956), .A2(new_n945), .A3(new_n954), .A4(new_n961), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT44), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n963), .A2(new_n968), .ZN(G397));
  INV_X1    g544(.A(G1384), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n858), .A2(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n470), .A2(new_n478), .A3(G40), .ZN(new_n974));
  NOR2_X1   g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(new_n821), .B(new_n823), .ZN(new_n976));
  INV_X1    g551(.A(G2067), .ZN(new_n977));
  XNOR2_X1  g552(.A(new_n766), .B(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(G1996), .ZN(new_n979));
  XNOR2_X1  g554(.A(new_n695), .B(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n976), .A2(new_n981), .ZN(new_n982));
  INV_X1    g557(.A(new_n982), .ZN(new_n983));
  XNOR2_X1  g558(.A(G290), .B(G1986), .ZN(new_n984));
  OAI21_X1  g559(.A(new_n975), .B1(new_n983), .B2(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n970), .B1(new_n501), .B2(new_n502), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(KEYINPUT50), .ZN(new_n987));
  INV_X1    g562(.A(G2090), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n481), .B1(new_n462), .B2(new_n463), .ZN(new_n989));
  INV_X1    g564(.A(G40), .ZN(new_n990));
  NOR3_X1   g565(.A1(new_n989), .A2(new_n477), .A3(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(G1384), .B1(new_n496), .B2(new_n500), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT50), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n992), .A2(new_n993), .ZN(new_n994));
  NAND4_X1  g569(.A1(new_n987), .A2(new_n988), .A3(new_n991), .A4(new_n994), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n974), .B1(KEYINPUT45), .B2(new_n992), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT71), .ZN(new_n997));
  INV_X1    g572(.A(G138), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n495), .B1(new_n475), .B2(new_n998), .ZN(new_n999));
  INV_X1    g574(.A(new_n492), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  INV_X1    g576(.A(new_n498), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n481), .A2(new_n1002), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n486), .B1(new_n1003), .B2(new_n497), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n997), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n496), .A2(new_n500), .A3(KEYINPUT71), .ZN(new_n1006));
  AOI21_X1  g581(.A(G1384), .B1(new_n1005), .B2(new_n1006), .ZN(new_n1007));
  OAI21_X1  g582(.A(new_n996), .B1(new_n1007), .B2(KEYINPUT45), .ZN(new_n1008));
  XNOR2_X1  g583(.A(KEYINPUT114), .B(G1971), .ZN(new_n1009));
  INV_X1    g584(.A(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1008), .A2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n995), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(G303), .A2(G8), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT55), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AND4_X1   g590(.A1(KEYINPUT115), .A2(new_n1012), .A3(G8), .A4(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(G8), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n995), .B2(new_n1011), .ZN(new_n1018));
  AOI21_X1  g593(.A(KEYINPUT115), .B1(new_n1018), .B2(new_n1015), .ZN(new_n1019));
  NOR2_X1   g594(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n788), .A2(G1976), .A3(new_n789), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1017), .B1(new_n992), .B2(new_n991), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1023), .A2(KEYINPUT52), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1021), .A2(new_n1022), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(new_n1022), .ZN(new_n1029));
  OAI21_X1  g604(.A(G1981), .B1(new_n888), .B2(KEYINPUT116), .ZN(new_n1030));
  XNOR2_X1  g605(.A(new_n1030), .B(new_n591), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT49), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  XNOR2_X1  g608(.A(G305), .B(new_n1030), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(KEYINPUT49), .ZN(new_n1035));
  AOI21_X1  g610(.A(new_n1028), .B1(new_n1033), .B2(new_n1035), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n974), .B1(new_n971), .B2(KEYINPUT50), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1037), .B1(new_n986), .B2(KEYINPUT50), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT117), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NAND2_X1  g615(.A1(new_n1007), .A2(new_n993), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1041), .A2(KEYINPUT117), .A3(new_n1037), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n988), .A3(new_n1042), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1017), .B1(new_n1043), .B2(new_n1011), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n1036), .B1(new_n1044), .B2(new_n1015), .ZN(new_n1045));
  NOR2_X1   g620(.A1(new_n1020), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(KEYINPUT45), .B(new_n970), .C1(new_n501), .C2(new_n502), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n974), .B1(new_n971), .B2(new_n972), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(KEYINPUT122), .B1(new_n1049), .B2(G2078), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT122), .ZN(new_n1051));
  NAND4_X1  g626(.A1(new_n1047), .A2(new_n1048), .A3(new_n1051), .A4(new_n735), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1052), .A3(KEYINPUT53), .ZN(new_n1053));
  INV_X1    g628(.A(KEYINPUT53), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n735), .B(new_n996), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n991), .B(new_n994), .C1(new_n1007), .C2(new_n993), .ZN(new_n1056));
  AOI22_X1  g631(.A1(new_n1054), .A2(new_n1055), .B1(new_n1056), .B2(new_n749), .ZN(new_n1057));
  AOI21_X1  g632(.A(G301), .B1(new_n1053), .B2(new_n1057), .ZN(new_n1058));
  INV_X1    g633(.A(G1966), .ZN(new_n1059));
  NAND2_X1  g634(.A1(new_n1049), .A2(new_n1059), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n974), .A2(G2084), .ZN(new_n1061));
  OAI211_X1 g636(.A(new_n994), .B(new_n1061), .C1(new_n1007), .C2(new_n993), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1060), .A2(G168), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(G8), .ZN(new_n1064));
  AOI21_X1  g639(.A(G168), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1065));
  OAI21_X1  g640(.A(KEYINPUT51), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT62), .ZN(new_n1067));
  INV_X1    g642(.A(new_n994), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1068), .B1(KEYINPUT50), .B2(new_n986), .ZN(new_n1069));
  AOI22_X1  g644(.A1(new_n1069), .A2(new_n1061), .B1(new_n1049), .B2(new_n1059), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n1017), .B1(new_n1070), .B2(G168), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT51), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g648(.A1(new_n1066), .A2(new_n1067), .A3(new_n1073), .ZN(new_n1074));
  INV_X1    g649(.A(new_n1065), .ZN(new_n1075));
  AOI21_X1  g650(.A(new_n1072), .B1(new_n1071), .B2(new_n1075), .ZN(new_n1076));
  NOR2_X1   g651(.A1(new_n1064), .A2(KEYINPUT51), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT62), .B1(new_n1076), .B2(new_n1077), .ZN(new_n1078));
  NAND4_X1  g653(.A1(new_n1046), .A2(new_n1058), .A3(new_n1074), .A4(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1033), .A2(new_n1035), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1080), .A2(new_n1025), .A3(new_n580), .A4(new_n579), .ZN(new_n1081));
  OAI21_X1  g656(.A(new_n1081), .B1(G1981), .B2(G305), .ZN(new_n1082));
  AOI22_X1  g657(.A1(new_n1082), .A2(new_n1022), .B1(new_n1020), .B2(new_n1036), .ZN(new_n1083));
  NAND2_X1  g658(.A1(G299), .A2(KEYINPUT57), .ZN(new_n1084));
  AOI21_X1  g659(.A(KEYINPUT57), .B1(new_n571), .B2(new_n565), .ZN(new_n1085));
  NAND2_X1  g660(.A1(new_n563), .A2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  OAI211_X1 g663(.A(new_n996), .B(new_n1088), .C1(new_n1007), .C2(KEYINPUT45), .ZN(new_n1089));
  INV_X1    g664(.A(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(G1956), .B1(new_n1041), .B2(new_n1037), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1087), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n992), .A2(new_n991), .A3(KEYINPUT118), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1093), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT118), .B1(new_n992), .B2(new_n991), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n977), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT119), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1096), .A2(new_n1097), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1056), .A2(new_n771), .ZN(new_n1099));
  OAI211_X1 g674(.A(KEYINPUT119), .B(new_n977), .C1(new_n1094), .C2(new_n1095), .ZN(new_n1100));
  NAND3_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1101), .A2(new_n606), .ZN(new_n1102));
  NOR3_X1   g677(.A1(new_n1090), .A2(new_n1091), .A3(new_n1087), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1092), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1038), .A2(new_n778), .ZN(new_n1105));
  AOI22_X1  g680(.A1(G299), .A2(KEYINPUT57), .B1(new_n563), .B2(new_n1085), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1105), .A2(new_n1106), .A3(new_n1089), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n1092), .A2(new_n1107), .A3(KEYINPUT61), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1095), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT58), .B(G1341), .Z(new_n1110));
  NAND3_X1  g685(.A1(new_n1109), .A2(new_n1093), .A3(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1111), .B1(new_n1008), .B2(G1996), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(new_n548), .ZN(new_n1113));
  XOR2_X1   g688(.A(KEYINPUT120), .B(KEYINPUT59), .Z(new_n1114));
  NAND2_X1  g689(.A1(new_n1113), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT60), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n606), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n1098), .A2(new_n1099), .A3(new_n1100), .A4(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1114), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1112), .A2(new_n548), .A3(new_n1120), .ZN(new_n1121));
  NAND4_X1  g696(.A1(new_n1108), .A2(new_n1115), .A3(new_n1119), .A4(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1098), .A2(new_n1099), .A3(new_n905), .A4(new_n1100), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1116), .B1(new_n1102), .B2(new_n1123), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1122), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT61), .ZN(new_n1126));
  AOI21_X1  g701(.A(new_n1106), .B1(new_n1105), .B2(new_n1089), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1126), .B1(new_n1103), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(KEYINPUT121), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  OAI211_X1 g705(.A(KEYINPUT121), .B(new_n1126), .C1(new_n1103), .C2(new_n1127), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1130), .A2(new_n1131), .ZN(new_n1132));
  AOI21_X1  g707(.A(new_n1104), .B1(new_n1125), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT54), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1055), .A2(new_n1054), .ZN(new_n1135));
  NAND2_X1  g710(.A1(new_n1056), .A2(new_n749), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n992), .A2(KEYINPUT45), .ZN(new_n1137));
  XOR2_X1   g712(.A(new_n477), .B(KEYINPUT123), .Z(new_n1138));
  OAI211_X1 g713(.A(KEYINPUT53), .B(G40), .C1(KEYINPUT124), .C2(G2078), .ZN(new_n1139));
  AOI211_X1 g714(.A(new_n1139), .B(new_n989), .C1(KEYINPUT124), .C2(G2078), .ZN(new_n1140));
  NAND4_X1  g715(.A1(new_n973), .A2(new_n1137), .A3(new_n1138), .A4(new_n1140), .ZN(new_n1141));
  NAND4_X1  g716(.A1(new_n1135), .A2(new_n1136), .A3(G301), .A4(new_n1141), .ZN(new_n1142));
  INV_X1    g717(.A(KEYINPUT125), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g719(.A1(new_n1057), .A2(KEYINPUT125), .A3(G301), .A4(new_n1141), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g721(.A(new_n1134), .B1(new_n1146), .B2(new_n1058), .ZN(new_n1147));
  NAND3_X1  g722(.A1(new_n1135), .A2(new_n1136), .A3(new_n1141), .ZN(new_n1148));
  AOI21_X1  g723(.A(new_n1134), .B1(new_n1148), .B2(G171), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1053), .A2(G301), .A3(new_n1057), .ZN(new_n1150));
  AOI22_X1  g725(.A1(new_n1066), .A2(new_n1073), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g726(.A(new_n1045), .ZN(new_n1152));
  OR2_X1    g727(.A1(new_n1016), .A2(new_n1019), .ZN(new_n1153));
  NAND4_X1  g728(.A1(new_n1147), .A2(new_n1151), .A3(new_n1152), .A4(new_n1153), .ZN(new_n1154));
  OAI211_X1 g729(.A(new_n1079), .B(new_n1083), .C1(new_n1133), .C2(new_n1154), .ZN(new_n1155));
  NOR3_X1   g730(.A1(new_n1070), .A2(new_n1017), .A3(G286), .ZN(new_n1156));
  NAND2_X1  g731(.A1(new_n1046), .A2(new_n1156), .ZN(new_n1157));
  INV_X1    g732(.A(KEYINPUT63), .ZN(new_n1158));
  NAND3_X1  g733(.A1(new_n1036), .A2(new_n1156), .A3(KEYINPUT63), .ZN(new_n1159));
  INV_X1    g734(.A(new_n1018), .ZN(new_n1160));
  AOI21_X1  g735(.A(new_n1159), .B1(new_n1014), .B2(new_n1160), .ZN(new_n1161));
  AOI22_X1  g736(.A1(new_n1157), .A2(new_n1158), .B1(new_n1153), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(new_n985), .B1(new_n1155), .B2(new_n1162), .ZN(new_n1163));
  INV_X1    g738(.A(new_n975), .ZN(new_n1164));
  OR3_X1    g739(.A1(new_n1164), .A2(G1986), .A3(G290), .ZN(new_n1165));
  INV_X1    g740(.A(KEYINPUT48), .ZN(new_n1166));
  OAI22_X1  g741(.A1(new_n982), .A2(new_n1164), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  AOI21_X1  g742(.A(new_n1167), .B1(new_n1166), .B2(new_n1165), .ZN(new_n1168));
  AOI21_X1  g743(.A(KEYINPUT46), .B1(new_n975), .B2(new_n979), .ZN(new_n1169));
  INV_X1    g744(.A(KEYINPUT126), .ZN(new_n1170));
  AND2_X1   g745(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1171));
  NOR2_X1   g746(.A1(new_n1169), .A2(new_n1170), .ZN(new_n1172));
  AOI21_X1  g747(.A(new_n695), .B1(KEYINPUT46), .B2(new_n979), .ZN(new_n1173));
  AND2_X1   g748(.A1(new_n978), .A2(new_n1173), .ZN(new_n1174));
  OAI22_X1  g749(.A1(new_n1171), .A2(new_n1172), .B1(new_n1164), .B2(new_n1174), .ZN(new_n1175));
  XOR2_X1   g750(.A(new_n1175), .B(KEYINPUT47), .Z(new_n1176));
  NAND2_X1  g751(.A1(new_n821), .A2(new_n823), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n981), .A2(new_n1177), .B1(G2067), .B2(new_n766), .ZN(new_n1178));
  AOI211_X1 g753(.A(new_n1168), .B(new_n1176), .C1(new_n975), .C2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g754(.A1(new_n1163), .A2(new_n1179), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g755(.A1(G227), .A2(G401), .A3(new_n459), .ZN(new_n1182));
  OAI21_X1  g756(.A(new_n1182), .B1(new_n688), .B2(new_n689), .ZN(new_n1183));
  NAND2_X1  g757(.A1(new_n1183), .A2(KEYINPUT127), .ZN(new_n1184));
  INV_X1    g758(.A(KEYINPUT127), .ZN(new_n1185));
  OAI211_X1 g759(.A(new_n1185), .B(new_n1182), .C1(new_n688), .C2(new_n689), .ZN(new_n1186));
  AOI22_X1  g760(.A1(new_n881), .A2(new_n883), .B1(new_n1184), .B2(new_n1186), .ZN(new_n1187));
  NAND2_X1  g761(.A1(new_n1187), .A2(new_n966), .ZN(G225));
  INV_X1    g762(.A(G225), .ZN(G308));
endmodule


