

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U546 ( .A1(G651), .A2(n562), .ZN(n787) );
  AND2_X1 U547 ( .A1(n522), .A2(G2105), .ZN(n881) );
  NAND2_X1 U548 ( .A1(n877), .A2(G101), .ZN(n526) );
  OR2_X1 U549 ( .A1(G301), .A2(n646), .ZN(n513) );
  XOR2_X1 U550 ( .A(KEYINPUT84), .B(n519), .Z(n514) );
  OR2_X1 U551 ( .A1(n689), .A2(n688), .ZN(n515) );
  XOR2_X1 U552 ( .A(n649), .B(KEYINPUT31), .Z(n516) );
  INV_X1 U553 ( .A(KEYINPUT29), .ZN(n636) );
  AND2_X1 U554 ( .A1(n690), .A2(n515), .ZN(n691) );
  NAND2_X1 U555 ( .A1(G160), .A2(G40), .ZN(n693) );
  NOR2_X1 U556 ( .A1(G164), .A2(G1384), .ZN(n694) );
  NOR2_X2 U557 ( .A1(G2105), .A2(n522), .ZN(n877) );
  XOR2_X1 U558 ( .A(KEYINPUT15), .B(n622), .Z(n894) );
  NOR2_X1 U559 ( .A1(n525), .A2(n524), .ZN(G164) );
  INV_X1 U560 ( .A(G2104), .ZN(n522) );
  NAND2_X1 U561 ( .A1(G126), .A2(n881), .ZN(n518) );
  AND2_X1 U562 ( .A1(G2104), .A2(G2105), .ZN(n882) );
  NAND2_X1 U563 ( .A1(G114), .A2(n882), .ZN(n517) );
  NAND2_X1 U564 ( .A1(n518), .A2(n517), .ZN(n519) );
  NOR2_X1 U565 ( .A1(G2104), .A2(G2105), .ZN(n520) );
  XOR2_X2 U566 ( .A(KEYINPUT17), .B(n520), .Z(n878) );
  NAND2_X1 U567 ( .A1(n878), .A2(G138), .ZN(n521) );
  NAND2_X1 U568 ( .A1(n514), .A2(n521), .ZN(n525) );
  NAND2_X1 U569 ( .A1(G102), .A2(n877), .ZN(n523) );
  XNOR2_X1 U570 ( .A(KEYINPUT85), .B(n523), .ZN(n524) );
  XOR2_X1 U571 ( .A(n526), .B(KEYINPUT23), .Z(n528) );
  NAND2_X1 U572 ( .A1(n881), .A2(G125), .ZN(n527) );
  NAND2_X1 U573 ( .A1(n528), .A2(n527), .ZN(n529) );
  XNOR2_X1 U574 ( .A(n529), .B(KEYINPUT64), .ZN(n533) );
  NAND2_X1 U575 ( .A1(G113), .A2(n882), .ZN(n531) );
  NAND2_X1 U576 ( .A1(G137), .A2(n878), .ZN(n530) );
  NAND2_X1 U577 ( .A1(n531), .A2(n530), .ZN(n532) );
  NOR2_X2 U578 ( .A1(n533), .A2(n532), .ZN(G160) );
  XOR2_X1 U579 ( .A(G543), .B(KEYINPUT0), .Z(n562) );
  NAND2_X1 U580 ( .A1(G52), .A2(n787), .ZN(n536) );
  INV_X1 U581 ( .A(G651), .ZN(n537) );
  NOR2_X1 U582 ( .A1(G543), .A2(n537), .ZN(n534) );
  XOR2_X1 U583 ( .A(KEYINPUT1), .B(n534), .Z(n789) );
  NAND2_X1 U584 ( .A1(G64), .A2(n789), .ZN(n535) );
  NAND2_X1 U585 ( .A1(n536), .A2(n535), .ZN(n543) );
  NOR2_X2 U586 ( .A1(n562), .A2(n537), .ZN(n783) );
  NAND2_X1 U587 ( .A1(n783), .A2(G77), .ZN(n538) );
  XNOR2_X1 U588 ( .A(n538), .B(KEYINPUT66), .ZN(n540) );
  NOR2_X1 U589 ( .A1(G651), .A2(G543), .ZN(n784) );
  NAND2_X1 U590 ( .A1(G90), .A2(n784), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XOR2_X1 U592 ( .A(KEYINPUT9), .B(n541), .Z(n542) );
  NOR2_X1 U593 ( .A1(n543), .A2(n542), .ZN(G171) );
  INV_X1 U594 ( .A(G171), .ZN(G301) );
  XNOR2_X1 U595 ( .A(KEYINPUT72), .B(KEYINPUT7), .ZN(n555) );
  NAND2_X1 U596 ( .A1(n784), .A2(G89), .ZN(n544) );
  XNOR2_X1 U597 ( .A(n544), .B(KEYINPUT4), .ZN(n546) );
  NAND2_X1 U598 ( .A1(G76), .A2(n783), .ZN(n545) );
  NAND2_X1 U599 ( .A1(n546), .A2(n545), .ZN(n547) );
  XNOR2_X1 U600 ( .A(KEYINPUT5), .B(n547), .ZN(n553) );
  NAND2_X1 U601 ( .A1(n787), .A2(G51), .ZN(n548) );
  XOR2_X1 U602 ( .A(KEYINPUT71), .B(n548), .Z(n550) );
  NAND2_X1 U603 ( .A1(n789), .A2(G63), .ZN(n549) );
  NAND2_X1 U604 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U605 ( .A(KEYINPUT6), .B(n551), .Z(n552) );
  NAND2_X1 U606 ( .A1(n553), .A2(n552), .ZN(n554) );
  XNOR2_X1 U607 ( .A(n555), .B(n554), .ZN(G168) );
  XOR2_X1 U608 ( .A(KEYINPUT8), .B(G168), .Z(G286) );
  NAND2_X1 U609 ( .A1(G75), .A2(n783), .ZN(n557) );
  NAND2_X1 U610 ( .A1(G88), .A2(n784), .ZN(n556) );
  NAND2_X1 U611 ( .A1(n557), .A2(n556), .ZN(n561) );
  NAND2_X1 U612 ( .A1(G50), .A2(n787), .ZN(n559) );
  NAND2_X1 U613 ( .A1(G62), .A2(n789), .ZN(n558) );
  NAND2_X1 U614 ( .A1(n559), .A2(n558), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n561), .A2(n560), .ZN(G166) );
  NAND2_X1 U616 ( .A1(n562), .A2(G87), .ZN(n567) );
  NAND2_X1 U617 ( .A1(G49), .A2(n787), .ZN(n564) );
  NAND2_X1 U618 ( .A1(G74), .A2(G651), .ZN(n563) );
  NAND2_X1 U619 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U620 ( .A1(n789), .A2(n565), .ZN(n566) );
  NAND2_X1 U621 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U622 ( .A(KEYINPUT75), .B(n568), .Z(G288) );
  INV_X1 U623 ( .A(G166), .ZN(G303) );
  NAND2_X1 U624 ( .A1(G48), .A2(n787), .ZN(n577) );
  XOR2_X1 U625 ( .A(KEYINPUT76), .B(KEYINPUT2), .Z(n570) );
  NAND2_X1 U626 ( .A1(G73), .A2(n783), .ZN(n569) );
  XNOR2_X1 U627 ( .A(n570), .B(n569), .ZN(n574) );
  NAND2_X1 U628 ( .A1(G86), .A2(n784), .ZN(n572) );
  NAND2_X1 U629 ( .A1(G61), .A2(n789), .ZN(n571) );
  NAND2_X1 U630 ( .A1(n572), .A2(n571), .ZN(n573) );
  NOR2_X1 U631 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U632 ( .A(KEYINPUT77), .B(n575), .Z(n576) );
  NAND2_X1 U633 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U634 ( .A(n578), .B(KEYINPUT78), .ZN(G305) );
  NAND2_X1 U635 ( .A1(G72), .A2(n783), .ZN(n580) );
  NAND2_X1 U636 ( .A1(G85), .A2(n784), .ZN(n579) );
  NAND2_X1 U637 ( .A1(n580), .A2(n579), .ZN(n583) );
  NAND2_X1 U638 ( .A1(G60), .A2(n789), .ZN(n581) );
  XNOR2_X1 U639 ( .A(KEYINPUT65), .B(n581), .ZN(n582) );
  NOR2_X1 U640 ( .A1(n583), .A2(n582), .ZN(n585) );
  NAND2_X1 U641 ( .A1(n787), .A2(G47), .ZN(n584) );
  NAND2_X1 U642 ( .A1(n585), .A2(n584), .ZN(G290) );
  INV_X1 U643 ( .A(n693), .ZN(n586) );
  NAND2_X2 U644 ( .A1(n586), .A2(n694), .ZN(n658) );
  NOR2_X1 U645 ( .A1(G2084), .A2(n658), .ZN(n642) );
  NAND2_X1 U646 ( .A1(n642), .A2(G8), .ZN(n655) );
  NAND2_X1 U647 ( .A1(G8), .A2(n658), .ZN(n689) );
  NOR2_X1 U648 ( .A1(G1966), .A2(n689), .ZN(n653) );
  INV_X1 U649 ( .A(KEYINPUT100), .ZN(n651) );
  NAND2_X1 U650 ( .A1(G53), .A2(n787), .ZN(n588) );
  NAND2_X1 U651 ( .A1(G65), .A2(n789), .ZN(n587) );
  NAND2_X1 U652 ( .A1(n588), .A2(n587), .ZN(n592) );
  NAND2_X1 U653 ( .A1(G78), .A2(n783), .ZN(n590) );
  NAND2_X1 U654 ( .A1(G91), .A2(n784), .ZN(n589) );
  NAND2_X1 U655 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U656 ( .A1(n592), .A2(n591), .ZN(n798) );
  INV_X1 U657 ( .A(n658), .ZN(n638) );
  NAND2_X1 U658 ( .A1(n638), .A2(G2072), .ZN(n593) );
  XNOR2_X1 U659 ( .A(n593), .B(KEYINPUT27), .ZN(n596) );
  NAND2_X1 U660 ( .A1(G1956), .A2(n658), .ZN(n594) );
  XNOR2_X1 U661 ( .A(KEYINPUT97), .B(n594), .ZN(n595) );
  NOR2_X1 U662 ( .A1(n596), .A2(n595), .ZN(n597) );
  XNOR2_X1 U663 ( .A(n597), .B(KEYINPUT98), .ZN(n631) );
  NOR2_X1 U664 ( .A1(n798), .A2(n631), .ZN(n599) );
  INV_X1 U665 ( .A(KEYINPUT28), .ZN(n598) );
  XNOR2_X1 U666 ( .A(n599), .B(n598), .ZN(n635) );
  INV_X1 U667 ( .A(G1996), .ZN(n741) );
  NOR2_X1 U668 ( .A1(n658), .A2(n741), .ZN(n600) );
  XNOR2_X1 U669 ( .A(n600), .B(KEYINPUT26), .ZN(n613) );
  NAND2_X1 U670 ( .A1(n658), .A2(G1341), .ZN(n611) );
  NAND2_X1 U671 ( .A1(G56), .A2(n789), .ZN(n601) );
  XOR2_X1 U672 ( .A(KEYINPUT14), .B(n601), .Z(n607) );
  NAND2_X1 U673 ( .A1(n784), .A2(G81), .ZN(n602) );
  XNOR2_X1 U674 ( .A(n602), .B(KEYINPUT12), .ZN(n604) );
  NAND2_X1 U675 ( .A1(G68), .A2(n783), .ZN(n603) );
  NAND2_X1 U676 ( .A1(n604), .A2(n603), .ZN(n605) );
  XOR2_X1 U677 ( .A(KEYINPUT13), .B(n605), .Z(n606) );
  NOR2_X1 U678 ( .A1(n607), .A2(n606), .ZN(n609) );
  NAND2_X1 U679 ( .A1(n787), .A2(G43), .ZN(n608) );
  NAND2_X1 U680 ( .A1(n609), .A2(n608), .ZN(n922) );
  INV_X1 U681 ( .A(n922), .ZN(n610) );
  NAND2_X1 U682 ( .A1(n611), .A2(n610), .ZN(n612) );
  NOR2_X1 U683 ( .A1(n613), .A2(n612), .ZN(n628) );
  NAND2_X1 U684 ( .A1(n783), .A2(G79), .ZN(n614) );
  XOR2_X1 U685 ( .A(KEYINPUT69), .B(n614), .Z(n616) );
  NAND2_X1 U686 ( .A1(n787), .A2(G54), .ZN(n615) );
  NAND2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n617) );
  XNOR2_X1 U688 ( .A(n617), .B(KEYINPUT70), .ZN(n621) );
  NAND2_X1 U689 ( .A1(G92), .A2(n784), .ZN(n619) );
  NAND2_X1 U690 ( .A1(G66), .A2(n789), .ZN(n618) );
  NAND2_X1 U691 ( .A1(n619), .A2(n618), .ZN(n620) );
  NOR2_X1 U692 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U693 ( .A1(n628), .A2(n894), .ZN(n626) );
  NOR2_X1 U694 ( .A1(n638), .A2(G1348), .ZN(n624) );
  NOR2_X1 U695 ( .A1(G2067), .A2(n658), .ZN(n623) );
  NOR2_X1 U696 ( .A1(n624), .A2(n623), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n626), .A2(n625), .ZN(n627) );
  XOR2_X1 U698 ( .A(KEYINPUT99), .B(n627), .Z(n630) );
  OR2_X1 U699 ( .A1(n894), .A2(n628), .ZN(n629) );
  NAND2_X1 U700 ( .A1(n630), .A2(n629), .ZN(n633) );
  NAND2_X1 U701 ( .A1(n798), .A2(n631), .ZN(n632) );
  NAND2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n634) );
  NAND2_X1 U703 ( .A1(n635), .A2(n634), .ZN(n637) );
  XNOR2_X1 U704 ( .A(n637), .B(n636), .ZN(n641) );
  XOR2_X1 U705 ( .A(KEYINPUT25), .B(G2078), .Z(n964) );
  NOR2_X1 U706 ( .A1(n964), .A2(n658), .ZN(n640) );
  NOR2_X1 U707 ( .A1(n638), .A2(G1961), .ZN(n639) );
  NOR2_X1 U708 ( .A1(n640), .A2(n639), .ZN(n646) );
  NAND2_X1 U709 ( .A1(n641), .A2(n513), .ZN(n650) );
  NOR2_X1 U710 ( .A1(n653), .A2(n642), .ZN(n643) );
  NAND2_X1 U711 ( .A1(G8), .A2(n643), .ZN(n644) );
  XNOR2_X1 U712 ( .A(KEYINPUT30), .B(n644), .ZN(n645) );
  NOR2_X1 U713 ( .A1(G168), .A2(n645), .ZN(n648) );
  AND2_X1 U714 ( .A1(G301), .A2(n646), .ZN(n647) );
  NOR2_X1 U715 ( .A1(n648), .A2(n647), .ZN(n649) );
  NAND2_X1 U716 ( .A1(n650), .A2(n516), .ZN(n656) );
  XNOR2_X1 U717 ( .A(n651), .B(n656), .ZN(n652) );
  NOR2_X1 U718 ( .A1(n653), .A2(n652), .ZN(n654) );
  NAND2_X1 U719 ( .A1(n655), .A2(n654), .ZN(n668) );
  NAND2_X1 U720 ( .A1(n656), .A2(G286), .ZN(n663) );
  NOR2_X1 U721 ( .A1(G1971), .A2(n689), .ZN(n657) );
  XNOR2_X1 U722 ( .A(KEYINPUT101), .B(n657), .ZN(n661) );
  NOR2_X1 U723 ( .A1(G2090), .A2(n658), .ZN(n659) );
  NOR2_X1 U724 ( .A1(G166), .A2(n659), .ZN(n660) );
  NAND2_X1 U725 ( .A1(n661), .A2(n660), .ZN(n662) );
  NAND2_X1 U726 ( .A1(n663), .A2(n662), .ZN(n664) );
  NAND2_X1 U727 ( .A1(n664), .A2(G8), .ZN(n666) );
  XNOR2_X1 U728 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n665) );
  XNOR2_X1 U729 ( .A(n666), .B(n665), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n668), .A2(n667), .ZN(n685) );
  NOR2_X1 U731 ( .A1(G1976), .A2(G288), .ZN(n908) );
  NOR2_X1 U732 ( .A1(G1971), .A2(G303), .ZN(n669) );
  XOR2_X1 U733 ( .A(n669), .B(KEYINPUT103), .Z(n670) );
  NOR2_X1 U734 ( .A1(n908), .A2(n670), .ZN(n671) );
  NAND2_X1 U735 ( .A1(n685), .A2(n671), .ZN(n674) );
  NAND2_X1 U736 ( .A1(G1976), .A2(G288), .ZN(n909) );
  INV_X1 U737 ( .A(n689), .ZN(n672) );
  AND2_X1 U738 ( .A1(n909), .A2(n672), .ZN(n673) );
  AND2_X1 U739 ( .A1(n674), .A2(n673), .ZN(n675) );
  NOR2_X1 U740 ( .A1(n675), .A2(KEYINPUT33), .ZN(n678) );
  NAND2_X1 U741 ( .A1(n908), .A2(KEYINPUT33), .ZN(n676) );
  NOR2_X1 U742 ( .A1(n676), .A2(n689), .ZN(n677) );
  NOR2_X1 U743 ( .A1(n678), .A2(n677), .ZN(n680) );
  XOR2_X1 U744 ( .A(G1981), .B(G305), .Z(n679) );
  XNOR2_X1 U745 ( .A(KEYINPUT104), .B(n679), .ZN(n917) );
  NAND2_X1 U746 ( .A1(n680), .A2(n917), .ZN(n681) );
  XNOR2_X1 U747 ( .A(n681), .B(KEYINPUT105), .ZN(n682) );
  INV_X1 U748 ( .A(n682), .ZN(n692) );
  NOR2_X1 U749 ( .A1(G2090), .A2(G303), .ZN(n683) );
  NAND2_X1 U750 ( .A1(G8), .A2(n683), .ZN(n684) );
  NAND2_X1 U751 ( .A1(n685), .A2(n684), .ZN(n686) );
  NAND2_X1 U752 ( .A1(n686), .A2(n689), .ZN(n690) );
  NOR2_X1 U753 ( .A1(G1981), .A2(G305), .ZN(n687) );
  XOR2_X1 U754 ( .A(n687), .B(KEYINPUT24), .Z(n688) );
  NAND2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n733) );
  NOR2_X1 U756 ( .A1(n694), .A2(n693), .ZN(n748) );
  XNOR2_X1 U757 ( .A(G2067), .B(KEYINPUT37), .ZN(n735) );
  NAND2_X1 U758 ( .A1(n881), .A2(G128), .ZN(n695) );
  XOR2_X1 U759 ( .A(KEYINPUT89), .B(n695), .Z(n697) );
  NAND2_X1 U760 ( .A1(n882), .A2(G116), .ZN(n696) );
  NAND2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  XOR2_X1 U762 ( .A(KEYINPUT35), .B(n698), .Z(n705) );
  XOR2_X1 U763 ( .A(KEYINPUT88), .B(KEYINPUT34), .Z(n703) );
  NAND2_X1 U764 ( .A1(n878), .A2(G140), .ZN(n699) );
  XOR2_X1 U765 ( .A(KEYINPUT87), .B(n699), .Z(n701) );
  NAND2_X1 U766 ( .A1(n877), .A2(G104), .ZN(n700) );
  NAND2_X1 U767 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U768 ( .A(n703), .B(n702), .Z(n704) );
  NOR2_X1 U769 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U770 ( .A(KEYINPUT36), .B(n706), .ZN(n890) );
  NOR2_X1 U771 ( .A1(n735), .A2(n890), .ZN(n988) );
  NAND2_X1 U772 ( .A1(n748), .A2(n988), .ZN(n744) );
  NAND2_X1 U773 ( .A1(n882), .A2(G117), .ZN(n707) );
  XNOR2_X1 U774 ( .A(KEYINPUT92), .B(n707), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n881), .A2(G129), .ZN(n708) );
  XOR2_X1 U776 ( .A(KEYINPUT91), .B(n708), .Z(n709) );
  NAND2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(KEYINPUT93), .ZN(n713) );
  NAND2_X1 U779 ( .A1(G141), .A2(n878), .ZN(n712) );
  NAND2_X1 U780 ( .A1(n713), .A2(n712), .ZN(n717) );
  XOR2_X1 U781 ( .A(KEYINPUT94), .B(KEYINPUT38), .Z(n715) );
  NAND2_X1 U782 ( .A1(G105), .A2(n877), .ZN(n714) );
  XNOR2_X1 U783 ( .A(n715), .B(n714), .ZN(n716) );
  NOR2_X1 U784 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U785 ( .A(n718), .B(KEYINPUT95), .Z(n873) );
  OR2_X1 U786 ( .A1(n741), .A2(n873), .ZN(n727) );
  NAND2_X1 U787 ( .A1(G95), .A2(n877), .ZN(n720) );
  NAND2_X1 U788 ( .A1(G131), .A2(n878), .ZN(n719) );
  NAND2_X1 U789 ( .A1(n720), .A2(n719), .ZN(n721) );
  XOR2_X1 U790 ( .A(KEYINPUT90), .B(n721), .Z(n725) );
  NAND2_X1 U791 ( .A1(G119), .A2(n881), .ZN(n723) );
  NAND2_X1 U792 ( .A1(G107), .A2(n882), .ZN(n722) );
  AND2_X1 U793 ( .A1(n723), .A2(n722), .ZN(n724) );
  NAND2_X1 U794 ( .A1(n725), .A2(n724), .ZN(n872) );
  NAND2_X1 U795 ( .A1(G1991), .A2(n872), .ZN(n726) );
  NAND2_X1 U796 ( .A1(n727), .A2(n726), .ZN(n1000) );
  NAND2_X1 U797 ( .A1(n748), .A2(n1000), .ZN(n739) );
  NAND2_X1 U798 ( .A1(n744), .A2(n739), .ZN(n728) );
  XNOR2_X1 U799 ( .A(KEYINPUT96), .B(n728), .ZN(n731) );
  XNOR2_X1 U800 ( .A(G1986), .B(G290), .ZN(n924) );
  NAND2_X1 U801 ( .A1(n748), .A2(n924), .ZN(n729) );
  XOR2_X1 U802 ( .A(KEYINPUT86), .B(n729), .Z(n730) );
  NOR2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U804 ( .A1(n733), .A2(n732), .ZN(n734) );
  XNOR2_X1 U805 ( .A(n734), .B(KEYINPUT106), .ZN(n750) );
  NAND2_X1 U806 ( .A1(n890), .A2(n735), .ZN(n736) );
  XNOR2_X1 U807 ( .A(n736), .B(KEYINPUT108), .ZN(n985) );
  NOR2_X1 U808 ( .A1(G1986), .A2(G290), .ZN(n737) );
  NOR2_X1 U809 ( .A1(G1991), .A2(n872), .ZN(n990) );
  NOR2_X1 U810 ( .A1(n737), .A2(n990), .ZN(n738) );
  XNOR2_X1 U811 ( .A(KEYINPUT107), .B(n738), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n740), .A2(n739), .ZN(n742) );
  NAND2_X1 U813 ( .A1(n873), .A2(n741), .ZN(n981) );
  NAND2_X1 U814 ( .A1(n742), .A2(n981), .ZN(n743) );
  XOR2_X1 U815 ( .A(KEYINPUT39), .B(n743), .Z(n745) );
  NAND2_X1 U816 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U817 ( .A1(n985), .A2(n746), .ZN(n747) );
  NAND2_X1 U818 ( .A1(n748), .A2(n747), .ZN(n749) );
  NAND2_X1 U819 ( .A1(n750), .A2(n749), .ZN(n751) );
  XNOR2_X1 U820 ( .A(n751), .B(KEYINPUT40), .ZN(G329) );
  XOR2_X1 U821 ( .A(G2427), .B(G2435), .Z(n753) );
  XNOR2_X1 U822 ( .A(G2454), .B(G2443), .ZN(n752) );
  XNOR2_X1 U823 ( .A(n753), .B(n752), .ZN(n760) );
  XOR2_X1 U824 ( .A(G2451), .B(KEYINPUT109), .Z(n755) );
  XNOR2_X1 U825 ( .A(G2430), .B(G2438), .ZN(n754) );
  XNOR2_X1 U826 ( .A(n755), .B(n754), .ZN(n756) );
  XOR2_X1 U827 ( .A(n756), .B(G2446), .Z(n758) );
  XNOR2_X1 U828 ( .A(G1341), .B(G1348), .ZN(n757) );
  XNOR2_X1 U829 ( .A(n758), .B(n757), .ZN(n759) );
  XNOR2_X1 U830 ( .A(n760), .B(n759), .ZN(n761) );
  AND2_X1 U831 ( .A1(n761), .A2(G14), .ZN(G401) );
  AND2_X1 U832 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U833 ( .A(n798), .ZN(G299) );
  NAND2_X1 U834 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U835 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U836 ( .A(G223), .ZN(n827) );
  NAND2_X1 U837 ( .A1(n827), .A2(G567), .ZN(n763) );
  XOR2_X1 U838 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  INV_X1 U839 ( .A(G860), .ZN(n795) );
  NOR2_X1 U840 ( .A1(n922), .A2(n795), .ZN(n764) );
  XOR2_X1 U841 ( .A(KEYINPUT68), .B(n764), .Z(G153) );
  NAND2_X1 U842 ( .A1(G868), .A2(G301), .ZN(n766) );
  INV_X1 U843 ( .A(n894), .ZN(n927) );
  INV_X1 U844 ( .A(G868), .ZN(n807) );
  NAND2_X1 U845 ( .A1(n927), .A2(n807), .ZN(n765) );
  NAND2_X1 U846 ( .A1(n766), .A2(n765), .ZN(G284) );
  NAND2_X1 U847 ( .A1(G868), .A2(G286), .ZN(n768) );
  NAND2_X1 U848 ( .A1(G299), .A2(n807), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U850 ( .A1(n795), .A2(G559), .ZN(n769) );
  NAND2_X1 U851 ( .A1(n769), .A2(n894), .ZN(n770) );
  XNOR2_X1 U852 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G868), .A2(n922), .ZN(n773) );
  NAND2_X1 U854 ( .A1(G868), .A2(n894), .ZN(n771) );
  NOR2_X1 U855 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U856 ( .A1(n773), .A2(n772), .ZN(G282) );
  NAND2_X1 U857 ( .A1(n881), .A2(G123), .ZN(n774) );
  XNOR2_X1 U858 ( .A(n774), .B(KEYINPUT18), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G111), .A2(n882), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n780) );
  NAND2_X1 U861 ( .A1(G99), .A2(n877), .ZN(n778) );
  NAND2_X1 U862 ( .A1(G135), .A2(n878), .ZN(n777) );
  NAND2_X1 U863 ( .A1(n778), .A2(n777), .ZN(n779) );
  NOR2_X1 U864 ( .A1(n780), .A2(n779), .ZN(n989) );
  XNOR2_X1 U865 ( .A(G2096), .B(n989), .ZN(n782) );
  INV_X1 U866 ( .A(G2100), .ZN(n781) );
  NAND2_X1 U867 ( .A1(n782), .A2(n781), .ZN(G156) );
  NAND2_X1 U868 ( .A1(G80), .A2(n783), .ZN(n786) );
  NAND2_X1 U869 ( .A1(G93), .A2(n784), .ZN(n785) );
  NAND2_X1 U870 ( .A1(n786), .A2(n785), .ZN(n793) );
  NAND2_X1 U871 ( .A1(n787), .A2(G55), .ZN(n788) );
  XNOR2_X1 U872 ( .A(n788), .B(KEYINPUT74), .ZN(n791) );
  NAND2_X1 U873 ( .A1(G67), .A2(n789), .ZN(n790) );
  NAND2_X1 U874 ( .A1(n791), .A2(n790), .ZN(n792) );
  OR2_X1 U875 ( .A1(n793), .A2(n792), .ZN(n808) );
  NAND2_X1 U876 ( .A1(G559), .A2(n894), .ZN(n794) );
  XOR2_X1 U877 ( .A(n922), .B(n794), .Z(n805) );
  NAND2_X1 U878 ( .A1(n795), .A2(n805), .ZN(n796) );
  XNOR2_X1 U879 ( .A(n796), .B(KEYINPUT73), .ZN(n797) );
  XOR2_X1 U880 ( .A(n808), .B(n797), .Z(G145) );
  XNOR2_X1 U881 ( .A(n798), .B(G290), .ZN(n804) );
  XOR2_X1 U882 ( .A(KEYINPUT19), .B(KEYINPUT79), .Z(n800) );
  XNOR2_X1 U883 ( .A(G166), .B(G305), .ZN(n799) );
  XNOR2_X1 U884 ( .A(n800), .B(n799), .ZN(n801) );
  XOR2_X1 U885 ( .A(n808), .B(n801), .Z(n802) );
  XNOR2_X1 U886 ( .A(n802), .B(G288), .ZN(n803) );
  XNOR2_X1 U887 ( .A(n804), .B(n803), .ZN(n893) );
  XOR2_X1 U888 ( .A(n893), .B(n805), .Z(n806) );
  NOR2_X1 U889 ( .A1(n807), .A2(n806), .ZN(n810) );
  NOR2_X1 U890 ( .A1(G868), .A2(n808), .ZN(n809) );
  NOR2_X1 U891 ( .A1(n810), .A2(n809), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n811) );
  XOR2_X1 U893 ( .A(KEYINPUT20), .B(n811), .Z(n812) );
  NAND2_X1 U894 ( .A1(G2090), .A2(n812), .ZN(n813) );
  XNOR2_X1 U895 ( .A(KEYINPUT21), .B(n813), .ZN(n814) );
  NAND2_X1 U896 ( .A1(n814), .A2(G2072), .ZN(n815) );
  XNOR2_X1 U897 ( .A(KEYINPUT80), .B(n815), .ZN(G158) );
  XNOR2_X1 U898 ( .A(KEYINPUT67), .B(G57), .ZN(G237) );
  XNOR2_X1 U899 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U900 ( .A1(G108), .A2(G120), .ZN(n816) );
  NOR2_X1 U901 ( .A1(G237), .A2(n816), .ZN(n817) );
  NAND2_X1 U902 ( .A1(G69), .A2(n817), .ZN(n831) );
  NAND2_X1 U903 ( .A1(n831), .A2(G567), .ZN(n824) );
  XOR2_X1 U904 ( .A(KEYINPUT22), .B(KEYINPUT82), .Z(n819) );
  NAND2_X1 U905 ( .A1(G132), .A2(G82), .ZN(n818) );
  XNOR2_X1 U906 ( .A(n819), .B(n818), .ZN(n820) );
  XNOR2_X1 U907 ( .A(n820), .B(KEYINPUT81), .ZN(n821) );
  NOR2_X1 U908 ( .A1(G218), .A2(n821), .ZN(n822) );
  NAND2_X1 U909 ( .A1(G96), .A2(n822), .ZN(n832) );
  NAND2_X1 U910 ( .A1(n832), .A2(G2106), .ZN(n823) );
  NAND2_X1 U911 ( .A1(n824), .A2(n823), .ZN(n906) );
  NAND2_X1 U912 ( .A1(G661), .A2(G483), .ZN(n825) );
  XOR2_X1 U913 ( .A(KEYINPUT83), .B(n825), .Z(n826) );
  NOR2_X1 U914 ( .A1(n906), .A2(n826), .ZN(n830) );
  NAND2_X1 U915 ( .A1(n830), .A2(G36), .ZN(G176) );
  NAND2_X1 U916 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U917 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U918 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U919 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U920 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U922 ( .A(G132), .ZN(G219) );
  INV_X1 U923 ( .A(G120), .ZN(G236) );
  INV_X1 U924 ( .A(G108), .ZN(G238) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G82), .ZN(G220) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  XOR2_X1 U930 ( .A(G2096), .B(KEYINPUT43), .Z(n834) );
  XNOR2_X1 U931 ( .A(G2090), .B(G2678), .ZN(n833) );
  XNOR2_X1 U932 ( .A(n834), .B(n833), .ZN(n835) );
  XOR2_X1 U933 ( .A(n835), .B(KEYINPUT110), .Z(n837) );
  XNOR2_X1 U934 ( .A(G2067), .B(G2072), .ZN(n836) );
  XNOR2_X1 U935 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U936 ( .A(KEYINPUT42), .B(G2100), .Z(n839) );
  XNOR2_X1 U937 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n840) );
  XNOR2_X1 U939 ( .A(n841), .B(n840), .ZN(G227) );
  XOR2_X1 U940 ( .A(KEYINPUT41), .B(G1976), .Z(n843) );
  XNOR2_X1 U941 ( .A(G1996), .B(G1991), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n843), .B(n842), .ZN(n844) );
  XOR2_X1 U943 ( .A(n844), .B(KEYINPUT112), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1981), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n850) );
  XOR2_X1 U946 ( .A(G1956), .B(G1961), .Z(n848) );
  XNOR2_X1 U947 ( .A(G1986), .B(G1971), .ZN(n847) );
  XNOR2_X1 U948 ( .A(n848), .B(n847), .ZN(n849) );
  XOR2_X1 U949 ( .A(n850), .B(n849), .Z(n852) );
  XNOR2_X1 U950 ( .A(G2474), .B(KEYINPUT111), .ZN(n851) );
  XNOR2_X1 U951 ( .A(n852), .B(n851), .ZN(G229) );
  NAND2_X1 U952 ( .A1(n881), .A2(G124), .ZN(n853) );
  XNOR2_X1 U953 ( .A(n853), .B(KEYINPUT44), .ZN(n855) );
  NAND2_X1 U954 ( .A1(G112), .A2(n882), .ZN(n854) );
  NAND2_X1 U955 ( .A1(n855), .A2(n854), .ZN(n859) );
  NAND2_X1 U956 ( .A1(G100), .A2(n877), .ZN(n857) );
  NAND2_X1 U957 ( .A1(G136), .A2(n878), .ZN(n856) );
  NAND2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n858) );
  NOR2_X1 U959 ( .A1(n859), .A2(n858), .ZN(G162) );
  XOR2_X1 U960 ( .A(KEYINPUT48), .B(KEYINPUT46), .Z(n870) );
  NAND2_X1 U961 ( .A1(G106), .A2(n877), .ZN(n861) );
  NAND2_X1 U962 ( .A1(G142), .A2(n878), .ZN(n860) );
  NAND2_X1 U963 ( .A1(n861), .A2(n860), .ZN(n862) );
  XNOR2_X1 U964 ( .A(n862), .B(KEYINPUT45), .ZN(n864) );
  NAND2_X1 U965 ( .A1(G118), .A2(n882), .ZN(n863) );
  NAND2_X1 U966 ( .A1(n864), .A2(n863), .ZN(n867) );
  NAND2_X1 U967 ( .A1(G130), .A2(n881), .ZN(n865) );
  XNOR2_X1 U968 ( .A(KEYINPUT113), .B(n865), .ZN(n866) );
  NOR2_X1 U969 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U970 ( .A(G162), .B(n868), .ZN(n869) );
  XNOR2_X1 U971 ( .A(n870), .B(n869), .ZN(n871) );
  XNOR2_X1 U972 ( .A(n872), .B(n871), .ZN(n875) );
  XNOR2_X1 U973 ( .A(G164), .B(n873), .ZN(n874) );
  XNOR2_X1 U974 ( .A(n875), .B(n874), .ZN(n876) );
  XOR2_X1 U975 ( .A(n876), .B(n989), .Z(n889) );
  NAND2_X1 U976 ( .A1(G103), .A2(n877), .ZN(n880) );
  NAND2_X1 U977 ( .A1(G139), .A2(n878), .ZN(n879) );
  NAND2_X1 U978 ( .A1(n880), .A2(n879), .ZN(n887) );
  NAND2_X1 U979 ( .A1(G127), .A2(n881), .ZN(n884) );
  NAND2_X1 U980 ( .A1(G115), .A2(n882), .ZN(n883) );
  NAND2_X1 U981 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U982 ( .A(KEYINPUT47), .B(n885), .Z(n886) );
  NOR2_X1 U983 ( .A1(n887), .A2(n886), .ZN(n991) );
  XNOR2_X1 U984 ( .A(G160), .B(n991), .ZN(n888) );
  XNOR2_X1 U985 ( .A(n889), .B(n888), .ZN(n891) );
  XOR2_X1 U986 ( .A(n891), .B(n890), .Z(n892) );
  NOR2_X1 U987 ( .A1(G37), .A2(n892), .ZN(G395) );
  XNOR2_X1 U988 ( .A(n922), .B(n893), .ZN(n896) );
  XNOR2_X1 U989 ( .A(G171), .B(n894), .ZN(n895) );
  XNOR2_X1 U990 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U991 ( .A(n897), .B(G286), .Z(n898) );
  NOR2_X1 U992 ( .A1(G37), .A2(n898), .ZN(G397) );
  NOR2_X1 U993 ( .A1(G227), .A2(G229), .ZN(n899) );
  XNOR2_X1 U994 ( .A(n899), .B(KEYINPUT49), .ZN(n902) );
  NOR2_X1 U995 ( .A1(G395), .A2(G397), .ZN(n900) );
  XNOR2_X1 U996 ( .A(n900), .B(KEYINPUT115), .ZN(n901) );
  NOR2_X1 U997 ( .A1(n902), .A2(n901), .ZN(n905) );
  NOR2_X1 U998 ( .A1(G401), .A2(n906), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n903), .B(KEYINPUT114), .ZN(n904) );
  NAND2_X1 U1000 ( .A1(n905), .A2(n904), .ZN(G225) );
  INV_X1 U1001 ( .A(G225), .ZN(G308) );
  INV_X1 U1002 ( .A(n906), .ZN(G319) );
  XNOR2_X1 U1003 ( .A(G16), .B(KEYINPUT56), .ZN(n934) );
  XNOR2_X1 U1004 ( .A(G166), .B(G1971), .ZN(n915) );
  XNOR2_X1 U1005 ( .A(G1956), .B(KEYINPUT122), .ZN(n907) );
  XNOR2_X1 U1006 ( .A(n907), .B(G299), .ZN(n913) );
  INV_X1 U1007 ( .A(n908), .ZN(n910) );
  NAND2_X1 U1008 ( .A1(n910), .A2(n909), .ZN(n911) );
  XOR2_X1 U1009 ( .A(KEYINPUT123), .B(n911), .Z(n912) );
  NOR2_X1 U1010 ( .A1(n913), .A2(n912), .ZN(n914) );
  NAND2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n916) );
  XNOR2_X1 U1012 ( .A(n916), .B(KEYINPUT124), .ZN(n921) );
  XNOR2_X1 U1013 ( .A(G168), .B(G1966), .ZN(n918) );
  NAND2_X1 U1014 ( .A1(n918), .A2(n917), .ZN(n919) );
  XOR2_X1 U1015 ( .A(KEYINPUT57), .B(n919), .Z(n920) );
  NOR2_X1 U1016 ( .A1(n921), .A2(n920), .ZN(n932) );
  XNOR2_X1 U1017 ( .A(G171), .B(G1961), .ZN(n926) );
  XNOR2_X1 U1018 ( .A(G1341), .B(n922), .ZN(n923) );
  NOR2_X1 U1019 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1020 ( .A1(n926), .A2(n925), .ZN(n930) );
  XOR2_X1 U1021 ( .A(G1348), .B(n927), .Z(n928) );
  XNOR2_X1 U1022 ( .A(KEYINPUT121), .B(n928), .ZN(n929) );
  NOR2_X1 U1023 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1024 ( .A1(n932), .A2(n931), .ZN(n933) );
  NAND2_X1 U1025 ( .A1(n934), .A2(n933), .ZN(n1011) );
  XOR2_X1 U1026 ( .A(G1348), .B(KEYINPUT59), .Z(n935) );
  XNOR2_X1 U1027 ( .A(G4), .B(n935), .ZN(n937) );
  XNOR2_X1 U1028 ( .A(G20), .B(G1956), .ZN(n936) );
  NOR2_X1 U1029 ( .A1(n937), .A2(n936), .ZN(n941) );
  XNOR2_X1 U1030 ( .A(G1341), .B(G19), .ZN(n939) );
  XNOR2_X1 U1031 ( .A(G6), .B(G1981), .ZN(n938) );
  NOR2_X1 U1032 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1033 ( .A1(n941), .A2(n940), .ZN(n942) );
  XNOR2_X1 U1034 ( .A(n942), .B(KEYINPUT60), .ZN(n950) );
  XNOR2_X1 U1035 ( .A(G1971), .B(G22), .ZN(n944) );
  XNOR2_X1 U1036 ( .A(G23), .B(G1976), .ZN(n943) );
  NOR2_X1 U1037 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1038 ( .A(G1986), .B(KEYINPUT126), .Z(n945) );
  XNOR2_X1 U1039 ( .A(G24), .B(n945), .ZN(n946) );
  NAND2_X1 U1040 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1041 ( .A(KEYINPUT58), .B(n948), .ZN(n949) );
  NOR2_X1 U1042 ( .A1(n950), .A2(n949), .ZN(n954) );
  XNOR2_X1 U1043 ( .A(G1961), .B(G5), .ZN(n952) );
  XNOR2_X1 U1044 ( .A(G1966), .B(G21), .ZN(n951) );
  NOR2_X1 U1045 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1046 ( .A1(n954), .A2(n953), .ZN(n955) );
  XNOR2_X1 U1047 ( .A(n955), .B(KEYINPUT127), .ZN(n956) );
  XNOR2_X1 U1048 ( .A(n956), .B(KEYINPUT61), .ZN(n958) );
  XNOR2_X1 U1049 ( .A(G16), .B(KEYINPUT125), .ZN(n957) );
  NAND2_X1 U1050 ( .A1(n958), .A2(n957), .ZN(n959) );
  NAND2_X1 U1051 ( .A1(G11), .A2(n959), .ZN(n1009) );
  XOR2_X1 U1052 ( .A(G2067), .B(G26), .Z(n960) );
  NAND2_X1 U1053 ( .A1(G28), .A2(n960), .ZN(n962) );
  XNOR2_X1 U1054 ( .A(G25), .B(G1991), .ZN(n961) );
  NOR2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n971) );
  XNOR2_X1 U1056 ( .A(G2072), .B(KEYINPUT118), .ZN(n963) );
  XNOR2_X1 U1057 ( .A(n963), .B(G33), .ZN(n969) );
  XNOR2_X1 U1058 ( .A(G1996), .B(G32), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(n964), .B(G27), .ZN(n965) );
  NOR2_X1 U1060 ( .A1(n966), .A2(n965), .ZN(n967) );
  XNOR2_X1 U1061 ( .A(KEYINPUT119), .B(n967), .ZN(n968) );
  NOR2_X1 U1062 ( .A1(n969), .A2(n968), .ZN(n970) );
  NAND2_X1 U1063 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1064 ( .A(n972), .B(KEYINPUT53), .ZN(n975) );
  XOR2_X1 U1065 ( .A(G2084), .B(G34), .Z(n973) );
  XNOR2_X1 U1066 ( .A(KEYINPUT54), .B(n973), .ZN(n974) );
  NAND2_X1 U1067 ( .A1(n975), .A2(n974), .ZN(n977) );
  XNOR2_X1 U1068 ( .A(G35), .B(G2090), .ZN(n976) );
  NOR2_X1 U1069 ( .A1(n977), .A2(n976), .ZN(n978) );
  XNOR2_X1 U1070 ( .A(KEYINPUT120), .B(n978), .ZN(n979) );
  NOR2_X1 U1071 ( .A1(G29), .A2(n979), .ZN(n980) );
  XNOR2_X1 U1072 ( .A(n980), .B(KEYINPUT55), .ZN(n1007) );
  XNOR2_X1 U1073 ( .A(G2090), .B(G162), .ZN(n982) );
  NAND2_X1 U1074 ( .A1(n982), .A2(n981), .ZN(n983) );
  XNOR2_X1 U1075 ( .A(n983), .B(KEYINPUT51), .ZN(n984) );
  XNOR2_X1 U1076 ( .A(KEYINPUT116), .B(n984), .ZN(n986) );
  NAND2_X1 U1077 ( .A1(n986), .A2(n985), .ZN(n987) );
  NOR2_X1 U1078 ( .A1(n988), .A2(n987), .ZN(n1002) );
  NOR2_X1 U1079 ( .A1(n990), .A2(n989), .ZN(n998) );
  XOR2_X1 U1080 ( .A(G2072), .B(n991), .Z(n993) );
  XOR2_X1 U1081 ( .A(G164), .B(G2078), .Z(n992) );
  NOR2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n994) );
  XOR2_X1 U1083 ( .A(KEYINPUT50), .B(n994), .Z(n996) );
  XOR2_X1 U1084 ( .A(G160), .B(G2084), .Z(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1086 ( .A1(n998), .A2(n997), .ZN(n999) );
  NOR2_X1 U1087 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1088 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XNOR2_X1 U1089 ( .A(KEYINPUT52), .B(n1003), .ZN(n1004) );
  XOR2_X1 U1090 ( .A(KEYINPUT117), .B(n1004), .Z(n1005) );
  NAND2_X1 U1091 ( .A1(G29), .A2(n1005), .ZN(n1006) );
  NAND2_X1 U1092 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1093 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1094 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1095 ( .A(KEYINPUT62), .B(n1012), .Z(G311) );
  INV_X1 U1096 ( .A(G311), .ZN(G150) );
endmodule

