//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 1 0 0 1 1 1 0 1 1 1 0 1 1 1 1 0 0 0 0 0 1 1 0 0 0 0 1 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:36:43 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n234, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n241, new_n242, new_n243, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1237,
    new_n1238, new_n1239, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0005(.A1(G1), .A2(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n206), .A2(G13), .ZN(new_n207));
  OAI211_X1 g0007(.A(new_n207), .B(G250), .C1(G257), .C2(G264), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT0), .ZN(new_n209));
  OAI21_X1  g0009(.A(G50), .B1(G58), .B2(G68), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT64), .ZN(new_n211));
  NAND2_X1  g0011(.A1(G1), .A2(G13), .ZN(new_n212));
  INV_X1    g0012(.A(G20), .ZN(new_n213));
  NOR2_X1   g0013(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n211), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(KEYINPUT65), .B(G77), .ZN(new_n216));
  AND2_X1   g0016(.A1(new_n216), .A2(G244), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n220));
  NAND2_X1  g0020(.A1(G58), .A2(G232), .ZN(new_n221));
  NAND4_X1  g0021(.A1(new_n218), .A2(new_n219), .A3(new_n220), .A4(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n206), .B1(new_n217), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n209), .B(new_n215), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XNOR2_X1  g0025(.A(G238), .B(G244), .ZN(new_n226));
  XNOR2_X1  g0026(.A(new_n226), .B(G232), .ZN(new_n227));
  XNOR2_X1  g0027(.A(KEYINPUT2), .B(G226), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n227), .B(new_n228), .ZN(new_n229));
  XOR2_X1   g0029(.A(G264), .B(G270), .Z(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n229), .B(new_n232), .ZN(G358));
  XNOR2_X1  g0033(.A(G50), .B(G68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G58), .B(G77), .ZN(new_n235));
  XOR2_X1   g0035(.A(new_n234), .B(new_n235), .Z(new_n236));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n236), .B(new_n239), .ZN(G351));
  NOR2_X1   g0040(.A1(G20), .A2(G33), .ZN(new_n241));
  AOI22_X1  g0041(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n241), .ZN(new_n242));
  INV_X1    g0042(.A(G33), .ZN(new_n243));
  NOR2_X1   g0043(.A1(new_n243), .A2(G20), .ZN(new_n244));
  XNOR2_X1  g0044(.A(new_n244), .B(KEYINPUT69), .ZN(new_n245));
  XNOR2_X1  g0045(.A(KEYINPUT8), .B(G58), .ZN(new_n246));
  OAI21_X1  g0046(.A(new_n242), .B1(new_n245), .B2(new_n246), .ZN(new_n247));
  NAND3_X1  g0047(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(new_n212), .ZN(new_n249));
  INV_X1    g0049(.A(KEYINPUT68), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND3_X1  g0051(.A1(new_n248), .A2(KEYINPUT68), .A3(new_n212), .ZN(new_n252));
  NAND2_X1  g0052(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n254), .A2(G1), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n255), .A2(G20), .ZN(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  AOI22_X1  g0057(.A1(new_n247), .A2(new_n253), .B1(new_n202), .B2(new_n257), .ZN(new_n258));
  NOR2_X1   g0058(.A1(new_n253), .A2(new_n257), .ZN(new_n259));
  OAI21_X1  g0059(.A(KEYINPUT70), .B1(new_n213), .B2(G1), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT70), .ZN(new_n261));
  INV_X1    g0061(.A(G1), .ZN(new_n262));
  NAND3_X1  g0062(.A1(new_n261), .A2(new_n262), .A3(G20), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n259), .A2(G50), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n258), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(new_n266), .ZN(new_n267));
  NAND2_X1  g0067(.A1(G33), .A2(G41), .ZN(new_n268));
  INV_X1    g0068(.A(KEYINPUT66), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n212), .ZN(new_n271));
  NAND3_X1  g0071(.A1(KEYINPUT66), .A2(G33), .A3(G41), .ZN(new_n272));
  NAND3_X1  g0072(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G45), .ZN(new_n275));
  AOI21_X1  g0075(.A(G1), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND3_X1  g0076(.A1(new_n273), .A2(G274), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n276), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G226), .ZN(new_n280));
  OAI21_X1  g0080(.A(new_n277), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n243), .A2(KEYINPUT3), .ZN(new_n282));
  INV_X1    g0082(.A(KEYINPUT3), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n283), .A2(G33), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n282), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n285), .A2(new_n216), .ZN(new_n286));
  OR2_X1    g0086(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n287));
  NAND2_X1  g0087(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n288));
  NAND4_X1  g0088(.A1(new_n287), .A2(new_n282), .A3(new_n284), .A4(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(G222), .ZN(new_n290));
  INV_X1    g0090(.A(G223), .ZN(new_n291));
  XNOR2_X1  g0091(.A(KEYINPUT3), .B(G33), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(G1698), .ZN(new_n293));
  OAI221_X1 g0093(.A(new_n286), .B1(new_n289), .B2(new_n290), .C1(new_n291), .C2(new_n293), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n271), .A2(new_n268), .ZN(new_n295));
  INV_X1    g0095(.A(new_n295), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n281), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G179), .ZN(new_n298));
  AND2_X1   g0098(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n297), .A2(G169), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n267), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  INV_X1    g0101(.A(G200), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n297), .A2(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT73), .ZN(new_n304));
  OAI21_X1  g0104(.A(KEYINPUT10), .B1(new_n303), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n297), .A2(G190), .ZN(new_n306));
  XNOR2_X1  g0106(.A(new_n306), .B(KEYINPUT72), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n266), .A2(KEYINPUT9), .ZN(new_n308));
  INV_X1    g0108(.A(KEYINPUT9), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n258), .A2(new_n309), .A3(new_n265), .ZN(new_n310));
  AOI21_X1  g0110(.A(new_n303), .B1(new_n308), .B2(new_n310), .ZN(new_n311));
  AOI21_X1  g0111(.A(new_n305), .B1(new_n307), .B2(new_n311), .ZN(new_n312));
  INV_X1    g0112(.A(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(new_n305), .A3(new_n311), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n301), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n273), .A2(new_n278), .A3(G238), .ZN(new_n316));
  AND2_X1   g0116(.A1(new_n277), .A2(new_n316), .ZN(new_n317));
  NAND3_X1  g0117(.A1(new_n287), .A2(G226), .A3(new_n288), .ZN(new_n318));
  NAND2_X1  g0118(.A1(G232), .A2(G1698), .ZN(new_n319));
  AOI21_X1  g0119(.A(new_n285), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND2_X1  g0120(.A1(G33), .A2(G97), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n296), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n317), .A2(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(KEYINPUT13), .ZN(new_n325));
  INV_X1    g0125(.A(KEYINPUT13), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n317), .B2(new_n323), .ZN(new_n327));
  OAI21_X1  g0127(.A(G169), .B1(new_n325), .B2(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(KEYINPUT14), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT14), .ZN(new_n330));
  OAI211_X1 g0130(.A(new_n330), .B(G169), .C1(new_n325), .C2(new_n327), .ZN(new_n331));
  INV_X1    g0131(.A(KEYINPUT74), .ZN(new_n332));
  AND2_X1   g0132(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n333));
  NOR2_X1   g0133(.A1(KEYINPUT67), .A2(G1698), .ZN(new_n334));
  NOR3_X1   g0134(.A1(new_n333), .A2(new_n334), .A3(new_n280), .ZN(new_n335));
  INV_X1    g0135(.A(new_n319), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n292), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n295), .B1(new_n337), .B2(new_n321), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n277), .A2(new_n316), .ZN(new_n339));
  OAI21_X1  g0139(.A(new_n332), .B1(new_n338), .B2(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n317), .A2(new_n323), .A3(KEYINPUT74), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(KEYINPUT13), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n338), .A2(new_n339), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n298), .B1(new_n343), .B2(new_n326), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT78), .ZN(new_n345));
  AND3_X1   g0145(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(new_n345), .B1(new_n342), .B2(new_n344), .ZN(new_n347));
  OAI211_X1 g0147(.A(new_n329), .B(new_n331), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G68), .ZN(new_n349));
  AOI21_X1  g0149(.A(KEYINPUT77), .B1(new_n257), .B2(new_n349), .ZN(new_n350));
  XOR2_X1   g0150(.A(new_n350), .B(KEYINPUT12), .Z(new_n351));
  INV_X1    g0151(.A(new_n249), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n352), .A2(new_n256), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  AOI21_X1  g0154(.A(new_n349), .B1(new_n260), .B2(new_n263), .ZN(new_n355));
  AOI21_X1  g0155(.A(new_n351), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  AOI22_X1  g0156(.A1(new_n241), .A2(G50), .B1(G20), .B2(new_n349), .ZN(new_n357));
  INV_X1    g0157(.A(G77), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n357), .B1(new_n245), .B2(new_n358), .ZN(new_n359));
  XNOR2_X1  g0159(.A(KEYINPUT75), .B(KEYINPUT11), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n359), .A2(new_n253), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n359), .B2(new_n253), .ZN(new_n362));
  OR3_X1    g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT76), .ZN(new_n363));
  OAI21_X1  g0163(.A(KEYINPUT76), .B1(new_n361), .B2(new_n362), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n356), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n348), .A2(new_n365), .ZN(new_n366));
  AND2_X1   g0166(.A1(new_n356), .A2(new_n364), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n342), .B(G190), .C1(KEYINPUT13), .C2(new_n324), .ZN(new_n368));
  OAI21_X1  g0168(.A(G200), .B1(new_n325), .B2(new_n327), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n367), .A2(new_n368), .A3(new_n363), .A4(new_n369), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n333), .A2(new_n334), .ZN(new_n371));
  NAND3_X1  g0171(.A1(new_n371), .A2(new_n292), .A3(G232), .ZN(new_n372));
  INV_X1    g0172(.A(G107), .ZN(new_n373));
  INV_X1    g0173(.A(G238), .ZN(new_n374));
  OAI221_X1 g0174(.A(new_n372), .B1(new_n373), .B2(new_n292), .C1(new_n374), .C2(new_n293), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(new_n296), .ZN(new_n376));
  NAND3_X1  g0176(.A1(new_n273), .A2(new_n278), .A3(G244), .ZN(new_n377));
  AND2_X1   g0177(.A1(new_n277), .A2(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(G169), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(KEYINPUT71), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n376), .A2(new_n378), .ZN(new_n381));
  OAI22_X1  g0181(.A1(new_n379), .A2(new_n380), .B1(new_n381), .B2(G179), .ZN(new_n382));
  NAND4_X1  g0182(.A1(new_n376), .A2(KEYINPUT71), .A3(new_n298), .A4(new_n378), .ZN(new_n383));
  XNOR2_X1  g0183(.A(KEYINPUT15), .B(G87), .ZN(new_n384));
  INV_X1    g0184(.A(new_n384), .ZN(new_n385));
  AOI22_X1  g0185(.A1(new_n385), .A2(new_n244), .B1(new_n216), .B2(G20), .ZN(new_n386));
  INV_X1    g0186(.A(new_n246), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n387), .A2(new_n241), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n352), .B1(new_n386), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n264), .A2(G77), .ZN(new_n390));
  OAI22_X1  g0190(.A1(new_n390), .A2(new_n353), .B1(new_n216), .B2(new_n256), .ZN(new_n391));
  OR2_X1    g0191(.A1(new_n389), .A2(new_n391), .ZN(new_n392));
  AND2_X1   g0192(.A1(new_n383), .A2(new_n392), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n381), .B2(G200), .ZN(new_n394));
  NAND3_X1  g0194(.A1(new_n376), .A2(G190), .A3(new_n378), .ZN(new_n395));
  AOI22_X1  g0195(.A1(new_n382), .A2(new_n393), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND4_X1  g0196(.A1(new_n315), .A2(new_n366), .A3(new_n370), .A4(new_n396), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT81), .ZN(new_n398));
  INV_X1    g0198(.A(G58), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n399), .A2(new_n349), .ZN(new_n400));
  OAI21_X1  g0200(.A(G20), .B1(new_n400), .B2(new_n201), .ZN(new_n401));
  NAND2_X1  g0201(.A1(new_n241), .A2(G159), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT7), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n292), .B2(G20), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n285), .A2(KEYINPUT7), .A3(new_n213), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n403), .B1(new_n407), .B2(G68), .ZN(new_n408));
  XNOR2_X1  g0208(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n409));
  OAI21_X1  g0209(.A(new_n249), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT79), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n408), .A2(new_n411), .A3(KEYINPUT16), .ZN(new_n412));
  AOI21_X1  g0212(.A(KEYINPUT7), .B1(new_n285), .B2(new_n213), .ZN(new_n413));
  AOI211_X1 g0213(.A(new_n404), .B(G20), .C1(new_n282), .C2(new_n284), .ZN(new_n414));
  OAI21_X1  g0214(.A(G68), .B1(new_n413), .B2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(new_n403), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n415), .A2(KEYINPUT16), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(KEYINPUT79), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n410), .B1(new_n412), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n387), .A2(new_n264), .ZN(new_n420));
  INV_X1    g0220(.A(new_n420), .ZN(new_n421));
  AOI22_X1  g0221(.A1(new_n259), .A2(new_n421), .B1(new_n257), .B2(new_n246), .ZN(new_n422));
  INV_X1    g0222(.A(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n398), .B1(new_n419), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n415), .A2(new_n416), .ZN(new_n425));
  INV_X1    g0225(.A(new_n409), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n352), .B1(new_n425), .B2(new_n426), .ZN(new_n427));
  AOI21_X1  g0227(.A(new_n411), .B1(new_n408), .B2(KEYINPUT16), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n349), .B1(new_n405), .B2(new_n406), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT16), .ZN(new_n430));
  NOR4_X1   g0230(.A1(new_n429), .A2(new_n403), .A3(KEYINPUT79), .A4(new_n430), .ZN(new_n431));
  OAI21_X1  g0231(.A(new_n427), .B1(new_n428), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n432), .A2(KEYINPUT81), .A3(new_n422), .ZN(new_n433));
  INV_X1    g0233(.A(G87), .ZN(new_n434));
  OAI22_X1  g0234(.A1(new_n289), .A2(new_n291), .B1(new_n243), .B2(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n293), .A2(new_n280), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n296), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n273), .A2(new_n278), .A3(G232), .ZN(new_n438));
  AND2_X1   g0238(.A1(new_n277), .A2(new_n438), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n437), .A2(G179), .A3(new_n439), .ZN(new_n440));
  AND2_X1   g0240(.A1(new_n437), .A2(new_n439), .ZN(new_n441));
  INV_X1    g0241(.A(G169), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n440), .B1(new_n441), .B2(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n424), .A2(new_n433), .A3(new_n443), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT18), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT18), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n424), .A2(new_n446), .A3(new_n433), .A4(new_n443), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n418), .A2(new_n412), .ZN(new_n448));
  AOI21_X1  g0248(.A(new_n423), .B1(new_n448), .B2(new_n427), .ZN(new_n449));
  INV_X1    g0249(.A(G190), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n437), .A2(new_n450), .A3(new_n439), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(new_n441), .B2(G200), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT17), .B1(new_n449), .B2(new_n452), .ZN(new_n453));
  AND4_X1   g0253(.A1(KEYINPUT17), .A2(new_n432), .A3(new_n452), .A4(new_n422), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND3_X1  g0255(.A1(new_n445), .A2(new_n447), .A3(new_n455), .ZN(new_n456));
  NOR2_X1   g0256(.A1(new_n397), .A2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT4), .ZN(new_n458));
  INV_X1    g0258(.A(G244), .ZN(new_n459));
  OAI21_X1  g0259(.A(new_n458), .B1(new_n289), .B2(new_n459), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n282), .A2(new_n284), .A3(G250), .A4(G1698), .ZN(new_n461));
  NAND2_X1  g0261(.A1(G33), .A2(G283), .ZN(new_n462));
  AND2_X1   g0262(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND4_X1  g0263(.A1(new_n371), .A2(new_n292), .A3(KEYINPUT4), .A4(G244), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n460), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  NAND2_X1  g0265(.A1(new_n465), .A2(new_n296), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT83), .ZN(new_n467));
  NOR2_X1   g0267(.A1(new_n275), .A2(G1), .ZN(new_n468));
  NAND2_X1  g0268(.A1(KEYINPUT5), .A2(G41), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NOR2_X1   g0270(.A1(KEYINPUT5), .A2(G41), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n468), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n273), .A2(new_n472), .ZN(new_n473));
  INV_X1    g0273(.A(G257), .ZN(new_n474));
  OAI21_X1  g0274(.A(new_n467), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  NAND4_X1  g0275(.A1(new_n273), .A2(new_n472), .A3(KEYINPUT83), .A4(G257), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g0277(.A1(new_n262), .A2(G45), .ZN(new_n478));
  INV_X1    g0278(.A(new_n471), .ZN(new_n479));
  AOI21_X1  g0279(.A(new_n478), .B1(new_n479), .B2(new_n469), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n480), .A2(G274), .A3(new_n273), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n466), .A2(new_n477), .A3(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT84), .ZN(new_n483));
  NAND2_X1  g0283(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n481), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n485), .B1(new_n465), .B2(new_n296), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n486), .A2(KEYINPUT84), .A3(new_n477), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g0288(.A(KEYINPUT85), .B1(new_n488), .B2(new_n450), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT85), .ZN(new_n490));
  NAND4_X1  g0290(.A1(new_n484), .A2(new_n490), .A3(G190), .A4(new_n487), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n241), .A2(G77), .ZN(new_n492));
  INV_X1    g0292(.A(KEYINPUT6), .ZN(new_n493));
  INV_X1    g0293(.A(G97), .ZN(new_n494));
  NOR3_X1   g0294(.A1(new_n493), .A2(new_n494), .A3(G107), .ZN(new_n495));
  XNOR2_X1  g0295(.A(G97), .B(G107), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n495), .B1(new_n493), .B2(new_n496), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n492), .B1(new_n497), .B2(new_n213), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n373), .B1(new_n405), .B2(new_n406), .ZN(new_n499));
  OAI21_X1  g0299(.A(new_n249), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n257), .A2(new_n494), .ZN(new_n501));
  INV_X1    g0301(.A(KEYINPUT82), .ZN(new_n502));
  OAI21_X1  g0302(.A(new_n502), .B1(new_n243), .B2(G1), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n262), .A2(KEYINPUT82), .A3(G33), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g0305(.A1(new_n251), .A2(new_n505), .A3(new_n256), .A4(new_n252), .ZN(new_n506));
  OAI211_X1 g0306(.A(new_n500), .B(new_n501), .C1(new_n494), .C2(new_n506), .ZN(new_n507));
  AOI21_X1  g0307(.A(new_n507), .B1(G200), .B2(new_n482), .ZN(new_n508));
  NAND3_X1  g0308(.A1(new_n489), .A2(new_n491), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n486), .A2(new_n298), .A3(new_n477), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  AOI21_X1  g0311(.A(new_n511), .B1(new_n488), .B2(new_n442), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n262), .A2(new_n373), .A3(G13), .A4(G20), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT25), .ZN(new_n515));
  XNOR2_X1  g0315(.A(new_n514), .B(new_n515), .ZN(new_n516));
  OAI21_X1  g0316(.A(new_n516), .B1(new_n506), .B2(new_n373), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(KEYINPUT91), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT91), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n519), .B(new_n516), .C1(new_n506), .C2(new_n373), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n518), .A2(new_n520), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n434), .A2(KEYINPUT90), .A3(G20), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n292), .A2(new_n522), .ZN(new_n523));
  INV_X1    g0323(.A(KEYINPUT22), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g0325(.A1(G33), .A2(G116), .ZN(new_n526));
  NOR2_X1   g0326(.A1(new_n526), .A2(G20), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT23), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n528), .B1(new_n213), .B2(G107), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n373), .A2(KEYINPUT23), .A3(G20), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n527), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n292), .A2(KEYINPUT22), .A3(new_n522), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n525), .A2(new_n531), .A3(new_n532), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT24), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  NAND4_X1  g0335(.A1(new_n525), .A2(new_n531), .A3(new_n532), .A4(KEYINPUT24), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n535), .A2(new_n249), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n521), .A2(new_n537), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n282), .A2(new_n284), .A3(G257), .A4(G1698), .ZN(new_n539));
  NAND2_X1  g0339(.A1(G33), .A2(G294), .ZN(new_n540));
  INV_X1    g0340(.A(G250), .ZN(new_n541));
  OAI211_X1 g0341(.A(new_n539), .B(new_n540), .C1(new_n289), .C2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n542), .A2(new_n296), .ZN(new_n543));
  NAND3_X1  g0343(.A1(new_n273), .A2(new_n472), .A3(G264), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n544), .A3(new_n481), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n442), .ZN(new_n546));
  NAND4_X1  g0346(.A1(new_n543), .A2(new_n544), .A3(new_n298), .A4(new_n481), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n538), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(KEYINPUT21), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n462), .B(new_n213), .C1(G33), .C2(new_n494), .ZN(new_n550));
  INV_X1    g0350(.A(G116), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n551), .A2(G20), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n550), .A2(new_n249), .A3(new_n552), .ZN(new_n553));
  OR2_X1    g0353(.A1(KEYINPUT89), .A2(KEYINPUT20), .ZN(new_n554));
  OR2_X1    g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(KEYINPUT89), .A2(KEYINPUT20), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n553), .A2(new_n554), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g0357(.A1(new_n255), .A2(G20), .A3(new_n551), .ZN(new_n558));
  NAND4_X1  g0358(.A1(new_n505), .A2(new_n352), .A3(new_n256), .A4(G116), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n555), .A2(new_n557), .A3(new_n558), .A4(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n560), .A2(G169), .ZN(new_n561));
  NAND3_X1  g0361(.A1(new_n273), .A2(new_n472), .A3(G270), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n481), .A2(new_n562), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n371), .A2(new_n292), .A3(G257), .ZN(new_n564));
  XNOR2_X1  g0364(.A(KEYINPUT88), .B(G303), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n285), .A2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(G264), .ZN(new_n567));
  OAI211_X1 g0367(.A(new_n564), .B(new_n566), .C1(new_n567), .C2(new_n293), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n563), .B1(new_n568), .B2(new_n296), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n549), .B1(new_n561), .B2(new_n569), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n569), .A2(G179), .A3(new_n560), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n568), .A2(new_n296), .ZN(new_n572));
  INV_X1    g0372(.A(new_n563), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND4_X1  g0374(.A1(new_n574), .A2(KEYINPUT21), .A3(G169), .A4(new_n560), .ZN(new_n575));
  NAND4_X1  g0375(.A1(new_n548), .A2(new_n570), .A3(new_n571), .A4(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n545), .A2(G200), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n543), .A2(new_n544), .A3(G190), .A4(new_n481), .ZN(new_n578));
  NAND4_X1  g0378(.A1(new_n577), .A2(new_n521), .A3(new_n537), .A4(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(KEYINPUT87), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n213), .A2(G68), .ZN(new_n581));
  OAI21_X1  g0381(.A(new_n580), .B1(new_n285), .B2(new_n581), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n292), .A2(KEYINPUT87), .A3(new_n213), .A4(G68), .ZN(new_n583));
  INV_X1    g0383(.A(KEYINPUT19), .ZN(new_n584));
  NOR2_X1   g0384(.A1(G97), .A2(G107), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(new_n434), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n321), .A2(new_n213), .ZN(new_n587));
  AOI21_X1  g0387(.A(new_n584), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NOR4_X1   g0388(.A1(new_n243), .A2(new_n494), .A3(KEYINPUT19), .A4(G20), .ZN(new_n589));
  OAI211_X1 g0389(.A(new_n582), .B(new_n583), .C1(new_n588), .C2(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n249), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n257), .A2(new_n384), .ZN(new_n592));
  OR2_X1    g0392(.A1(new_n506), .A2(new_n434), .ZN(new_n593));
  AND3_X1   g0393(.A1(new_n591), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT86), .ZN(new_n595));
  AND3_X1   g0395(.A1(new_n270), .A2(new_n271), .A3(new_n272), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n478), .A2(G250), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n595), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n273), .A2(KEYINPUT86), .A3(G250), .A4(new_n478), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  NAND4_X1  g0400(.A1(new_n282), .A2(new_n284), .A3(G244), .A4(G1698), .ZN(new_n601));
  OAI211_X1 g0401(.A(new_n526), .B(new_n601), .C1(new_n289), .C2(new_n374), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n602), .A2(new_n296), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n273), .A2(G274), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n604), .A2(new_n468), .ZN(new_n605));
  NAND3_X1  g0405(.A1(new_n600), .A2(new_n603), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(G200), .ZN(new_n607));
  AOI22_X1  g0407(.A1(new_n602), .A2(new_n296), .B1(new_n604), .B2(new_n468), .ZN(new_n608));
  NAND3_X1  g0408(.A1(new_n608), .A2(G190), .A3(new_n600), .ZN(new_n609));
  NAND3_X1  g0409(.A1(new_n594), .A2(new_n607), .A3(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n606), .A2(new_n442), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n608), .A2(new_n298), .A3(new_n600), .ZN(new_n612));
  OR2_X1    g0412(.A1(new_n506), .A2(new_n384), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n591), .A2(new_n592), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n612), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n572), .A2(new_n573), .A3(G190), .ZN(new_n616));
  INV_X1    g0416(.A(new_n560), .ZN(new_n617));
  OAI211_X1 g0417(.A(new_n616), .B(new_n617), .C1(new_n569), .C2(new_n302), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n579), .A2(new_n610), .A3(new_n615), .A4(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(new_n576), .A2(new_n619), .ZN(new_n620));
  AND4_X1   g0420(.A1(new_n457), .A2(new_n509), .A3(new_n513), .A4(new_n620), .ZN(G372));
  NAND3_X1  g0421(.A1(new_n579), .A2(new_n610), .A3(new_n615), .ZN(new_n622));
  NAND3_X1  g0422(.A1(new_n570), .A2(new_n571), .A3(new_n575), .ZN(new_n623));
  INV_X1    g0423(.A(new_n623), .ZN(new_n624));
  AOI21_X1  g0424(.A(new_n622), .B1(new_n624), .B2(new_n548), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n509), .A2(new_n625), .A3(new_n513), .ZN(new_n626));
  AND4_X1   g0426(.A1(KEYINPUT84), .A2(new_n466), .A3(new_n477), .A4(new_n481), .ZN(new_n627));
  AOI21_X1  g0427(.A(KEYINPUT84), .B1(new_n486), .B2(new_n477), .ZN(new_n628));
  OAI21_X1  g0428(.A(new_n442), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n507), .A2(new_n510), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n629), .A2(new_n630), .A3(new_n615), .A4(new_n610), .ZN(new_n631));
  INV_X1    g0431(.A(KEYINPUT26), .ZN(new_n632));
  NOR2_X1   g0432(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n610), .A2(new_n615), .ZN(new_n634));
  INV_X1    g0434(.A(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(KEYINPUT26), .B1(new_n512), .B2(new_n635), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n615), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g0437(.A(new_n457), .B1(new_n626), .B2(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n442), .B1(new_n437), .B2(new_n439), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(G179), .B2(new_n441), .ZN(new_n640));
  OAI21_X1  g0440(.A(KEYINPUT18), .B1(new_n449), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n432), .A2(new_n422), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n642), .A2(new_n446), .A3(new_n443), .ZN(new_n643));
  AND2_X1   g0443(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n382), .A2(new_n393), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n348), .A2(new_n365), .B1(new_n370), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n432), .A2(new_n452), .A3(new_n422), .ZN(new_n647));
  INV_X1    g0447(.A(KEYINPUT17), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND3_X1  g0449(.A1(new_n449), .A2(KEYINPUT17), .A3(new_n452), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g0451(.A(new_n644), .B1(new_n646), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n313), .A2(new_n314), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n301), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n638), .A2(new_n654), .ZN(G369));
  NAND2_X1  g0455(.A1(new_n255), .A2(new_n213), .ZN(new_n656));
  OR2_X1    g0456(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n656), .A2(KEYINPUT27), .ZN(new_n658));
  NAND3_X1  g0458(.A1(new_n657), .A2(G213), .A3(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(G343), .ZN(new_n660));
  NOR2_X1   g0460(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(new_n661), .ZN(new_n662));
  NOR2_X1   g0462(.A1(new_n617), .A2(new_n662), .ZN(new_n663));
  XNOR2_X1  g0463(.A(new_n623), .B(new_n663), .ZN(new_n664));
  AND2_X1   g0464(.A1(new_n664), .A2(new_n618), .ZN(new_n665));
  XNOR2_X1  g0465(.A(KEYINPUT92), .B(G330), .ZN(new_n666));
  INV_X1    g0466(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n538), .A2(new_n661), .ZN(new_n670));
  AND2_X1   g0470(.A1(new_n546), .A2(new_n547), .ZN(new_n671));
  AOI22_X1  g0471(.A1(new_n670), .A2(new_n579), .B1(new_n671), .B2(new_n538), .ZN(new_n672));
  NOR2_X1   g0472(.A1(new_n548), .A2(new_n661), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n623), .A2(new_n662), .ZN(new_n676));
  OAI22_X1  g0476(.A1(new_n672), .A2(new_n676), .B1(new_n548), .B2(new_n661), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n675), .A2(new_n678), .ZN(G399));
  NOR2_X1   g0479(.A1(new_n586), .A2(G116), .ZN(new_n680));
  XOR2_X1   g0480(.A(new_n680), .B(KEYINPUT93), .Z(new_n681));
  INV_X1    g0481(.A(new_n207), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n682), .A2(G41), .ZN(new_n683));
  NOR3_X1   g0483(.A1(new_n681), .A2(new_n262), .A3(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n210), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n684), .B1(new_n685), .B2(new_n683), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT28), .Z(new_n687));
  OAI21_X1  g0487(.A(new_n662), .B1(new_n637), .B2(new_n626), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT29), .ZN(new_n689));
  NAND3_X1  g0489(.A1(new_n688), .A2(KEYINPUT95), .A3(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT95), .ZN(new_n691));
  INV_X1    g0491(.A(new_n615), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n631), .A2(new_n632), .ZN(new_n693));
  NAND3_X1  g0493(.A1(new_n512), .A2(KEYINPUT26), .A3(new_n635), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n509), .A2(new_n625), .A3(new_n513), .ZN(new_n696));
  AOI21_X1  g0496(.A(new_n661), .B1(new_n695), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n691), .B1(new_n697), .B2(KEYINPUT29), .ZN(new_n698));
  NAND2_X1  g0498(.A1(new_n509), .A2(new_n513), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n624), .A2(KEYINPUT96), .A3(new_n548), .ZN(new_n700));
  INV_X1    g0500(.A(new_n622), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  AOI21_X1  g0502(.A(KEYINPUT96), .B1(new_n624), .B2(new_n548), .ZN(new_n703));
  NOR3_X1   g0503(.A1(new_n699), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  OAI211_X1 g0504(.A(KEYINPUT29), .B(new_n662), .C1(new_n704), .C2(new_n637), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n690), .A2(new_n698), .A3(new_n705), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n620), .A2(new_n509), .A3(new_n513), .A4(new_n662), .ZN(new_n707));
  INV_X1    g0507(.A(KEYINPUT30), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n708), .A2(KEYINPUT94), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n627), .A2(new_n628), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n572), .A2(new_n573), .A3(G179), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n543), .A2(new_n544), .ZN(new_n712));
  NOR3_X1   g0512(.A1(new_n711), .A2(new_n606), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n710), .B2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n713), .A2(new_n484), .A3(new_n487), .A4(new_n709), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n569), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n716), .A2(new_n482), .A3(new_n545), .A4(new_n606), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n717), .ZN(new_n718));
  OAI21_X1  g0518(.A(new_n661), .B1(new_n714), .B2(new_n718), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  OAI211_X1 g0521(.A(KEYINPUT31), .B(new_n661), .C1(new_n714), .C2(new_n718), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n707), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(new_n667), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n706), .A2(new_n724), .ZN(new_n725));
  OAI21_X1  g0525(.A(new_n687), .B1(new_n725), .B2(G1), .ZN(G364));
  NOR2_X1   g0526(.A1(new_n254), .A2(G20), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n262), .B1(new_n727), .B2(G45), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n683), .A2(new_n729), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n669), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n665), .A2(new_n667), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(G13), .A2(G33), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(G20), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  OR2_X1    g0537(.A1(new_n665), .A2(new_n737), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n212), .B1(G20), .B2(new_n442), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  NAND2_X1  g0540(.A1(G20), .A2(G179), .ZN(new_n741));
  NOR3_X1   g0541(.A1(new_n741), .A2(new_n450), .A3(G200), .ZN(new_n742));
  INV_X1    g0542(.A(new_n742), .ZN(new_n743));
  INV_X1    g0543(.A(G322), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR3_X1   g0545(.A1(new_n741), .A2(G190), .A3(G200), .ZN(new_n746));
  INV_X1    g0546(.A(new_n746), .ZN(new_n747));
  INV_X1    g0547(.A(G311), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n285), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n213), .A2(G179), .ZN(new_n750));
  NAND3_X1  g0550(.A1(new_n750), .A2(new_n450), .A3(new_n302), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  AOI211_X1 g0552(.A(new_n745), .B(new_n749), .C1(G329), .C2(new_n752), .ZN(new_n753));
  INV_X1    g0553(.A(new_n741), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G200), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(new_n450), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n756), .A2(G326), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n750), .A2(G190), .A3(G200), .ZN(new_n758));
  INV_X1    g0558(.A(new_n758), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n754), .A2(new_n450), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  XNOR2_X1  g0561(.A(KEYINPUT33), .B(G317), .ZN(new_n762));
  AOI22_X1  g0562(.A1(G303), .A2(new_n759), .B1(new_n761), .B2(new_n762), .ZN(new_n763));
  NOR3_X1   g0563(.A1(new_n450), .A2(G179), .A3(G200), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n764), .A2(new_n213), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g0566(.A1(new_n750), .A2(new_n450), .A3(G200), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  AOI22_X1  g0568(.A1(new_n766), .A2(G294), .B1(new_n768), .B2(G283), .ZN(new_n769));
  NAND4_X1  g0569(.A1(new_n753), .A2(new_n757), .A3(new_n763), .A4(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n743), .A2(new_n399), .ZN(new_n771));
  AOI211_X1 g0571(.A(new_n285), .B(new_n771), .C1(new_n216), .C2(new_n746), .ZN(new_n772));
  INV_X1    g0572(.A(new_n756), .ZN(new_n773));
  OAI22_X1  g0573(.A1(new_n773), .A2(new_n202), .B1(new_n767), .B2(new_n373), .ZN(new_n774));
  OAI22_X1  g0574(.A1(new_n765), .A2(new_n494), .B1(new_n760), .B2(new_n349), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n752), .A2(G159), .ZN(new_n777));
  OR2_X1    g0577(.A1(new_n777), .A2(KEYINPUT32), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n758), .A2(new_n434), .ZN(new_n779));
  AOI21_X1  g0579(.A(new_n779), .B1(new_n777), .B2(KEYINPUT32), .ZN(new_n780));
  NAND4_X1  g0580(.A1(new_n772), .A2(new_n776), .A3(new_n778), .A4(new_n780), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n740), .B1(new_n770), .B2(new_n781), .ZN(new_n782));
  NAND3_X1  g0582(.A1(new_n292), .A2(G355), .A3(new_n207), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n783), .B1(G116), .B2(new_n207), .ZN(new_n784));
  OR2_X1    g0584(.A1(new_n236), .A2(new_n275), .ZN(new_n785));
  NOR2_X1   g0585(.A1(new_n682), .A2(new_n292), .ZN(new_n786));
  INV_X1    g0586(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n211), .B2(new_n275), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n784), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n736), .A2(new_n739), .ZN(new_n790));
  INV_X1    g0590(.A(new_n790), .ZN(new_n791));
  OAI21_X1  g0591(.A(new_n730), .B1(new_n789), .B2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n782), .A2(new_n792), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n731), .A2(new_n733), .B1(new_n738), .B2(new_n793), .ZN(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(G396));
  NAND3_X1  g0595(.A1(new_n382), .A2(new_n393), .A3(new_n661), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n796), .A2(KEYINPUT99), .ZN(new_n797));
  INV_X1    g0597(.A(KEYINPUT99), .ZN(new_n798));
  NAND4_X1  g0598(.A1(new_n382), .A2(new_n393), .A3(new_n798), .A4(new_n661), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n392), .A2(new_n661), .ZN(new_n800));
  AOI22_X1  g0600(.A1(new_n797), .A2(new_n799), .B1(new_n396), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n697), .B(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n730), .B1(new_n803), .B2(new_n724), .ZN(new_n804));
  OAI21_X1  g0604(.A(new_n804), .B1(new_n724), .B2(new_n803), .ZN(new_n805));
  INV_X1    g0605(.A(new_n730), .ZN(new_n806));
  NOR2_X1   g0606(.A1(new_n739), .A2(new_n734), .ZN(new_n807));
  AOI21_X1  g0607(.A(new_n806), .B1(new_n358), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(G283), .ZN(new_n809));
  OAI22_X1  g0609(.A1(new_n758), .A2(new_n373), .B1(new_n760), .B2(new_n809), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n766), .A2(G97), .B1(new_n756), .B2(G303), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n292), .B1(new_n746), .B2(G116), .ZN(new_n812));
  AOI22_X1  g0612(.A1(new_n752), .A2(G311), .B1(new_n742), .B2(G294), .ZN(new_n813));
  NAND3_X1  g0613(.A1(new_n811), .A2(new_n812), .A3(new_n813), .ZN(new_n814));
  AOI211_X1 g0614(.A(new_n810), .B(new_n814), .C1(G87), .C2(new_n768), .ZN(new_n815));
  XNOR2_X1  g0615(.A(new_n815), .B(KEYINPUT97), .ZN(new_n816));
  AOI22_X1  g0616(.A1(G143), .A2(new_n742), .B1(new_n746), .B2(G159), .ZN(new_n817));
  INV_X1    g0617(.A(G150), .ZN(new_n818));
  INV_X1    g0618(.A(G137), .ZN(new_n819));
  OAI221_X1 g0619(.A(new_n817), .B1(new_n818), .B2(new_n760), .C1(new_n773), .C2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n820), .B(KEYINPUT34), .ZN(new_n821));
  INV_X1    g0621(.A(KEYINPUT98), .ZN(new_n822));
  OR2_X1    g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(G132), .ZN(new_n824));
  OAI221_X1 g0624(.A(new_n292), .B1(new_n751), .B2(new_n824), .C1(new_n202), .C2(new_n758), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n768), .A2(G68), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n826), .B1(new_n399), .B2(new_n765), .ZN(new_n827));
  AOI211_X1 g0627(.A(new_n825), .B(new_n827), .C1(new_n821), .C2(new_n822), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n816), .B1(new_n823), .B2(new_n828), .ZN(new_n829));
  OAI221_X1 g0629(.A(new_n808), .B1(new_n829), .B2(new_n740), .C1(new_n802), .C2(new_n735), .ZN(new_n830));
  NAND2_X1  g0630(.A1(new_n805), .A2(new_n830), .ZN(G384));
  INV_X1    g0631(.A(new_n497), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n832), .A2(KEYINPUT35), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n832), .A2(KEYINPUT35), .ZN(new_n834));
  NAND4_X1  g0634(.A1(new_n833), .A2(G116), .A3(new_n214), .A4(new_n834), .ZN(new_n835));
  XOR2_X1   g0635(.A(new_n835), .B(KEYINPUT36), .Z(new_n836));
  OAI211_X1 g0636(.A(new_n216), .B(new_n685), .C1(new_n399), .C2(new_n349), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n202), .A2(G68), .ZN(new_n838));
  AOI211_X1 g0638(.A(new_n262), .B(G13), .C1(new_n837), .C2(new_n838), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n836), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g0640(.A1(new_n690), .A2(new_n698), .A3(new_n457), .A4(new_n705), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n841), .A2(new_n654), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT101), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n645), .A2(new_n662), .ZN(new_n844));
  INV_X1    g0644(.A(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(new_n845), .B1(new_n697), .B2(new_n802), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n365), .A2(new_n661), .ZN(new_n847));
  NAND3_X1  g0647(.A1(new_n366), .A2(new_n370), .A3(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n348), .A2(new_n365), .A3(new_n661), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n846), .A2(new_n851), .ZN(new_n852));
  INV_X1    g0652(.A(KEYINPUT38), .ZN(new_n853));
  INV_X1    g0653(.A(new_n659), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n253), .B1(new_n408), .B2(new_n409), .ZN(new_n855));
  AOI21_X1  g0655(.A(new_n855), .B1(new_n412), .B2(new_n418), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n854), .B1(new_n856), .B2(new_n423), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n651), .B1(KEYINPUT18), .B2(new_n444), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n857), .B1(new_n858), .B2(new_n447), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n424), .A2(new_n433), .A3(new_n854), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT37), .B1(new_n449), .B2(new_n452), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n444), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n443), .B1(new_n856), .B2(new_n423), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n863), .A2(new_n857), .A3(new_n647), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g0665(.A1(new_n862), .A2(new_n865), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI21_X1  g0667(.A(new_n853), .B1(new_n859), .B2(new_n867), .ZN(new_n868));
  INV_X1    g0668(.A(new_n857), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n456), .A2(new_n869), .ZN(new_n870));
  NAND3_X1  g0670(.A1(new_n870), .A2(KEYINPUT38), .A3(new_n866), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n641), .A2(new_n643), .ZN(new_n873));
  AOI22_X1  g0673(.A1(new_n852), .A2(new_n872), .B1(new_n873), .B2(new_n659), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  AND3_X1   g0675(.A1(new_n424), .A2(new_n433), .A3(new_n854), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n649), .A2(new_n650), .A3(KEYINPUT100), .ZN(new_n877));
  NAND2_X1  g0677(.A1(new_n644), .A2(new_n877), .ZN(new_n878));
  AOI21_X1  g0678(.A(KEYINPUT100), .B1(new_n649), .B2(new_n650), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n876), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n647), .B1(new_n449), .B2(new_n640), .ZN(new_n881));
  OAI21_X1  g0681(.A(KEYINPUT37), .B1(new_n876), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g0682(.A1(new_n882), .A2(new_n862), .ZN(new_n883));
  AOI21_X1  g0683(.A(KEYINPUT38), .B1(new_n880), .B2(new_n883), .ZN(new_n884));
  AOI221_X4 g0684(.A(new_n853), .B1(new_n862), .B2(new_n865), .C1(new_n456), .C2(new_n869), .ZN(new_n885));
  OAI21_X1  g0685(.A(new_n875), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  NAND3_X1  g0686(.A1(new_n868), .A2(KEYINPUT39), .A3(new_n871), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n366), .A2(new_n661), .ZN(new_n888));
  NAND3_X1  g0688(.A1(new_n886), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n874), .A2(new_n889), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n843), .B(new_n890), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT40), .ZN(new_n892));
  INV_X1    g0692(.A(KEYINPUT100), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n651), .A2(new_n893), .ZN(new_n894));
  NAND3_X1  g0694(.A1(new_n894), .A2(new_n644), .A3(new_n877), .ZN(new_n895));
  AOI22_X1  g0695(.A1(new_n895), .A2(new_n876), .B1(new_n862), .B2(new_n882), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n871), .B1(new_n896), .B2(KEYINPUT38), .ZN(new_n897));
  AOI21_X1  g0697(.A(new_n801), .B1(new_n848), .B2(new_n849), .ZN(new_n898));
  AND2_X1   g0698(.A1(new_n898), .A2(new_n723), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n892), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NAND3_X1  g0700(.A1(new_n898), .A2(new_n723), .A3(new_n892), .ZN(new_n901));
  AOI21_X1  g0701(.A(new_n901), .B1(new_n868), .B2(new_n871), .ZN(new_n902));
  NOR2_X1   g0702(.A1(new_n900), .A2(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n457), .A2(new_n723), .ZN(new_n904));
  XNOR2_X1  g0704(.A(new_n903), .B(new_n904), .ZN(new_n905));
  NOR2_X1   g0705(.A1(new_n905), .A2(new_n666), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n891), .A2(new_n906), .B1(new_n262), .B2(new_n727), .ZN(new_n907));
  AND2_X1   g0707(.A1(new_n891), .A2(new_n906), .ZN(new_n908));
  OAI21_X1  g0708(.A(new_n840), .B1(new_n907), .B2(new_n908), .ZN(G367));
  OAI221_X1 g0709(.A(new_n790), .B1(new_n207), .B2(new_n384), .C1(new_n232), .C2(new_n787), .ZN(new_n910));
  AND2_X1   g0710(.A1(new_n910), .A2(new_n730), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n594), .A2(new_n662), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n692), .A2(new_n912), .ZN(new_n913));
  OAI21_X1  g0713(.A(new_n913), .B1(new_n634), .B2(new_n912), .ZN(new_n914));
  AOI22_X1  g0714(.A1(new_n768), .A2(G97), .B1(new_n761), .B2(G294), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n915), .B1(new_n373), .B2(new_n765), .C1(new_n748), .C2(new_n773), .ZN(new_n916));
  AOI22_X1  g0716(.A1(new_n752), .A2(G317), .B1(G283), .B2(new_n746), .ZN(new_n917));
  NAND3_X1  g0717(.A1(new_n759), .A2(KEYINPUT46), .A3(G116), .ZN(new_n918));
  INV_X1    g0718(.A(KEYINPUT46), .ZN(new_n919));
  OAI21_X1  g0719(.A(new_n919), .B1(new_n758), .B2(new_n551), .ZN(new_n920));
  AOI21_X1  g0720(.A(new_n292), .B1(new_n565), .B2(new_n742), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n917), .A2(new_n918), .A3(new_n920), .A4(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n292), .B1(new_n743), .B2(new_n818), .ZN(new_n923));
  AOI21_X1  g0723(.A(new_n923), .B1(G137), .B2(new_n752), .ZN(new_n924));
  AOI22_X1  g0724(.A1(G143), .A2(new_n756), .B1(new_n759), .B2(G58), .ZN(new_n925));
  AOI22_X1  g0725(.A1(new_n766), .A2(G68), .B1(new_n768), .B2(new_n216), .ZN(new_n926));
  NAND3_X1  g0726(.A1(new_n924), .A2(new_n925), .A3(new_n926), .ZN(new_n927));
  INV_X1    g0727(.A(G159), .ZN(new_n928));
  OAI22_X1  g0728(.A1(new_n747), .A2(new_n202), .B1(new_n760), .B2(new_n928), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(KEYINPUT105), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n916), .A2(new_n922), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  XOR2_X1   g0731(.A(new_n931), .B(KEYINPUT47), .Z(new_n932));
  OAI221_X1 g0732(.A(new_n911), .B1(new_n914), .B2(new_n737), .C1(new_n740), .C2(new_n932), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n507), .A2(new_n661), .ZN(new_n934));
  NAND3_X1  g0734(.A1(new_n509), .A2(new_n513), .A3(new_n934), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n512), .A2(new_n661), .ZN(new_n936));
  NAND3_X1  g0736(.A1(new_n935), .A2(new_n936), .A3(new_n677), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  AND2_X1   g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NOR2_X1   g0739(.A1(new_n937), .A2(new_n938), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n935), .A2(new_n936), .ZN(new_n941));
  AOI21_X1  g0741(.A(KEYINPUT45), .B1(new_n941), .B2(new_n678), .ZN(new_n942));
  INV_X1    g0742(.A(KEYINPUT45), .ZN(new_n943));
  AOI211_X1 g0743(.A(new_n943), .B(new_n677), .C1(new_n935), .C2(new_n936), .ZN(new_n944));
  OAI22_X1  g0744(.A1(new_n939), .A2(new_n940), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  INV_X1    g0745(.A(new_n674), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n668), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  OAI221_X1 g0748(.A(new_n675), .B1(new_n942), .B2(new_n944), .C1(new_n939), .C2(new_n940), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT104), .ZN(new_n951));
  INV_X1    g0751(.A(new_n676), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n674), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n946), .A2(new_n676), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n669), .A2(new_n951), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n954), .A2(new_n953), .ZN(new_n956));
  OAI21_X1  g0756(.A(KEYINPUT104), .B1(new_n668), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n955), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n668), .A2(new_n956), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n959), .A2(KEYINPUT103), .ZN(new_n960));
  INV_X1    g0760(.A(KEYINPUT103), .ZN(new_n961));
  NAND3_X1  g0761(.A1(new_n668), .A2(new_n956), .A3(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n960), .A2(new_n962), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n958), .A2(new_n963), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n725), .B1(new_n950), .B2(new_n964), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n683), .B(KEYINPUT41), .Z(new_n966));
  INV_X1    g0766(.A(new_n966), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n729), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n947), .A2(new_n941), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT102), .ZN(new_n970));
  XNOR2_X1  g0770(.A(new_n969), .B(new_n970), .ZN(new_n971));
  AND2_X1   g0771(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT42), .ZN(new_n973));
  INV_X1    g0773(.A(new_n953), .ZN(new_n974));
  AOI21_X1  g0774(.A(new_n973), .B1(new_n941), .B2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n548), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n509), .A2(new_n513), .A3(new_n976), .A4(new_n934), .ZN(new_n977));
  AOI21_X1  g0777(.A(new_n661), .B1(new_n977), .B2(new_n513), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n975), .A2(new_n978), .ZN(new_n979));
  NAND3_X1  g0779(.A1(new_n941), .A2(new_n973), .A3(new_n974), .ZN(new_n980));
  AOI21_X1  g0780(.A(new_n972), .B1(new_n979), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g0781(.A1(new_n914), .A2(KEYINPUT43), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n982), .ZN(new_n984));
  INV_X1    g0784(.A(new_n980), .ZN(new_n985));
  NOR3_X1   g0785(.A1(new_n985), .A2(new_n975), .A3(new_n978), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n984), .B1(new_n986), .B2(new_n972), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n971), .A2(new_n983), .A3(new_n987), .ZN(new_n988));
  AND2_X1   g0788(.A1(new_n983), .A2(new_n987), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT102), .B1(new_n947), .B2(new_n941), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n933), .B1(new_n968), .B2(new_n991), .ZN(G387));
  NAND3_X1  g0792(.A1(new_n681), .A2(new_n207), .A3(new_n292), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n993), .B1(G107), .B2(new_n207), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT106), .Z(new_n995));
  NAND2_X1  g0795(.A1(new_n387), .A2(new_n202), .ZN(new_n996));
  XNOR2_X1  g0796(.A(new_n996), .B(KEYINPUT50), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n275), .B1(new_n349), .B2(new_n358), .ZN(new_n998));
  NOR3_X1   g0798(.A1(new_n997), .A2(new_n681), .A3(new_n998), .ZN(new_n999));
  OAI21_X1  g0799(.A(new_n786), .B1(new_n229), .B2(new_n275), .ZN(new_n1000));
  OAI21_X1  g0800(.A(new_n995), .B1(new_n999), .B2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g0801(.A(new_n806), .B1(new_n1001), .B2(new_n790), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(G159), .A2(new_n756), .B1(new_n759), .B2(new_n216), .ZN(new_n1003));
  OAI221_X1 g0803(.A(new_n1003), .B1(new_n494), .B2(new_n767), .C1(new_n246), .C2(new_n760), .ZN(new_n1004));
  OAI22_X1  g0804(.A1(new_n765), .A2(new_n384), .B1(new_n743), .B2(new_n202), .ZN(new_n1005));
  XNOR2_X1  g0805(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n292), .B1(new_n751), .B2(new_n818), .C1(new_n747), .C2(new_n349), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n1004), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(new_n766), .A2(G283), .B1(new_n759), .B2(G294), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(new_n565), .A2(new_n746), .B1(new_n742), .B2(G317), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1010), .B1(new_n748), .B2(new_n760), .C1(new_n773), .C2(new_n744), .ZN(new_n1011));
  INV_X1    g0811(.A(KEYINPUT48), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1009), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT108), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n1014), .B1(new_n1012), .B2(new_n1011), .ZN(new_n1015));
  OR2_X1    g0815(.A1(new_n1015), .A2(KEYINPUT49), .ZN(new_n1016));
  AOI21_X1  g0816(.A(new_n292), .B1(new_n752), .B2(G326), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1017), .B1(new_n551), .B2(new_n767), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n1015), .B2(KEYINPUT49), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1008), .B1(new_n1016), .B2(new_n1019), .ZN(new_n1020));
  OAI221_X1 g0820(.A(new_n1002), .B1(new_n674), .B2(new_n737), .C1(new_n1020), .C2(new_n740), .ZN(new_n1021));
  AOI22_X1  g0821(.A1(new_n955), .A2(new_n957), .B1(new_n960), .B2(new_n962), .ZN(new_n1022));
  NAND3_X1  g0822(.A1(new_n1022), .A2(new_n706), .A3(new_n724), .ZN(new_n1023));
  NAND2_X1  g0823(.A1(new_n1023), .A2(new_n683), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n725), .A2(new_n1022), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n1021), .B1(new_n728), .B2(new_n964), .C1(new_n1024), .C2(new_n1025), .ZN(G393));
  NAND3_X1  g0826(.A1(new_n948), .A2(new_n949), .A3(new_n729), .ZN(new_n1027));
  OAI221_X1 g0827(.A(new_n790), .B1(new_n494), .B2(new_n207), .C1(new_n239), .C2(new_n787), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n1028), .A2(new_n730), .ZN(new_n1029));
  AOI22_X1  g0829(.A1(new_n756), .A2(G150), .B1(G159), .B2(new_n742), .ZN(new_n1030));
  XNOR2_X1  g0830(.A(new_n1030), .B(KEYINPUT51), .ZN(new_n1031));
  AOI22_X1  g0831(.A1(G68), .A2(new_n759), .B1(new_n752), .B2(G143), .ZN(new_n1032));
  XOR2_X1   g0832(.A(new_n1032), .B(KEYINPUT109), .Z(new_n1033));
  OAI221_X1 g0833(.A(new_n292), .B1(new_n767), .B2(new_n434), .C1(new_n747), .C2(new_n246), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n765), .A2(new_n358), .B1(new_n760), .B2(new_n202), .ZN(new_n1035));
  OR4_X1    g0835(.A1(new_n1031), .A2(new_n1033), .A3(new_n1034), .A4(new_n1035), .ZN(new_n1036));
  OR2_X1    g0836(.A1(new_n1036), .A2(KEYINPUT110), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(new_n756), .A2(G317), .B1(G311), .B2(new_n742), .ZN(new_n1038));
  XOR2_X1   g0838(.A(new_n1038), .B(KEYINPUT52), .Z(new_n1039));
  OAI21_X1  g0839(.A(new_n285), .B1(new_n751), .B2(new_n744), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n1040), .B1(G294), .B2(new_n746), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G107), .A2(new_n768), .B1(new_n761), .B2(new_n565), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(new_n766), .A2(G116), .B1(new_n759), .B2(G283), .ZN(new_n1043));
  NAND4_X1  g0843(.A1(new_n1039), .A2(new_n1041), .A3(new_n1042), .A4(new_n1043), .ZN(new_n1044));
  NAND2_X1  g0844(.A1(new_n1036), .A2(KEYINPUT110), .ZN(new_n1045));
  NAND3_X1  g0845(.A1(new_n1037), .A2(new_n1044), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1029), .B1(new_n1046), .B2(new_n739), .ZN(new_n1047));
  OAI21_X1  g0847(.A(new_n1047), .B1(new_n941), .B2(new_n737), .ZN(new_n1048));
  NAND3_X1  g0848(.A1(new_n1027), .A2(KEYINPUT111), .A3(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  AOI21_X1  g0850(.A(KEYINPUT111), .B1(new_n1027), .B2(new_n1048), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1023), .A2(new_n950), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n683), .B1(new_n1023), .B2(new_n950), .ZN(new_n1054));
  OAI22_X1  g0854(.A1(new_n1050), .A2(new_n1051), .B1(new_n1053), .B2(new_n1054), .ZN(G390));
  NAND2_X1  g0855(.A1(new_n886), .A2(new_n887), .ZN(new_n1056));
  AOI211_X1 g0856(.A(new_n661), .B(new_n801), .C1(new_n695), .C2(new_n696), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n850), .B1(new_n1057), .B2(new_n845), .ZN(new_n1058));
  INV_X1    g0858(.A(new_n888), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  OAI211_X1 g0861(.A(new_n662), .B(new_n802), .C1(new_n704), .C2(new_n637), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1062), .A2(new_n844), .ZN(new_n1063));
  OAI211_X1 g0863(.A(new_n1059), .B(new_n897), .C1(new_n1063), .C2(new_n851), .ZN(new_n1064));
  NAND3_X1  g0864(.A1(new_n723), .A2(new_n667), .A3(new_n802), .ZN(new_n1065));
  OR2_X1    g0865(.A1(new_n1065), .A2(new_n851), .ZN(new_n1066));
  NAND3_X1  g0866(.A1(new_n1061), .A2(new_n1064), .A3(new_n1066), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n898), .A2(new_n723), .A3(G330), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1068), .A2(KEYINPUT112), .ZN(new_n1069));
  INV_X1    g0869(.A(KEYINPUT112), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n898), .A2(new_n723), .A3(new_n1070), .A4(G330), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  AOI22_X1  g0872(.A1(new_n886), .A2(new_n887), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1059), .B1(new_n884), .B2(new_n885), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n851), .B1(new_n1062), .B2(new_n844), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n1072), .B1(new_n1073), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n1067), .A2(new_n1077), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1078), .A2(new_n728), .ZN(new_n1079));
  NAND2_X1  g0879(.A1(new_n1056), .A2(new_n734), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n807), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n730), .B1(new_n1081), .B2(new_n387), .ZN(new_n1082));
  INV_X1    g0882(.A(G294), .ZN(new_n1083));
  OAI21_X1  g0883(.A(new_n826), .B1(new_n1083), .B2(new_n751), .ZN(new_n1084));
  XOR2_X1   g0884(.A(new_n1084), .B(KEYINPUT114), .Z(new_n1085));
  OAI22_X1  g0885(.A1(new_n773), .A2(new_n809), .B1(new_n373), .B2(new_n760), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n779), .B(new_n1086), .C1(G77), .C2(new_n766), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n285), .B1(new_n743), .B2(new_n551), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n1088), .B1(G97), .B2(new_n746), .ZN(new_n1089));
  NAND3_X1  g0889(.A1(new_n1085), .A2(new_n1087), .A3(new_n1089), .ZN(new_n1090));
  XNOR2_X1  g0890(.A(KEYINPUT54), .B(G143), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  AOI22_X1  g0892(.A1(new_n761), .A2(G137), .B1(new_n1092), .B2(new_n746), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(new_n1093), .B(KEYINPUT113), .ZN(new_n1094));
  INV_X1    g0894(.A(G125), .ZN(new_n1095));
  OAI221_X1 g0895(.A(new_n292), .B1(new_n751), .B2(new_n1095), .C1(new_n743), .C2(new_n824), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n759), .A2(G150), .ZN(new_n1097));
  AOI21_X1  g0897(.A(new_n1096), .B1(KEYINPUT53), .B2(new_n1097), .ZN(new_n1098));
  OAI22_X1  g0898(.A1(new_n765), .A2(new_n928), .B1(new_n767), .B2(new_n202), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n1099), .B1(G128), .B2(new_n756), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n1098), .B(new_n1100), .C1(KEYINPUT53), .C2(new_n1097), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1090), .B1(new_n1094), .B2(new_n1101), .ZN(new_n1102));
  AOI21_X1  g0902(.A(new_n1082), .B1(new_n1102), .B2(new_n739), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1079), .B1(new_n1080), .B2(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n723), .A2(G330), .ZN(new_n1105));
  INV_X1    g0905(.A(new_n1105), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n1106), .A2(new_n457), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n841), .A2(new_n654), .A3(new_n1107), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n1065), .A2(new_n851), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1069), .A2(new_n1109), .A3(new_n1071), .ZN(new_n1110));
  INV_X1    g0910(.A(new_n846), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1110), .A2(new_n1111), .ZN(new_n1112));
  OAI21_X1  g0912(.A(new_n851), .B1(new_n1105), .B2(new_n801), .ZN(new_n1113));
  NAND3_X1  g0913(.A1(new_n1066), .A2(new_n1063), .A3(new_n1113), .ZN(new_n1114));
  NAND2_X1  g0914(.A1(new_n1112), .A2(new_n1114), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n1115), .ZN(new_n1116));
  OAI21_X1  g0916(.A(new_n1078), .B1(new_n1108), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1108), .B1(new_n1112), .B2(new_n1114), .ZN(new_n1118));
  NAND3_X1  g0918(.A1(new_n1118), .A2(new_n1067), .A3(new_n1077), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n1117), .A2(new_n683), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1104), .A2(new_n1120), .ZN(G378));
  INV_X1    g0921(.A(KEYINPUT117), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n267), .A2(new_n659), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n315), .A2(new_n1124), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n301), .ZN(new_n1126));
  INV_X1    g0926(.A(new_n314), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1126), .B1(new_n1127), .B2(new_n312), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1129));
  XNOR2_X1  g0929(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1130));
  AND3_X1   g0930(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1130), .B1(new_n1125), .B2(new_n1129), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1122), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1130), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n315), .A2(new_n1124), .ZN(new_n1135));
  NOR2_X1   g0935(.A1(new_n1128), .A2(new_n1123), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1134), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND3_X1  g0937(.A1(new_n1125), .A2(new_n1129), .A3(new_n1130), .ZN(new_n1138));
  NAND3_X1  g0938(.A1(new_n1137), .A2(KEYINPUT117), .A3(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1133), .A2(new_n1139), .ZN(new_n1140));
  OAI211_X1 g0940(.A(new_n1140), .B(G330), .C1(new_n900), .C2(new_n902), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  NOR2_X1   g0942(.A1(new_n1131), .A2(new_n1132), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(KEYINPUT38), .B1(new_n870), .B2(new_n866), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n899), .B(new_n892), .C1(new_n885), .C2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n898), .A2(new_n723), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n873), .B1(new_n455), .B2(KEYINPUT100), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n860), .B1(new_n1148), .B2(new_n894), .ZN(new_n1149));
  AND2_X1   g0949(.A1(new_n882), .A2(new_n862), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n853), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1147), .B1(new_n1151), .B2(new_n871), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1146), .B1(new_n1152), .B2(new_n892), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1144), .B1(new_n1153), .B2(G330), .ZN(new_n1154));
  OAI21_X1  g0954(.A(new_n890), .B1(new_n1142), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT119), .ZN(new_n1156));
  INV_X1    g0956(.A(G330), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1143), .B1(new_n903), .B2(new_n1157), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n890), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1158), .A2(new_n1159), .A3(new_n1141), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1155), .A2(new_n1156), .A3(new_n1160), .ZN(new_n1161));
  INV_X1    g0961(.A(KEYINPUT57), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n1108), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1162), .B1(new_n1119), .B2(new_n1163), .ZN(new_n1164));
  OAI211_X1 g0964(.A(KEYINPUT119), .B(new_n890), .C1(new_n1142), .C2(new_n1154), .ZN(new_n1165));
  NAND3_X1  g0965(.A1(new_n1161), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(KEYINPUT120), .ZN(new_n1167));
  INV_X1    g0967(.A(KEYINPUT120), .ZN(new_n1168));
  NAND4_X1  g0968(.A1(new_n1161), .A2(new_n1164), .A3(new_n1168), .A4(new_n1165), .ZN(new_n1169));
  NAND2_X1  g0969(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1170));
  AOI22_X1  g0970(.A1(new_n1155), .A2(new_n1160), .B1(new_n1119), .B2(new_n1163), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n683), .B1(new_n1171), .B2(KEYINPUT57), .ZN(new_n1172));
  INV_X1    g0972(.A(new_n1172), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1170), .A2(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n728), .B1(new_n1155), .B2(new_n1160), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n806), .B1(new_n202), .B2(new_n807), .ZN(new_n1176));
  NOR2_X1   g0976(.A1(new_n292), .A2(G41), .ZN(new_n1177));
  OAI21_X1  g0977(.A(new_n1177), .B1(new_n809), .B2(new_n751), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n767), .A2(new_n399), .ZN(new_n1179));
  XNOR2_X1  g0979(.A(new_n1179), .B(KEYINPUT115), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1178), .B(new_n1180), .C1(new_n216), .C2(new_n759), .ZN(new_n1181));
  XNOR2_X1  g0981(.A(new_n1181), .B(KEYINPUT116), .ZN(new_n1182));
  OAI22_X1  g0982(.A1(new_n373), .A2(new_n743), .B1(new_n747), .B2(new_n384), .ZN(new_n1183));
  AOI21_X1  g0983(.A(new_n1183), .B1(G68), .B2(new_n766), .ZN(new_n1184));
  AOI22_X1  g0984(.A1(G116), .A2(new_n756), .B1(new_n761), .B2(G97), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n1182), .A2(new_n1184), .A3(new_n1185), .ZN(new_n1186));
  INV_X1    g0986(.A(KEYINPUT58), .ZN(new_n1187));
  OR2_X1    g0987(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(G33), .A2(G41), .ZN(new_n1190));
  NOR3_X1   g0990(.A1(new_n1177), .A2(G50), .A3(new_n1190), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n773), .A2(new_n1095), .B1(new_n824), .B2(new_n760), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n1192), .B1(G150), .B2(new_n766), .ZN(new_n1193));
  AOI22_X1  g0993(.A1(G128), .A2(new_n742), .B1(new_n746), .B2(G137), .ZN(new_n1194));
  OAI211_X1 g0994(.A(new_n1193), .B(new_n1194), .C1(new_n758), .C2(new_n1091), .ZN(new_n1195));
  OR2_X1    g0995(.A1(new_n1195), .A2(KEYINPUT59), .ZN(new_n1196));
  INV_X1    g0996(.A(G124), .ZN(new_n1197));
  OAI221_X1 g0997(.A(new_n1190), .B1(new_n751), .B2(new_n1197), .C1(new_n928), .C2(new_n767), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(new_n1195), .B2(KEYINPUT59), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n1191), .B1(new_n1196), .B2(new_n1199), .ZN(new_n1200));
  AND3_X1   g1000(.A1(new_n1188), .A2(new_n1189), .A3(new_n1200), .ZN(new_n1201));
  OAI221_X1 g1001(.A(new_n1176), .B1(new_n740), .B2(new_n1201), .C1(new_n1140), .C2(new_n735), .ZN(new_n1202));
  XNOR2_X1  g1002(.A(new_n1202), .B(KEYINPUT118), .ZN(new_n1203));
  NOR2_X1   g1003(.A1(new_n1175), .A2(new_n1203), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1174), .A2(new_n1204), .ZN(G375));
  AOI21_X1  g1005(.A(new_n806), .B1(new_n349), .B2(new_n807), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n752), .A2(G303), .B1(new_n742), .B2(G283), .ZN(new_n1207));
  OAI211_X1 g1007(.A(new_n1207), .B(new_n285), .C1(new_n373), .C2(new_n747), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n773), .A2(new_n1083), .B1(new_n767), .B2(new_n358), .ZN(new_n1209));
  NOR2_X1   g1009(.A1(new_n758), .A2(new_n494), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n765), .A2(new_n384), .B1(new_n760), .B2(new_n551), .ZN(new_n1211));
  NOR4_X1   g1011(.A1(new_n1208), .A2(new_n1209), .A3(new_n1210), .A4(new_n1211), .ZN(new_n1212));
  AOI22_X1  g1012(.A1(G128), .A2(new_n752), .B1(new_n759), .B2(G159), .ZN(new_n1213));
  XNOR2_X1  g1013(.A(new_n1213), .B(KEYINPUT121), .ZN(new_n1214));
  AOI22_X1  g1014(.A1(new_n766), .A2(G50), .B1(new_n761), .B2(new_n1092), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n824), .B2(new_n773), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n292), .B1(new_n747), .B2(new_n818), .C1(new_n819), .C2(new_n743), .ZN(new_n1217));
  NOR3_X1   g1017(.A1(new_n1216), .A2(new_n1180), .A3(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1212), .B1(new_n1214), .B2(new_n1218), .ZN(new_n1219));
  OAI221_X1 g1019(.A(new_n1206), .B1(new_n740), .B2(new_n1219), .C1(new_n850), .C2(new_n735), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1220), .B1(new_n1116), .B2(new_n728), .ZN(new_n1221));
  NOR2_X1   g1021(.A1(new_n1118), .A2(new_n966), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1116), .A2(new_n1108), .ZN(new_n1223));
  AOI21_X1  g1023(.A(new_n1221), .B1(new_n1222), .B2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n1224), .ZN(G381));
  INV_X1    g1025(.A(new_n1051), .ZN(new_n1226));
  INV_X1    g1026(.A(new_n683), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n950), .ZN(new_n1228));
  AND4_X1   g1028(.A1(new_n724), .A2(new_n706), .A3(new_n958), .A4(new_n963), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1227), .B1(new_n1228), .B2(new_n1229), .ZN(new_n1230));
  AOI22_X1  g1030(.A1(new_n1226), .A2(new_n1049), .B1(new_n1230), .B2(new_n1052), .ZN(new_n1231));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G396), .A2(G381), .A3(new_n1233), .A4(G393), .ZN(new_n1234));
  NOR4_X1   g1034(.A1(G375), .A2(G387), .A3(new_n1234), .A4(G378), .ZN(new_n1235));
  XNOR2_X1  g1035(.A(new_n1235), .B(KEYINPUT122), .ZN(G407));
  NAND2_X1  g1036(.A1(new_n660), .A2(G213), .ZN(new_n1237));
  NOR3_X1   g1037(.A1(G375), .A2(G378), .A3(new_n1237), .ZN(new_n1238));
  XOR2_X1   g1038(.A(new_n1238), .B(KEYINPUT123), .Z(new_n1239));
  NAND3_X1  g1039(.A1(new_n1239), .A2(G407), .A3(G213), .ZN(G409));
  XNOR2_X1  g1040(.A(G393), .B(new_n794), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n988), .ZN(new_n1242));
  AOI22_X1  g1042(.A1(new_n983), .A2(new_n987), .B1(new_n970), .B2(new_n969), .ZN(new_n1243));
  NOR2_X1   g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n725), .A2(new_n1022), .A3(new_n949), .A4(new_n948), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n966), .B1(new_n1245), .B2(new_n725), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1244), .B1(new_n1246), .B2(new_n729), .ZN(new_n1247));
  AOI21_X1  g1047(.A(G390), .B1(new_n1247), .B2(new_n933), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(G387), .A2(new_n1231), .ZN(new_n1249));
  NOR3_X1   g1049(.A1(new_n1241), .A2(new_n1248), .A3(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(KEYINPUT126), .B1(G387), .B2(new_n1231), .ZN(new_n1251));
  INV_X1    g1051(.A(KEYINPUT126), .ZN(new_n1252));
  NAND4_X1  g1052(.A1(new_n1247), .A2(new_n1252), .A3(new_n933), .A4(G390), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(G387), .A2(new_n1231), .ZN(new_n1254));
  NAND3_X1  g1054(.A1(new_n1251), .A2(new_n1253), .A3(new_n1254), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1241), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(KEYINPUT127), .ZN(new_n1257));
  INV_X1    g1057(.A(KEYINPUT127), .ZN(new_n1258));
  NAND3_X1  g1058(.A1(new_n1255), .A2(new_n1258), .A3(new_n1241), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1250), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n1172), .B1(new_n1167), .B2(new_n1169), .ZN(new_n1261));
  INV_X1    g1061(.A(G378), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n1204), .ZN(new_n1263));
  NOR3_X1   g1063(.A1(new_n1261), .A2(new_n1262), .A3(new_n1263), .ZN(new_n1264));
  INV_X1    g1064(.A(new_n1202), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1265), .B1(new_n1171), .B2(new_n967), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n1161), .A2(new_n729), .A3(new_n1165), .ZN(new_n1267));
  AOI21_X1  g1067(.A(G378), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1237), .B1(new_n1264), .B2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT60), .ZN(new_n1270));
  OAI21_X1  g1070(.A(new_n1223), .B1(new_n1270), .B2(new_n1118), .ZN(new_n1271));
  NOR3_X1   g1071(.A1(new_n1115), .A2(new_n1163), .A3(new_n1270), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1272), .A2(new_n1227), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1221), .B1(new_n1271), .B2(new_n1273), .ZN(new_n1274));
  NOR2_X1   g1074(.A1(new_n1274), .A2(G384), .ZN(new_n1275));
  AOI211_X1 g1075(.A(new_n1232), .B(new_n1221), .C1(new_n1271), .C2(new_n1273), .ZN(new_n1276));
  NOR3_X1   g1076(.A1(new_n1275), .A2(new_n1276), .A3(KEYINPUT125), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1237), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1275), .A2(new_n1276), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT125), .ZN(new_n1280));
  OAI211_X1 g1080(.A(G2897), .B(new_n1278), .C1(new_n1279), .C2(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1278), .A2(G2897), .ZN(new_n1282));
  OAI211_X1 g1082(.A(KEYINPUT125), .B(new_n1282), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1277), .B1(new_n1281), .B2(new_n1283), .ZN(new_n1284));
  AOI211_X1 g1084(.A(KEYINPUT61), .B(new_n1260), .C1(new_n1269), .C2(new_n1284), .ZN(new_n1285));
  OAI211_X1 g1085(.A(new_n1237), .B(new_n1279), .C1(new_n1264), .C2(new_n1268), .ZN(new_n1286));
  INV_X1    g1086(.A(KEYINPUT63), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1286), .A2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1288), .A2(KEYINPUT124), .ZN(new_n1289));
  NAND3_X1  g1089(.A1(new_n1174), .A2(G378), .A3(new_n1204), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1268), .ZN(new_n1291));
  AOI21_X1  g1091(.A(new_n1278), .B1(new_n1290), .B2(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(new_n1292), .A2(KEYINPUT63), .A3(new_n1279), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT124), .ZN(new_n1294));
  NAND3_X1  g1094(.A1(new_n1286), .A2(new_n1294), .A3(new_n1287), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1285), .A2(new_n1289), .A3(new_n1293), .A4(new_n1295), .ZN(new_n1296));
  AOI21_X1  g1096(.A(KEYINPUT61), .B1(new_n1269), .B2(new_n1284), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT62), .ZN(new_n1298));
  NAND3_X1  g1098(.A1(new_n1292), .A2(new_n1298), .A3(new_n1279), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1286), .A2(KEYINPUT62), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1297), .A2(new_n1299), .A3(new_n1300), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n1260), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1296), .A2(new_n1302), .ZN(G405));
  NAND2_X1  g1103(.A1(G375), .A2(new_n1262), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n1290), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1305), .A2(new_n1279), .ZN(new_n1306));
  OAI211_X1 g1106(.A(new_n1304), .B(new_n1290), .C1(new_n1275), .C2(new_n1276), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1306), .A2(new_n1307), .ZN(new_n1308));
  XNOR2_X1  g1108(.A(new_n1308), .B(new_n1260), .ZN(G402));
endmodule


