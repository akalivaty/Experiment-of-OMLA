

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599,
         n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
         n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, n654,
         n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665,
         n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
         n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687,
         n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698,
         n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
         n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720,
         n721, n722, n723, n724, n725, n726, n727, n728, n729, n730, n731,
         n732, n733, n734, n735, n736, n737, n738, n739, n740, n741, n742,
         n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
         n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764,
         n765, n766, n767, n768, n769;

  INV_X1 U368 ( .A(n581), .ZN(n407) );
  INV_X1 U369 ( .A(n655), .ZN(n686) );
  XNOR2_X2 U370 ( .A(n568), .B(n567), .ZN(n696) );
  XNOR2_X2 U371 ( .A(n603), .B(KEYINPUT45), .ZN(n665) );
  OR2_X1 U372 ( .A1(n486), .A2(n434), .ZN(n435) );
  AND2_X1 U373 ( .A1(n367), .A2(n382), .ZN(n360) );
  NOR2_X1 U374 ( .A1(n602), .A2(n601), .ZN(n603) );
  NAND2_X1 U375 ( .A1(n664), .A2(n663), .ZN(n734) );
  XNOR2_X1 U376 ( .A(n400), .B(n355), .ZN(n664) );
  OR2_X1 U377 ( .A1(n594), .A2(n593), .ZN(n597) );
  NOR2_X1 U378 ( .A1(n641), .A2(n640), .ZN(n693) );
  XNOR2_X1 U379 ( .A(n363), .B(n564), .ZN(n572) );
  NAND2_X1 U380 ( .A1(n408), .A2(n405), .ZN(n675) );
  NAND2_X1 U381 ( .A1(n413), .A2(n415), .ZN(n617) );
  AND2_X2 U382 ( .A1(n562), .A2(n561), .ZN(n575) );
  INV_X1 U383 ( .A(n417), .ZN(n413) );
  BUF_X1 U384 ( .A(n541), .Z(n638) );
  XNOR2_X1 U385 ( .A(n453), .B(n452), .ZN(n541) );
  XNOR2_X1 U386 ( .A(n361), .B(n503), .ZN(n752) );
  XNOR2_X1 U387 ( .A(n435), .B(n436), .ZN(n439) );
  NAND2_X1 U388 ( .A1(n666), .A2(KEYINPUT86), .ZN(n382) );
  XNOR2_X1 U389 ( .A(n440), .B(G128), .ZN(n484) );
  XNOR2_X2 U390 ( .A(KEYINPUT64), .B(G953), .ZN(n486) );
  XNOR2_X1 U391 ( .A(KEYINPUT82), .B(G143), .ZN(n440) );
  INV_X1 U392 ( .A(G237), .ZN(n450) );
  NAND2_X1 U393 ( .A1(n410), .A2(n349), .ZN(n565) );
  NAND2_X1 U394 ( .A1(n413), .A2(n411), .ZN(n410) );
  XOR2_X1 U395 ( .A(KEYINPUT84), .B(KEYINPUT8), .Z(n488) );
  NAND2_X1 U396 ( .A1(n750), .A2(G475), .ZN(n389) );
  AND2_X1 U397 ( .A1(n523), .A2(n420), .ZN(n416) );
  NOR2_X1 U398 ( .A1(n763), .A2(G237), .ZN(n512) );
  XNOR2_X1 U399 ( .A(G146), .B(G125), .ZN(n476) );
  XNOR2_X1 U400 ( .A(n458), .B(n457), .ZN(n648) );
  XNOR2_X1 U401 ( .A(n481), .B(n480), .ZN(n569) );
  XNOR2_X1 U402 ( .A(n527), .B(n526), .ZN(n756) );
  NOR2_X1 U403 ( .A1(n486), .A2(n528), .ZN(n372) );
  AND2_X1 U404 ( .A1(n643), .A2(n362), .ZN(n624) );
  INV_X1 U405 ( .A(KEYINPUT110), .ZN(n428) );
  NAND2_X1 U406 ( .A1(n565), .A2(n675), .ZN(n552) );
  NAND2_X1 U407 ( .A1(n642), .A2(n714), .ZN(n426) );
  INV_X1 U408 ( .A(n569), .ZN(n582) );
  XNOR2_X1 U409 ( .A(n498), .B(n497), .ZN(n536) );
  XNOR2_X1 U410 ( .A(n530), .B(n576), .ZN(n531) );
  XNOR2_X1 U411 ( .A(n422), .B(n421), .ZN(n431) );
  AND2_X2 U412 ( .A1(n398), .A2(n381), .ZN(n750) );
  NOR2_X1 U413 ( .A1(n369), .A2(n364), .ZN(n381) );
  NAND2_X1 U414 ( .A1(n750), .A2(G210), .ZN(n394) );
  NAND2_X1 U415 ( .A1(n419), .A2(n418), .ZN(n417) );
  NAND2_X1 U416 ( .A1(G902), .A2(G472), .ZN(n418) );
  OR2_X1 U417 ( .A1(n674), .A2(n420), .ZN(n419) );
  NOR2_X1 U418 ( .A1(n412), .A2(n534), .ZN(n411) );
  XNOR2_X1 U419 ( .A(G113), .B(G122), .ZN(n472) );
  XNOR2_X1 U420 ( .A(G143), .B(G131), .ZN(n470) );
  XOR2_X1 U421 ( .A(G104), .B(G140), .Z(n471) );
  INV_X1 U422 ( .A(KEYINPUT86), .ZN(n383) );
  NAND2_X1 U423 ( .A1(n734), .A2(n354), .ZN(n367) );
  XNOR2_X1 U424 ( .A(KEYINPUT79), .B(KEYINPUT18), .ZN(n437) );
  NAND2_X1 U425 ( .A1(G234), .A2(G237), .ZN(n459) );
  OR2_X1 U426 ( .A1(n569), .A2(n581), .ZN(n433) );
  NAND2_X1 U427 ( .A1(n563), .A2(n575), .ZN(n363) );
  XNOR2_X1 U428 ( .A(G134), .B(G131), .ZN(n524) );
  XOR2_X1 U429 ( .A(KEYINPUT5), .B(G116), .Z(n514) );
  XNOR2_X1 U430 ( .A(G137), .B(G101), .ZN(n515) );
  XOR2_X1 U431 ( .A(KEYINPUT76), .B(G146), .Z(n516) );
  XNOR2_X1 U432 ( .A(G113), .B(KEYINPUT70), .ZN(n446) );
  XNOR2_X1 U433 ( .A(n423), .B(KEYINPUT7), .ZN(n422) );
  XNOR2_X1 U434 ( .A(KEYINPUT9), .B(KEYINPUT102), .ZN(n423) );
  XNOR2_X1 U435 ( .A(G134), .B(G107), .ZN(n421) );
  INV_X1 U436 ( .A(n734), .ZN(n366) );
  INV_X1 U437 ( .A(KEYINPUT2), .ZN(n399) );
  BUF_X1 U438 ( .A(n696), .Z(n724) );
  INV_X1 U439 ( .A(n714), .ZN(n425) );
  NAND2_X1 U440 ( .A1(n648), .A2(n465), .ZN(n466) );
  NOR2_X1 U441 ( .A1(n622), .A2(n621), .ZN(n643) );
  NAND2_X1 U442 ( .A1(n575), .A2(n620), .ZN(n621) );
  XNOR2_X1 U443 ( .A(n502), .B(n505), .ZN(n361) );
  XNOR2_X1 U444 ( .A(n501), .B(n432), .ZN(n502) );
  XNOR2_X1 U445 ( .A(n756), .B(n370), .ZN(n670) );
  XNOR2_X1 U446 ( .A(n372), .B(n350), .ZN(n371) );
  BUF_X1 U447 ( .A(G953), .Z(n763) );
  INV_X1 U448 ( .A(n639), .ZN(n640) );
  XNOR2_X1 U449 ( .A(n424), .B(KEYINPUT36), .ZN(n641) );
  OR2_X1 U450 ( .A1(n427), .A2(n426), .ZN(n424) );
  INV_X1 U451 ( .A(n644), .ZN(n571) );
  AND2_X1 U452 ( .A1(n538), .A2(n535), .ZN(n430) );
  AND2_X1 U453 ( .A1(n409), .A2(n406), .ZN(n405) );
  NAND2_X1 U454 ( .A1(n582), .A2(KEYINPUT109), .ZN(n409) );
  NAND2_X1 U455 ( .A1(n396), .A2(n392), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n397), .B(n357), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n386), .B(n385), .ZN(n749) );
  XNOR2_X1 U458 ( .A(n748), .B(n747), .ZN(n385) );
  NAND2_X1 U459 ( .A1(n750), .A2(G478), .ZN(n386) );
  NAND2_X1 U460 ( .A1(n388), .A2(n392), .ZN(n387) );
  XNOR2_X1 U461 ( .A(n389), .B(n356), .ZN(n388) );
  INV_X1 U462 ( .A(KEYINPUT56), .ZN(n390) );
  NAND2_X1 U463 ( .A1(n393), .A2(n392), .ZN(n391) );
  XNOR2_X1 U464 ( .A(n394), .B(n348), .ZN(n393) );
  NAND2_X1 U465 ( .A1(n674), .A2(n353), .ZN(n347) );
  XOR2_X1 U466 ( .A(n744), .B(n746), .Z(n348) );
  AND2_X1 U467 ( .A1(n414), .A2(n347), .ZN(n349) );
  XOR2_X1 U468 ( .A(G146), .B(KEYINPUT78), .Z(n350) );
  AND2_X1 U469 ( .A1(n569), .A2(n551), .ZN(n351) );
  NOR2_X1 U470 ( .A1(n427), .A2(n425), .ZN(n352) );
  AND2_X1 U471 ( .A1(n534), .A2(n416), .ZN(n353) );
  INV_X1 U472 ( .A(KEYINPUT109), .ZN(n551) );
  INV_X1 U473 ( .A(G902), .ZN(n523) );
  AND2_X1 U474 ( .A1(n384), .A2(n383), .ZN(n354) );
  XOR2_X1 U475 ( .A(KEYINPUT48), .B(KEYINPUT68), .Z(n355) );
  XNOR2_X1 U476 ( .A(KEYINPUT59), .B(n667), .ZN(n356) );
  XNOR2_X1 U477 ( .A(KEYINPUT62), .B(n674), .ZN(n357) );
  XOR2_X1 U478 ( .A(n636), .B(n635), .Z(n358) );
  INV_X1 U479 ( .A(n666), .ZN(n384) );
  XOR2_X1 U480 ( .A(KEYINPUT118), .B(KEYINPUT60), .Z(n359) );
  AND2_X1 U481 ( .A1(n486), .A2(n668), .ZN(n754) );
  INV_X1 U482 ( .A(n754), .ZN(n392) );
  NAND2_X1 U483 ( .A1(n360), .A2(n368), .ZN(n369) );
  XNOR2_X1 U484 ( .A(n637), .B(n358), .ZN(n401) );
  NOR2_X1 U485 ( .A1(n626), .A2(n631), .ZN(n362) );
  XNOR2_X2 U486 ( .A(n492), .B(n491), .ZN(n581) );
  NOR2_X1 U487 ( .A1(n628), .A2(n552), .ZN(n553) );
  XOR2_X1 U488 ( .A(n490), .B(n489), .Z(n748) );
  NAND2_X1 U489 ( .A1(n366), .A2(n666), .ZN(n365) );
  XNOR2_X1 U490 ( .A(n572), .B(KEYINPUT107), .ZN(n566) );
  NOR2_X2 U491 ( .A1(n665), .A2(n734), .ZN(n730) );
  NOR2_X1 U492 ( .A1(n665), .A2(n365), .ZN(n364) );
  NAND2_X1 U493 ( .A1(n665), .A2(n354), .ZN(n368) );
  XNOR2_X1 U494 ( .A(n371), .B(n529), .ZN(n370) );
  XNOR2_X2 U495 ( .A(n484), .B(KEYINPUT4), .ZN(n527) );
  NAND2_X1 U496 ( .A1(n373), .A2(n580), .ZN(n377) );
  NOR2_X1 U497 ( .A1(n696), .A2(n378), .ZN(n373) );
  NAND2_X1 U498 ( .A1(n374), .A2(n378), .ZN(n376) );
  NAND2_X1 U499 ( .A1(n375), .A2(n580), .ZN(n374) );
  INV_X1 U500 ( .A(n696), .ZN(n375) );
  NAND2_X1 U501 ( .A1(n377), .A2(n376), .ZN(n380) );
  INV_X1 U502 ( .A(KEYINPUT34), .ZN(n378) );
  XNOR2_X2 U503 ( .A(n379), .B(KEYINPUT35), .ZN(n595) );
  NAND2_X1 U504 ( .A1(n380), .A2(n571), .ZN(n379) );
  XNOR2_X1 U505 ( .A(n387), .B(n359), .ZN(G60) );
  XNOR2_X1 U506 ( .A(n391), .B(n390), .ZN(G51) );
  XNOR2_X1 U507 ( .A(n395), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U508 ( .A1(n750), .A2(G472), .ZN(n397) );
  XNOR2_X1 U509 ( .A(n730), .B(n399), .ZN(n398) );
  NAND2_X1 U510 ( .A1(n402), .A2(n401), .ZN(n400) );
  AND2_X1 U511 ( .A1(n403), .A2(n660), .ZN(n402) );
  XNOR2_X1 U512 ( .A(n693), .B(n404), .ZN(n403) );
  INV_X1 U513 ( .A(KEYINPUT88), .ZN(n404) );
  NAND2_X1 U514 ( .A1(n407), .A2(n351), .ZN(n406) );
  NAND2_X1 U515 ( .A1(n674), .A2(n416), .ZN(n415) );
  NAND2_X1 U516 ( .A1(n581), .A2(KEYINPUT109), .ZN(n408) );
  NOR2_X1 U517 ( .A1(n581), .A2(n582), .ZN(n584) );
  INV_X1 U518 ( .A(n415), .ZN(n412) );
  NAND2_X1 U519 ( .A1(n417), .A2(n534), .ZN(n414) );
  INV_X1 U520 ( .A(G472), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n553), .B(n428), .ZN(n427) );
  AND2_X1 U522 ( .A1(n536), .A2(n535), .ZN(n558) );
  NAND2_X1 U523 ( .A1(n536), .A2(n430), .ZN(n429) );
  XNOR2_X1 U524 ( .A(n429), .B(n539), .ZN(n594) );
  XOR2_X1 U525 ( .A(n500), .B(n499), .Z(n432) );
  INV_X1 U526 ( .A(KEYINPUT65), .ZN(n635) );
  INV_X1 U527 ( .A(n619), .ZN(n620) );
  XNOR2_X1 U528 ( .A(KEYINPUT13), .B(G475), .ZN(n480) );
  XNOR2_X1 U529 ( .A(n525), .B(n524), .ZN(n526) );
  BUF_X1 U530 ( .A(n665), .Z(n731) );
  INV_X1 U531 ( .A(KEYINPUT39), .ZN(n623) );
  NOR2_X1 U532 ( .A1(n560), .A2(n559), .ZN(n588) );
  XOR2_X1 U533 ( .A(KEYINPUT80), .B(KEYINPUT17), .Z(n436) );
  INV_X1 U534 ( .A(G224), .ZN(n434) );
  XNOR2_X1 U535 ( .A(n476), .B(n437), .ZN(n438) );
  XNOR2_X1 U536 ( .A(n439), .B(n438), .ZN(n441) );
  XNOR2_X1 U537 ( .A(n441), .B(n527), .ZN(n449) );
  XNOR2_X1 U538 ( .A(G104), .B(G101), .ZN(n443) );
  XNOR2_X1 U539 ( .A(G110), .B(G107), .ZN(n442) );
  XNOR2_X1 U540 ( .A(n443), .B(n442), .ZN(n529) );
  XNOR2_X1 U541 ( .A(G122), .B(G116), .ZN(n482) );
  XNOR2_X1 U542 ( .A(n482), .B(KEYINPUT16), .ZN(n444) );
  XNOR2_X1 U543 ( .A(n529), .B(n444), .ZN(n448) );
  XNOR2_X1 U544 ( .A(KEYINPUT3), .B(G119), .ZN(n445) );
  XNOR2_X1 U545 ( .A(n445), .B(KEYINPUT93), .ZN(n447) );
  XNOR2_X1 U546 ( .A(n447), .B(n446), .ZN(n519) );
  XNOR2_X1 U547 ( .A(n448), .B(n519), .ZN(n613) );
  XNOR2_X1 U548 ( .A(n449), .B(n613), .ZN(n744) );
  XNOR2_X2 U549 ( .A(KEYINPUT15), .B(G902), .ZN(n666) );
  NAND2_X1 U550 ( .A1(n744), .A2(n666), .ZN(n453) );
  NAND2_X1 U551 ( .A1(n523), .A2(n450), .ZN(n454) );
  NAND2_X1 U552 ( .A1(n454), .A2(G210), .ZN(n451) );
  XNOR2_X1 U553 ( .A(n451), .B(KEYINPUT94), .ZN(n452) );
  INV_X1 U554 ( .A(n541), .ZN(n455) );
  NAND2_X1 U555 ( .A1(n454), .A2(G214), .ZN(n714) );
  NAND2_X1 U556 ( .A1(n455), .A2(n714), .ZN(n458) );
  XNOR2_X1 U557 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n456) );
  XNOR2_X1 U558 ( .A(n456), .B(KEYINPUT67), .ZN(n457) );
  XNOR2_X1 U559 ( .A(n459), .B(KEYINPUT14), .ZN(n460) );
  XNOR2_X1 U560 ( .A(KEYINPUT74), .B(n460), .ZN(n461) );
  NAND2_X1 U561 ( .A1(G952), .A2(n461), .ZN(n729) );
  NOR2_X1 U562 ( .A1(n763), .A2(n729), .ZN(n546) );
  NAND2_X1 U563 ( .A1(n461), .A2(G902), .ZN(n543) );
  INV_X1 U564 ( .A(n763), .ZN(n604) );
  NOR2_X1 U565 ( .A1(n604), .A2(G898), .ZN(n462) );
  XNOR2_X1 U566 ( .A(n462), .B(KEYINPUT95), .ZN(n612) );
  NOR2_X1 U567 ( .A1(n543), .A2(n612), .ZN(n463) );
  OR2_X1 U568 ( .A1(n546), .A2(n463), .ZN(n464) );
  XNOR2_X1 U569 ( .A(n464), .B(KEYINPUT96), .ZN(n465) );
  XNOR2_X2 U570 ( .A(n466), .B(KEYINPUT0), .ZN(n573) );
  INV_X1 U571 ( .A(n573), .ZN(n495) );
  NAND2_X1 U572 ( .A1(n666), .A2(G234), .ZN(n467) );
  XNOR2_X1 U573 ( .A(n467), .B(KEYINPUT20), .ZN(n506) );
  NAND2_X1 U574 ( .A1(n506), .A2(G221), .ZN(n468) );
  XOR2_X1 U575 ( .A(KEYINPUT21), .B(n468), .Z(n698) );
  INV_X1 U576 ( .A(KEYINPUT101), .ZN(n469) );
  XNOR2_X1 U577 ( .A(n698), .B(n469), .ZN(n561) );
  INV_X1 U578 ( .A(n561), .ZN(n493) );
  XNOR2_X1 U579 ( .A(n471), .B(n470), .ZN(n475) );
  XOR2_X1 U580 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n473) );
  XNOR2_X1 U581 ( .A(n473), .B(n472), .ZN(n474) );
  XOR2_X1 U582 ( .A(n475), .B(n474), .Z(n479) );
  XNOR2_X1 U583 ( .A(n476), .B(KEYINPUT10), .ZN(n755) );
  NAND2_X1 U584 ( .A1(G214), .A2(n512), .ZN(n477) );
  XNOR2_X1 U585 ( .A(n755), .B(n477), .ZN(n478) );
  XNOR2_X1 U586 ( .A(n479), .B(n478), .ZN(n667) );
  NOR2_X1 U587 ( .A1(G902), .A2(n667), .ZN(n481) );
  INV_X1 U588 ( .A(n482), .ZN(n483) );
  XNOR2_X1 U589 ( .A(n484), .B(n483), .ZN(n485) );
  XNOR2_X1 U590 ( .A(n431), .B(n485), .ZN(n490) );
  INV_X1 U591 ( .A(n486), .ZN(n542) );
  NAND2_X1 U592 ( .A1(G234), .A2(n542), .ZN(n487) );
  XNOR2_X1 U593 ( .A(n488), .B(n487), .ZN(n504) );
  NAND2_X1 U594 ( .A1(G217), .A2(n504), .ZN(n489) );
  NOR2_X1 U595 ( .A1(G902), .A2(n748), .ZN(n492) );
  XNOR2_X1 U596 ( .A(KEYINPUT103), .B(G478), .ZN(n491) );
  XNOR2_X1 U597 ( .A(KEYINPUT106), .B(n433), .ZN(n717) );
  NOR2_X1 U598 ( .A1(n493), .A2(n717), .ZN(n494) );
  NAND2_X1 U599 ( .A1(n495), .A2(n494), .ZN(n498) );
  INV_X1 U600 ( .A(KEYINPUT72), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n496), .B(KEYINPUT22), .ZN(n497) );
  XOR2_X1 U602 ( .A(n755), .B(G110), .Z(n503) );
  INV_X1 U603 ( .A(G140), .ZN(n557) );
  XNOR2_X1 U604 ( .A(n557), .B(G137), .ZN(n525) );
  XNOR2_X1 U605 ( .A(G128), .B(n525), .ZN(n501) );
  XOR2_X1 U606 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n500) );
  XNOR2_X1 U607 ( .A(G119), .B(KEYINPUT98), .ZN(n499) );
  NAND2_X1 U608 ( .A1(n504), .A2(G221), .ZN(n505) );
  NOR2_X1 U609 ( .A1(n752), .A2(G902), .ZN(n511) );
  XOR2_X1 U610 ( .A(KEYINPUT100), .B(KEYINPUT25), .Z(n508) );
  NAND2_X1 U611 ( .A1(G217), .A2(n506), .ZN(n507) );
  XNOR2_X1 U612 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U613 ( .A(n509), .B(KEYINPUT99), .ZN(n510) );
  XNOR2_X1 U614 ( .A(n511), .B(n510), .ZN(n562) );
  INV_X1 U615 ( .A(n562), .ZN(n549) );
  INV_X1 U616 ( .A(n549), .ZN(n699) );
  NAND2_X1 U617 ( .A1(n512), .A2(G210), .ZN(n513) );
  XNOR2_X1 U618 ( .A(n514), .B(n513), .ZN(n518) );
  XNOR2_X1 U619 ( .A(n516), .B(n515), .ZN(n517) );
  XNOR2_X1 U620 ( .A(n518), .B(n517), .ZN(n520) );
  XNOR2_X1 U621 ( .A(n520), .B(n519), .ZN(n522) );
  XNOR2_X1 U622 ( .A(n527), .B(n524), .ZN(n521) );
  XNOR2_X1 U623 ( .A(n522), .B(n521), .ZN(n674) );
  NOR2_X1 U624 ( .A1(n699), .A2(n617), .ZN(n532) );
  INV_X1 U625 ( .A(G227), .ZN(n528) );
  OR2_X2 U626 ( .A1(n670), .A2(G902), .ZN(n577) );
  XNOR2_X1 U627 ( .A(KEYINPUT66), .B(KEYINPUT1), .ZN(n530) );
  INV_X1 U628 ( .A(G469), .ZN(n576) );
  XNOR2_X2 U629 ( .A(n577), .B(n531), .ZN(n702) );
  AND2_X1 U630 ( .A1(n532), .A2(n702), .ZN(n533) );
  AND2_X1 U631 ( .A1(n536), .A2(n533), .ZN(n593) );
  XOR2_X1 U632 ( .A(G110), .B(n593), .Z(G12) );
  INV_X1 U633 ( .A(KEYINPUT6), .ZN(n534) );
  INV_X1 U634 ( .A(n565), .ZN(n535) );
  INV_X1 U635 ( .A(KEYINPUT92), .ZN(n537) );
  XNOR2_X1 U636 ( .A(n702), .B(n537), .ZN(n639) );
  AND2_X1 U637 ( .A1(n639), .A2(n549), .ZN(n538) );
  XNOR2_X1 U638 ( .A(KEYINPUT81), .B(KEYINPUT32), .ZN(n539) );
  XNOR2_X1 U639 ( .A(G119), .B(KEYINPUT127), .ZN(n540) );
  XNOR2_X1 U640 ( .A(n594), .B(n540), .ZN(G21) );
  OR2_X1 U641 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U642 ( .A1(G900), .A2(n544), .ZN(n545) );
  NOR2_X1 U643 ( .A1(n546), .A2(n545), .ZN(n619) );
  INV_X1 U644 ( .A(n698), .ZN(n547) );
  NOR2_X1 U645 ( .A1(n619), .A2(n547), .ZN(n548) );
  NAND2_X1 U646 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U647 ( .A(n550), .B(KEYINPUT69), .Z(n628) );
  NAND2_X1 U648 ( .A1(n352), .A2(n702), .ZN(n555) );
  XOR2_X1 U649 ( .A(KEYINPUT43), .B(KEYINPUT111), .Z(n554) );
  XNOR2_X1 U650 ( .A(n555), .B(n554), .ZN(n556) );
  AND2_X1 U651 ( .A1(n638), .A2(n556), .ZN(n662) );
  XNOR2_X1 U652 ( .A(n662), .B(n557), .ZN(G42) );
  XNOR2_X1 U653 ( .A(n558), .B(KEYINPUT89), .ZN(n560) );
  NAND2_X1 U654 ( .A1(n702), .A2(n699), .ZN(n559) );
  XOR2_X1 U655 ( .A(G101), .B(n588), .Z(G3) );
  INV_X1 U656 ( .A(n702), .ZN(n563) );
  INV_X1 U657 ( .A(KEYINPUT75), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n566), .A2(n565), .ZN(n568) );
  XNOR2_X1 U659 ( .A(KEYINPUT71), .B(KEYINPUT33), .ZN(n567) );
  XNOR2_X1 U660 ( .A(n573), .B(KEYINPUT97), .ZN(n580) );
  NAND2_X1 U661 ( .A1(n569), .A2(n581), .ZN(n570) );
  XNOR2_X1 U662 ( .A(n570), .B(KEYINPUT108), .ZN(n644) );
  XOR2_X1 U663 ( .A(n595), .B(G122), .Z(G24) );
  NAND2_X1 U664 ( .A1(n595), .A2(KEYINPUT44), .ZN(n591) );
  INV_X1 U665 ( .A(n617), .ZN(n629) );
  OR2_X1 U666 ( .A1(n572), .A2(n629), .ZN(n709) );
  NOR2_X1 U667 ( .A1(n709), .A2(n573), .ZN(n574) );
  XNOR2_X1 U668 ( .A(n574), .B(KEYINPUT31), .ZN(n690) );
  NAND2_X1 U669 ( .A1(n575), .A2(n629), .ZN(n578) );
  XNOR2_X1 U670 ( .A(n577), .B(n576), .ZN(n631) );
  NOR2_X1 U671 ( .A1(n578), .A2(n631), .ZN(n579) );
  NAND2_X1 U672 ( .A1(n580), .A2(n579), .ZN(n679) );
  AND2_X1 U673 ( .A1(n690), .A2(n679), .ZN(n587) );
  NAND2_X1 U674 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U675 ( .A(n583), .B(KEYINPUT104), .Z(n683) );
  NOR2_X1 U676 ( .A1(n683), .A2(n584), .ZN(n586) );
  INV_X1 U677 ( .A(KEYINPUT105), .ZN(n585) );
  XNOR2_X1 U678 ( .A(n586), .B(n585), .ZN(n720) );
  NOR2_X1 U679 ( .A1(n587), .A2(n720), .ZN(n589) );
  NOR2_X1 U680 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U681 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U682 ( .A(n592), .B(KEYINPUT90), .ZN(n602) );
  NOR2_X1 U683 ( .A1(n595), .A2(n597), .ZN(n596) );
  NOR2_X1 U684 ( .A1(n596), .A2(KEYINPUT44), .ZN(n600) );
  INV_X1 U685 ( .A(n597), .ZN(n598) );
  AND2_X1 U686 ( .A1(n598), .A2(KEYINPUT44), .ZN(n599) );
  NOR2_X1 U687 ( .A1(n600), .A2(n599), .ZN(n601) );
  INV_X1 U688 ( .A(n731), .ZN(n605) );
  NAND2_X1 U689 ( .A1(n605), .A2(n604), .ZN(n611) );
  XOR2_X1 U690 ( .A(KEYINPUT61), .B(KEYINPUT122), .Z(n607) );
  NAND2_X1 U691 ( .A1(G224), .A2(n763), .ZN(n606) );
  XNOR2_X1 U692 ( .A(n607), .B(n606), .ZN(n608) );
  XNOR2_X1 U693 ( .A(KEYINPUT121), .B(n608), .ZN(n609) );
  NAND2_X1 U694 ( .A1(n609), .A2(G898), .ZN(n610) );
  NAND2_X1 U695 ( .A1(n611), .A2(n610), .ZN(n616) );
  NAND2_X1 U696 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U697 ( .A(n614), .B(KEYINPUT123), .ZN(n615) );
  XNOR2_X1 U698 ( .A(n616), .B(n615), .ZN(G69) );
  NAND2_X1 U699 ( .A1(n617), .A2(n714), .ZN(n618) );
  XNOR2_X1 U700 ( .A(KEYINPUT30), .B(n618), .ZN(n622) );
  INV_X1 U701 ( .A(n631), .ZN(n649) );
  XOR2_X1 U702 ( .A(KEYINPUT38), .B(n638), .Z(n626) );
  XNOR2_X1 U703 ( .A(n624), .B(n623), .ZN(n661) );
  NAND2_X1 U704 ( .A1(n661), .A2(n584), .ZN(n625) );
  XNOR2_X1 U705 ( .A(n625), .B(KEYINPUT40), .ZN(n768) );
  INV_X1 U706 ( .A(n626), .ZN(n715) );
  NAND2_X1 U707 ( .A1(n715), .A2(n714), .ZN(n719) );
  NOR2_X1 U708 ( .A1(n717), .A2(n719), .ZN(n627) );
  XNOR2_X1 U709 ( .A(KEYINPUT41), .B(n627), .ZN(n712) );
  INV_X1 U710 ( .A(n712), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n629), .A2(n628), .ZN(n630) );
  XOR2_X1 U712 ( .A(KEYINPUT28), .B(n630), .Z(n651) );
  NOR2_X1 U713 ( .A1(n651), .A2(n631), .ZN(n632) );
  NAND2_X1 U714 ( .A1(n633), .A2(n632), .ZN(n634) );
  XNOR2_X1 U715 ( .A(n634), .B(KEYINPUT42), .ZN(n767) );
  NAND2_X1 U716 ( .A1(n768), .A2(n767), .ZN(n637) );
  XOR2_X1 U717 ( .A(KEYINPUT46), .B(KEYINPUT87), .Z(n636) );
  INV_X1 U718 ( .A(n638), .ZN(n642) );
  NAND2_X1 U719 ( .A1(n643), .A2(n642), .ZN(n645) );
  NOR2_X1 U720 ( .A1(n645), .A2(n644), .ZN(n646) );
  NAND2_X1 U721 ( .A1(n646), .A2(n649), .ZN(n647) );
  XNOR2_X1 U722 ( .A(KEYINPUT112), .B(n647), .ZN(n769) );
  NAND2_X1 U723 ( .A1(n649), .A2(n648), .ZN(n650) );
  OR2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n655) );
  INV_X1 U725 ( .A(n720), .ZN(n652) );
  NOR2_X1 U726 ( .A1(n655), .A2(n652), .ZN(n653) );
  NAND2_X1 U727 ( .A1(KEYINPUT73), .A2(n653), .ZN(n654) );
  NAND2_X1 U728 ( .A1(n769), .A2(n654), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n720), .A2(KEYINPUT73), .ZN(n656) );
  NAND2_X1 U730 ( .A1(n686), .A2(n656), .ZN(n657) );
  XNOR2_X1 U731 ( .A(KEYINPUT47), .B(n657), .ZN(n658) );
  NOR2_X1 U732 ( .A1(n659), .A2(n658), .ZN(n660) );
  AND2_X1 U733 ( .A1(n683), .A2(n661), .ZN(n695) );
  NOR2_X1 U734 ( .A1(n662), .A2(n695), .ZN(n663) );
  INV_X1 U735 ( .A(G952), .ZN(n668) );
  NAND2_X1 U736 ( .A1(n750), .A2(G469), .ZN(n672) );
  XOR2_X1 U737 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n669) );
  XNOR2_X1 U738 ( .A(n670), .B(n669), .ZN(n671) );
  XNOR2_X1 U739 ( .A(n672), .B(n671), .ZN(n673) );
  NOR2_X1 U740 ( .A1(n673), .A2(n754), .ZN(G54) );
  INV_X1 U741 ( .A(n675), .ZN(n688) );
  NOR2_X1 U742 ( .A1(n688), .A2(n679), .ZN(n677) );
  XNOR2_X1 U743 ( .A(KEYINPUT113), .B(KEYINPUT114), .ZN(n676) );
  XNOR2_X1 U744 ( .A(n677), .B(n676), .ZN(n678) );
  XNOR2_X1 U745 ( .A(G104), .B(n678), .ZN(G6) );
  INV_X1 U746 ( .A(n683), .ZN(n691) );
  NOR2_X1 U747 ( .A1(n691), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n680) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(n682) );
  XNOR2_X1 U750 ( .A(G107), .B(n682), .ZN(G9) );
  XOR2_X1 U751 ( .A(G128), .B(KEYINPUT29), .Z(n685) );
  NAND2_X1 U752 ( .A1(n686), .A2(n683), .ZN(n684) );
  XNOR2_X1 U753 ( .A(n685), .B(n684), .ZN(G30) );
  NAND2_X1 U754 ( .A1(n686), .A2(n675), .ZN(n687) );
  XNOR2_X1 U755 ( .A(n687), .B(G146), .ZN(G48) );
  NOR2_X1 U756 ( .A1(n688), .A2(n690), .ZN(n689) );
  XOR2_X1 U757 ( .A(G113), .B(n689), .Z(G15) );
  NOR2_X1 U758 ( .A1(n691), .A2(n690), .ZN(n692) );
  XOR2_X1 U759 ( .A(G116), .B(n692), .Z(G18) );
  XNOR2_X1 U760 ( .A(n693), .B(G125), .ZN(n694) );
  XNOR2_X1 U761 ( .A(n694), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U762 ( .A(G134), .B(n695), .Z(G36) );
  NOR2_X1 U763 ( .A1(n712), .A2(n724), .ZN(n697) );
  NOR2_X1 U764 ( .A1(n697), .A2(n763), .ZN(n742) );
  NOR2_X1 U765 ( .A1(n699), .A2(n698), .ZN(n700) );
  XOR2_X1 U766 ( .A(KEYINPUT115), .B(n700), .Z(n701) );
  XNOR2_X1 U767 ( .A(KEYINPUT49), .B(n701), .ZN(n708) );
  INV_X1 U768 ( .A(n575), .ZN(n703) );
  NAND2_X1 U769 ( .A1(n703), .A2(n702), .ZN(n705) );
  XOR2_X1 U770 ( .A(KEYINPUT50), .B(KEYINPUT116), .Z(n704) );
  XNOR2_X1 U771 ( .A(n705), .B(n704), .ZN(n706) );
  NOR2_X1 U772 ( .A1(n706), .A2(n617), .ZN(n707) );
  NAND2_X1 U773 ( .A1(n708), .A2(n707), .ZN(n710) );
  NAND2_X1 U774 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U775 ( .A(KEYINPUT51), .B(n711), .ZN(n713) );
  NOR2_X1 U776 ( .A1(n713), .A2(n712), .ZN(n726) );
  NOR2_X1 U777 ( .A1(n715), .A2(n714), .ZN(n716) );
  NOR2_X1 U778 ( .A1(n717), .A2(n716), .ZN(n718) );
  XOR2_X1 U779 ( .A(KEYINPUT117), .B(n718), .Z(n722) );
  NOR2_X1 U780 ( .A1(n720), .A2(n719), .ZN(n721) );
  NOR2_X1 U781 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U782 ( .A1(n724), .A2(n723), .ZN(n725) );
  NOR2_X1 U783 ( .A1(n726), .A2(n725), .ZN(n727) );
  XNOR2_X1 U784 ( .A(n727), .B(KEYINPUT52), .ZN(n728) );
  NOR2_X1 U785 ( .A1(n729), .A2(n728), .ZN(n740) );
  NAND2_X1 U786 ( .A1(n730), .A2(KEYINPUT2), .ZN(n733) );
  XNOR2_X1 U787 ( .A(KEYINPUT83), .B(KEYINPUT2), .ZN(n735) );
  NAND2_X1 U788 ( .A1(n731), .A2(n735), .ZN(n732) );
  NAND2_X1 U789 ( .A1(n733), .A2(n732), .ZN(n738) );
  NAND2_X1 U790 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U791 ( .A(KEYINPUT85), .B(n736), .ZN(n737) );
  NOR2_X1 U792 ( .A1(n738), .A2(n737), .ZN(n739) );
  NOR2_X1 U793 ( .A1(n740), .A2(n739), .ZN(n741) );
  NAND2_X1 U794 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U795 ( .A(KEYINPUT53), .B(n743), .Z(G75) );
  XOR2_X1 U796 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n745) );
  XNOR2_X1 U797 ( .A(n745), .B(KEYINPUT91), .ZN(n746) );
  XOR2_X1 U798 ( .A(KEYINPUT119), .B(KEYINPUT120), .Z(n747) );
  NOR2_X1 U799 ( .A1(n754), .A2(n749), .ZN(G63) );
  NAND2_X1 U800 ( .A1(n750), .A2(G217), .ZN(n751) );
  XNOR2_X1 U801 ( .A(n752), .B(n751), .ZN(n753) );
  NOR2_X1 U802 ( .A1(n754), .A2(n753), .ZN(G66) );
  XNOR2_X1 U803 ( .A(n756), .B(n755), .ZN(n761) );
  XOR2_X1 U804 ( .A(KEYINPUT124), .B(n761), .Z(n757) );
  XNOR2_X1 U805 ( .A(n757), .B(n734), .ZN(n758) );
  NOR2_X1 U806 ( .A1(n486), .A2(n758), .ZN(n759) );
  XNOR2_X1 U807 ( .A(n759), .B(KEYINPUT125), .ZN(n766) );
  XNOR2_X1 U808 ( .A(G227), .B(KEYINPUT126), .ZN(n760) );
  XNOR2_X1 U809 ( .A(n761), .B(n760), .ZN(n762) );
  NAND2_X1 U810 ( .A1(n762), .A2(G900), .ZN(n764) );
  NAND2_X1 U811 ( .A1(n764), .A2(n763), .ZN(n765) );
  NAND2_X1 U812 ( .A1(n766), .A2(n765), .ZN(G72) );
  XNOR2_X1 U813 ( .A(G137), .B(n767), .ZN(G39) );
  XNOR2_X1 U814 ( .A(G131), .B(n768), .ZN(G33) );
  XNOR2_X1 U815 ( .A(G143), .B(n769), .ZN(G45) );
endmodule

