//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 1 0 0 1 0 1 0 1 1 1 1 0 0 1 0 1 0 1 0 1 1 0 0 0 0 0 1 1 1 0 1 1 0 0 1 1 1 1 0 1 0 1 1 0 0 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:38 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n658, new_n659, new_n660, new_n661, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n699, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n732, new_n733, new_n735,
    new_n736, new_n738, new_n739, new_n740, new_n742, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n824, new_n825, new_n826, new_n828,
    new_n830, new_n831, new_n832, new_n833, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n902, new_n903, new_n904, new_n906,
    new_n907, new_n908, new_n909, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(G1gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(KEYINPUT16), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  OAI21_X1  g004(.A(new_n205), .B1(G1gat), .B2(new_n202), .ZN(new_n206));
  INV_X1    g005(.A(G8gat), .ZN(new_n207));
  XNOR2_X1  g006(.A(new_n206), .B(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT14), .ZN(new_n209));
  INV_X1    g008(.A(G29gat), .ZN(new_n210));
  INV_X1    g009(.A(G36gat), .ZN(new_n211));
  NAND3_X1  g010(.A1(new_n209), .A2(new_n210), .A3(new_n211), .ZN(new_n212));
  OAI21_X1  g011(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n213));
  AOI22_X1  g012(.A1(new_n212), .A2(new_n213), .B1(G29gat), .B2(G36gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(G43gat), .B(G50gat), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n214), .B1(KEYINPUT15), .B2(new_n215), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n216), .A2(new_n218), .ZN(new_n219));
  OR2_X1    g018(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n220));
  NAND3_X1  g019(.A1(new_n220), .A2(new_n217), .A3(new_n214), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n219), .A2(new_n221), .ZN(new_n222));
  AND3_X1   g021(.A1(new_n222), .A2(KEYINPUT88), .A3(KEYINPUT17), .ZN(new_n223));
  AOI21_X1  g022(.A(KEYINPUT17), .B1(new_n222), .B2(KEYINPUT88), .ZN(new_n224));
  OAI21_X1  g023(.A(new_n208), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(new_n206), .B(G8gat), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n226), .A2(new_n222), .ZN(new_n227));
  AND2_X1   g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NAND2_X1  g027(.A1(G229gat), .A2(G233gat), .ZN(new_n229));
  AOI21_X1  g028(.A(KEYINPUT18), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OR3_X1    g029(.A1(new_n226), .A2(KEYINPUT90), .A3(new_n222), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT90), .B1(new_n226), .B2(new_n222), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n231), .A2(new_n227), .A3(new_n232), .ZN(new_n233));
  XOR2_X1   g032(.A(new_n229), .B(KEYINPUT13), .Z(new_n234));
  NAND2_X1  g033(.A1(new_n233), .A2(new_n234), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n225), .A2(KEYINPUT18), .A3(new_n229), .A4(new_n227), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n230), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g037(.A(KEYINPUT11), .B(G169gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n239), .B(G197gat), .ZN(new_n240));
  XOR2_X1   g039(.A(G113gat), .B(G141gat), .Z(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(KEYINPUT12), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(KEYINPUT89), .ZN(new_n245));
  OAI21_X1  g044(.A(new_n244), .B1(new_n237), .B2(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(new_n238), .B(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT85), .ZN(new_n249));
  NAND2_X1  g048(.A1(G225gat), .A2(G233gat), .ZN(new_n250));
  INV_X1    g049(.A(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT69), .ZN(new_n252));
  AND2_X1   g051(.A1(G127gat), .A2(G134gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(G127gat), .A2(G134gat), .ZN(new_n254));
  OAI21_X1  g053(.A(new_n252), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G134gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g057(.A1(G127gat), .A2(G134gat), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n258), .A2(KEYINPUT69), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT70), .ZN(new_n262));
  INV_X1    g061(.A(KEYINPUT1), .ZN(new_n263));
  INV_X1    g062(.A(G113gat), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n264), .A2(G120gat), .ZN(new_n265));
  INV_X1    g064(.A(G120gat), .ZN(new_n266));
  NOR2_X1   g065(.A1(new_n266), .A2(G113gat), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n263), .B1(new_n265), .B2(new_n267), .ZN(new_n268));
  AND3_X1   g067(.A1(new_n261), .A2(new_n262), .A3(new_n268), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n262), .B1(new_n261), .B2(new_n268), .ZN(new_n270));
  INV_X1    g069(.A(new_n267), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT71), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(G113gat), .B2(new_n266), .ZN(new_n273));
  NOR3_X1   g072(.A1(new_n264), .A2(KEYINPUT71), .A3(G120gat), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n271), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  OAI22_X1  g074(.A1(new_n275), .A2(KEYINPUT72), .B1(new_n254), .B2(new_n253), .ZN(new_n276));
  OAI21_X1  g075(.A(KEYINPUT71), .B1(new_n264), .B2(G120gat), .ZN(new_n277));
  NAND3_X1  g076(.A1(new_n272), .A2(new_n266), .A3(G113gat), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n267), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(KEYINPUT72), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n263), .B1(new_n279), .B2(new_n280), .ZN(new_n281));
  OAI22_X1  g080(.A1(new_n269), .A2(new_n270), .B1(new_n276), .B2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(KEYINPUT80), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT78), .ZN(new_n284));
  INV_X1    g083(.A(G148gat), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n284), .B1(new_n285), .B2(G141gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(G141gat), .ZN(new_n287));
  INV_X1    g086(.A(G141gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n288), .A2(KEYINPUT78), .A3(G148gat), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G155gat), .A2(G162gat), .ZN(new_n291));
  OR2_X1    g090(.A1(G155gat), .A2(G162gat), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n291), .B1(new_n292), .B2(KEYINPUT2), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n290), .A2(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(G155gat), .A2(G162gat), .ZN(new_n295));
  NOR2_X1   g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n295), .A2(new_n296), .ZN(new_n297));
  XNOR2_X1  g096(.A(G141gat), .B(G148gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n297), .B1(new_n298), .B2(KEYINPUT2), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n294), .A2(new_n299), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n282), .A2(new_n283), .A3(new_n300), .ZN(new_n301));
  NOR3_X1   g100(.A1(new_n253), .A2(new_n254), .A3(new_n252), .ZN(new_n302));
  AOI21_X1  g101(.A(KEYINPUT69), .B1(new_n258), .B2(new_n259), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n268), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(KEYINPUT70), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n261), .A2(new_n262), .A3(new_n268), .ZN(new_n306));
  AOI21_X1  g105(.A(KEYINPUT1), .B1(new_n275), .B2(KEYINPUT72), .ZN(new_n307));
  AOI22_X1  g106(.A1(new_n279), .A2(new_n280), .B1(new_n258), .B2(new_n259), .ZN(new_n308));
  AOI22_X1  g107(.A1(new_n305), .A2(new_n306), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n300), .ZN(new_n310));
  AOI21_X1  g109(.A(KEYINPUT80), .B1(new_n309), .B2(new_n310), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n301), .A2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT81), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n313), .B1(new_n309), .B2(new_n310), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n282), .A2(KEYINPUT81), .A3(new_n300), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n251), .B1(new_n312), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT4), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n318), .B1(new_n301), .B2(new_n311), .ZN(new_n319));
  AND3_X1   g118(.A1(new_n294), .A2(KEYINPUT79), .A3(new_n299), .ZN(new_n320));
  AOI21_X1  g119(.A(KEYINPUT79), .B1(new_n294), .B2(new_n299), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n309), .A2(new_n322), .A3(KEYINPUT4), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT3), .ZN(new_n324));
  NAND3_X1  g123(.A1(new_n294), .A2(new_n299), .A3(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n324), .B1(new_n294), .B2(new_n299), .ZN(new_n327));
  NOR2_X1   g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(new_n282), .ZN(new_n329));
  AND3_X1   g128(.A1(new_n323), .A2(new_n329), .A3(new_n250), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n319), .A2(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n317), .A2(new_n331), .A3(KEYINPUT5), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n309), .A2(new_n322), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n300), .A2(KEYINPUT3), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n325), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n309), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n333), .B1(new_n336), .B2(new_n318), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n283), .B1(new_n282), .B2(new_n300), .ZN(new_n338));
  NAND3_X1  g137(.A1(new_n309), .A2(KEYINPUT80), .A3(new_n310), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT4), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n251), .A2(KEYINPUT5), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n332), .A2(new_n342), .ZN(new_n343));
  XNOR2_X1  g142(.A(KEYINPUT0), .B(G57gat), .ZN(new_n344));
  XNOR2_X1  g143(.A(new_n344), .B(G85gat), .ZN(new_n345));
  XNOR2_X1  g144(.A(G1gat), .B(G29gat), .ZN(new_n346));
  XOR2_X1   g145(.A(new_n345), .B(new_n346), .Z(new_n347));
  INV_X1    g146(.A(new_n347), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n343), .A2(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT82), .B(KEYINPUT6), .Z(new_n350));
  INV_X1    g149(.A(new_n350), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n332), .A2(new_n342), .A3(new_n347), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n349), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n343), .A2(new_n348), .A3(new_n350), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(KEYINPUT84), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n347), .B1(new_n332), .B2(new_n342), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT84), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n356), .A2(new_n357), .A3(new_n350), .ZN(new_n358));
  NAND3_X1  g157(.A1(new_n353), .A2(new_n355), .A3(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(G226gat), .ZN(new_n360));
  INV_X1    g159(.A(G233gat), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n360), .A2(new_n361), .ZN(new_n362));
  OAI21_X1  g161(.A(KEYINPUT67), .B1(G169gat), .B2(G176gat), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n363), .A2(KEYINPUT23), .ZN(new_n364));
  NAND2_X1  g163(.A1(G169gat), .A2(G176gat), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT23), .ZN(new_n366));
  OAI211_X1 g165(.A(new_n366), .B(KEYINPUT67), .C1(G169gat), .C2(G176gat), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n364), .A2(new_n365), .A3(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT68), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g169(.A1(new_n364), .A2(KEYINPUT68), .A3(new_n367), .A4(new_n365), .ZN(new_n371));
  INV_X1    g170(.A(G183gat), .ZN(new_n372));
  INV_X1    g171(.A(G190gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(G183gat), .A2(G190gat), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n374), .A2(KEYINPUT24), .A3(new_n375), .ZN(new_n376));
  OR2_X1    g175(.A1(new_n375), .A2(KEYINPUT24), .ZN(new_n377));
  INV_X1    g176(.A(KEYINPUT66), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n378), .A2(KEYINPUT25), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n376), .A2(new_n377), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(KEYINPUT66), .B1(new_n376), .B2(new_n377), .ZN(new_n381));
  OAI211_X1 g180(.A(new_n370), .B(new_n371), .C1(new_n380), .C2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n376), .A2(new_n377), .ZN(new_n383));
  OAI21_X1  g182(.A(KEYINPUT25), .B1(new_n383), .B2(new_n368), .ZN(new_n384));
  AND2_X1   g183(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n385));
  NOR2_X1   g184(.A1(KEYINPUT27), .A2(G183gat), .ZN(new_n386));
  OAI21_X1  g185(.A(new_n373), .B1(new_n385), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(KEYINPUT28), .ZN(new_n388));
  AOI21_X1  g187(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n389));
  OAI21_X1  g188(.A(new_n389), .B1(G169gat), .B2(G176gat), .ZN(new_n390));
  NOR2_X1   g189(.A1(G169gat), .A2(G176gat), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n391), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT28), .ZN(new_n393));
  OAI211_X1 g192(.A(new_n393), .B(new_n373), .C1(new_n385), .C2(new_n386), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n388), .A2(new_n390), .A3(new_n392), .A4(new_n394), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n382), .A2(new_n384), .A3(new_n395), .ZN(new_n396));
  INV_X1    g195(.A(KEYINPUT29), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n362), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n396), .A2(new_n362), .ZN(new_n400));
  INV_X1    g199(.A(KEYINPUT76), .ZN(new_n401));
  NAND2_X1  g200(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(new_n362), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n384), .A2(new_n395), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n403), .B1(new_n404), .B2(new_n382), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT76), .ZN(new_n406));
  NAND3_X1  g205(.A1(new_n399), .A2(new_n402), .A3(new_n406), .ZN(new_n407));
  XNOR2_X1  g206(.A(G197gat), .B(G204gat), .ZN(new_n408));
  INV_X1    g207(.A(G211gat), .ZN(new_n409));
  INV_X1    g208(.A(G218gat), .ZN(new_n410));
  NOR2_X1   g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n408), .B1(KEYINPUT22), .B2(new_n411), .ZN(new_n412));
  XOR2_X1   g211(.A(G211gat), .B(G218gat), .Z(new_n413));
  INV_X1    g212(.A(new_n413), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n412), .B(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(KEYINPUT75), .ZN(new_n416));
  XNOR2_X1  g215(.A(new_n412), .B(new_n413), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT75), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n416), .A2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n407), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT37), .ZN(new_n422));
  NOR3_X1   g221(.A1(new_n398), .A2(new_n420), .A3(new_n405), .ZN(new_n423));
  INV_X1    g222(.A(new_n423), .ZN(new_n424));
  NAND3_X1  g223(.A1(new_n421), .A2(new_n422), .A3(new_n424), .ZN(new_n425));
  XNOR2_X1  g224(.A(G8gat), .B(G36gat), .ZN(new_n426));
  INV_X1    g225(.A(G64gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(G92gat), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n428), .B(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n425), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n423), .B1(new_n407), .B2(new_n420), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n432), .A2(new_n422), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT38), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  OAI21_X1  g233(.A(new_n420), .B1(new_n398), .B2(new_n405), .ZN(new_n435));
  INV_X1    g234(.A(KEYINPUT83), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  OAI211_X1 g236(.A(KEYINPUT83), .B(new_n420), .C1(new_n398), .C2(new_n405), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n437), .B(new_n438), .C1(new_n420), .C2(new_n407), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n439), .A2(KEYINPUT37), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT38), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n440), .A2(new_n441), .A3(new_n430), .A4(new_n425), .ZN(new_n442));
  INV_X1    g241(.A(new_n430), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n421), .A2(new_n424), .A3(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n434), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n359), .A2(new_n445), .ZN(new_n446));
  XNOR2_X1  g245(.A(KEYINPUT31), .B(G50gat), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n324), .B1(new_n415), .B2(KEYINPUT29), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n321), .B2(new_n320), .ZN(new_n449));
  NAND2_X1  g248(.A1(G228gat), .A2(G233gat), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n325), .A2(new_n397), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n416), .A2(new_n419), .A3(new_n451), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n449), .A2(new_n450), .A3(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n448), .A2(new_n300), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n450), .B1(new_n455), .B2(new_n452), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n447), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(G78gat), .B(G106gat), .ZN(new_n458));
  XOR2_X1   g257(.A(new_n458), .B(G22gat), .Z(new_n459));
  INV_X1    g258(.A(new_n456), .ZN(new_n460));
  INV_X1    g259(.A(new_n447), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(new_n461), .A3(new_n453), .ZN(new_n462));
  AND3_X1   g261(.A1(new_n457), .A2(new_n459), .A3(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n459), .B1(new_n457), .B2(new_n462), .ZN(new_n464));
  OR2_X1    g263(.A1(new_n463), .A2(new_n464), .ZN(new_n465));
  OR2_X1    g264(.A1(new_n432), .A2(new_n443), .ZN(new_n466));
  NAND4_X1  g265(.A1(new_n421), .A2(new_n424), .A3(KEYINPUT30), .A4(new_n443), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT77), .ZN(new_n468));
  NAND2_X1  g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(KEYINPUT30), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n444), .A2(new_n470), .ZN(new_n471));
  NAND4_X1  g270(.A1(new_n432), .A2(KEYINPUT77), .A3(KEYINPUT30), .A4(new_n443), .ZN(new_n472));
  AND4_X1   g271(.A1(new_n466), .A2(new_n469), .A3(new_n471), .A4(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n338), .A2(new_n339), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n474), .A2(new_n250), .A3(new_n314), .A4(new_n315), .ZN(new_n475));
  AND2_X1   g274(.A1(new_n337), .A2(new_n340), .ZN(new_n476));
  OAI211_X1 g275(.A(KEYINPUT39), .B(new_n475), .C1(new_n476), .C2(new_n250), .ZN(new_n477));
  AOI21_X1  g276(.A(new_n250), .B1(new_n337), .B2(new_n340), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT39), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n348), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n477), .A2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT40), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n477), .A2(KEYINPUT40), .A3(new_n480), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n349), .A3(new_n484), .ZN(new_n485));
  OAI21_X1  g284(.A(new_n465), .B1(new_n473), .B2(new_n485), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n249), .B1(new_n446), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n353), .A2(new_n354), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n465), .B1(new_n488), .B2(new_n473), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n396), .A2(new_n282), .ZN(new_n490));
  NAND2_X1  g289(.A1(new_n305), .A2(new_n306), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n307), .A2(new_n308), .ZN(new_n492));
  NAND4_X1  g291(.A1(new_n404), .A2(new_n491), .A3(new_n492), .A4(new_n382), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  NAND2_X1  g293(.A1(G227gat), .A2(G233gat), .ZN(new_n495));
  XNOR2_X1  g294(.A(new_n495), .B(KEYINPUT64), .ZN(new_n496));
  XNOR2_X1  g295(.A(new_n496), .B(KEYINPUT65), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n494), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT33), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  XNOR2_X1  g300(.A(G15gat), .B(G43gat), .ZN(new_n502));
  XNOR2_X1  g301(.A(G71gat), .B(G99gat), .ZN(new_n503));
  XOR2_X1   g302(.A(new_n502), .B(new_n503), .Z(new_n504));
  NAND2_X1  g303(.A1(new_n501), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n490), .A2(new_n493), .A3(new_n496), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n506), .A2(KEYINPUT73), .ZN(new_n507));
  INV_X1    g306(.A(KEYINPUT34), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n490), .A2(new_n493), .A3(new_n497), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n507), .A2(new_n508), .A3(new_n509), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n499), .A2(KEYINPUT32), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT73), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n513), .A2(KEYINPUT34), .ZN(new_n514));
  AND3_X1   g313(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n511), .B1(new_n510), .B2(new_n514), .ZN(new_n516));
  OAI21_X1  g315(.A(new_n505), .B1(new_n515), .B2(new_n516), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n510), .A2(new_n514), .ZN(new_n518));
  INV_X1    g317(.A(new_n511), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g319(.A(new_n505), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n510), .A2(new_n511), .A3(new_n514), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n520), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT74), .ZN(new_n524));
  NAND3_X1  g323(.A1(new_n517), .A2(new_n523), .A3(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT36), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n517), .A2(new_n523), .A3(new_n524), .A4(KEYINPUT36), .ZN(new_n528));
  NAND2_X1  g327(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NOR2_X1   g328(.A1(new_n489), .A2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n434), .A2(new_n442), .A3(new_n444), .ZN(new_n531));
  AND4_X1   g330(.A1(new_n357), .A2(new_n343), .A3(new_n348), .A4(new_n350), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n357), .B1(new_n356), .B2(new_n350), .ZN(new_n533));
  NOR2_X1   g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n534), .A3(new_n353), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n463), .A2(new_n464), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n483), .A2(new_n349), .A3(new_n484), .ZN(new_n537));
  NAND4_X1  g336(.A1(new_n466), .A2(new_n469), .A3(new_n471), .A4(new_n472), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n536), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n535), .A2(new_n539), .A3(KEYINPUT85), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n487), .A2(new_n530), .A3(new_n540), .ZN(new_n541));
  AND2_X1   g340(.A1(new_n517), .A2(new_n523), .ZN(new_n542));
  NOR3_X1   g341(.A1(new_n542), .A2(new_n536), .A3(new_n538), .ZN(new_n543));
  XOR2_X1   g342(.A(KEYINPUT86), .B(KEYINPUT35), .Z(new_n544));
  NAND4_X1  g343(.A1(new_n543), .A2(KEYINPUT87), .A3(new_n359), .A4(new_n544), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT87), .ZN(new_n546));
  INV_X1    g345(.A(new_n359), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n517), .A2(new_n523), .ZN(new_n548));
  NAND4_X1  g347(.A1(new_n473), .A2(new_n548), .A3(new_n465), .A4(new_n544), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n546), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n536), .B1(new_n523), .B2(new_n517), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n551), .A2(new_n488), .A3(new_n473), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT35), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n545), .A2(new_n550), .A3(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n248), .B1(new_n541), .B2(new_n554), .ZN(new_n555));
  INV_X1    g354(.A(KEYINPUT21), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n427), .A2(G57gat), .ZN(new_n557));
  INV_X1    g356(.A(G57gat), .ZN(new_n558));
  NOR2_X1   g357(.A1(new_n558), .A2(G64gat), .ZN(new_n559));
  OAI21_X1  g358(.A(KEYINPUT9), .B1(new_n557), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(G71gat), .A2(G78gat), .ZN(new_n561));
  OR2_X1    g360(.A1(G71gat), .A2(G78gat), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n560), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT9), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n561), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT91), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(new_n558), .B2(G64gat), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n427), .A2(KEYINPUT91), .A3(G57gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n565), .B1(new_n569), .B2(new_n557), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n563), .A2(new_n570), .ZN(new_n571));
  OAI21_X1  g370(.A(new_n208), .B1(new_n556), .B2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(G183gat), .ZN(new_n573));
  INV_X1    g372(.A(G231gat), .ZN(new_n574));
  OAI21_X1  g373(.A(new_n573), .B1(new_n574), .B2(new_n361), .ZN(new_n575));
  OR2_X1    g374(.A1(new_n572), .A2(G183gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n572), .A2(G183gat), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n576), .A2(G231gat), .A3(G233gat), .A4(new_n577), .ZN(new_n578));
  XNOR2_X1  g377(.A(G127gat), .B(G155gat), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n579), .B(KEYINPUT92), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND3_X1   g380(.A1(new_n575), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(new_n581), .B1(new_n575), .B2(new_n578), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n571), .A2(new_n556), .ZN(new_n584));
  XNOR2_X1  g383(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n585));
  XNOR2_X1  g384(.A(new_n585), .B(new_n409), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n584), .B(new_n586), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  OR3_X1    g387(.A1(new_n582), .A2(new_n583), .A3(new_n588), .ZN(new_n589));
  OAI21_X1  g388(.A(new_n588), .B1(new_n582), .B2(new_n583), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(G99gat), .A2(G106gat), .ZN(new_n592));
  INV_X1    g391(.A(G85gat), .ZN(new_n593));
  AOI22_X1  g392(.A1(KEYINPUT8), .A2(new_n592), .B1(new_n593), .B2(new_n429), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n594), .B(KEYINPUT95), .ZN(new_n595));
  XNOR2_X1  g394(.A(KEYINPUT94), .B(KEYINPUT7), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n593), .A2(new_n429), .ZN(new_n597));
  XNOR2_X1  g396(.A(new_n596), .B(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  XOR2_X1   g398(.A(G99gat), .B(G106gat), .Z(new_n600));
  XNOR2_X1  g399(.A(new_n599), .B(new_n600), .ZN(new_n601));
  OAI21_X1  g400(.A(new_n601), .B1(new_n223), .B2(new_n224), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n602), .A2(KEYINPUT96), .ZN(new_n603));
  AND3_X1   g402(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n604));
  AND2_X1   g403(.A1(new_n595), .A2(new_n598), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n600), .ZN(new_n606));
  INV_X1    g405(.A(new_n600), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n599), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n606), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n604), .B1(new_n609), .B2(new_n222), .ZN(new_n610));
  INV_X1    g409(.A(KEYINPUT96), .ZN(new_n611));
  OAI211_X1 g410(.A(new_n601), .B(new_n611), .C1(new_n223), .C2(new_n224), .ZN(new_n612));
  NAND3_X1  g411(.A1(new_n603), .A2(new_n610), .A3(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(G190gat), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n603), .A2(new_n373), .A3(new_n610), .A4(new_n612), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n616), .A2(new_n410), .ZN(new_n617));
  NAND3_X1  g416(.A1(new_n614), .A2(G218gat), .A3(new_n615), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  AOI21_X1  g418(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  NAND4_X1  g420(.A1(new_n617), .A2(KEYINPUT93), .A3(new_n618), .A4(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n617), .A2(KEYINPUT93), .A3(new_n618), .ZN(new_n623));
  INV_X1    g422(.A(new_n621), .ZN(new_n624));
  NAND2_X1  g423(.A1(new_n623), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n591), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(G230gat), .A2(G233gat), .ZN(new_n628));
  INV_X1    g427(.A(new_n571), .ZN(new_n629));
  OAI21_X1  g428(.A(new_n629), .B1(new_n605), .B2(KEYINPUT97), .ZN(new_n630));
  INV_X1    g429(.A(new_n608), .ZN(new_n631));
  NOR2_X1   g430(.A1(new_n599), .A2(new_n607), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(KEYINPUT97), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n571), .B1(new_n599), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g434(.A1(new_n606), .A2(new_n635), .A3(new_n608), .ZN(new_n636));
  AOI21_X1  g435(.A(KEYINPUT10), .B1(new_n633), .B2(new_n636), .ZN(new_n637));
  INV_X1    g436(.A(KEYINPUT10), .ZN(new_n638));
  NOR3_X1   g437(.A1(new_n601), .A2(new_n638), .A3(new_n571), .ZN(new_n639));
  OAI21_X1  g438(.A(new_n628), .B1(new_n637), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(G120gat), .B(G148gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(G176gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(G204gat), .ZN(new_n643));
  INV_X1    g442(.A(new_n643), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n633), .A2(new_n636), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n640), .B(new_n644), .C1(new_n628), .C2(new_n645), .ZN(new_n646));
  AOI21_X1  g445(.A(new_n639), .B1(new_n645), .B2(new_n638), .ZN(new_n647));
  XNOR2_X1  g446(.A(new_n628), .B(KEYINPUT98), .ZN(new_n648));
  INV_X1    g447(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n647), .A2(new_n649), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n645), .A2(new_n628), .ZN(new_n651));
  NOR2_X1   g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  OAI21_X1  g451(.A(new_n646), .B1(new_n652), .B2(new_n644), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n627), .A2(new_n653), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n555), .A2(new_n654), .ZN(new_n655));
  NOR2_X1   g454(.A1(new_n655), .A2(new_n488), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(new_n203), .ZN(G1324gat));
  NOR2_X1   g456(.A1(new_n655), .A2(new_n473), .ZN(new_n658));
  OAI21_X1  g457(.A(new_n658), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n659), .B1(KEYINPUT16), .B2(G8gat), .ZN(new_n660));
  XOR2_X1   g459(.A(new_n660), .B(KEYINPUT42), .Z(new_n661));
  OAI21_X1  g460(.A(new_n661), .B1(new_n207), .B2(new_n658), .ZN(G1325gat));
  INV_X1    g461(.A(new_n655), .ZN(new_n663));
  AOI21_X1  g462(.A(G15gat), .B1(new_n663), .B2(new_n548), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n529), .A2(G15gat), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n665), .B(KEYINPUT99), .ZN(new_n666));
  AOI21_X1  g465(.A(new_n664), .B1(new_n663), .B2(new_n666), .ZN(G1326gat));
  NOR2_X1   g466(.A1(new_n655), .A2(new_n465), .ZN(new_n668));
  XOR2_X1   g467(.A(KEYINPUT43), .B(G22gat), .Z(new_n669));
  XNOR2_X1  g468(.A(new_n668), .B(new_n669), .ZN(G1327gat));
  NAND2_X1  g469(.A1(new_n625), .A2(new_n622), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(new_n653), .ZN(new_n673));
  NAND3_X1  g472(.A1(new_n672), .A2(new_n591), .A3(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(KEYINPUT100), .ZN(new_n675));
  OR2_X1    g474(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  AND2_X1   g475(.A1(new_n555), .A2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n675), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  NOR3_X1   g478(.A1(new_n679), .A2(G29gat), .A3(new_n488), .ZN(new_n680));
  XOR2_X1   g479(.A(new_n680), .B(KEYINPUT45), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n541), .A2(new_n554), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n682), .A2(new_n672), .ZN(new_n683));
  INV_X1    g482(.A(KEYINPUT44), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n653), .B(KEYINPUT101), .Z(new_n686));
  NOR2_X1   g485(.A1(new_n686), .A2(new_n248), .ZN(new_n687));
  AOI21_X1  g486(.A(new_n671), .B1(new_n541), .B2(new_n554), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n688), .A2(KEYINPUT44), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n685), .A2(new_n591), .A3(new_n687), .A4(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT102), .ZN(new_n691));
  AOI21_X1  g490(.A(KEYINPUT44), .B1(new_n682), .B2(new_n672), .ZN(new_n692));
  AOI211_X1 g491(.A(new_n684), .B(new_n671), .C1(new_n541), .C2(new_n554), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(KEYINPUT102), .ZN(new_n695));
  NAND4_X1  g494(.A1(new_n694), .A2(new_n695), .A3(new_n591), .A4(new_n687), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n488), .B1(new_n691), .B2(new_n696), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n681), .B1(new_n210), .B2(new_n697), .ZN(G1328gat));
  NOR3_X1   g497(.A1(new_n679), .A2(G36gat), .A3(new_n473), .ZN(new_n699));
  XNOR2_X1  g498(.A(new_n699), .B(KEYINPUT46), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n473), .B1(new_n691), .B2(new_n696), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n700), .B1(new_n211), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  OAI211_X1 g503(.A(new_n700), .B(KEYINPUT103), .C1(new_n211), .C2(new_n701), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n704), .A2(new_n705), .ZN(G1329gat));
  NOR3_X1   g505(.A1(new_n679), .A2(G43gat), .A3(new_n542), .ZN(new_n707));
  INV_X1    g506(.A(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n529), .ZN(new_n709));
  OAI21_X1  g508(.A(G43gat), .B1(new_n690), .B2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n708), .A2(KEYINPUT47), .A3(new_n710), .ZN(new_n711));
  INV_X1    g510(.A(new_n687), .ZN(new_n712));
  NOR3_X1   g511(.A1(new_n692), .A2(new_n693), .A3(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n695), .B1(new_n713), .B2(new_n591), .ZN(new_n714));
  NOR2_X1   g513(.A1(new_n690), .A2(KEYINPUT102), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n529), .B1(new_n714), .B2(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n707), .B1(new_n716), .B2(G43gat), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n711), .B1(new_n717), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g517(.A(new_n536), .B1(new_n714), .B2(new_n715), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n719), .A2(KEYINPUT104), .A3(G50gat), .ZN(new_n720));
  INV_X1    g519(.A(G50gat), .ZN(new_n721));
  NAND4_X1  g520(.A1(new_n677), .A2(new_n721), .A3(new_n536), .A4(new_n678), .ZN(new_n722));
  INV_X1    g521(.A(KEYINPUT104), .ZN(new_n723));
  AOI21_X1  g522(.A(new_n465), .B1(new_n691), .B2(new_n696), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n723), .B1(new_n724), .B2(new_n721), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n720), .A2(new_n722), .A3(new_n725), .ZN(new_n726));
  INV_X1    g525(.A(KEYINPUT48), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OAI21_X1  g527(.A(G50gat), .B1(new_n690), .B2(new_n465), .ZN(new_n729));
  NAND3_X1  g528(.A1(new_n729), .A2(KEYINPUT48), .A3(new_n722), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n728), .A2(new_n730), .ZN(G1331gat));
  NAND4_X1  g530(.A1(new_n682), .A2(new_n248), .A3(new_n626), .A4(new_n686), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n732), .A2(new_n488), .ZN(new_n733));
  XNOR2_X1  g532(.A(new_n733), .B(new_n558), .ZN(G1332gat));
  AOI211_X1 g533(.A(new_n473), .B(new_n732), .C1(KEYINPUT49), .C2(G64gat), .ZN(new_n735));
  NOR2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  XNOR2_X1  g535(.A(new_n735), .B(new_n736), .ZN(G1333gat));
  OAI21_X1  g536(.A(G71gat), .B1(new_n732), .B2(new_n709), .ZN(new_n738));
  OR2_X1    g537(.A1(new_n732), .A2(G71gat), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n738), .B1(new_n739), .B2(new_n542), .ZN(new_n740));
  XOR2_X1   g539(.A(new_n740), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g540(.A1(new_n732), .A2(new_n465), .ZN(new_n742));
  XOR2_X1   g541(.A(new_n742), .B(G78gat), .Z(G1335gat));
  INV_X1    g542(.A(new_n591), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n744), .A2(new_n247), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n688), .A2(new_n745), .ZN(new_n746));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n688), .A2(KEYINPUT51), .A3(new_n745), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n751), .A2(KEYINPUT105), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n748), .A2(KEYINPUT105), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NOR2_X1   g553(.A1(new_n754), .A2(new_n673), .ZN(new_n755));
  INV_X1    g554(.A(new_n488), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n755), .A2(new_n593), .A3(new_n756), .ZN(new_n757));
  NOR3_X1   g556(.A1(new_n692), .A2(new_n693), .A3(new_n673), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n758), .A2(new_n745), .ZN(new_n759));
  OAI21_X1  g558(.A(G85gat), .B1(new_n759), .B2(new_n488), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n757), .A2(new_n760), .ZN(G1336gat));
  INV_X1    g560(.A(KEYINPUT106), .ZN(new_n762));
  OAI21_X1  g561(.A(new_n762), .B1(new_n759), .B2(new_n473), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n758), .A2(KEYINPUT106), .A3(new_n538), .A4(new_n745), .ZN(new_n764));
  NAND3_X1  g563(.A1(new_n763), .A2(G92gat), .A3(new_n764), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT52), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n686), .A2(new_n429), .A3(new_n538), .ZN(new_n767));
  OAI211_X1 g566(.A(new_n765), .B(new_n766), .C1(new_n754), .C2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G92gat), .B1(new_n759), .B2(new_n473), .ZN(new_n769));
  OAI21_X1  g568(.A(new_n769), .B1(new_n751), .B2(new_n767), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n768), .A2(new_n771), .ZN(G1337gat));
  XOR2_X1   g571(.A(KEYINPUT107), .B(G99gat), .Z(new_n773));
  NOR2_X1   g572(.A1(new_n542), .A2(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n755), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g574(.A(new_n773), .B1(new_n759), .B2(new_n709), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n775), .A2(new_n776), .ZN(G1338gat));
  NAND3_X1  g576(.A1(new_n758), .A2(new_n536), .A3(new_n745), .ZN(new_n778));
  AND2_X1   g577(.A1(new_n778), .A2(G106gat), .ZN(new_n779));
  NOR2_X1   g578(.A1(new_n779), .A2(KEYINPUT53), .ZN(new_n780));
  INV_X1    g579(.A(new_n686), .ZN(new_n781));
  NOR3_X1   g580(.A1(new_n781), .A2(G106gat), .A3(new_n465), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n752), .A2(new_n753), .A3(new_n782), .ZN(new_n783));
  AND2_X1   g582(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(KEYINPUT108), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n780), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n750), .A2(new_n782), .ZN(new_n787));
  OAI21_X1  g586(.A(KEYINPUT53), .B1(new_n779), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n786), .A2(new_n788), .ZN(G1339gat));
  INV_X1    g588(.A(KEYINPUT54), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n644), .B1(new_n650), .B2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT109), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n790), .B1(new_n647), .B2(new_n649), .ZN(new_n793));
  AOI21_X1  g592(.A(new_n792), .B1(new_n793), .B2(new_n640), .ZN(new_n794));
  INV_X1    g593(.A(new_n636), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n635), .B1(new_n608), .B2(new_n606), .ZN(new_n796));
  OAI21_X1  g595(.A(new_n638), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(new_n639), .ZN(new_n798));
  NAND3_X1  g597(.A1(new_n797), .A2(new_n798), .A3(new_n649), .ZN(new_n799));
  AND4_X1   g598(.A1(new_n792), .A2(new_n799), .A3(new_n640), .A4(KEYINPUT54), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n791), .B1(new_n794), .B2(new_n800), .ZN(new_n801));
  INV_X1    g600(.A(KEYINPUT55), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g602(.A(KEYINPUT55), .B(new_n791), .C1(new_n794), .C2(new_n800), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n803), .A2(new_n247), .A3(new_n646), .A4(new_n804), .ZN(new_n805));
  OR3_X1    g604(.A1(new_n228), .A2(KEYINPUT110), .A3(new_n229), .ZN(new_n806));
  OAI21_X1  g605(.A(KEYINPUT110), .B1(new_n228), .B2(new_n229), .ZN(new_n807));
  OAI211_X1 g606(.A(new_n806), .B(new_n807), .C1(new_n234), .C2(new_n233), .ZN(new_n808));
  AOI22_X1  g607(.A1(new_n808), .A2(new_n242), .B1(new_n238), .B2(new_n243), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n809), .A2(new_n653), .ZN(new_n810));
  AOI22_X1  g609(.A1(new_n805), .A2(new_n810), .B1(new_n622), .B2(new_n625), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n803), .A2(new_n646), .A3(new_n804), .ZN(new_n812));
  NAND3_X1  g611(.A1(new_n625), .A2(new_n622), .A3(new_n809), .ZN(new_n813));
  NOR2_X1   g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n591), .B1(new_n811), .B2(new_n814), .ZN(new_n815));
  NAND4_X1  g614(.A1(new_n671), .A2(new_n744), .A3(new_n248), .A4(new_n673), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g616(.A1(new_n817), .A2(new_n551), .ZN(new_n818));
  NOR2_X1   g617(.A1(new_n488), .A2(new_n538), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR2_X1   g619(.A1(new_n820), .A2(new_n248), .ZN(new_n821));
  XNOR2_X1  g620(.A(KEYINPUT111), .B(G113gat), .ZN(new_n822));
  XNOR2_X1  g621(.A(new_n821), .B(new_n822), .ZN(G1340gat));
  INV_X1    g622(.A(new_n820), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n824), .A2(new_n266), .A3(new_n653), .ZN(new_n825));
  OAI21_X1  g624(.A(G120gat), .B1(new_n820), .B2(new_n781), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(G1341gat));
  NOR2_X1   g626(.A1(new_n820), .A2(new_n591), .ZN(new_n828));
  XNOR2_X1  g627(.A(new_n828), .B(new_n256), .ZN(G1342gat));
  NAND2_X1  g628(.A1(new_n824), .A2(new_n672), .ZN(new_n830));
  NOR2_X1   g629(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n831));
  AND2_X1   g630(.A1(KEYINPUT56), .A2(G134gat), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n830), .A2(new_n831), .A3(new_n832), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n830), .B2(new_n831), .ZN(G1343gat));
  NAND2_X1  g633(.A1(new_n709), .A2(new_n819), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n817), .A2(new_n536), .ZN(new_n836));
  XNOR2_X1  g635(.A(KEYINPUT112), .B(KEYINPUT57), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n465), .B1(new_n815), .B2(new_n816), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT57), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  OAI21_X1  g641(.A(G141gat), .B1(new_n842), .B2(new_n248), .ZN(new_n843));
  INV_X1    g642(.A(new_n835), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n839), .A2(new_n844), .ZN(new_n845));
  INV_X1    g644(.A(new_n845), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n846), .A2(new_n288), .A3(new_n247), .ZN(new_n847));
  XOR2_X1   g646(.A(KEYINPUT114), .B(KEYINPUT58), .Z(new_n848));
  NAND3_X1  g647(.A1(new_n843), .A2(new_n847), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n849), .A2(new_n850), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n849), .A2(new_n850), .ZN(new_n852));
  INV_X1    g651(.A(new_n847), .ZN(new_n853));
  AOI21_X1  g652(.A(KEYINPUT113), .B1(new_n838), .B2(new_n841), .ZN(new_n854));
  INV_X1    g653(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n838), .A2(KEYINPUT113), .A3(new_n841), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(new_n247), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n853), .B1(new_n858), .B2(G141gat), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT58), .ZN(new_n860));
  OAI211_X1 g659(.A(new_n851), .B(new_n852), .C1(new_n859), .C2(new_n860), .ZN(G1344gat));
  NAND2_X1  g660(.A1(new_n805), .A2(new_n810), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n671), .ZN(new_n863));
  OR2_X1    g662(.A1(new_n812), .A2(new_n813), .ZN(new_n864));
  AOI21_X1  g663(.A(new_n744), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT117), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n816), .A2(new_n866), .ZN(new_n867));
  NAND4_X1  g666(.A1(new_n626), .A2(KEYINPUT117), .A3(new_n248), .A4(new_n673), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  OAI21_X1  g668(.A(KEYINPUT118), .B1(new_n865), .B2(new_n869), .ZN(new_n870));
  INV_X1    g669(.A(KEYINPUT118), .ZN(new_n871));
  NAND4_X1  g670(.A1(new_n815), .A2(new_n871), .A3(new_n867), .A4(new_n868), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n870), .A2(new_n536), .A3(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n840), .ZN(new_n874));
  INV_X1    g673(.A(new_n837), .ZN(new_n875));
  AOI211_X1 g674(.A(new_n465), .B(new_n875), .C1(new_n815), .C2(new_n816), .ZN(new_n876));
  INV_X1    g675(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n874), .A2(new_n877), .ZN(new_n878));
  XOR2_X1   g677(.A(KEYINPUT116), .B(KEYINPUT59), .Z(new_n879));
  NAND4_X1  g678(.A1(new_n878), .A2(new_n653), .A3(new_n844), .A4(new_n879), .ZN(new_n880));
  INV_X1    g679(.A(new_n856), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n881), .A2(new_n854), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n882), .A2(new_n673), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n880), .B1(new_n883), .B2(KEYINPUT59), .ZN(new_n884));
  AOI21_X1  g683(.A(G148gat), .B1(new_n846), .B2(new_n653), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n884), .A2(G148gat), .B1(new_n879), .B2(new_n885), .ZN(G1345gat));
  AOI21_X1  g685(.A(G155gat), .B1(new_n846), .B2(new_n744), .ZN(new_n887));
  NAND2_X1  g686(.A1(new_n744), .A2(G155gat), .ZN(new_n888));
  XOR2_X1   g687(.A(new_n888), .B(KEYINPUT119), .Z(new_n889));
  AOI21_X1  g688(.A(new_n887), .B1(new_n857), .B2(new_n889), .ZN(G1346gat));
  AOI21_X1  g689(.A(G162gat), .B1(new_n846), .B2(new_n672), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n882), .A2(new_n671), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n891), .B1(new_n892), .B2(G162gat), .ZN(G1347gat));
  INV_X1    g692(.A(G169gat), .ZN(new_n894));
  NOR2_X1   g693(.A1(new_n756), .A2(new_n473), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n818), .A2(new_n896), .ZN(new_n897));
  AOI21_X1  g696(.A(new_n894), .B1(new_n897), .B2(new_n247), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n818), .A2(new_n895), .ZN(new_n899));
  NOR3_X1   g698(.A1(new_n899), .A2(G169gat), .A3(new_n248), .ZN(new_n900));
  OR2_X1    g699(.A1(new_n898), .A2(new_n900), .ZN(G1348gat));
  NAND3_X1  g700(.A1(new_n897), .A2(G176gat), .A3(new_n686), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n899), .A2(new_n673), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n902), .B1(G176gat), .B2(new_n903), .ZN(new_n904));
  XNOR2_X1  g703(.A(new_n904), .B(KEYINPUT121), .ZN(G1349gat));
  AOI21_X1  g704(.A(new_n372), .B1(new_n897), .B2(new_n744), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n385), .A2(new_n386), .ZN(new_n907));
  NOR3_X1   g706(.A1(new_n899), .A2(new_n907), .A3(new_n591), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n906), .A2(new_n908), .ZN(new_n909));
  XOR2_X1   g708(.A(new_n909), .B(KEYINPUT60), .Z(G1350gat));
  NAND2_X1  g709(.A1(new_n897), .A2(new_n672), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(G190gat), .ZN(new_n912));
  INV_X1    g711(.A(KEYINPUT122), .ZN(new_n913));
  OAI21_X1  g712(.A(KEYINPUT61), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n912), .A2(new_n913), .ZN(new_n915));
  XNOR2_X1  g714(.A(new_n914), .B(new_n915), .ZN(new_n916));
  NAND4_X1  g715(.A1(new_n818), .A2(new_n373), .A3(new_n672), .A4(new_n895), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1351gat));
  NOR2_X1   g717(.A1(new_n836), .A2(new_n529), .ZN(new_n919));
  NAND2_X1  g718(.A1(new_n919), .A2(new_n895), .ZN(new_n920));
  INV_X1    g719(.A(new_n920), .ZN(new_n921));
  INV_X1    g720(.A(G197gat), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n921), .A2(new_n922), .A3(new_n247), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n896), .A2(new_n709), .ZN(new_n924));
  INV_X1    g723(.A(new_n924), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n876), .B1(new_n873), .B2(new_n840), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n925), .B1(new_n926), .B2(KEYINPUT123), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT123), .ZN(new_n928));
  AOI211_X1 g727(.A(new_n928), .B(new_n876), .C1(new_n873), .C2(new_n840), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n927), .A2(new_n248), .A3(new_n929), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n923), .B1(new_n930), .B2(new_n922), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n931), .A2(KEYINPUT124), .ZN(new_n932));
  INV_X1    g731(.A(KEYINPUT124), .ZN(new_n933));
  OAI211_X1 g732(.A(new_n933), .B(new_n923), .C1(new_n930), .C2(new_n922), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n932), .A2(new_n934), .ZN(G1352gat));
  INV_X1    g734(.A(KEYINPUT126), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n924), .B1(new_n878), .B2(new_n928), .ZN(new_n937));
  INV_X1    g736(.A(new_n929), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n936), .B1(new_n939), .B2(new_n781), .ZN(new_n940));
  NAND4_X1  g739(.A1(new_n937), .A2(KEYINPUT126), .A3(new_n686), .A4(new_n938), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n940), .A2(G204gat), .A3(new_n941), .ZN(new_n942));
  NOR3_X1   g741(.A1(new_n920), .A2(G204gat), .A3(new_n673), .ZN(new_n943));
  XNOR2_X1  g742(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n943), .B(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n942), .A2(new_n945), .ZN(G1353gat));
  NAND3_X1  g745(.A1(new_n921), .A2(new_n409), .A3(new_n744), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT127), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n924), .B1(new_n874), .B2(new_n877), .ZN(new_n949));
  AOI21_X1  g748(.A(new_n948), .B1(new_n949), .B2(new_n744), .ZN(new_n950));
  NOR4_X1   g749(.A1(new_n926), .A2(KEYINPUT127), .A3(new_n591), .A4(new_n924), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(KEYINPUT63), .B1(new_n952), .B2(G211gat), .ZN(new_n953));
  INV_X1    g752(.A(KEYINPUT63), .ZN(new_n954));
  NOR4_X1   g753(.A1(new_n950), .A2(new_n951), .A3(new_n954), .A4(new_n409), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n947), .B1(new_n953), .B2(new_n955), .ZN(G1354gat));
  OAI21_X1  g755(.A(G218gat), .B1(new_n939), .B2(new_n671), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n921), .A2(new_n410), .A3(new_n672), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1355gat));
endmodule


