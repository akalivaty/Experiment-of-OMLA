//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 0 1 1 0 1 1 0 1 0 1 0 1 0 0 0 0 1 1 0 1 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 0 0 0 0 1 0 0 0 0 1 1 1 0 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n713, new_n714, new_n715, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n724, new_n726, new_n727,
    new_n728, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n755, new_n756, new_n757,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n788, new_n789, new_n790, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n813, new_n814, new_n815, new_n816, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n928, new_n929, new_n930, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n991, new_n992, new_n993, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008;
  INV_X1    g000(.A(KEYINPUT70), .ZN(new_n187));
  INV_X1    g001(.A(G128), .ZN(new_n188));
  OAI21_X1  g002(.A(new_n187), .B1(new_n188), .B2(G119), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n188), .A2(G119), .ZN(new_n190));
  INV_X1    g004(.A(G119), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n191), .A2(KEYINPUT70), .A3(G128), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n189), .A2(new_n190), .A3(new_n192), .ZN(new_n193));
  XNOR2_X1  g007(.A(KEYINPUT24), .B(G110), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(KEYINPUT23), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n190), .A2(new_n196), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n188), .A2(KEYINPUT23), .A3(G119), .ZN(new_n198));
  INV_X1    g012(.A(G110), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n191), .A2(G128), .ZN(new_n200));
  NAND4_X1  g014(.A1(new_n197), .A2(new_n198), .A3(new_n199), .A4(new_n200), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n195), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(KEYINPUT71), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT71), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n204), .A3(new_n201), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G140), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G125), .ZN(new_n208));
  INV_X1    g022(.A(G125), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G140), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n208), .A2(new_n210), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G146), .ZN(new_n212));
  NOR3_X1   g026(.A1(new_n209), .A2(KEYINPUT16), .A3(G140), .ZN(new_n213));
  XNOR2_X1  g027(.A(G125), .B(G140), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n213), .B1(new_n214), .B2(KEYINPUT16), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n212), .B1(new_n215), .B2(G146), .ZN(new_n216));
  AOI21_X1  g030(.A(KEYINPUT72), .B1(new_n206), .B2(new_n216), .ZN(new_n217));
  AND3_X1   g031(.A1(new_n195), .A2(new_n204), .A3(new_n201), .ZN(new_n218));
  AOI21_X1  g032(.A(new_n204), .B1(new_n195), .B2(new_n201), .ZN(new_n219));
  OAI211_X1 g033(.A(KEYINPUT72), .B(new_n216), .C1(new_n218), .C2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(new_n220), .ZN(new_n221));
  INV_X1    g035(.A(new_n213), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT16), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n222), .B1(new_n211), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G146), .ZN(new_n225));
  NOR2_X1   g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n215), .A2(G146), .ZN(new_n227));
  NOR2_X1   g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  AND3_X1   g042(.A1(new_n197), .A2(new_n200), .A3(new_n198), .ZN(new_n229));
  OAI22_X1  g043(.A1(new_n229), .A2(new_n199), .B1(new_n194), .B2(new_n193), .ZN(new_n230));
  OAI22_X1  g044(.A1(new_n217), .A2(new_n221), .B1(new_n228), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT22), .B(G137), .ZN(new_n232));
  INV_X1    g046(.A(G953), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n233), .A2(G221), .A3(G234), .ZN(new_n234));
  XNOR2_X1  g048(.A(new_n232), .B(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n231), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n228), .A2(new_n230), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n216), .B1(new_n218), .B2(new_n219), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT72), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n239), .A2(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n238), .B1(new_n241), .B2(new_n220), .ZN(new_n242));
  INV_X1    g056(.A(new_n235), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n237), .A3(new_n244), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n236), .A2(new_n244), .A3(KEYINPUT25), .A4(new_n237), .ZN(new_n248));
  AND3_X1   g062(.A1(new_n247), .A2(KEYINPUT73), .A3(new_n248), .ZN(new_n249));
  INV_X1    g063(.A(G217), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n250), .B1(G234), .B2(new_n237), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n251), .B1(new_n247), .B2(KEYINPUT73), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT74), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n242), .A2(new_n243), .ZN(new_n254));
  AOI211_X1 g068(.A(new_n235), .B(new_n238), .C1(new_n241), .C2(new_n220), .ZN(new_n255));
  OAI21_X1  g069(.A(new_n253), .B1(new_n254), .B2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n254), .A2(new_n255), .A3(new_n253), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n251), .A2(G902), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  OAI22_X1  g075(.A1(new_n249), .A2(new_n252), .B1(new_n259), .B2(new_n261), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n225), .A2(G143), .ZN(new_n263));
  INV_X1    g077(.A(G143), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n264), .A2(G146), .ZN(new_n265));
  AND2_X1   g079(.A1(KEYINPUT0), .A2(G128), .ZN(new_n266));
  NAND3_X1  g080(.A1(new_n263), .A2(new_n265), .A3(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(KEYINPUT65), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT65), .ZN(new_n269));
  NAND4_X1  g083(.A1(new_n263), .A2(new_n265), .A3(new_n266), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n264), .A2(G146), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT64), .B1(new_n225), .B2(G143), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT64), .ZN(new_n274));
  NAND3_X1  g088(.A1(new_n274), .A2(new_n264), .A3(G146), .ZN(new_n275));
  AOI21_X1  g089(.A(new_n272), .B1(new_n273), .B2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(KEYINPUT0), .B(G128), .ZN(new_n277));
  NOR2_X1   g091(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g092(.A1(new_n271), .A2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT11), .ZN(new_n280));
  INV_X1    g094(.A(G134), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n280), .B1(new_n281), .B2(G137), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(G137), .ZN(new_n283));
  INV_X1    g097(.A(G137), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n284), .A2(KEYINPUT11), .A3(G134), .ZN(new_n285));
  NAND3_X1  g099(.A1(new_n282), .A2(new_n283), .A3(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(G131), .ZN(new_n287));
  INV_X1    g101(.A(G131), .ZN(new_n288));
  NAND4_X1  g102(.A1(new_n282), .A2(new_n285), .A3(new_n288), .A4(new_n283), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND3_X1  g104(.A1(new_n279), .A2(KEYINPUT67), .A3(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(KEYINPUT67), .ZN(new_n292));
  AND2_X1   g106(.A1(new_n287), .A2(new_n289), .ZN(new_n293));
  OAI211_X1 g107(.A(new_n268), .B(new_n270), .C1(new_n276), .C2(new_n277), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n291), .A2(new_n295), .ZN(new_n296));
  NOR2_X1   g110(.A1(new_n281), .A2(G137), .ZN(new_n297));
  NOR2_X1   g111(.A1(new_n284), .A2(G134), .ZN(new_n298));
  OAI21_X1  g112(.A(G131), .B1(new_n297), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g113(.A1(new_n289), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(KEYINPUT1), .ZN(new_n301));
  NAND4_X1  g115(.A1(new_n263), .A2(new_n265), .A3(new_n301), .A4(G128), .ZN(new_n302));
  AOI21_X1  g116(.A(new_n188), .B1(new_n263), .B2(KEYINPUT1), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n302), .B1(new_n276), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n300), .A2(new_n304), .A3(KEYINPUT68), .ZN(new_n305));
  AOI21_X1  g119(.A(KEYINPUT68), .B1(new_n300), .B2(new_n304), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n296), .A2(new_n307), .A3(KEYINPUT30), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n279), .A2(new_n290), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n300), .A2(new_n304), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n310), .A2(KEYINPUT66), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n300), .A2(new_n304), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n309), .A2(new_n311), .A3(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT30), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n191), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(G116), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G119), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n320), .ZN(new_n321));
  XNOR2_X1  g135(.A(KEYINPUT2), .B(G113), .ZN(new_n322));
  INV_X1    g136(.A(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n320), .A2(new_n322), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n308), .A2(new_n316), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n326), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n296), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT69), .B(KEYINPUT27), .Z(new_n330));
  INV_X1    g144(.A(G237), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n331), .A2(new_n233), .A3(G210), .ZN(new_n332));
  XNOR2_X1  g146(.A(new_n330), .B(new_n332), .ZN(new_n333));
  XNOR2_X1  g147(.A(KEYINPUT26), .B(G101), .ZN(new_n334));
  XNOR2_X1  g148(.A(new_n333), .B(new_n334), .ZN(new_n335));
  NAND3_X1  g149(.A1(new_n327), .A2(new_n329), .A3(new_n335), .ZN(new_n336));
  INV_X1    g150(.A(KEYINPUT31), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NAND4_X1  g152(.A1(new_n327), .A2(KEYINPUT31), .A3(new_n329), .A4(new_n335), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n326), .B1(new_n304), .B2(new_n300), .ZN(new_n341));
  AOI21_X1  g155(.A(KEYINPUT28), .B1(new_n309), .B2(new_n341), .ZN(new_n342));
  INV_X1    g156(.A(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n314), .A2(new_n326), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n329), .A2(new_n344), .ZN(new_n345));
  INV_X1    g159(.A(KEYINPUT28), .ZN(new_n346));
  OAI21_X1  g160(.A(new_n343), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g161(.A(new_n335), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n340), .A2(new_n349), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT32), .ZN(new_n351));
  NOR2_X1   g165(.A1(G472), .A2(G902), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n350), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  AOI22_X1  g167(.A1(new_n338), .A2(new_n339), .B1(new_n347), .B2(new_n348), .ZN(new_n354));
  INV_X1    g168(.A(new_n352), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT32), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n353), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G472), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n296), .A2(new_n307), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n326), .ZN(new_n360));
  AOI21_X1  g174(.A(new_n346), .B1(new_n360), .B2(new_n329), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n361), .A2(new_n342), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT29), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n348), .A2(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n327), .A2(new_n329), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n366), .A2(new_n348), .ZN(new_n367));
  OAI211_X1 g181(.A(new_n367), .B(new_n363), .C1(new_n347), .C2(new_n348), .ZN(new_n368));
  AOI21_X1  g182(.A(new_n358), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  AOI21_X1  g184(.A(new_n262), .B1(new_n357), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(G469), .ZN(new_n372));
  XNOR2_X1  g186(.A(G110), .B(G140), .ZN(new_n373));
  INV_X1    g187(.A(G227), .ZN(new_n374));
  NOR2_X1   g188(.A1(new_n374), .A2(G953), .ZN(new_n375));
  XNOR2_X1  g189(.A(new_n373), .B(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G104), .ZN(new_n378));
  NOR2_X1   g192(.A1(new_n378), .A2(KEYINPUT3), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT76), .ZN(new_n380));
  INV_X1    g194(.A(G107), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT76), .A2(G107), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n379), .A2(new_n382), .A3(new_n383), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n385));
  INV_X1    g199(.A(KEYINPUT75), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G104), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n385), .A2(new_n387), .A3(G107), .ZN(new_n388));
  AOI21_X1  g202(.A(G107), .B1(new_n385), .B2(new_n387), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT3), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n384), .B(new_n388), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT4), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n391), .A2(new_n392), .A3(G101), .ZN(new_n393));
  AND2_X1   g207(.A1(new_n279), .A2(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n386), .A2(G104), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n396));
  OAI21_X1  g210(.A(new_n381), .B1(new_n395), .B2(new_n396), .ZN(new_n397));
  AND2_X1   g211(.A1(KEYINPUT76), .A2(G107), .ZN(new_n398));
  NOR2_X1   g212(.A1(KEYINPUT76), .A2(G107), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n397), .A2(KEYINPUT3), .B1(new_n400), .B2(new_n379), .ZN(new_n401));
  INV_X1    g215(.A(G101), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n388), .A2(new_n402), .ZN(new_n403));
  INV_X1    g217(.A(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n391), .A2(G101), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(KEYINPUT4), .ZN(new_n407));
  AOI21_X1  g221(.A(G104), .B1(new_n382), .B2(new_n383), .ZN(new_n408));
  OAI21_X1  g222(.A(G101), .B1(new_n389), .B2(new_n408), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT77), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n378), .B1(new_n398), .B2(new_n399), .ZN(new_n412));
  XNOR2_X1  g226(.A(KEYINPUT75), .B(G104), .ZN(new_n413));
  OAI21_X1  g227(.A(new_n412), .B1(new_n413), .B2(G107), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n414), .A2(KEYINPUT77), .A3(G101), .ZN(new_n415));
  AOI22_X1  g229(.A1(new_n411), .A2(new_n415), .B1(new_n401), .B2(new_n404), .ZN(new_n416));
  INV_X1    g230(.A(new_n304), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT10), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AOI22_X1  g233(.A1(new_n394), .A2(new_n407), .B1(new_n416), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n411), .A2(new_n415), .ZN(new_n421));
  OAI21_X1  g235(.A(G128), .B1(new_n272), .B2(new_n301), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n263), .A2(new_n265), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI22_X1  g238(.A1(new_n401), .A2(new_n404), .B1(new_n302), .B2(new_n424), .ZN(new_n425));
  AOI211_X1 g239(.A(KEYINPUT78), .B(KEYINPUT10), .C1(new_n421), .C2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(KEYINPUT78), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n424), .A2(new_n302), .ZN(new_n428));
  AOI211_X1 g242(.A(new_n410), .B(new_n402), .C1(new_n397), .C2(new_n412), .ZN(new_n429));
  AOI21_X1  g243(.A(KEYINPUT77), .B1(new_n414), .B2(G101), .ZN(new_n430));
  OAI211_X1 g244(.A(new_n405), .B(new_n428), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n427), .B1(new_n431), .B2(new_n418), .ZN(new_n432));
  OAI21_X1  g246(.A(new_n420), .B1(new_n426), .B2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n290), .ZN(new_n434));
  OAI211_X1 g248(.A(new_n293), .B(new_n420), .C1(new_n426), .C2(new_n432), .ZN(new_n435));
  AOI21_X1  g249(.A(new_n377), .B1(new_n434), .B2(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT12), .ZN(new_n437));
  OAI21_X1  g251(.A(new_n405), .B1(new_n429), .B2(new_n430), .ZN(new_n438));
  AOI22_X1  g252(.A1(new_n438), .A2(new_n417), .B1(new_n421), .B2(new_n425), .ZN(new_n439));
  OAI21_X1  g253(.A(new_n437), .B1(new_n439), .B2(new_n293), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n431), .B1(new_n416), .B2(new_n304), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n441), .A2(KEYINPUT12), .A3(new_n290), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  AND3_X1   g257(.A1(new_n443), .A2(new_n435), .A3(new_n377), .ZN(new_n444));
  OAI211_X1 g258(.A(new_n372), .B(new_n237), .C1(new_n436), .C2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n443), .A2(new_n435), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n446), .A2(new_n376), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n435), .A2(KEYINPUT79), .A3(new_n377), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n448), .A2(new_n434), .ZN(new_n449));
  AOI21_X1  g263(.A(KEYINPUT79), .B1(new_n435), .B2(new_n377), .ZN(new_n450));
  OAI211_X1 g264(.A(new_n447), .B(G469), .C1(new_n449), .C2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(G469), .A2(G902), .ZN(new_n452));
  NAND3_X1  g266(.A1(new_n445), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  XNOR2_X1  g267(.A(KEYINPUT9), .B(G234), .ZN(new_n454));
  OAI21_X1  g268(.A(G221), .B1(new_n454), .B2(G902), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n453), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT96), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n264), .A2(G128), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n188), .A2(G143), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n460), .A2(G134), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n458), .A2(new_n459), .A3(new_n281), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n318), .A2(G122), .ZN(new_n464));
  INV_X1    g278(.A(G122), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n465), .A2(G116), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n400), .A2(new_n464), .A3(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(KEYINPUT14), .B1(new_n465), .B2(G116), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT14), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n318), .A3(G122), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n468), .A2(new_n470), .A3(new_n466), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G107), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n463), .A2(new_n467), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(KEYINPUT95), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT95), .ZN(new_n475));
  NAND4_X1  g289(.A1(new_n463), .A2(new_n475), .A3(new_n472), .A4(new_n467), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  AND4_X1   g291(.A1(new_n382), .A2(new_n464), .A3(new_n466), .A4(new_n383), .ZN(new_n478));
  AOI22_X1  g292(.A1(new_n464), .A2(new_n466), .B1(new_n382), .B2(new_n383), .ZN(new_n479));
  OAI21_X1  g293(.A(new_n462), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  INV_X1    g294(.A(KEYINPUT13), .ZN(new_n481));
  AOI21_X1  g295(.A(new_n481), .B1(new_n188), .B2(G143), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n188), .A2(G143), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT93), .B1(new_n482), .B2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n459), .A2(KEYINPUT13), .ZN(new_n485));
  INV_X1    g299(.A(KEYINPUT93), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n485), .A2(new_n486), .A3(new_n458), .ZN(new_n487));
  INV_X1    g301(.A(KEYINPUT94), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n483), .A2(new_n488), .A3(KEYINPUT13), .ZN(new_n489));
  OAI21_X1  g303(.A(KEYINPUT94), .B1(new_n458), .B2(new_n481), .ZN(new_n490));
  NAND4_X1  g304(.A1(new_n484), .A2(new_n487), .A3(new_n489), .A4(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n480), .B1(G134), .B2(new_n491), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n457), .B1(new_n477), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n491), .A2(G134), .ZN(new_n494));
  OR2_X1    g308(.A1(new_n478), .A2(new_n479), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n494), .A2(new_n495), .A3(new_n462), .ZN(new_n496));
  NAND4_X1  g310(.A1(new_n496), .A2(KEYINPUT96), .A3(new_n474), .A4(new_n476), .ZN(new_n497));
  NOR3_X1   g311(.A1(new_n454), .A2(new_n250), .A3(G953), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n493), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n496), .A2(new_n474), .A3(new_n476), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n457), .A3(new_n498), .ZN(new_n502));
  NAND4_X1  g316(.A1(new_n500), .A2(KEYINPUT98), .A3(new_n237), .A4(new_n502), .ZN(new_n503));
  INV_X1    g317(.A(KEYINPUT97), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g319(.A1(new_n500), .A2(KEYINPUT97), .A3(new_n237), .A4(new_n502), .ZN(new_n506));
  INV_X1    g320(.A(G478), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n507), .A2(KEYINPUT15), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n506), .A3(new_n508), .ZN(new_n509));
  NAND3_X1  g323(.A1(new_n500), .A2(new_n237), .A3(new_n502), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n511));
  OAI221_X1 g325(.A(new_n504), .B1(KEYINPUT15), .B2(new_n507), .C1(new_n510), .C2(new_n511), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n509), .A2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(G113), .B(G122), .ZN(new_n514));
  XNOR2_X1  g328(.A(new_n514), .B(new_n378), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT89), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT90), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n516), .B(KEYINPUT19), .C1(new_n211), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(KEYINPUT89), .B1(new_n214), .B2(KEYINPUT90), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT19), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n520), .B1(new_n214), .B2(KEYINPUT89), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n518), .B(new_n225), .C1(new_n519), .C2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n215), .A2(G146), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n524), .A2(KEYINPUT91), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n331), .A2(new_n233), .A3(G214), .ZN(new_n526));
  OR2_X1    g340(.A1(new_n526), .A2(new_n264), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n264), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n529), .A2(G131), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n288), .A3(new_n528), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n530), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT91), .ZN(new_n533));
  NAND3_X1  g347(.A1(new_n522), .A2(new_n533), .A3(new_n523), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n525), .A2(new_n532), .A3(new_n534), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n529), .A2(KEYINPUT18), .A3(G131), .ZN(new_n536));
  XNOR2_X1  g350(.A(new_n214), .B(new_n225), .ZN(new_n537));
  NAND2_X1  g351(.A1(KEYINPUT18), .A2(G131), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n527), .A2(new_n528), .A3(new_n538), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  AOI21_X1  g354(.A(new_n515), .B1(new_n535), .B2(new_n540), .ZN(new_n541));
  OAI21_X1  g355(.A(KEYINPUT92), .B1(new_n226), .B2(new_n227), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT17), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n530), .A2(new_n543), .A3(new_n531), .ZN(new_n544));
  NAND3_X1  g358(.A1(new_n529), .A2(KEYINPUT17), .A3(G131), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n224), .A2(new_n225), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT92), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n523), .A3(new_n547), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n542), .A2(new_n544), .A3(new_n545), .A4(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n549), .A2(new_n515), .A3(new_n540), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n541), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(G475), .A2(G902), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(KEYINPUT20), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(new_n540), .ZN(new_n556));
  AOI22_X1  g370(.A1(new_n524), .A2(KEYINPUT91), .B1(new_n530), .B2(new_n531), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n556), .B1(new_n557), .B2(new_n534), .ZN(new_n558));
  OAI21_X1  g372(.A(new_n550), .B1(new_n558), .B2(new_n515), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT20), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n559), .A2(new_n560), .A3(new_n553), .ZN(new_n561));
  AOI21_X1  g375(.A(new_n515), .B1(new_n549), .B2(new_n540), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n237), .B1(new_n551), .B2(new_n562), .ZN(new_n563));
  AOI22_X1  g377(.A1(new_n555), .A2(new_n561), .B1(G475), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n233), .A2(G952), .ZN(new_n565));
  AOI21_X1  g379(.A(new_n565), .B1(G234), .B2(G237), .ZN(new_n566));
  AOI211_X1 g380(.A(new_n237), .B(new_n233), .C1(G234), .C2(G237), .ZN(new_n567));
  XNOR2_X1  g381(.A(KEYINPUT21), .B(G898), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n566), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n513), .A2(new_n564), .A3(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(new_n456), .A2(new_n571), .ZN(new_n572));
  OAI21_X1  g386(.A(G214), .B1(G237), .B2(G902), .ZN(new_n573));
  INV_X1    g387(.A(new_n573), .ZN(new_n574));
  AND2_X1   g388(.A1(new_n391), .A2(G101), .ZN(new_n575));
  OAI21_X1  g389(.A(new_n384), .B1(new_n389), .B2(new_n390), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT4), .B1(new_n576), .B2(new_n403), .ZN(new_n577));
  OAI211_X1 g391(.A(new_n326), .B(new_n393), .C1(new_n575), .C2(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n579));
  NOR2_X1   g393(.A1(new_n317), .A2(KEYINPUT5), .ZN(new_n580));
  INV_X1    g394(.A(G113), .ZN(new_n581));
  NOR2_X1   g395(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  AOI22_X1  g396(.A1(new_n579), .A2(new_n582), .B1(new_n321), .B2(new_n323), .ZN(new_n583));
  OAI211_X1 g397(.A(new_n405), .B(new_n583), .C1(new_n429), .C2(new_n430), .ZN(new_n584));
  AOI21_X1  g398(.A(KEYINPUT80), .B1(new_n578), .B2(new_n584), .ZN(new_n585));
  INV_X1    g399(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n578), .A2(KEYINPUT80), .A3(new_n584), .ZN(new_n587));
  XNOR2_X1  g401(.A(G110), .B(G122), .ZN(new_n588));
  XOR2_X1   g402(.A(new_n588), .B(KEYINPUT81), .Z(new_n589));
  INV_X1    g403(.A(new_n589), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n586), .A2(KEYINPUT6), .A3(new_n587), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(KEYINPUT6), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n578), .A2(new_n584), .A3(new_n589), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT82), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n578), .A2(KEYINPUT82), .A3(new_n584), .A4(new_n589), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n592), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  AND3_X1   g411(.A1(new_n578), .A2(KEYINPUT80), .A3(new_n584), .ZN(new_n598));
  NOR3_X1   g412(.A1(new_n598), .A2(new_n585), .A3(new_n589), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n591), .B1(new_n597), .B2(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n294), .A2(G125), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n601), .B1(G125), .B2(new_n304), .ZN(new_n602));
  INV_X1    g416(.A(KEYINPUT83), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(KEYINPUT83), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT84), .B(G224), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT85), .ZN(new_n608));
  OR3_X1    g422(.A1(new_n607), .A2(new_n608), .A3(G953), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n608), .B1(new_n607), .B2(G953), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(new_n611), .B(KEYINPUT86), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n606), .B(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n600), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(new_n583), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n438), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n584), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n589), .B(KEYINPUT8), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT87), .ZN(new_n620));
  OAI21_X1  g434(.A(KEYINPUT7), .B1(new_n611), .B2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n621), .B1(new_n620), .B2(new_n611), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n622), .A2(new_n604), .A3(new_n605), .ZN(new_n623));
  INV_X1    g437(.A(KEYINPUT7), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n602), .B1(new_n624), .B2(new_n611), .ZN(new_n625));
  NAND3_X1  g439(.A1(new_n619), .A2(new_n623), .A3(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n595), .A2(new_n596), .ZN(new_n628));
  AOI21_X1  g442(.A(G902), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n614), .A2(new_n629), .ZN(new_n630));
  OAI21_X1  g444(.A(G210), .B1(G237), .B2(G902), .ZN(new_n631));
  XOR2_X1   g445(.A(new_n631), .B(KEYINPUT88), .Z(new_n632));
  NAND2_X1  g446(.A1(new_n630), .A2(new_n632), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n614), .A2(new_n631), .A3(new_n629), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n574), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n371), .A2(new_n572), .A3(new_n635), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(G101), .ZN(G3));
  OAI21_X1  g451(.A(G472), .B1(new_n354), .B2(G902), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n350), .A2(new_n352), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  NOR3_X1   g454(.A1(new_n456), .A2(new_n640), .A3(new_n262), .ZN(new_n641));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n642));
  AND3_X1   g456(.A1(new_n501), .A2(new_n642), .A3(new_n498), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n498), .B1(new_n501), .B2(new_n642), .ZN(new_n644));
  OAI21_X1  g458(.A(KEYINPUT33), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g459(.A(KEYINPUT33), .ZN(new_n646));
  NAND3_X1  g460(.A1(new_n500), .A2(new_n646), .A3(new_n502), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n507), .A2(G902), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n645), .A2(new_n647), .A3(new_n648), .ZN(new_n649));
  AND3_X1   g463(.A1(new_n510), .A2(KEYINPUT100), .A3(new_n507), .ZN(new_n650));
  AOI21_X1  g464(.A(KEYINPUT100), .B1(new_n510), .B2(new_n507), .ZN(new_n651));
  OAI21_X1  g465(.A(new_n649), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n563), .A2(G475), .ZN(new_n653));
  INV_X1    g467(.A(new_n561), .ZN(new_n654));
  AOI21_X1  g468(.A(new_n560), .B1(new_n559), .B2(new_n553), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n653), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n652), .A2(new_n656), .ZN(new_n657));
  INV_X1    g471(.A(new_n657), .ZN(new_n658));
  INV_X1    g472(.A(new_n631), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n630), .A2(new_n659), .ZN(new_n660));
  AOI211_X1 g474(.A(new_n574), .B(new_n569), .C1(new_n660), .C2(new_n634), .ZN(new_n661));
  NAND3_X1  g475(.A1(new_n641), .A2(new_n658), .A3(new_n661), .ZN(new_n662));
  XOR2_X1   g476(.A(KEYINPUT34), .B(G104), .Z(new_n663));
  XNOR2_X1  g477(.A(new_n662), .B(new_n663), .ZN(G6));
  NOR2_X1   g478(.A1(new_n513), .A2(new_n656), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n641), .A2(new_n661), .A3(new_n665), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(KEYINPUT101), .ZN(new_n667));
  XNOR2_X1  g481(.A(KEYINPUT35), .B(G107), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n667), .B(new_n668), .ZN(G9));
  NAND2_X1  g483(.A1(new_n231), .A2(KEYINPUT102), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n235), .A2(KEYINPUT36), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT102), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n242), .A2(new_n672), .ZN(new_n673));
  AND3_X1   g487(.A1(new_n670), .A2(new_n671), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n671), .B1(new_n670), .B2(new_n673), .ZN(new_n675));
  OAI21_X1  g489(.A(new_n260), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(new_n676), .B1(new_n249), .B2(new_n252), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n677), .A2(KEYINPUT103), .ZN(new_n678));
  INV_X1    g492(.A(KEYINPUT103), .ZN(new_n679));
  OAI211_X1 g493(.A(new_n679), .B(new_n676), .C1(new_n249), .C2(new_n252), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n678), .A2(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n640), .ZN(new_n682));
  NAND4_X1  g496(.A1(new_n681), .A2(new_n572), .A3(new_n635), .A4(new_n682), .ZN(new_n683));
  XOR2_X1   g497(.A(KEYINPUT37), .B(G110), .Z(new_n684));
  XNOR2_X1  g498(.A(new_n683), .B(new_n684), .ZN(G12));
  AOI21_X1  g499(.A(new_n369), .B1(new_n353), .B2(new_n356), .ZN(new_n686));
  AND3_X1   g500(.A1(new_n614), .A2(new_n631), .A3(new_n629), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n631), .B1(new_n614), .B2(new_n629), .ZN(new_n688));
  OAI21_X1  g502(.A(new_n573), .B1(new_n687), .B2(new_n688), .ZN(new_n689));
  NOR3_X1   g503(.A1(new_n686), .A2(new_n689), .A3(new_n456), .ZN(new_n690));
  INV_X1    g504(.A(G900), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n566), .B1(new_n567), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n665), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n694), .B1(new_n678), .B2(new_n680), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n696), .B(G128), .ZN(G30));
  NOR4_X1   g511(.A1(new_n681), .A2(new_n574), .A3(new_n564), .A4(new_n513), .ZN(new_n698));
  XOR2_X1   g512(.A(KEYINPUT105), .B(KEYINPUT39), .Z(new_n699));
  XNOR2_X1  g513(.A(new_n692), .B(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n453), .A2(new_n455), .A3(new_n700), .ZN(new_n701));
  XOR2_X1   g515(.A(new_n701), .B(KEYINPUT40), .Z(new_n702));
  NAND2_X1  g516(.A1(new_n633), .A2(new_n634), .ZN(new_n703));
  XNOR2_X1  g517(.A(KEYINPUT104), .B(KEYINPUT38), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n703), .B(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n336), .ZN(new_n706));
  NAND2_X1  g520(.A1(new_n360), .A2(new_n329), .ZN(new_n707));
  AOI21_X1  g521(.A(new_n706), .B1(new_n348), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g522(.A(G472), .B1(new_n708), .B2(G902), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n357), .A2(new_n709), .ZN(new_n710));
  NAND4_X1  g524(.A1(new_n698), .A2(new_n702), .A3(new_n705), .A4(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G143), .ZN(G45));
  NAND3_X1  g526(.A1(new_n652), .A2(new_n656), .A3(new_n693), .ZN(new_n713));
  AOI21_X1  g527(.A(new_n713), .B1(new_n678), .B2(new_n680), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n690), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G146), .ZN(G48));
  NOR2_X1   g530(.A1(new_n436), .A2(new_n444), .ZN(new_n717));
  OAI21_X1  g531(.A(G469), .B1(new_n717), .B2(G902), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n718), .A2(new_n455), .A3(new_n445), .ZN(new_n719));
  INV_X1    g533(.A(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n371), .A2(new_n661), .A3(new_n658), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(KEYINPUT41), .B(G113), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n721), .B(new_n722), .ZN(G15));
  NAND4_X1  g537(.A1(new_n371), .A2(new_n661), .A3(new_n665), .A4(new_n720), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G116), .ZN(G18));
  NOR2_X1   g539(.A1(new_n689), .A2(new_n719), .ZN(new_n726));
  AOI21_X1  g540(.A(new_n571), .B1(new_n357), .B2(new_n370), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n681), .ZN(new_n728));
  XNOR2_X1  g542(.A(new_n728), .B(G119), .ZN(G21));
  NOR2_X1   g543(.A1(new_n513), .A2(new_n564), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n573), .C1(new_n687), .C2(new_n688), .ZN(new_n731));
  INV_X1    g545(.A(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n258), .ZN(new_n733));
  AOI21_X1  g547(.A(new_n261), .B1(new_n733), .B2(new_n256), .ZN(new_n734));
  INV_X1    g548(.A(new_n251), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n254), .A2(new_n255), .ZN(new_n736));
  AOI21_X1  g550(.A(KEYINPUT25), .B1(new_n736), .B2(new_n237), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT73), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n735), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n247), .A2(KEYINPUT73), .A3(new_n248), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n734), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g555(.A(KEYINPUT106), .B1(new_n361), .B2(new_n342), .ZN(new_n742));
  INV_X1    g556(.A(new_n329), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n328), .B1(new_n296), .B2(new_n307), .ZN(new_n744));
  OAI21_X1  g558(.A(KEYINPUT28), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  INV_X1    g559(.A(KEYINPUT106), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n746), .A3(new_n343), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n742), .A2(new_n747), .A3(new_n348), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(new_n340), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(new_n352), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n741), .A2(new_n638), .A3(new_n750), .ZN(new_n751));
  AND4_X1   g565(.A1(new_n570), .A2(new_n718), .A3(new_n455), .A4(new_n445), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n732), .A2(new_n751), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G122), .ZN(G24));
  XNOR2_X1  g568(.A(new_n713), .B(KEYINPUT107), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n750), .A2(new_n638), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n755), .A2(new_n726), .A3(new_n681), .A4(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G125), .ZN(G27));
  INV_X1    g572(.A(KEYINPUT108), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n456), .A2(new_n759), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n453), .A2(KEYINPUT108), .A3(new_n455), .ZN(new_n761));
  INV_X1    g575(.A(new_n632), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n595), .A2(new_n596), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n237), .B1(new_n763), .B2(new_n626), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n764), .B1(new_n613), .B2(new_n600), .ZN(new_n765));
  OAI211_X1 g579(.A(new_n634), .B(new_n573), .C1(new_n762), .C2(new_n765), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n760), .A2(new_n761), .A3(new_n767), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n768), .A2(KEYINPUT109), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n766), .B1(new_n456), .B2(new_n759), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n770), .A2(new_n771), .A3(new_n761), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n769), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n371), .A2(KEYINPUT110), .ZN(new_n774));
  INV_X1    g588(.A(KEYINPUT110), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n775), .B1(new_n686), .B2(new_n262), .ZN(new_n776));
  AND2_X1   g590(.A1(new_n774), .A2(new_n776), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n773), .A2(new_n755), .A3(new_n777), .ZN(new_n778));
  INV_X1    g592(.A(new_n371), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n779), .B1(new_n769), .B2(new_n772), .ZN(new_n780));
  XOR2_X1   g594(.A(new_n713), .B(KEYINPUT107), .Z(new_n781));
  NOR2_X1   g595(.A1(new_n781), .A2(KEYINPUT42), .ZN(new_n782));
  AOI22_X1  g596(.A1(new_n778), .A2(KEYINPUT42), .B1(new_n780), .B2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  INV_X1    g598(.A(new_n694), .ZN(new_n785));
  INV_X1    g599(.A(new_n761), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT108), .B1(new_n453), .B2(new_n455), .ZN(new_n787));
  NOR4_X1   g601(.A1(new_n786), .A2(new_n787), .A3(KEYINPUT109), .A4(new_n766), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n771), .B1(new_n770), .B2(new_n761), .ZN(new_n789));
  OAI211_X1 g603(.A(new_n371), .B(new_n785), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(G134), .ZN(G36));
  NAND2_X1  g605(.A1(new_n652), .A2(new_n564), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT43), .Z(new_n793));
  NAND3_X1  g607(.A1(new_n793), .A2(new_n640), .A3(new_n681), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT44), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n767), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  AOI21_X1  g610(.A(new_n796), .B1(new_n795), .B2(new_n794), .ZN(new_n797));
  INV_X1    g611(.A(new_n455), .ZN(new_n798));
  OAI21_X1  g612(.A(new_n447), .B1(new_n449), .B2(new_n450), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT45), .ZN(new_n800));
  OR2_X1    g614(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  AOI21_X1  g615(.A(new_n372), .B1(new_n799), .B2(new_n800), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  AOI21_X1  g617(.A(KEYINPUT46), .B1(new_n803), .B2(new_n452), .ZN(new_n804));
  INV_X1    g618(.A(new_n445), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n803), .A2(KEYINPUT46), .A3(new_n452), .ZN(new_n807));
  AOI21_X1  g621(.A(new_n798), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(new_n700), .ZN(new_n809));
  INV_X1    g623(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n797), .A2(new_n810), .ZN(new_n811));
  XNOR2_X1  g625(.A(new_n811), .B(G137), .ZN(G39));
  XNOR2_X1  g626(.A(new_n808), .B(KEYINPUT47), .ZN(new_n813));
  INV_X1    g627(.A(new_n686), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n814), .A2(new_n741), .A3(new_n713), .A4(new_n766), .ZN(new_n815));
  NAND2_X1  g629(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g630(.A(new_n816), .B(G140), .ZN(G42));
  INV_X1    g631(.A(new_n705), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n718), .A2(new_n445), .ZN(new_n819));
  XOR2_X1   g633(.A(new_n819), .B(KEYINPUT49), .Z(new_n820));
  NOR2_X1   g634(.A1(new_n710), .A2(new_n262), .ZN(new_n821));
  NOR3_X1   g635(.A1(new_n792), .A2(new_n574), .A3(new_n798), .ZN(new_n822));
  NAND4_X1  g636(.A1(new_n818), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n793), .A2(new_n566), .A3(new_n751), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n574), .A3(new_n818), .A4(new_n720), .ZN(new_n825));
  XNOR2_X1  g639(.A(new_n825), .B(KEYINPUT50), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n819), .A2(new_n455), .ZN(new_n827));
  OR2_X1    g641(.A1(new_n813), .A2(new_n827), .ZN(new_n828));
  AND2_X1   g642(.A1(new_n824), .A2(new_n767), .ZN(new_n829));
  AOI21_X1  g643(.A(new_n826), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n681), .A2(new_n756), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n720), .A2(new_n566), .A3(new_n767), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(new_n793), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(new_n821), .ZN(new_n834));
  INV_X1    g648(.A(new_n651), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n510), .A2(KEYINPUT100), .A3(new_n507), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n645), .A2(new_n647), .ZN(new_n837));
  AOI22_X1  g651(.A1(new_n835), .A2(new_n836), .B1(new_n837), .B2(new_n648), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n838), .A2(new_n564), .ZN(new_n839));
  OAI22_X1  g653(.A1(new_n831), .A2(new_n833), .B1(new_n834), .B2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT112), .ZN(new_n841));
  OAI21_X1  g655(.A(KEYINPUT51), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  AOI21_X1  g656(.A(new_n842), .B1(new_n841), .B2(new_n840), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n830), .A2(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n777), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n833), .ZN(new_n846));
  XNOR2_X1  g660(.A(new_n846), .B(KEYINPUT48), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n824), .A2(new_n726), .ZN(new_n848));
  XNOR2_X1  g662(.A(new_n565), .B(KEYINPUT113), .ZN(new_n849));
  OAI211_X1 g663(.A(new_n848), .B(new_n849), .C1(new_n834), .C2(new_n657), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n847), .A2(new_n850), .ZN(new_n851));
  AOI211_X1 g665(.A(new_n840), .B(new_n826), .C1(new_n828), .C2(new_n829), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n844), .B(new_n851), .C1(new_n852), .C2(KEYINPUT51), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT54), .ZN(new_n854));
  NOR2_X1   g668(.A1(new_n831), .A2(new_n781), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n788), .B2(new_n789), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n686), .A2(new_n456), .ZN(new_n857));
  AND3_X1   g671(.A1(new_n513), .A2(new_n564), .A3(new_n693), .ZN(new_n858));
  NAND4_X1  g672(.A1(new_n857), .A2(new_n681), .A3(new_n767), .A4(new_n858), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n790), .A2(new_n856), .A3(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n860), .A2(KEYINPUT111), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n456), .A2(new_n262), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n564), .A2(new_n512), .A3(new_n509), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n569), .B1(new_n863), .B2(new_n657), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n862), .A2(new_n635), .A3(new_n682), .A4(new_n864), .ZN(new_n865));
  NAND4_X1  g679(.A1(new_n683), .A2(new_n865), .A3(new_n636), .A4(new_n753), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n721), .A2(new_n724), .A3(new_n728), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n861), .A2(new_n783), .A3(new_n868), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n690), .B1(new_n695), .B2(new_n714), .ZN(new_n870));
  NOR3_X1   g684(.A1(new_n456), .A2(new_n677), .A3(new_n692), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n871), .A2(new_n710), .A3(new_n732), .ZN(new_n872));
  NAND3_X1  g686(.A1(new_n870), .A2(new_n757), .A3(new_n872), .ZN(new_n873));
  INV_X1    g687(.A(KEYINPUT52), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n870), .A2(KEYINPUT52), .A3(new_n757), .A4(new_n872), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g691(.A(KEYINPUT111), .ZN(new_n878));
  NAND4_X1  g692(.A1(new_n790), .A2(new_n856), .A3(new_n878), .A4(new_n859), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n877), .A2(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NOR3_X1   g695(.A1(new_n869), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(new_n859), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n883), .B1(new_n773), .B2(new_n855), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n878), .B1(new_n884), .B2(new_n790), .ZN(new_n885));
  NOR2_X1   g699(.A1(new_n788), .A2(new_n789), .ZN(new_n886));
  NAND3_X1  g700(.A1(new_n774), .A2(new_n755), .A3(new_n776), .ZN(new_n887));
  OAI21_X1  g701(.A(KEYINPUT42), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n780), .A2(new_n782), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(new_n889), .A3(new_n868), .ZN(new_n890));
  NOR2_X1   g704(.A1(new_n885), .A2(new_n890), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n877), .A2(new_n879), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT53), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n854), .B1(new_n882), .B2(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n881), .B1(new_n869), .B2(new_n880), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n891), .A2(KEYINPUT53), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n896), .A3(KEYINPUT54), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n853), .B1(new_n894), .B2(new_n897), .ZN(new_n898));
  NOR2_X1   g712(.A1(G952), .A2(G953), .ZN(new_n899));
  OAI21_X1  g713(.A(new_n823), .B1(new_n898), .B2(new_n899), .ZN(G75));
  NOR2_X1   g714(.A1(new_n233), .A2(G952), .ZN(new_n901));
  INV_X1    g715(.A(new_n901), .ZN(new_n902));
  AOI21_X1  g716(.A(new_n237), .B1(new_n895), .B2(new_n896), .ZN(new_n903));
  AOI21_X1  g717(.A(KEYINPUT56), .B1(new_n903), .B2(G210), .ZN(new_n904));
  INV_X1    g718(.A(new_n600), .ZN(new_n905));
  OR2_X1    g719(.A1(new_n905), .A2(KEYINPUT114), .ZN(new_n906));
  NAND2_X1  g720(.A1(new_n905), .A2(KEYINPUT114), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT55), .Z(new_n909));
  XNOR2_X1  g723(.A(new_n909), .B(new_n613), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n902), .B1(new_n904), .B2(new_n910), .ZN(new_n911));
  AND2_X1   g725(.A1(new_n903), .A2(new_n632), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT115), .ZN(new_n913));
  INV_X1    g727(.A(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n910), .A2(new_n914), .ZN(new_n915));
  OR3_X1    g729(.A1(new_n912), .A2(new_n913), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n913), .B1(new_n912), .B2(new_n915), .ZN(new_n917));
  AOI21_X1  g731(.A(new_n911), .B1(new_n916), .B2(new_n917), .ZN(G51));
  XOR2_X1   g732(.A(new_n452), .B(KEYINPUT57), .Z(new_n919));
  NAND3_X1  g733(.A1(new_n894), .A2(new_n897), .A3(new_n919), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT116), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  INV_X1    g736(.A(new_n717), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n894), .A2(KEYINPUT116), .A3(new_n897), .A4(new_n919), .ZN(new_n924));
  NAND3_X1  g738(.A1(new_n922), .A2(new_n923), .A3(new_n924), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n903), .A2(new_n801), .A3(new_n802), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n901), .B1(new_n925), .B2(new_n926), .ZN(G54));
  NAND3_X1  g741(.A1(new_n903), .A2(KEYINPUT58), .A3(G475), .ZN(new_n928));
  AND2_X1   g742(.A1(new_n928), .A2(new_n552), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n552), .ZN(new_n930));
  NOR3_X1   g744(.A1(new_n929), .A2(new_n930), .A3(new_n901), .ZN(G60));
  AND3_X1   g745(.A1(new_n895), .A2(KEYINPUT54), .A3(new_n896), .ZN(new_n932));
  AOI21_X1  g746(.A(KEYINPUT54), .B1(new_n895), .B2(new_n896), .ZN(new_n933));
  NAND2_X1  g747(.A1(G478), .A2(G902), .ZN(new_n934));
  XOR2_X1   g748(.A(new_n934), .B(KEYINPUT59), .Z(new_n935));
  NOR3_X1   g749(.A1(new_n932), .A2(new_n933), .A3(new_n935), .ZN(new_n936));
  OAI21_X1  g750(.A(new_n902), .B1(new_n936), .B2(new_n837), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n894), .A2(new_n837), .A3(new_n897), .A4(new_n938), .ZN(new_n939));
  OR2_X1    g753(.A1(new_n939), .A2(KEYINPUT117), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n939), .A2(KEYINPUT117), .ZN(new_n941));
  AOI21_X1  g755(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G63));
  NAND2_X1  g756(.A1(G217), .A2(G902), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(KEYINPUT60), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n944), .B1(new_n895), .B2(new_n896), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n674), .A2(new_n675), .ZN(new_n946));
  XNOR2_X1  g760(.A(new_n946), .B(KEYINPUT118), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n945), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n259), .ZN(new_n949));
  OAI21_X1  g763(.A(new_n902), .B1(new_n945), .B2(new_n949), .ZN(new_n950));
  NOR2_X1   g764(.A1(new_n948), .A2(new_n950), .ZN(new_n951));
  OAI211_X1 g765(.A(KEYINPUT119), .B(new_n902), .C1(new_n945), .C2(new_n949), .ZN(new_n952));
  INV_X1    g766(.A(new_n952), .ZN(new_n953));
  OAI21_X1  g767(.A(new_n951), .B1(KEYINPUT61), .B2(new_n953), .ZN(new_n954));
  INV_X1    g768(.A(KEYINPUT61), .ZN(new_n955));
  OAI211_X1 g769(.A(new_n955), .B(new_n952), .C1(new_n948), .C2(new_n950), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n954), .A2(new_n956), .ZN(G66));
  OAI21_X1  g771(.A(G953), .B1(new_n607), .B2(new_n568), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n958), .B1(new_n868), .B2(G953), .ZN(new_n959));
  OAI211_X1 g773(.A(new_n906), .B(new_n907), .C1(G898), .C2(new_n233), .ZN(new_n960));
  XNOR2_X1  g774(.A(new_n960), .B(KEYINPUT120), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n959), .B(new_n961), .ZN(G69));
  NAND2_X1  g776(.A1(new_n308), .A2(new_n316), .ZN(new_n963));
  OAI21_X1  g777(.A(new_n518), .B1(new_n519), .B2(new_n521), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n964), .B(KEYINPUT121), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n963), .B(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n691), .B1(new_n966), .B2(new_n374), .ZN(new_n967));
  OAI21_X1  g781(.A(new_n967), .B1(new_n374), .B2(new_n966), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n968), .A2(G953), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n783), .A2(new_n790), .ZN(new_n970));
  INV_X1    g784(.A(KEYINPUT123), .ZN(new_n971));
  XNOR2_X1  g785(.A(new_n970), .B(new_n971), .ZN(new_n972));
  AOI22_X1  g786(.A1(new_n813), .A2(new_n815), .B1(new_n797), .B2(new_n810), .ZN(new_n973));
  NAND3_X1  g787(.A1(new_n810), .A2(new_n732), .A3(new_n777), .ZN(new_n974));
  NAND4_X1  g788(.A1(new_n973), .A2(new_n757), .A3(new_n870), .A4(new_n974), .ZN(new_n975));
  NOR2_X1   g789(.A1(new_n972), .A2(new_n975), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n233), .B1(new_n976), .B2(new_n966), .ZN(new_n977));
  NOR2_X1   g791(.A1(new_n658), .A2(new_n665), .ZN(new_n978));
  NOR4_X1   g792(.A1(new_n779), .A2(new_n701), .A3(new_n766), .A4(new_n978), .ZN(new_n979));
  AND3_X1   g793(.A1(new_n711), .A2(new_n757), .A3(new_n870), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT62), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n979), .B1(new_n980), .B2(new_n981), .ZN(new_n982));
  NAND3_X1  g796(.A1(new_n711), .A2(new_n757), .A3(new_n870), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n983), .A2(KEYINPUT62), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n973), .A2(new_n982), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT122), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  NAND4_X1  g801(.A1(new_n973), .A2(new_n982), .A3(KEYINPUT122), .A4(new_n984), .ZN(new_n988));
  AND3_X1   g802(.A1(new_n987), .A2(new_n966), .A3(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n969), .B1(new_n977), .B2(new_n989), .ZN(G72));
  XNOR2_X1  g804(.A(new_n366), .B(KEYINPUT125), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n991), .A2(new_n335), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n987), .A2(new_n868), .A3(new_n988), .ZN(new_n993));
  NAND2_X1  g807(.A1(G472), .A2(G902), .ZN(new_n994));
  XOR2_X1   g808(.A(new_n994), .B(KEYINPUT63), .Z(new_n995));
  NAND2_X1  g809(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n996), .A2(KEYINPUT124), .ZN(new_n997));
  INV_X1    g811(.A(KEYINPUT124), .ZN(new_n998));
  NAND3_X1  g812(.A1(new_n993), .A2(new_n998), .A3(new_n995), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n992), .B1(new_n997), .B2(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n895), .A2(new_n896), .ZN(new_n1001));
  INV_X1    g815(.A(new_n995), .ZN(new_n1002));
  AOI21_X1  g816(.A(new_n1002), .B1(new_n367), .B2(new_n336), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT126), .Z(new_n1004));
  AOI21_X1  g818(.A(new_n901), .B1(new_n1001), .B2(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n976), .B2(new_n868), .ZN(new_n1006));
  OR2_X1    g820(.A1(new_n991), .A2(new_n335), .ZN(new_n1007));
  OAI21_X1  g821(.A(new_n1005), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g822(.A1(new_n1000), .A2(new_n1008), .ZN(G57));
endmodule


