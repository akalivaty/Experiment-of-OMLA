//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 1 1 0 0 0 1 0 1 1 0 0 1 1 1 0 1 1 1 0 0 0 1 1 0 1 1 1 1 1 1 0 1 0 1 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:30 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n721, new_n722, new_n724, new_n725, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n738, new_n739, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n902, new_n903,
    new_n904, new_n905, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n949, new_n950, new_n951, new_n952, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n994,
    new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  AND2_X1   g001(.A1(new_n187), .A2(KEYINPUT32), .ZN(new_n188));
  XNOR2_X1  g002(.A(KEYINPUT26), .B(G101), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT69), .B(KEYINPUT27), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  NOR2_X1   g005(.A1(G237), .A2(G953), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G210), .ZN(new_n193));
  XNOR2_X1  g007(.A(new_n193), .B(KEYINPUT70), .ZN(new_n194));
  XNOR2_X1  g008(.A(new_n191), .B(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G143), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n196), .A2(G146), .ZN(new_n197));
  INV_X1    g011(.A(G146), .ZN(new_n198));
  OAI21_X1  g012(.A(KEYINPUT64), .B1(new_n198), .B2(G143), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT64), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n200), .A2(new_n196), .A3(G146), .ZN(new_n201));
  AOI21_X1  g015(.A(new_n197), .B1(new_n199), .B2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(KEYINPUT0), .A2(G128), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  OR2_X1    g018(.A1(KEYINPUT0), .A2(G128), .ZN(new_n205));
  AND2_X1   g019(.A1(new_n205), .A2(new_n203), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n198), .A2(G143), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n196), .A2(G146), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g023(.A1(new_n202), .A2(new_n204), .B1(new_n206), .B2(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G131), .ZN(new_n211));
  INV_X1    g025(.A(G137), .ZN(new_n212));
  OAI21_X1  g026(.A(KEYINPUT66), .B1(new_n212), .B2(G134), .ZN(new_n213));
  INV_X1    g027(.A(KEYINPUT66), .ZN(new_n214));
  INV_X1    g028(.A(G134), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n214), .A2(new_n215), .A3(G137), .ZN(new_n216));
  INV_X1    g030(.A(KEYINPUT65), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n217), .B1(new_n215), .B2(G137), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n213), .A2(new_n216), .B1(new_n218), .B2(KEYINPUT11), .ZN(new_n219));
  INV_X1    g033(.A(KEYINPUT11), .ZN(new_n220));
  OAI211_X1 g034(.A(new_n217), .B(new_n220), .C1(new_n215), .C2(G137), .ZN(new_n221));
  AOI21_X1  g035(.A(new_n211), .B1(new_n219), .B2(new_n221), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n213), .A2(new_n216), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n218), .A2(KEYINPUT11), .ZN(new_n224));
  AND4_X1   g038(.A1(new_n211), .A2(new_n223), .A3(new_n224), .A4(new_n221), .ZN(new_n225));
  OAI21_X1  g039(.A(new_n210), .B1(new_n222), .B2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT67), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n226), .A2(new_n227), .ZN(new_n228));
  NAND4_X1  g042(.A1(new_n223), .A2(new_n224), .A3(new_n211), .A4(new_n221), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n215), .A2(G137), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n212), .A2(G134), .ZN(new_n231));
  OAI21_X1  g045(.A(G131), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  AND2_X1   g046(.A1(new_n229), .A2(new_n232), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT1), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G128), .ZN(new_n235));
  INV_X1    g049(.A(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n200), .B1(new_n196), .B2(G146), .ZN(new_n237));
  NOR3_X1   g051(.A1(new_n198), .A2(KEYINPUT64), .A3(G143), .ZN(new_n238));
  OAI211_X1 g052(.A(new_n207), .B(new_n236), .C1(new_n237), .C2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT1), .B1(new_n196), .B2(G146), .ZN(new_n240));
  NAND2_X1  g054(.A1(new_n240), .A2(G128), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(new_n209), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n239), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G119), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G116), .ZN(new_n245));
  INV_X1    g059(.A(G116), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G119), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT2), .ZN(new_n248));
  NOR2_X1   g062(.A1(new_n248), .A2(G113), .ZN(new_n249));
  INV_X1    g063(.A(G113), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n250), .A2(KEYINPUT2), .ZN(new_n251));
  OAI211_X1 g065(.A(new_n245), .B(new_n247), .C1(new_n249), .C2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n245), .A2(new_n247), .ZN(new_n253));
  XNOR2_X1  g067(.A(KEYINPUT2), .B(G113), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n252), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(KEYINPUT68), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  NAND3_X1  g072(.A1(new_n252), .A2(new_n255), .A3(KEYINPUT68), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n233), .A2(new_n243), .B1(new_n258), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n223), .A2(new_n224), .A3(new_n221), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n261), .A2(G131), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n229), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n263), .A2(KEYINPUT67), .A3(new_n210), .ZN(new_n264));
  NAND3_X1  g078(.A1(new_n228), .A2(new_n260), .A3(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n206), .A2(new_n209), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n207), .B(new_n204), .C1(new_n237), .C2(new_n238), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  AOI21_X1  g082(.A(new_n268), .B1(new_n262), .B2(new_n229), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n229), .A2(new_n232), .ZN(new_n270));
  AOI22_X1  g084(.A1(new_n202), .A2(new_n236), .B1(new_n241), .B2(new_n209), .ZN(new_n271));
  NOR2_X1   g085(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  OAI21_X1  g086(.A(new_n256), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  INV_X1    g089(.A(KEYINPUT73), .ZN(new_n276));
  OAI21_X1  g090(.A(new_n276), .B1(new_n269), .B2(new_n272), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n258), .A2(new_n259), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n243), .A2(new_n229), .A3(new_n232), .ZN(new_n279));
  NAND3_X1  g093(.A1(new_n226), .A2(KEYINPUT73), .A3(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT28), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n281), .A2(new_n282), .ZN(new_n283));
  AOI21_X1  g097(.A(new_n195), .B1(new_n275), .B2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT30), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n233), .B2(new_n243), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n228), .A2(new_n264), .A3(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n285), .B1(new_n269), .B2(new_n272), .ZN(new_n288));
  NAND3_X1  g102(.A1(new_n287), .A2(new_n256), .A3(new_n288), .ZN(new_n289));
  XOR2_X1   g103(.A(KEYINPUT72), .B(KEYINPUT31), .Z(new_n290));
  AND4_X1   g104(.A1(new_n289), .A2(new_n265), .A3(new_n195), .A4(new_n290), .ZN(new_n291));
  NOR2_X1   g105(.A1(new_n284), .A2(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(KEYINPUT71), .ZN(new_n293));
  AND3_X1   g107(.A1(new_n228), .A2(new_n264), .A3(new_n286), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n288), .A2(new_n256), .ZN(new_n295));
  NOR2_X1   g109(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g110(.A1(new_n265), .A2(new_n195), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n293), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n297), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n299), .A2(KEYINPUT71), .A3(new_n289), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n301));
  AND3_X1   g115(.A1(new_n292), .A2(KEYINPUT74), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g116(.A(KEYINPUT74), .B1(new_n292), .B2(new_n301), .ZN(new_n303));
  OAI21_X1  g117(.A(new_n188), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND3_X1   g118(.A1(new_n228), .A2(new_n264), .A3(new_n279), .ZN(new_n305));
  OAI21_X1  g119(.A(new_n265), .B1(new_n305), .B2(new_n278), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(KEYINPUT28), .ZN(new_n307));
  INV_X1    g121(.A(new_n195), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n309));
  NOR2_X1   g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n307), .A2(new_n283), .A3(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n312));
  INV_X1    g126(.A(G902), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n275), .A2(new_n195), .A3(new_n283), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n289), .A2(new_n265), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(new_n308), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n314), .A2(new_n316), .A3(new_n309), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n312), .A2(new_n313), .A3(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n311), .A2(KEYINPUT75), .ZN(new_n319));
  OAI21_X1  g133(.A(G472), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(new_n187), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT74), .ZN(new_n322));
  AND3_X1   g136(.A1(new_n298), .A2(KEYINPUT31), .A3(new_n300), .ZN(new_n323));
  INV_X1    g137(.A(new_n283), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n282), .B1(new_n265), .B2(new_n273), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n308), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n299), .A2(new_n289), .A3(new_n290), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(new_n322), .B1(new_n323), .B2(new_n328), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n292), .A2(new_n301), .A3(KEYINPUT74), .ZN(new_n330));
  AOI21_X1  g144(.A(new_n321), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n304), .B(new_n320), .C1(new_n331), .C2(KEYINPUT32), .ZN(new_n332));
  AOI21_X1  g146(.A(G125), .B1(new_n241), .B2(new_n209), .ZN(new_n333));
  AND3_X1   g147(.A1(new_n333), .A2(KEYINPUT84), .A3(new_n239), .ZN(new_n334));
  AOI21_X1  g148(.A(KEYINPUT84), .B1(new_n333), .B2(new_n239), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  AOI21_X1  g150(.A(new_n336), .B1(new_n266), .B2(new_n267), .ZN(new_n337));
  NOR3_X1   g151(.A1(new_n334), .A2(new_n335), .A3(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G953), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G224), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(KEYINPUT7), .ZN(new_n341));
  INV_X1    g155(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(KEYINPUT85), .B1(new_n338), .B2(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(KEYINPUT79), .ZN(new_n344));
  INV_X1    g158(.A(G107), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(KEYINPUT79), .A2(G107), .ZN(new_n347));
  AOI21_X1  g161(.A(G104), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G104), .ZN(new_n349));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n349), .B2(G107), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT80), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n345), .A3(G104), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  OAI21_X1  g167(.A(G101), .B1(new_n348), .B2(new_n353), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n349), .A2(KEYINPUT3), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n355), .A2(new_n346), .A3(new_n347), .ZN(new_n356));
  OAI21_X1  g170(.A(KEYINPUT3), .B1(new_n349), .B2(G107), .ZN(new_n357));
  AOI21_X1  g171(.A(G101), .B1(new_n349), .B2(G107), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n354), .A2(new_n359), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n245), .A2(new_n247), .A3(KEYINPUT5), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n361), .B(G113), .C1(KEYINPUT5), .C2(new_n245), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n362), .A2(new_n252), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n354), .A2(new_n362), .A3(new_n252), .A4(new_n359), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G122), .ZN(new_n367));
  XNOR2_X1  g181(.A(new_n367), .B(KEYINPUT8), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n268), .A2(G125), .B1(new_n239), .B2(new_n333), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n366), .A2(new_n368), .B1(new_n369), .B2(new_n342), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT85), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n333), .A2(new_n239), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT84), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n268), .A2(G125), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OAI211_X1 g190(.A(new_n371), .B(new_n341), .C1(new_n376), .C2(new_n334), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n349), .A2(G107), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n356), .A2(new_n357), .A3(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT4), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n379), .A2(new_n380), .A3(G101), .ZN(new_n381));
  INV_X1    g195(.A(G101), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT3), .ZN(new_n383));
  AOI21_X1  g197(.A(new_n383), .B1(G104), .B2(new_n345), .ZN(new_n384));
  AND2_X1   g198(.A1(KEYINPUT79), .A2(G107), .ZN(new_n385));
  NOR2_X1   g199(.A1(KEYINPUT79), .A2(G107), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  AOI21_X1  g201(.A(new_n384), .B1(new_n387), .B2(new_n355), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n382), .B1(new_n388), .B2(new_n378), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n359), .A2(KEYINPUT4), .ZN(new_n390));
  OAI211_X1 g204(.A(new_n256), .B(new_n381), .C1(new_n389), .C2(new_n390), .ZN(new_n391));
  NAND3_X1  g205(.A1(new_n391), .A2(new_n367), .A3(new_n365), .ZN(new_n392));
  NAND4_X1  g206(.A1(new_n343), .A2(new_n370), .A3(new_n377), .A4(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n393), .A2(new_n313), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n394), .A2(KEYINPUT86), .ZN(new_n395));
  OAI21_X1  g209(.A(G210), .B1(G237), .B2(G902), .ZN(new_n396));
  INV_X1    g210(.A(KEYINPUT86), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n393), .A2(new_n397), .A3(new_n313), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n391), .A2(new_n365), .ZN(new_n399));
  INV_X1    g213(.A(new_n367), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n401), .A2(KEYINPUT6), .A3(new_n392), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n399), .A2(new_n403), .A3(new_n400), .ZN(new_n404));
  XNOR2_X1  g218(.A(new_n369), .B(new_n340), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n402), .A2(new_n404), .A3(new_n405), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n395), .A2(new_n396), .A3(new_n398), .A4(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(new_n407), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n395), .A2(new_n398), .A3(new_n406), .ZN(new_n409));
  INV_X1    g223(.A(KEYINPUT87), .ZN(new_n410));
  AOI21_X1  g224(.A(new_n396), .B1(new_n409), .B2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n395), .A2(KEYINPUT87), .A3(new_n398), .A4(new_n406), .ZN(new_n412));
  AOI21_X1  g226(.A(new_n408), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G469), .ZN(new_n414));
  INV_X1    g228(.A(G128), .ZN(new_n415));
  AOI21_X1  g229(.A(new_n234), .B1(G143), .B2(new_n198), .ZN(new_n416));
  INV_X1    g230(.A(KEYINPUT81), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n415), .B1(new_n416), .B2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n240), .A2(KEYINPUT81), .ZN(new_n419));
  AOI21_X1  g233(.A(new_n202), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(new_n235), .B(new_n197), .C1(new_n199), .C2(new_n201), .ZN(new_n421));
  OAI211_X1 g235(.A(new_n359), .B(new_n354), .C1(new_n420), .C2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT10), .ZN(new_n423));
  NAND4_X1  g237(.A1(new_n243), .A2(KEYINPUT10), .A3(new_n359), .A4(new_n354), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT82), .ZN(new_n425));
  AOI22_X1  g239(.A1(new_n422), .A2(new_n423), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n263), .ZN(new_n427));
  OAI21_X1  g241(.A(new_n349), .B1(new_n385), .B2(new_n386), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n428), .A2(new_n350), .A3(new_n352), .ZN(new_n429));
  AOI22_X1  g243(.A1(new_n429), .A2(G101), .B1(new_n388), .B2(new_n358), .ZN(new_n430));
  NAND4_X1  g244(.A1(new_n430), .A2(KEYINPUT82), .A3(KEYINPUT10), .A4(new_n243), .ZN(new_n431));
  OAI211_X1 g245(.A(new_n210), .B(new_n381), .C1(new_n389), .C2(new_n390), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n426), .A2(new_n427), .A3(new_n431), .A4(new_n432), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G140), .ZN(new_n434));
  AND2_X1   g248(.A1(new_n339), .A2(G227), .ZN(new_n435));
  XNOR2_X1  g249(.A(new_n434), .B(new_n435), .ZN(new_n436));
  INV_X1    g250(.A(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n433), .A2(new_n437), .ZN(new_n438));
  AND2_X1   g252(.A1(new_n350), .A2(new_n352), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n382), .B1(new_n439), .B2(new_n428), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n356), .A2(new_n357), .A3(new_n358), .ZN(new_n441));
  OAI21_X1  g255(.A(new_n271), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT83), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n360), .A2(KEYINPUT83), .A3(new_n271), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n422), .A3(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(KEYINPUT12), .A3(new_n263), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n263), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT12), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n438), .B1(new_n447), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n202), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n418), .A2(new_n419), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n421), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  OAI21_X1  g268(.A(new_n423), .B1(new_n454), .B2(new_n360), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n424), .A2(new_n425), .ZN(new_n456));
  NAND4_X1  g270(.A1(new_n455), .A2(new_n456), .A3(new_n431), .A4(new_n432), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(new_n263), .ZN(new_n458));
  AOI21_X1  g272(.A(new_n437), .B1(new_n458), .B2(new_n433), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n414), .B(new_n313), .C1(new_n451), .C2(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(new_n457), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n436), .B1(new_n461), .B2(new_n427), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(new_n458), .ZN(new_n463));
  AOI22_X1  g277(.A1(new_n450), .A2(new_n447), .B1(new_n427), .B2(new_n461), .ZN(new_n464));
  XNOR2_X1  g278(.A(new_n436), .B(KEYINPUT78), .ZN(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  OAI211_X1 g280(.A(new_n463), .B(G469), .C1(new_n464), .C2(new_n466), .ZN(new_n467));
  NOR2_X1   g281(.A1(new_n414), .A2(new_n313), .ZN(new_n468));
  INV_X1    g282(.A(new_n468), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n460), .A2(new_n467), .A3(new_n469), .ZN(new_n470));
  XNOR2_X1  g284(.A(KEYINPUT9), .B(G234), .ZN(new_n471));
  OAI21_X1  g285(.A(G221), .B1(new_n471), .B2(G902), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  OAI21_X1  g287(.A(G214), .B1(G237), .B2(G902), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NOR2_X1   g289(.A1(new_n473), .A2(new_n475), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(KEYINPUT90), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n336), .A2(KEYINPUT16), .A3(G140), .ZN(new_n479));
  XNOR2_X1  g293(.A(G125), .B(G140), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n480), .B2(KEYINPUT16), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n481), .A2(G146), .ZN(new_n482));
  INV_X1    g296(.A(G140), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n483), .A2(G125), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n336), .A2(G140), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT19), .ZN(new_n486));
  AOI21_X1  g300(.A(KEYINPUT19), .B1(new_n484), .B2(new_n485), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n198), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n192), .A2(G143), .A3(G214), .ZN(new_n489));
  INV_X1    g303(.A(new_n489), .ZN(new_n490));
  AOI21_X1  g304(.A(G143), .B1(new_n192), .B2(G214), .ZN(new_n491));
  NOR3_X1   g305(.A1(new_n490), .A2(new_n491), .A3(G131), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n192), .A2(G214), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(new_n196), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n211), .B1(new_n494), .B2(new_n489), .ZN(new_n495));
  OAI211_X1 g309(.A(new_n482), .B(new_n488), .C1(new_n492), .C2(new_n495), .ZN(new_n496));
  OAI211_X1 g310(.A(KEYINPUT18), .B(G131), .C1(new_n490), .C2(new_n491), .ZN(new_n497));
  NAND2_X1  g311(.A1(KEYINPUT18), .A2(G131), .ZN(new_n498));
  NAND3_X1  g312(.A1(new_n494), .A2(new_n489), .A3(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n480), .A2(new_n198), .ZN(new_n500));
  NOR2_X1   g314(.A1(new_n480), .A2(new_n198), .ZN(new_n501));
  OAI211_X1 g315(.A(new_n497), .B(new_n499), .C1(new_n500), .C2(new_n501), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n496), .A2(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(G113), .B(G122), .ZN(new_n504));
  XNOR2_X1  g318(.A(new_n504), .B(new_n349), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n503), .A2(new_n506), .ZN(new_n507));
  NOR3_X1   g321(.A1(new_n492), .A2(new_n495), .A3(KEYINPUT17), .ZN(new_n508));
  OAI211_X1 g322(.A(KEYINPUT17), .B(G131), .C1(new_n490), .C2(new_n491), .ZN(new_n509));
  AND3_X1   g323(.A1(new_n484), .A2(new_n485), .A3(KEYINPUT16), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n198), .B1(new_n510), .B2(new_n479), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n482), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  OAI211_X1 g326(.A(new_n505), .B(new_n502), .C1(new_n508), .C2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n507), .A2(new_n513), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT88), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  NOR2_X1   g330(.A1(G475), .A2(G902), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n507), .A2(new_n513), .A3(KEYINPUT88), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n516), .A2(new_n517), .A3(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n517), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n520), .A2(KEYINPUT20), .ZN(new_n521));
  AOI22_X1  g335(.A1(new_n519), .A2(KEYINPUT20), .B1(new_n514), .B2(new_n521), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n502), .B1(new_n508), .B2(new_n512), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n506), .ZN(new_n524));
  AOI21_X1  g338(.A(G902), .B1(new_n524), .B2(new_n513), .ZN(new_n525));
  XNOR2_X1  g339(.A(KEYINPUT89), .B(G475), .ZN(new_n526));
  NOR2_X1   g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  OAI21_X1  g341(.A(new_n478), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n514), .A2(new_n521), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n507), .A2(new_n513), .A3(KEYINPUT88), .ZN(new_n530));
  AOI21_X1  g344(.A(KEYINPUT88), .B1(new_n507), .B2(new_n513), .ZN(new_n531));
  NOR3_X1   g345(.A1(new_n530), .A2(new_n531), .A3(new_n520), .ZN(new_n532));
  INV_X1    g346(.A(KEYINPUT20), .ZN(new_n533));
  OAI21_X1  g347(.A(new_n529), .B1(new_n532), .B2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n527), .ZN(new_n535));
  NAND3_X1  g349(.A1(new_n534), .A2(KEYINPUT90), .A3(new_n535), .ZN(new_n536));
  NOR2_X1   g350(.A1(KEYINPUT93), .A2(G952), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(KEYINPUT93), .A2(G952), .ZN(new_n539));
  AOI21_X1  g353(.A(G953), .B1(new_n538), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(G234), .A2(G237), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g356(.A(KEYINPUT21), .B(G898), .ZN(new_n543));
  NAND4_X1  g357(.A1(new_n543), .A2(G902), .A3(G953), .A4(new_n541), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT91), .ZN(new_n546));
  INV_X1    g360(.A(G122), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n547), .A2(G116), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n246), .A2(G122), .ZN(new_n549));
  AOI21_X1  g363(.A(new_n546), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n550), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n549), .A3(new_n546), .ZN(new_n552));
  OAI211_X1 g366(.A(new_n551), .B(new_n552), .C1(new_n386), .C2(new_n385), .ZN(new_n553));
  INV_X1    g367(.A(new_n552), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n387), .B1(new_n554), .B2(new_n550), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n196), .A2(G128), .ZN(new_n557));
  INV_X1    g371(.A(new_n557), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n196), .A2(G128), .ZN(new_n559));
  NOR3_X1   g373(.A1(new_n558), .A2(new_n559), .A3(G134), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n558), .A2(KEYINPUT92), .A3(KEYINPUT13), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT13), .ZN(new_n562));
  OAI21_X1  g376(.A(new_n557), .B1(new_n559), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT92), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n564), .B1(new_n557), .B2(new_n562), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n561), .A2(new_n563), .A3(new_n565), .ZN(new_n566));
  AOI21_X1  g380(.A(new_n560), .B1(new_n566), .B2(G134), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n556), .A2(new_n567), .ZN(new_n568));
  NOR2_X1   g382(.A1(new_n558), .A2(new_n559), .ZN(new_n569));
  NOR2_X1   g383(.A1(new_n569), .A2(new_n215), .ZN(new_n570));
  OR2_X1    g384(.A1(new_n549), .A2(KEYINPUT14), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n549), .A2(KEYINPUT14), .ZN(new_n572));
  AND3_X1   g386(.A1(new_n571), .A2(new_n548), .A3(new_n572), .ZN(new_n573));
  OAI221_X1 g387(.A(new_n555), .B1(new_n570), .B2(new_n560), .C1(new_n573), .C2(new_n345), .ZN(new_n574));
  INV_X1    g388(.A(G217), .ZN(new_n575));
  NOR3_X1   g389(.A1(new_n471), .A2(new_n575), .A3(G953), .ZN(new_n576));
  AND3_X1   g390(.A1(new_n568), .A2(new_n574), .A3(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n576), .B1(new_n568), .B2(new_n574), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n313), .B1(new_n577), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(G478), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n580), .A2(KEYINPUT15), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  OAI221_X1 g396(.A(new_n313), .B1(KEYINPUT15), .B2(new_n580), .C1(new_n577), .C2(new_n578), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n582), .A2(new_n583), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  NAND4_X1  g399(.A1(new_n528), .A2(new_n536), .A3(new_n545), .A4(new_n585), .ZN(new_n586));
  NOR3_X1   g400(.A1(new_n413), .A2(new_n477), .A3(new_n586), .ZN(new_n587));
  AOI21_X1  g401(.A(new_n575), .B1(G234), .B2(new_n313), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n482), .A2(new_n511), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n244), .A2(G128), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n415), .A2(KEYINPUT23), .A3(G119), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n415), .A2(G119), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  OAI211_X1 g408(.A(new_n591), .B(new_n592), .C1(new_n594), .C2(KEYINPUT23), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(G110), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n593), .A2(new_n591), .ZN(new_n597));
  XNOR2_X1  g411(.A(KEYINPUT24), .B(G110), .ZN(new_n598));
  OAI211_X1 g412(.A(new_n590), .B(new_n596), .C1(new_n597), .C2(new_n598), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n500), .B1(new_n481), .B2(G146), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT76), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n597), .A2(new_n598), .ZN(new_n602));
  OAI21_X1  g416(.A(new_n602), .B1(new_n595), .B2(G110), .ZN(new_n603));
  AND3_X1   g417(.A1(new_n600), .A2(new_n601), .A3(new_n603), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n601), .B1(new_n600), .B2(new_n603), .ZN(new_n605));
  OAI21_X1  g419(.A(new_n599), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  XNOR2_X1  g420(.A(KEYINPUT22), .B(G137), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n339), .A2(G221), .A3(G234), .ZN(new_n608));
  XNOR2_X1  g422(.A(new_n607), .B(new_n608), .ZN(new_n609));
  INV_X1    g423(.A(new_n609), .ZN(new_n610));
  NAND2_X1  g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  OAI211_X1 g425(.A(new_n599), .B(new_n609), .C1(new_n604), .C2(new_n605), .ZN(new_n612));
  NAND3_X1  g426(.A1(new_n611), .A2(new_n313), .A3(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT25), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n611), .A2(KEYINPUT25), .A3(new_n313), .A4(new_n612), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n589), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AND2_X1   g431(.A1(new_n611), .A2(new_n612), .ZN(new_n618));
  NOR2_X1   g432(.A1(new_n588), .A2(G902), .ZN(new_n619));
  AOI21_X1  g433(.A(new_n617), .B1(new_n618), .B2(new_n619), .ZN(new_n620));
  XOR2_X1   g434(.A(new_n620), .B(KEYINPUT77), .Z(new_n621));
  NAND3_X1  g435(.A1(new_n332), .A2(new_n587), .A3(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n622), .B(G101), .ZN(G3));
  OAI21_X1  g437(.A(new_n313), .B1(new_n302), .B2(new_n303), .ZN(new_n624));
  AOI21_X1  g438(.A(new_n331), .B1(G472), .B2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n470), .A2(new_n472), .ZN(new_n626));
  NAND3_X1  g440(.A1(new_n625), .A2(new_n621), .A3(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n396), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n409), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n475), .B1(new_n629), .B2(new_n407), .ZN(new_n630));
  OR2_X1    g444(.A1(new_n577), .A2(new_n578), .ZN(new_n631));
  NAND2_X1  g445(.A1(new_n631), .A2(KEYINPUT33), .ZN(new_n632));
  OR3_X1    g446(.A1(new_n577), .A2(new_n578), .A3(KEYINPUT33), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n632), .A2(G478), .A3(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n631), .A2(new_n580), .A3(new_n313), .ZN(new_n635));
  NOR2_X1   g449(.A1(new_n580), .A2(new_n313), .ZN(new_n636));
  INV_X1    g450(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n634), .A2(new_n635), .A3(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(new_n638), .B1(new_n528), .B2(new_n536), .ZN(new_n639));
  AND3_X1   g453(.A1(new_n630), .A2(new_n639), .A3(new_n545), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NOR2_X1   g455(.A1(new_n627), .A2(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT34), .B(G104), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  INV_X1    g458(.A(KEYINPUT96), .ZN(new_n645));
  AND2_X1   g459(.A1(new_n402), .A2(new_n404), .ZN(new_n646));
  AOI22_X1  g460(.A1(new_n646), .A2(new_n405), .B1(new_n394), .B2(KEYINPUT86), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n396), .B1(new_n647), .B2(new_n398), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n474), .B1(new_n648), .B2(new_n408), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n516), .A2(new_n518), .A3(new_n521), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n650), .B1(new_n532), .B2(new_n533), .ZN(new_n651));
  INV_X1    g465(.A(new_n525), .ZN(new_n652));
  INV_X1    g466(.A(new_n526), .ZN(new_n653));
  AOI22_X1  g467(.A1(new_n582), .A2(new_n583), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g468(.A(new_n545), .B(KEYINPUT94), .Z(new_n655));
  NAND3_X1  g469(.A1(new_n651), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n656), .A2(KEYINPUT95), .ZN(new_n657));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n658));
  NAND4_X1  g472(.A1(new_n651), .A2(new_n654), .A3(new_n658), .A4(new_n655), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  OAI21_X1  g474(.A(new_n645), .B1(new_n649), .B2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n630), .A2(KEYINPUT96), .A3(new_n657), .A4(new_n659), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n627), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  XNOR2_X1  g477(.A(KEYINPUT35), .B(G107), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  NOR2_X1   g479(.A1(new_n413), .A2(new_n477), .ZN(new_n666));
  OR2_X1    g480(.A1(new_n610), .A2(KEYINPUT36), .ZN(new_n667));
  AND2_X1   g481(.A1(new_n606), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n606), .A2(new_n667), .ZN(new_n669));
  NOR4_X1   g483(.A1(new_n668), .A2(new_n669), .A3(G902), .A4(new_n588), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n617), .A2(new_n670), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n586), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n625), .A2(new_n666), .A3(new_n672), .ZN(new_n673));
  XOR2_X1   g487(.A(KEYINPUT37), .B(G110), .Z(new_n674));
  XNOR2_X1  g488(.A(new_n673), .B(new_n674), .ZN(G12));
  NAND2_X1  g489(.A1(new_n470), .A2(new_n472), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n649), .A2(new_n676), .A3(new_n671), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n541), .A2(G902), .A3(G953), .ZN(new_n678));
  OAI21_X1  g492(.A(new_n542), .B1(G900), .B2(new_n678), .ZN(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT97), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n651), .A2(new_n654), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND3_X1  g496(.A1(new_n332), .A2(new_n677), .A3(new_n682), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G128), .ZN(G30));
  AND2_X1   g498(.A1(new_n298), .A2(new_n300), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n306), .A2(new_n308), .ZN(new_n686));
  AOI21_X1  g500(.A(KEYINPUT98), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n298), .A2(new_n686), .A3(new_n300), .A4(KEYINPUT98), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n688), .A2(new_n313), .ZN(new_n689));
  OAI21_X1  g503(.A(G472), .B1(new_n687), .B2(new_n689), .ZN(new_n690));
  OAI211_X1 g504(.A(new_n304), .B(new_n690), .C1(new_n331), .C2(KEYINPUT32), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(KEYINPUT99), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n528), .A2(new_n536), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n694), .A2(new_n584), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n671), .A2(new_n474), .ZN(new_n696));
  XNOR2_X1  g510(.A(new_n680), .B(KEYINPUT39), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n626), .A2(new_n697), .ZN(new_n698));
  AOI211_X1 g512(.A(new_n695), .B(new_n696), .C1(new_n698), .C2(KEYINPUT40), .ZN(new_n699));
  OAI21_X1  g513(.A(new_n699), .B1(KEYINPUT40), .B2(new_n698), .ZN(new_n700));
  XNOR2_X1  g514(.A(new_n413), .B(KEYINPUT38), .ZN(new_n701));
  NOR3_X1   g515(.A1(new_n693), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(new_n196), .ZN(G45));
  INV_X1    g517(.A(new_n638), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n694), .A2(new_n704), .A3(new_n680), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n332), .A2(new_n677), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(G146), .ZN(G48));
  NAND2_X1  g522(.A1(new_n450), .A2(new_n447), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n458), .A2(new_n433), .ZN(new_n710));
  AOI22_X1  g524(.A1(new_n709), .A2(new_n462), .B1(new_n710), .B2(new_n436), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(G902), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n712), .A2(new_n460), .A3(new_n472), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n713), .A2(KEYINPUT100), .ZN(new_n714));
  INV_X1    g528(.A(KEYINPUT100), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n712), .A2(new_n460), .A3(new_n715), .A4(new_n472), .ZN(new_n716));
  AND2_X1   g530(.A1(new_n714), .A2(new_n716), .ZN(new_n717));
  NAND4_X1  g531(.A1(new_n332), .A2(new_n621), .A3(new_n717), .A4(new_n640), .ZN(new_n718));
  XNOR2_X1  g532(.A(KEYINPUT41), .B(G113), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n718), .B(new_n719), .ZN(G15));
  NAND2_X1  g534(.A1(new_n661), .A2(new_n662), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n721), .A2(new_n332), .A3(new_n621), .A4(new_n717), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G116), .ZN(G18));
  AND3_X1   g537(.A1(new_n714), .A2(new_n630), .A3(new_n716), .ZN(new_n724));
  NAND3_X1  g538(.A1(new_n332), .A2(new_n724), .A3(new_n672), .ZN(new_n725));
  XNOR2_X1  g539(.A(new_n725), .B(G119), .ZN(G21));
  INV_X1    g540(.A(KEYINPUT101), .ZN(new_n727));
  AOI21_X1  g541(.A(new_n195), .B1(new_n307), .B2(new_n283), .ZN(new_n728));
  OAI21_X1  g542(.A(new_n727), .B1(new_n323), .B2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n324), .B1(KEYINPUT28), .B2(new_n306), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n301), .B(KEYINPUT101), .C1(new_n195), .C2(new_n730), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n729), .A2(new_n327), .A3(new_n731), .ZN(new_n732));
  AOI22_X1  g546(.A1(G472), .A2(new_n624), .B1(new_n732), .B2(new_n187), .ZN(new_n733));
  AND3_X1   g547(.A1(new_n714), .A2(new_n655), .A3(new_n716), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n695), .A2(new_n649), .ZN(new_n735));
  NAND4_X1  g549(.A1(new_n733), .A2(new_n734), .A3(new_n620), .A4(new_n735), .ZN(new_n736));
  XNOR2_X1  g550(.A(new_n736), .B(G122), .ZN(G24));
  OR2_X1    g551(.A1(new_n617), .A2(new_n670), .ZN(new_n738));
  NAND4_X1  g552(.A1(new_n733), .A2(new_n724), .A3(new_n738), .A4(new_n706), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G125), .ZN(G27));
  XOR2_X1   g554(.A(KEYINPUT102), .B(KEYINPUT42), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n409), .A2(new_n410), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n742), .A2(new_n628), .A3(new_n412), .ZN(new_n743));
  NAND2_X1  g557(.A1(new_n407), .A2(new_n474), .ZN(new_n744));
  INV_X1    g558(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n743), .A2(new_n745), .ZN(new_n746));
  NOR2_X1   g560(.A1(new_n746), .A2(new_n676), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n332), .A2(new_n621), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n741), .B1(new_n748), .B2(new_n705), .ZN(new_n749));
  AOI21_X1  g563(.A(new_n744), .B1(new_n411), .B2(new_n412), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n706), .A2(new_n626), .A3(new_n750), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n332), .A2(KEYINPUT42), .A3(new_n620), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n749), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  NAND4_X1  g568(.A1(new_n332), .A2(new_n621), .A3(new_n747), .A4(new_n682), .ZN(new_n755));
  XOR2_X1   g569(.A(KEYINPUT103), .B(G134), .Z(new_n756));
  XNOR2_X1  g570(.A(new_n755), .B(new_n756), .ZN(G36));
  NOR2_X1   g571(.A1(new_n464), .A2(new_n466), .ZN(new_n758));
  AOI21_X1  g572(.A(new_n758), .B1(new_n458), .B2(new_n462), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n759), .B2(KEYINPUT45), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n760), .B1(KEYINPUT45), .B2(new_n759), .ZN(new_n761));
  OR2_X1    g575(.A1(new_n761), .A2(new_n468), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT46), .ZN(new_n763));
  OR2_X1    g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g578(.A(new_n460), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n765), .B1(new_n762), .B2(new_n763), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n473), .B1(new_n764), .B2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n767), .A2(new_n697), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT44), .ZN(new_n769));
  XOR2_X1   g583(.A(new_n694), .B(KEYINPUT104), .Z(new_n770));
  NAND3_X1  g584(.A1(new_n770), .A2(KEYINPUT43), .A3(new_n704), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n694), .A2(new_n638), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n771), .B1(KEYINPUT43), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(new_n625), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n773), .A2(new_n774), .A3(new_n738), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n768), .B1(new_n769), .B2(new_n775), .ZN(new_n776));
  OR2_X1    g590(.A1(new_n775), .A2(new_n769), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n777), .A2(KEYINPUT105), .A3(new_n750), .ZN(new_n778));
  NAND2_X1  g592(.A1(new_n776), .A2(new_n778), .ZN(new_n779));
  INV_X1    g593(.A(new_n779), .ZN(new_n780));
  AOI21_X1  g594(.A(KEYINPUT105), .B1(new_n777), .B2(new_n750), .ZN(new_n781));
  INV_X1    g595(.A(new_n781), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n780), .A2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G137), .ZN(G39));
  OR2_X1    g598(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n785));
  NAND2_X1  g599(.A1(KEYINPUT106), .A2(KEYINPUT47), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n767), .B1(new_n785), .B2(new_n786), .ZN(new_n787));
  AND2_X1   g601(.A1(new_n767), .A2(new_n786), .ZN(new_n788));
  OR4_X1    g602(.A1(new_n332), .A2(new_n621), .A3(new_n705), .A4(new_n746), .ZN(new_n789));
  NOR3_X1   g603(.A1(new_n787), .A2(new_n788), .A3(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n483), .ZN(G42));
  NAND2_X1  g605(.A1(new_n712), .A2(new_n460), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT49), .Z(new_n793));
  AND4_X1   g607(.A1(new_n620), .A2(new_n793), .A3(new_n476), .A4(new_n704), .ZN(new_n794));
  NAND4_X1  g608(.A1(new_n693), .A2(new_n701), .A3(new_n770), .A4(new_n794), .ZN(new_n795));
  XOR2_X1   g609(.A(KEYINPUT113), .B(KEYINPUT54), .Z(new_n796));
  OAI211_X1 g610(.A(new_n332), .B(new_n677), .C1(new_n682), .C2(new_n706), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n671), .A2(new_n680), .ZN(new_n798));
  INV_X1    g612(.A(new_n798), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n626), .A2(KEYINPUT110), .A3(new_n799), .ZN(new_n800));
  INV_X1    g614(.A(KEYINPUT110), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n801), .B1(new_n676), .B2(new_n798), .ZN(new_n802));
  NAND4_X1  g616(.A1(new_n691), .A2(new_n735), .A3(new_n800), .A4(new_n802), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n797), .A2(new_n739), .A3(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT52), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n797), .A2(new_n739), .A3(new_n803), .A4(KEYINPUT52), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n808), .A2(KEYINPUT111), .ZN(new_n809));
  INV_X1    g623(.A(KEYINPUT111), .ZN(new_n810));
  NAND3_X1  g624(.A1(new_n806), .A2(new_n810), .A3(new_n807), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n809), .A2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n624), .A2(G472), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n732), .A2(new_n187), .ZN(new_n814));
  NAND3_X1  g628(.A1(new_n813), .A2(new_n814), .A3(new_n738), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT109), .B1(new_n815), .B2(new_n751), .ZN(new_n816));
  NOR3_X1   g630(.A1(new_n746), .A2(new_n705), .A3(new_n676), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT109), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n817), .A2(new_n733), .A3(new_n818), .A4(new_n738), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  INV_X1    g634(.A(KEYINPUT108), .ZN(new_n821));
  INV_X1    g635(.A(new_n680), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n527), .A2(new_n822), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n651), .A2(new_n585), .A3(new_n823), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n470), .A2(new_n824), .A3(new_n738), .A4(new_n472), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n746), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n332), .A2(new_n821), .A3(new_n826), .ZN(new_n827));
  AOI21_X1  g641(.A(new_n821), .B1(new_n332), .B2(new_n826), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n755), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n820), .A2(new_n829), .ZN(new_n830));
  AND3_X1   g644(.A1(new_n528), .A2(new_n536), .A3(new_n584), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT107), .B1(new_n831), .B2(new_n639), .ZN(new_n832));
  INV_X1    g646(.A(KEYINPUT107), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n833), .B1(new_n694), .B2(new_n585), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  INV_X1    g649(.A(new_n655), .ZN(new_n836));
  NOR3_X1   g650(.A1(new_n413), .A2(new_n477), .A3(new_n836), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n835), .A2(new_n625), .A3(new_n621), .A4(new_n837), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n722), .A2(new_n718), .A3(new_n838), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n736), .A2(new_n673), .A3(new_n725), .A4(new_n622), .ZN(new_n840));
  NOR2_X1   g654(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  AND3_X1   g655(.A1(new_n830), .A2(new_n841), .A3(new_n753), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n812), .A2(KEYINPUT53), .A3(new_n842), .ZN(new_n843));
  NAND4_X1  g657(.A1(new_n808), .A2(new_n830), .A3(new_n753), .A4(new_n841), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT53), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n844), .A2(KEYINPUT112), .A3(new_n845), .ZN(new_n846));
  AOI21_X1  g660(.A(KEYINPUT112), .B1(new_n844), .B2(new_n845), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n796), .B(new_n843), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT53), .B1(new_n812), .B2(new_n842), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n844), .A2(new_n845), .ZN(new_n850));
  OAI21_X1  g664(.A(KEYINPUT54), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n848), .A2(new_n851), .ZN(new_n852));
  INV_X1    g666(.A(KEYINPUT114), .ZN(new_n853));
  NAND2_X1  g667(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n848), .A2(new_n851), .A3(KEYINPUT114), .ZN(new_n855));
  NAND2_X1  g669(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI22_X1  g670(.A1(new_n787), .A2(new_n788), .B1(new_n472), .B2(new_n792), .ZN(new_n857));
  INV_X1    g671(.A(new_n542), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n773), .A2(new_n858), .ZN(new_n859));
  AND2_X1   g673(.A1(new_n733), .A2(new_n620), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  INV_X1    g675(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n857), .A2(new_n750), .A3(new_n862), .ZN(new_n863));
  INV_X1    g677(.A(new_n717), .ZN(new_n864));
  NOR2_X1   g678(.A1(new_n864), .A2(new_n746), .ZN(new_n865));
  OR2_X1    g679(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n865), .A2(KEYINPUT115), .ZN(new_n867));
  NAND2_X1  g681(.A1(new_n866), .A2(new_n867), .ZN(new_n868));
  INV_X1    g682(.A(new_n868), .ZN(new_n869));
  NAND2_X1  g683(.A1(new_n869), .A2(new_n859), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n870), .A2(new_n815), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT50), .ZN(new_n872));
  INV_X1    g686(.A(new_n701), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n873), .A2(new_n474), .A3(new_n864), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n872), .B1(new_n861), .B2(new_n875), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n862), .A2(KEYINPUT50), .A3(new_n874), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n871), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n621), .A2(new_n858), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n869), .A2(KEYINPUT116), .A3(new_n693), .A4(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT116), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n693), .A2(new_n879), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n881), .B1(new_n868), .B2(new_n882), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n694), .A2(new_n704), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n880), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g699(.A1(new_n863), .A2(new_n878), .A3(new_n885), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT51), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n880), .A2(new_n639), .A3(new_n883), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n540), .B(KEYINPUT117), .ZN(new_n890));
  INV_X1    g704(.A(new_n724), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n890), .B1(new_n861), .B2(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n332), .A2(new_n620), .ZN(new_n893));
  OR3_X1    g707(.A1(new_n870), .A2(KEYINPUT48), .A3(new_n893), .ZN(new_n894));
  OAI21_X1  g708(.A(KEYINPUT48), .B1(new_n870), .B2(new_n893), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n892), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n888), .A2(new_n889), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n886), .A2(new_n887), .ZN(new_n898));
  NOR3_X1   g712(.A1(new_n856), .A2(new_n897), .A3(new_n898), .ZN(new_n899));
  NOR2_X1   g713(.A1(G952), .A2(G953), .ZN(new_n900));
  OAI21_X1  g714(.A(new_n795), .B1(new_n899), .B2(new_n900), .ZN(G75));
  NOR2_X1   g715(.A1(new_n339), .A2(G952), .ZN(new_n902));
  INV_X1    g716(.A(KEYINPUT56), .ZN(new_n903));
  OAI21_X1  g717(.A(new_n843), .B1(new_n846), .B2(new_n847), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(G902), .ZN(new_n905));
  INV_X1    g719(.A(G210), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n903), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  XNOR2_X1  g721(.A(new_n646), .B(new_n405), .ZN(new_n908));
  XNOR2_X1  g722(.A(KEYINPUT118), .B(KEYINPUT55), .ZN(new_n909));
  XNOR2_X1  g723(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n907), .A2(new_n910), .ZN(new_n911));
  XNOR2_X1  g725(.A(new_n905), .B(KEYINPUT119), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(new_n628), .ZN(new_n913));
  NOR2_X1   g727(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n914));
  AOI211_X1 g728(.A(new_n902), .B(new_n911), .C1(new_n913), .C2(new_n914), .ZN(G51));
  INV_X1    g729(.A(KEYINPUT120), .ZN(new_n916));
  INV_X1    g730(.A(new_n796), .ZN(new_n917));
  AND3_X1   g731(.A1(new_n904), .A2(new_n916), .A3(new_n917), .ZN(new_n918));
  AOI21_X1  g732(.A(new_n916), .B1(new_n904), .B2(new_n917), .ZN(new_n919));
  INV_X1    g733(.A(new_n848), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n918), .A2(new_n919), .A3(new_n920), .ZN(new_n921));
  XOR2_X1   g735(.A(new_n468), .B(KEYINPUT57), .Z(new_n922));
  OAI22_X1  g736(.A1(new_n921), .A2(new_n922), .B1(new_n459), .B2(new_n451), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n912), .A2(new_n761), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n902), .B1(new_n923), .B2(new_n924), .ZN(G54));
  AND2_X1   g739(.A1(KEYINPUT58), .A2(G475), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n912), .A2(new_n926), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n516), .A2(new_n518), .ZN(new_n928));
  NAND2_X1  g742(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  INV_X1    g743(.A(new_n902), .ZN(new_n930));
  NAND4_X1  g744(.A1(new_n912), .A2(new_n516), .A3(new_n518), .A4(new_n926), .ZN(new_n931));
  AND3_X1   g745(.A1(new_n929), .A2(new_n930), .A3(new_n931), .ZN(G60));
  AND2_X1   g746(.A1(new_n632), .A2(new_n633), .ZN(new_n933));
  INV_X1    g747(.A(new_n933), .ZN(new_n934));
  XNOR2_X1  g748(.A(KEYINPUT121), .B(KEYINPUT59), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n935), .B(new_n636), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n934), .A2(new_n936), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n930), .B1(new_n921), .B2(new_n937), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n934), .B1(new_n856), .B2(new_n936), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT122), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  INV_X1    g754(.A(new_n855), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT114), .B1(new_n848), .B2(new_n851), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n936), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n933), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n904), .A2(new_n917), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n945), .A2(KEYINPUT120), .ZN(new_n946));
  NAND3_X1  g760(.A1(new_n904), .A2(new_n916), .A3(new_n917), .ZN(new_n947));
  NAND3_X1  g761(.A1(new_n946), .A2(new_n848), .A3(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n937), .ZN(new_n949));
  AOI21_X1  g763(.A(new_n902), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g764(.A(KEYINPUT122), .ZN(new_n951));
  NAND3_X1  g765(.A1(new_n944), .A2(new_n950), .A3(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n940), .A2(new_n952), .ZN(G63));
  NAND2_X1  g767(.A1(G217), .A2(G902), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n954), .B(KEYINPUT60), .Z(new_n955));
  NAND2_X1  g769(.A1(new_n904), .A2(new_n955), .ZN(new_n956));
  OR3_X1    g770(.A1(new_n956), .A2(new_n669), .A3(new_n668), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n618), .B(KEYINPUT124), .ZN(new_n958));
  AOI21_X1  g772(.A(new_n902), .B1(new_n956), .B2(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n957), .A2(new_n959), .ZN(new_n960));
  AOI21_X1  g774(.A(KEYINPUT61), .B1(new_n959), .B2(KEYINPUT123), .ZN(new_n961));
  XNOR2_X1  g775(.A(new_n960), .B(new_n961), .ZN(G66));
  INV_X1    g776(.A(G224), .ZN(new_n963));
  OAI21_X1  g777(.A(G953), .B1(new_n543), .B2(new_n963), .ZN(new_n964));
  XOR2_X1   g778(.A(new_n964), .B(KEYINPUT125), .Z(new_n965));
  OAI21_X1  g779(.A(new_n965), .B1(new_n841), .B2(G953), .ZN(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT126), .Z(new_n967));
  INV_X1    g781(.A(G898), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n646), .B1(new_n968), .B2(G953), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n967), .B(new_n969), .ZN(G69));
  AOI21_X1  g784(.A(new_n339), .B1(G227), .B2(G900), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n287), .A2(new_n288), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n486), .A2(new_n487), .ZN(new_n973));
  XNOR2_X1  g787(.A(new_n972), .B(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n790), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n975), .B1(new_n779), .B2(new_n781), .ZN(new_n976));
  OR4_X1    g790(.A1(new_n649), .A2(new_n768), .A3(new_n695), .A4(new_n893), .ZN(new_n977));
  NAND2_X1  g791(.A1(new_n797), .A2(new_n739), .ZN(new_n978));
  INV_X1    g792(.A(new_n978), .ZN(new_n979));
  NAND4_X1  g793(.A1(new_n977), .A2(new_n753), .A3(new_n755), .A4(new_n979), .ZN(new_n980));
  OAI211_X1 g794(.A(new_n339), .B(new_n974), .C1(new_n976), .C2(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(new_n976), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n835), .A2(new_n697), .ZN(new_n983));
  NOR2_X1   g797(.A1(new_n983), .A2(new_n748), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT62), .ZN(new_n985));
  OR3_X1    g799(.A1(new_n702), .A2(new_n985), .A3(new_n978), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n985), .B1(new_n702), .B2(new_n978), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n984), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  AOI21_X1  g802(.A(G953), .B1(new_n982), .B2(new_n988), .ZN(new_n989));
  OAI21_X1  g803(.A(new_n981), .B1(new_n989), .B2(new_n974), .ZN(new_n990));
  INV_X1    g804(.A(G900), .ZN(new_n991));
  OAI21_X1  g805(.A(new_n971), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n992), .B1(new_n971), .B2(new_n990), .ZN(G72));
  XNOR2_X1  g807(.A(new_n315), .B(KEYINPUT127), .ZN(new_n994));
  NOR4_X1   g808(.A1(new_n976), .A2(new_n980), .A3(new_n840), .A4(new_n839), .ZN(new_n995));
  NAND2_X1  g809(.A1(G472), .A2(G902), .ZN(new_n996));
  XOR2_X1   g810(.A(new_n996), .B(KEYINPUT63), .Z(new_n997));
  INV_X1    g811(.A(new_n997), .ZN(new_n998));
  OAI211_X1 g812(.A(new_n308), .B(new_n994), .C1(new_n995), .C2(new_n998), .ZN(new_n999));
  AOI21_X1  g813(.A(new_n998), .B1(new_n685), .B2(new_n316), .ZN(new_n1000));
  OAI21_X1  g814(.A(new_n1000), .B1(new_n849), .B2(new_n850), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n994), .A2(new_n308), .ZN(new_n1002));
  AND3_X1   g816(.A1(new_n982), .A2(new_n841), .A3(new_n988), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n1002), .B1(new_n1003), .B2(new_n998), .ZN(new_n1004));
  AND4_X1   g818(.A1(new_n930), .A2(new_n999), .A3(new_n1001), .A4(new_n1004), .ZN(G57));
endmodule


