//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 1 0 1 0 0 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 1 0 0 1 0 1 1 0 0 0 1 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:54 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n446, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n561, new_n563, new_n564, new_n566, new_n567, new_n568,
    new_n569, new_n570, new_n571, new_n572, new_n573, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n605, new_n606, new_n609, new_n610, new_n612,
    new_n613, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n894, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1106,
    new_n1107;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT64), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  NAND2_X1  g020(.A1(G94), .A2(G452), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT65), .Z(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT66), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  OR4_X1    g029(.A1(G237), .A2(G236), .A3(G235), .A4(G238), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n454), .A2(new_n455), .ZN(G325));
  XNOR2_X1  g031(.A(G325), .B(KEYINPUT67), .ZN(G261));
  NAND2_X1  g032(.A1(new_n454), .A2(G2106), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n455), .A2(G567), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  INV_X1    g035(.A(new_n460), .ZN(G319));
  INV_X1    g036(.A(G2105), .ZN(new_n462));
  XNOR2_X1  g037(.A(KEYINPUT3), .B(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G125), .ZN(new_n464));
  NAND2_X1  g039(.A1(G113), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(new_n462), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(G101), .A2(G2104), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  OAI21_X1  g043(.A(KEYINPUT69), .B1(new_n468), .B2(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n468), .A2(KEYINPUT68), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT68), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(KEYINPUT3), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  AOI21_X1  g048(.A(new_n469), .B1(new_n473), .B2(G2104), .ZN(new_n474));
  INV_X1    g049(.A(G2104), .ZN(new_n475));
  AOI211_X1 g050(.A(KEYINPUT69), .B(new_n475), .C1(new_n470), .C2(new_n472), .ZN(new_n476));
  NOR2_X1   g051(.A1(new_n474), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(G137), .ZN(new_n478));
  OAI21_X1  g053(.A(new_n467), .B1(new_n477), .B2(new_n478), .ZN(new_n479));
  AOI21_X1  g054(.A(new_n466), .B1(new_n479), .B2(new_n462), .ZN(G160));
  NOR2_X1   g055(.A1(new_n477), .A2(new_n462), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G124), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n477), .A2(G2105), .ZN(new_n483));
  NAND2_X1  g058(.A1(new_n483), .A2(G136), .ZN(new_n484));
  NOR2_X1   g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT70), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G112), .C2(new_n462), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n482), .A2(new_n484), .A3(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(new_n488), .ZN(G162));
  XNOR2_X1  g064(.A(KEYINPUT71), .B(G114), .ZN(new_n490));
  OAI21_X1  g065(.A(KEYINPUT72), .B1(new_n490), .B2(new_n462), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT72), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT71), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G114), .ZN(new_n494));
  INV_X1    g069(.A(G114), .ZN(new_n495));
  NOR2_X1   g070(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n496));
  OAI211_X1 g071(.A(new_n492), .B(G2105), .C1(new_n494), .C2(new_n496), .ZN(new_n497));
  NAND2_X1  g072(.A1(new_n491), .A2(new_n497), .ZN(new_n498));
  OAI21_X1  g073(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  AOI21_X1  g075(.A(KEYINPUT73), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT73), .ZN(new_n502));
  AOI211_X1 g077(.A(new_n502), .B(new_n499), .C1(new_n491), .C2(new_n497), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n501), .A2(new_n503), .ZN(new_n504));
  OAI211_X1 g079(.A(G126), .B(G2105), .C1(new_n474), .C2(new_n476), .ZN(new_n505));
  AND2_X1   g080(.A1(KEYINPUT4), .A2(G138), .ZN(new_n506));
  OAI211_X1 g081(.A(new_n462), .B(new_n506), .C1(new_n474), .C2(new_n476), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n463), .A2(G138), .A3(new_n462), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT4), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n504), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(G543), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(KEYINPUT5), .ZN(new_n514));
  INV_X1    g089(.A(KEYINPUT5), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G543), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n514), .A2(new_n516), .ZN(new_n517));
  INV_X1    g092(.A(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n518), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AND2_X1   g096(.A1(KEYINPUT6), .A2(G651), .ZN(new_n522));
  NOR2_X1   g097(.A1(KEYINPUT6), .A2(G651), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n518), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G88), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(G543), .ZN(new_n527));
  INV_X1    g102(.A(G50), .ZN(new_n528));
  OAI22_X1  g103(.A1(new_n525), .A2(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OR2_X1    g104(.A1(new_n521), .A2(new_n529), .ZN(G303));
  INV_X1    g105(.A(G303), .ZN(G166));
  AOI22_X1  g106(.A1(new_n524), .A2(G89), .B1(G63), .B2(G651), .ZN(new_n532));
  INV_X1    g107(.A(new_n532), .ZN(new_n533));
  NOR2_X1   g108(.A1(new_n522), .A2(new_n523), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n534), .A2(new_n513), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n533), .A2(new_n518), .B1(new_n535), .B2(G51), .ZN(new_n536));
  NAND3_X1  g111(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT7), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n536), .A2(new_n538), .ZN(G286));
  INV_X1    g114(.A(G286), .ZN(G168));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  XNOR2_X1  g116(.A(KEYINPUT74), .B(G52), .ZN(new_n542));
  OAI22_X1  g117(.A1(new_n525), .A2(new_n541), .B1(new_n527), .B2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT75), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(new_n545));
  AOI22_X1  g120(.A1(new_n518), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n546));
  OR2_X1    g121(.A1(new_n546), .A2(new_n520), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n545), .A2(new_n547), .ZN(G301));
  INV_X1    g123(.A(G301), .ZN(G171));
  NAND2_X1  g124(.A1(G68), .A2(G543), .ZN(new_n550));
  INV_X1    g125(.A(G56), .ZN(new_n551));
  OAI21_X1  g126(.A(new_n550), .B1(new_n517), .B2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT76), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G651), .ZN(new_n554));
  INV_X1    g129(.A(new_n525), .ZN(new_n555));
  XNOR2_X1  g130(.A(KEYINPUT77), .B(G43), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n555), .A2(G81), .B1(new_n535), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n554), .A2(new_n557), .ZN(new_n558));
  INV_X1    g133(.A(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(G153));
  AND3_X1   g135(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G36), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n561), .A2(new_n564), .ZN(G188));
  NAND2_X1  g140(.A1(new_n535), .A2(G53), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  INV_X1    g142(.A(G78), .ZN(new_n568));
  OR3_X1    g143(.A1(new_n568), .A2(new_n513), .A3(KEYINPUT78), .ZN(new_n569));
  OAI21_X1  g144(.A(KEYINPUT78), .B1(new_n568), .B2(new_n513), .ZN(new_n570));
  INV_X1    g145(.A(G65), .ZN(new_n571));
  OAI211_X1 g146(.A(new_n569), .B(new_n570), .C1(new_n571), .C2(new_n517), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n555), .A2(G91), .B1(new_n572), .B2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n567), .A2(new_n573), .ZN(G299));
  OAI21_X1  g149(.A(G651), .B1(new_n518), .B2(G74), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n535), .A2(G49), .ZN(new_n576));
  INV_X1    g151(.A(G87), .ZN(new_n577));
  OAI211_X1 g152(.A(new_n575), .B(new_n576), .C1(new_n577), .C2(new_n525), .ZN(G288));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(new_n579), .B1(new_n517), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(new_n581), .A2(G651), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n535), .A2(G48), .ZN(new_n583));
  INV_X1    g158(.A(G86), .ZN(new_n584));
  OAI211_X1 g159(.A(new_n582), .B(new_n583), .C1(new_n584), .C2(new_n525), .ZN(G305));
  AOI22_X1  g160(.A1(new_n518), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n586), .A2(new_n520), .ZN(new_n587));
  INV_X1    g162(.A(G85), .ZN(new_n588));
  INV_X1    g163(.A(G47), .ZN(new_n589));
  OAI22_X1  g164(.A1(new_n525), .A2(new_n588), .B1(new_n527), .B2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n587), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  OR3_X1    g168(.A1(new_n525), .A2(KEYINPUT10), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g169(.A1(G79), .A2(G543), .ZN(new_n595));
  INV_X1    g170(.A(G66), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n517), .B2(new_n596), .ZN(new_n597));
  AOI22_X1  g172(.A1(new_n597), .A2(G651), .B1(new_n535), .B2(G54), .ZN(new_n598));
  OAI21_X1  g173(.A(KEYINPUT10), .B1(new_n525), .B2(new_n593), .ZN(new_n599));
  NAND3_X1  g174(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G284));
  OAI21_X1  g178(.A(new_n602), .B1(G171), .B2(new_n601), .ZN(G321));
  NOR2_X1   g179(.A1(G168), .A2(new_n601), .ZN(new_n605));
  AOI21_X1  g180(.A(new_n605), .B1(new_n601), .B2(G299), .ZN(new_n606));
  XOR2_X1   g181(.A(new_n606), .B(KEYINPUT79), .Z(G297));
  XNOR2_X1  g182(.A(new_n606), .B(KEYINPUT80), .ZN(G280));
  AND3_X1   g183(.A1(new_n594), .A2(new_n598), .A3(new_n599), .ZN(new_n609));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n609), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n558), .A2(new_n601), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n600), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n601), .B2(new_n613), .ZN(G323));
  XNOR2_X1  g189(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g190(.A1(new_n481), .A2(G123), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n483), .A2(G135), .ZN(new_n617));
  NOR2_X1   g192(.A1(G99), .A2(G2105), .ZN(new_n618));
  OAI21_X1  g193(.A(G2104), .B1(new_n462), .B2(G111), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n616), .B(new_n617), .C1(new_n618), .C2(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND3_X1  g196(.A1(new_n462), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XOR2_X1   g206(.A(G2451), .B(G2454), .Z(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT16), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n631), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(G1341), .B(G1348), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n634), .B(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2443), .B(G2446), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n636), .B(new_n637), .Z(new_n638));
  AND2_X1   g213(.A1(new_n638), .A2(G14), .ZN(G401));
  XNOR2_X1  g214(.A(G2072), .B(G2078), .ZN(new_n640));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT81), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  AND2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(KEYINPUT82), .B(KEYINPUT18), .ZN(new_n646));
  OAI21_X1  g221(.A(new_n640), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2096), .B(G2100), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  OAI21_X1  g224(.A(KEYINPUT17), .B1(new_n643), .B2(new_n644), .ZN(new_n650));
  OAI21_X1  g225(.A(new_n646), .B1(new_n645), .B2(new_n650), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n649), .B(new_n651), .ZN(G227));
  XNOR2_X1  g227(.A(G1971), .B(G1976), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT83), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n654), .B(KEYINPUT19), .Z(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G1956), .B(G2474), .Z(new_n657));
  XOR2_X1   g232(.A(G1961), .B(G1966), .Z(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NOR2_X1   g234(.A1(new_n656), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g235(.A(KEYINPUT84), .B(KEYINPUT20), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n660), .B(new_n661), .ZN(new_n662));
  NOR2_X1   g237(.A1(new_n657), .A2(new_n658), .ZN(new_n663));
  INV_X1    g238(.A(new_n663), .ZN(new_n664));
  NAND3_X1  g239(.A1(new_n656), .A2(new_n664), .A3(new_n659), .ZN(new_n665));
  OAI211_X1 g240(.A(new_n662), .B(new_n665), .C1(new_n664), .C2(new_n656), .ZN(new_n666));
  XOR2_X1   g241(.A(KEYINPUT21), .B(G1986), .Z(new_n667));
  XNOR2_X1  g242(.A(new_n666), .B(new_n667), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(KEYINPUT22), .B(G1981), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(G229));
  NOR2_X1   g247(.A1(G29), .A2(G33), .ZN(new_n673));
  AOI22_X1  g248(.A1(new_n463), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n674), .A2(new_n462), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n462), .A2(G103), .A3(G2104), .ZN(new_n676));
  XOR2_X1   g251(.A(new_n676), .B(KEYINPUT25), .Z(new_n677));
  OR2_X1    g252(.A1(new_n474), .A2(new_n476), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n678), .A2(new_n462), .ZN(new_n679));
  INV_X1    g254(.A(G139), .ZN(new_n680));
  OAI211_X1 g255(.A(new_n675), .B(new_n677), .C1(new_n679), .C2(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT91), .ZN(new_n682));
  INV_X1    g257(.A(KEYINPUT92), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n673), .B1(new_n684), .B2(G29), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n685), .B(G2072), .ZN(new_n686));
  INV_X1    g261(.A(G29), .ZN(new_n687));
  INV_X1    g262(.A(G34), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(KEYINPUT24), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(KEYINPUT24), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n687), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g266(.A(new_n691), .B1(G160), .B2(new_n687), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n686), .B1(G2084), .B2(new_n692), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n687), .A2(G26), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n481), .A2(G128), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n483), .A2(G140), .ZN(new_n696));
  OR2_X1    g271(.A1(G104), .A2(G2105), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n697), .B(G2104), .C1(G116), .C2(new_n462), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n695), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  OAI21_X1  g275(.A(new_n694), .B1(new_n700), .B2(new_n687), .ZN(new_n701));
  MUX2_X1   g276(.A(new_n694), .B(new_n701), .S(KEYINPUT28), .Z(new_n702));
  INV_X1    g277(.A(G2067), .ZN(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(G16), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(G19), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n706), .B1(new_n559), .B2(new_n705), .ZN(new_n707));
  XOR2_X1   g282(.A(new_n707), .B(G1341), .Z(new_n708));
  NAND2_X1  g283(.A1(new_n705), .A2(G20), .ZN(new_n709));
  XOR2_X1   g284(.A(new_n709), .B(KEYINPUT96), .Z(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(KEYINPUT23), .ZN(new_n711));
  AOI21_X1  g286(.A(new_n711), .B1(G299), .B2(G16), .ZN(new_n712));
  INV_X1    g287(.A(G1956), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n712), .B(new_n713), .ZN(new_n714));
  NAND2_X1  g289(.A1(G171), .A2(G16), .ZN(new_n715));
  OAI21_X1  g290(.A(new_n715), .B1(G5), .B2(G16), .ZN(new_n716));
  INV_X1    g291(.A(G1961), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(new_n716), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g293(.A1(new_n704), .A2(new_n708), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n687), .A2(G27), .ZN(new_n720));
  OAI21_X1  g295(.A(new_n720), .B1(G164), .B2(new_n687), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G2078), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n687), .A2(G35), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(G162), .B2(new_n687), .ZN(new_n724));
  XNOR2_X1  g299(.A(new_n724), .B(G2090), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR3_X1   g302(.A1(new_n719), .A2(new_n722), .A3(new_n727), .ZN(new_n728));
  OAI211_X1 g303(.A(new_n693), .B(new_n728), .C1(G2084), .C2(new_n692), .ZN(new_n729));
  NOR2_X1   g304(.A1(G16), .A2(G23), .ZN(new_n730));
  XNOR2_X1  g305(.A(G288), .B(KEYINPUT87), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n730), .B1(new_n731), .B2(G16), .ZN(new_n732));
  INV_X1    g307(.A(KEYINPUT88), .ZN(new_n733));
  AND2_X1   g308(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n732), .A2(new_n733), .ZN(new_n735));
  XNOR2_X1  g310(.A(KEYINPUT33), .B(G1976), .ZN(new_n736));
  INV_X1    g311(.A(new_n736), .ZN(new_n737));
  OR3_X1    g312(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n705), .A2(G22), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G166), .B2(new_n705), .ZN(new_n740));
  INV_X1    g315(.A(G1971), .ZN(new_n741));
  XNOR2_X1  g316(.A(new_n740), .B(new_n741), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(new_n743));
  MUX2_X1   g318(.A(G6), .B(G305), .S(G16), .Z(new_n744));
  XOR2_X1   g319(.A(KEYINPUT32), .B(G1981), .Z(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  NAND4_X1  g321(.A1(new_n738), .A2(new_n742), .A3(new_n743), .A4(new_n746), .ZN(new_n747));
  AND2_X1   g322(.A1(new_n747), .A2(KEYINPUT89), .ZN(new_n748));
  NOR2_X1   g323(.A1(new_n747), .A2(KEYINPUT89), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT34), .ZN(new_n750));
  OR3_X1    g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G16), .A2(G24), .ZN(new_n752));
  XOR2_X1   g327(.A(new_n591), .B(KEYINPUT86), .Z(new_n753));
  AOI21_X1  g328(.A(new_n752), .B1(new_n753), .B2(G16), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n754), .B(G1986), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n481), .A2(G119), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n483), .A2(G131), .ZN(new_n757));
  NOR2_X1   g332(.A1(G95), .A2(G2105), .ZN(new_n758));
  OAI21_X1  g333(.A(G2104), .B1(new_n462), .B2(G107), .ZN(new_n759));
  OAI211_X1 g334(.A(new_n756), .B(new_n757), .C1(new_n758), .C2(new_n759), .ZN(new_n760));
  MUX2_X1   g335(.A(G25), .B(new_n760), .S(G29), .Z(new_n761));
  XOR2_X1   g336(.A(KEYINPUT35), .B(G1991), .Z(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT85), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n761), .B(new_n763), .ZN(new_n764));
  NOR2_X1   g339(.A1(new_n755), .A2(new_n764), .ZN(new_n765));
  OAI21_X1  g340(.A(new_n750), .B1(new_n748), .B2(new_n749), .ZN(new_n766));
  NAND3_X1  g341(.A1(new_n751), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n767), .A2(KEYINPUT36), .ZN(new_n768));
  INV_X1    g343(.A(KEYINPUT36), .ZN(new_n769));
  NAND4_X1  g344(.A1(new_n751), .A2(new_n769), .A3(new_n765), .A4(new_n766), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n729), .B1(new_n768), .B2(new_n770), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT31), .B(G11), .Z(new_n772));
  INV_X1    g347(.A(KEYINPUT30), .ZN(new_n773));
  AND2_X1   g348(.A1(new_n773), .A2(G28), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n773), .A2(G28), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n774), .A2(new_n775), .A3(G29), .ZN(new_n776));
  OR3_X1    g351(.A1(new_n716), .A2(KEYINPUT93), .A3(new_n717), .ZN(new_n777));
  OAI21_X1  g352(.A(KEYINPUT93), .B1(new_n716), .B2(new_n717), .ZN(new_n778));
  AOI211_X1 g353(.A(new_n772), .B(new_n776), .C1(new_n777), .C2(new_n778), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n705), .A2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(G168), .B2(new_n705), .ZN(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n781), .B(new_n782), .ZN(new_n783));
  OAI211_X1 g358(.A(new_n779), .B(new_n783), .C1(new_n687), .C2(new_n620), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT94), .Z(new_n785));
  NOR2_X1   g360(.A1(G29), .A2(G32), .ZN(new_n786));
  AOI22_X1  g361(.A1(new_n678), .A2(G141), .B1(G105), .B2(G2104), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(G2105), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n481), .A2(G129), .ZN(new_n789));
  NAND3_X1  g364(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n790));
  XOR2_X1   g365(.A(new_n790), .B(KEYINPUT26), .Z(new_n791));
  NAND3_X1  g366(.A1(new_n788), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  INV_X1    g367(.A(new_n792), .ZN(new_n793));
  AOI21_X1  g368(.A(new_n786), .B1(new_n793), .B2(G29), .ZN(new_n794));
  XNOR2_X1  g369(.A(KEYINPUT27), .B(G1996), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  OAI21_X1  g371(.A(KEYINPUT90), .B1(G4), .B2(G16), .ZN(new_n797));
  OR3_X1    g372(.A1(KEYINPUT90), .A2(G4), .A3(G16), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n797), .B(new_n798), .C1(new_n600), .C2(new_n705), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1348), .Z(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  NAND4_X1  g376(.A1(new_n771), .A2(new_n785), .A3(new_n796), .A4(new_n801), .ZN(G150));
  INV_X1    g377(.A(KEYINPUT97), .ZN(new_n803));
  NAND2_X1  g378(.A1(G150), .A2(new_n803), .ZN(new_n804));
  AOI211_X1 g379(.A(new_n800), .B(new_n729), .C1(new_n768), .C2(new_n770), .ZN(new_n805));
  NAND4_X1  g380(.A1(new_n805), .A2(KEYINPUT97), .A3(new_n785), .A4(new_n796), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n804), .A2(new_n806), .ZN(G311));
  AOI22_X1  g382(.A1(new_n518), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n808), .A2(new_n520), .ZN(new_n809));
  XNOR2_X1  g384(.A(KEYINPUT98), .B(G93), .ZN(new_n810));
  INV_X1    g385(.A(G55), .ZN(new_n811));
  OAI22_X1  g386(.A1(new_n525), .A2(new_n810), .B1(new_n527), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G860), .ZN(new_n814));
  NOR2_X1   g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT37), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n558), .B1(KEYINPUT99), .B2(new_n813), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n813), .A2(KEYINPUT99), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n817), .B(new_n818), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n819), .B(KEYINPUT38), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n609), .A2(G559), .ZN(new_n821));
  XNOR2_X1  g396(.A(new_n820), .B(new_n821), .ZN(new_n822));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(KEYINPUT100), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n814), .B1(new_n822), .B2(new_n823), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n816), .B1(new_n825), .B2(new_n826), .ZN(G145));
  INV_X1    g402(.A(KEYINPUT101), .ZN(new_n828));
  INV_X1    g403(.A(G142), .ZN(new_n829));
  OAI21_X1  g404(.A(new_n828), .B1(new_n679), .B2(new_n829), .ZN(new_n830));
  OAI21_X1  g405(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n831));
  INV_X1    g406(.A(new_n831), .ZN(new_n832));
  NOR2_X1   g407(.A1(new_n462), .A2(G118), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT102), .ZN(new_n834));
  AOI22_X1  g409(.A1(new_n481), .A2(G130), .B1(new_n832), .B2(new_n834), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n483), .A2(KEYINPUT101), .A3(G142), .ZN(new_n836));
  NAND3_X1  g411(.A1(new_n830), .A2(new_n835), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g412(.A(new_n837), .B(new_n760), .Z(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT103), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(new_n623), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n505), .A2(new_n507), .A3(new_n510), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n495), .A2(KEYINPUT71), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n493), .A2(G114), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n492), .B1(new_n844), .B2(G2105), .ZN(new_n845));
  AOI211_X1 g420(.A(KEYINPUT72), .B(new_n462), .C1(new_n842), .C2(new_n843), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n500), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(new_n502), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n498), .A2(KEYINPUT73), .A3(new_n500), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n841), .A2(new_n850), .ZN(new_n851));
  XNOR2_X1  g426(.A(new_n699), .B(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(new_n792), .ZN(new_n853));
  MUX2_X1   g428(.A(new_n684), .B(new_n682), .S(new_n853), .Z(new_n854));
  XNOR2_X1  g429(.A(new_n840), .B(new_n854), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT104), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g432(.A(new_n620), .B(G160), .ZN(new_n858));
  XNOR2_X1  g433(.A(new_n858), .B(G162), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AND2_X1   g435(.A1(new_n840), .A2(new_n854), .ZN(new_n861));
  OAI211_X1 g436(.A(new_n857), .B(new_n860), .C1(new_n856), .C2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G37), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n855), .A2(new_n859), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n862), .A2(new_n863), .A3(new_n864), .ZN(new_n865));
  XNOR2_X1  g440(.A(new_n865), .B(KEYINPUT40), .ZN(G395));
  NAND3_X1  g441(.A1(new_n600), .A2(new_n573), .A3(new_n567), .ZN(new_n867));
  INV_X1    g442(.A(KEYINPUT105), .ZN(new_n868));
  NOR2_X1   g443(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g444(.A1(G299), .A2(new_n609), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n867), .ZN(new_n871));
  INV_X1    g446(.A(new_n871), .ZN(new_n872));
  AOI21_X1  g447(.A(new_n869), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  INV_X1    g448(.A(new_n873), .ZN(new_n874));
  OR2_X1    g449(.A1(new_n874), .A2(KEYINPUT41), .ZN(new_n875));
  NAND2_X1  g450(.A1(new_n872), .A2(KEYINPUT41), .ZN(new_n876));
  NAND2_X1  g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  XNOR2_X1  g452(.A(new_n819), .B(new_n613), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI21_X1  g454(.A(new_n879), .B1(new_n878), .B2(new_n872), .ZN(new_n880));
  OR2_X1    g455(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n881));
  XNOR2_X1  g456(.A(G303), .B(G305), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n731), .B(new_n591), .ZN(new_n883));
  INV_X1    g458(.A(KEYINPUT106), .ZN(new_n884));
  OAI21_X1  g459(.A(new_n882), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n883), .A2(new_n884), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n885), .B(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n880), .A2(KEYINPUT42), .ZN(new_n888));
  AND3_X1   g463(.A1(new_n881), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n887), .B1(new_n881), .B2(new_n888), .ZN(new_n890));
  OAI21_X1  g465(.A(G868), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n601), .B1(new_n809), .B2(new_n812), .ZN(new_n892));
  NAND2_X1  g467(.A1(new_n891), .A2(new_n892), .ZN(G295));
  INV_X1    g468(.A(KEYINPUT107), .ZN(new_n894));
  XNOR2_X1  g469(.A(G295), .B(new_n894), .ZN(G331));
  INV_X1    g470(.A(KEYINPUT109), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n887), .B(KEYINPUT108), .Z(new_n897));
  XNOR2_X1  g472(.A(G301), .B(G286), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n819), .B(new_n898), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n899), .A2(new_n876), .A3(new_n875), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n900), .B1(new_n871), .B2(new_n899), .ZN(new_n901));
  OR2_X1    g476(.A1(new_n897), .A2(new_n901), .ZN(new_n902));
  AOI21_X1  g477(.A(G37), .B1(new_n901), .B2(new_n887), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n896), .B1(new_n904), .B2(KEYINPUT43), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n899), .A2(KEYINPUT41), .A3(new_n873), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n871), .B1(new_n899), .B2(KEYINPUT41), .ZN(new_n907));
  OR3_X1    g482(.A1(new_n897), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n903), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(KEYINPUT43), .ZN(new_n910));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND4_X1  g486(.A1(new_n902), .A2(new_n903), .A3(KEYINPUT109), .A4(new_n911), .ZN(new_n912));
  NAND4_X1  g487(.A1(new_n905), .A2(new_n910), .A3(KEYINPUT44), .A4(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n908), .A2(new_n903), .A3(new_n911), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n914), .A2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n913), .B1(KEYINPUT44), .B2(new_n916), .ZN(G397));
  INV_X1    g492(.A(G1384), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n918), .B1(new_n504), .B2(new_n511), .ZN(new_n919));
  INV_X1    g494(.A(KEYINPUT45), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  INV_X1    g496(.A(new_n921), .ZN(new_n922));
  AND2_X1   g497(.A1(G160), .A2(G40), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(new_n924), .ZN(new_n925));
  INV_X1    g500(.A(G1996), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT46), .ZN(new_n928));
  NAND2_X1  g503(.A1(new_n928), .A2(KEYINPUT125), .ZN(new_n929));
  XNOR2_X1  g504(.A(new_n927), .B(new_n929), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n699), .B(new_n703), .ZN(new_n931));
  AND2_X1   g506(.A1(new_n931), .A2(new_n793), .ZN(new_n932));
  OAI221_X1 g507(.A(new_n930), .B1(KEYINPUT125), .B2(new_n928), .C1(new_n924), .C2(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(KEYINPUT47), .ZN(new_n934));
  NAND3_X1  g509(.A1(new_n925), .A2(G1996), .A3(new_n792), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n935), .B(KEYINPUT110), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n931), .B1(G1996), .B2(new_n792), .ZN(new_n937));
  AOI21_X1  g512(.A(new_n936), .B1(new_n925), .B2(new_n937), .ZN(new_n938));
  XOR2_X1   g513(.A(new_n760), .B(new_n763), .Z(new_n939));
  OAI21_X1  g514(.A(new_n938), .B1(new_n924), .B2(new_n939), .ZN(new_n940));
  NOR3_X1   g515(.A1(new_n924), .A2(G1986), .A3(G290), .ZN(new_n941));
  XOR2_X1   g516(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n942));
  XNOR2_X1  g517(.A(new_n941), .B(new_n942), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n940), .A2(new_n943), .ZN(new_n944));
  NOR2_X1   g519(.A1(new_n760), .A2(new_n763), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n938), .A2(new_n945), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n700), .A2(new_n703), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n924), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  INV_X1    g524(.A(KEYINPUT124), .ZN(new_n950));
  INV_X1    g525(.A(new_n919), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(new_n923), .A3(new_n703), .ZN(new_n952));
  NAND2_X1  g527(.A1(G160), .A2(G40), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT50), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n919), .A2(new_n954), .ZN(new_n955));
  OAI211_X1 g530(.A(KEYINPUT50), .B(new_n918), .C1(new_n504), .C2(new_n511), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n953), .B1(new_n955), .B2(new_n956), .ZN(new_n957));
  OAI21_X1  g532(.A(new_n952), .B1(new_n957), .B2(G1348), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n958), .A2(KEYINPUT116), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT116), .ZN(new_n960));
  OAI211_X1 g535(.A(new_n960), .B(new_n952), .C1(new_n957), .C2(G1348), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT60), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n600), .B1(new_n962), .B2(KEYINPUT60), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n964), .B(new_n609), .C1(new_n959), .C2(new_n961), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n965), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT61), .ZN(new_n969));
  NAND3_X1  g544(.A1(G299), .A2(KEYINPUT115), .A3(KEYINPUT57), .ZN(new_n970));
  NAND2_X1  g545(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n971));
  OR2_X1    g546(.A1(KEYINPUT115), .A2(KEYINPUT57), .ZN(new_n972));
  NAND4_X1  g547(.A1(new_n567), .A2(new_n573), .A3(new_n971), .A4(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n970), .A2(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT50), .B1(new_n851), .B2(new_n918), .ZN(new_n976));
  INV_X1    g551(.A(new_n956), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n923), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n978), .A2(new_n713), .ZN(new_n979));
  OAI211_X1 g554(.A(KEYINPUT45), .B(new_n918), .C1(new_n504), .C2(new_n511), .ZN(new_n980));
  XNOR2_X1  g555(.A(KEYINPUT56), .B(G2072), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n921), .A2(new_n923), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI21_X1  g557(.A(new_n975), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  OAI211_X1 g558(.A(new_n975), .B(new_n982), .C1(new_n957), .C2(G1956), .ZN(new_n984));
  INV_X1    g559(.A(new_n984), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n969), .B1(new_n983), .B2(new_n985), .ZN(new_n986));
  OAI21_X1  g561(.A(new_n982), .B1(new_n957), .B2(G1956), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(new_n974), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n988), .A2(KEYINPUT61), .A3(new_n984), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT117), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n990), .A2(KEYINPUT59), .ZN(new_n991));
  XNOR2_X1  g566(.A(new_n991), .B(KEYINPUT118), .ZN(new_n992));
  NAND4_X1  g567(.A1(new_n921), .A2(new_n923), .A3(new_n926), .A4(new_n980), .ZN(new_n993));
  XOR2_X1   g568(.A(KEYINPUT58), .B(G1341), .Z(new_n994));
  OAI21_X1  g569(.A(new_n994), .B1(new_n953), .B2(new_n919), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n992), .B1(new_n996), .B2(new_n559), .ZN(new_n997));
  INV_X1    g572(.A(new_n992), .ZN(new_n998));
  AOI211_X1 g573(.A(new_n558), .B(new_n998), .C1(new_n993), .C2(new_n995), .ZN(new_n999));
  NOR2_X1   g574(.A1(new_n997), .A2(new_n999), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n986), .A2(new_n989), .A3(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT119), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT119), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n986), .A2(new_n1000), .A3(new_n989), .A4(new_n1003), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n968), .A2(new_n1002), .A3(new_n1004), .ZN(new_n1005));
  NOR2_X1   g580(.A1(new_n985), .A2(new_n600), .ZN(new_n1006));
  AOI21_X1  g581(.A(new_n983), .B1(new_n963), .B2(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1008), .A2(KEYINPUT120), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT123), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G286), .A2(G8), .ZN(new_n1011));
  INV_X1    g586(.A(KEYINPUT121), .ZN(new_n1012));
  INV_X1    g587(.A(G2084), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n921), .A2(new_n923), .A3(new_n980), .ZN(new_n1014));
  AOI22_X1  g589(.A1(new_n1013), .A2(new_n957), .B1(new_n1014), .B2(new_n782), .ZN(new_n1015));
  INV_X1    g590(.A(G8), .ZN(new_n1016));
  OAI221_X1 g591(.A(new_n1011), .B1(new_n1012), .B2(KEYINPUT51), .C1(new_n1015), .C2(new_n1016), .ZN(new_n1017));
  AOI21_X1  g592(.A(KEYINPUT51), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1014), .A2(new_n782), .ZN(new_n1019));
  OAI21_X1  g594(.A(new_n1019), .B1(G2084), .B2(new_n978), .ZN(new_n1020));
  OAI211_X1 g595(.A(G8), .B(new_n1018), .C1(new_n1020), .C2(G286), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(G8), .A3(G286), .ZN(new_n1022));
  NAND3_X1  g597(.A1(new_n1017), .A2(new_n1021), .A3(new_n1022), .ZN(new_n1023));
  INV_X1    g598(.A(G2078), .ZN(new_n1024));
  NAND4_X1  g599(.A1(new_n921), .A2(new_n923), .A3(new_n1024), .A4(new_n980), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  AOI22_X1  g601(.A1(new_n978), .A2(new_n717), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT122), .ZN(new_n1028));
  AND2_X1   g603(.A1(new_n1025), .A2(new_n1028), .ZN(new_n1029));
  OAI21_X1  g604(.A(KEYINPUT53), .B1(new_n1025), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(G301), .B(KEYINPUT54), .Z(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  AND2_X1   g609(.A1(new_n1023), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n957), .A2(new_n1036), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1037), .A2(KEYINPUT111), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1014), .A2(new_n741), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT111), .ZN(new_n1040));
  NAND3_X1  g615(.A1(new_n957), .A2(new_n1040), .A3(new_n1036), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1038), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  NAND2_X1  g617(.A1(G303), .A2(G8), .ZN(new_n1043));
  XOR2_X1   g618(.A(new_n1043), .B(KEYINPUT55), .Z(new_n1044));
  XNOR2_X1  g619(.A(new_n1044), .B(KEYINPUT112), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1042), .A2(G8), .A3(new_n1045), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1016), .B1(new_n951), .B2(new_n923), .ZN(new_n1047));
  XNOR2_X1  g622(.A(G305), .B(KEYINPUT49), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n582), .A2(KEYINPUT113), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(G1981), .ZN(new_n1050));
  OR2_X1    g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1047), .A2(new_n1051), .A3(new_n1052), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n731), .A2(G1976), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1054), .B(G8), .C1(new_n953), .C2(new_n919), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1055), .A2(KEYINPUT52), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n951), .A2(new_n923), .ZN(new_n1057));
  INV_X1    g632(.A(G1976), .ZN(new_n1058));
  AOI21_X1  g633(.A(KEYINPUT52), .B1(G288), .B2(new_n1058), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1057), .A2(G8), .A3(new_n1054), .A4(new_n1059), .ZN(new_n1060));
  NAND3_X1  g635(.A1(new_n1053), .A2(new_n1056), .A3(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(KEYINPUT114), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NAND4_X1  g638(.A1(new_n1053), .A2(new_n1056), .A3(new_n1060), .A4(KEYINPUT114), .ZN(new_n1064));
  NAND2_X1  g639(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g640(.A(new_n1044), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1037), .A2(new_n1039), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1066), .B1(new_n1067), .B2(new_n1016), .ZN(new_n1068));
  OAI211_X1 g643(.A(new_n1027), .B(new_n1032), .C1(new_n1026), .C2(new_n1025), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1046), .A2(new_n1065), .A3(new_n1068), .A4(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1010), .B1(new_n1035), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1023), .A2(new_n1034), .ZN(new_n1073));
  NOR3_X1   g648(.A1(new_n1073), .A2(new_n1070), .A3(KEYINPUT123), .ZN(new_n1074));
  NOR2_X1   g649(.A1(new_n1072), .A2(new_n1074), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT120), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1005), .A2(new_n1076), .A3(new_n1007), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1009), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  OR2_X1    g653(.A1(new_n1046), .A2(new_n1061), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1053), .A2(new_n1058), .ZN(new_n1080));
  OAI22_X1  g655(.A1(new_n1080), .A2(G288), .B1(G1981), .B2(G305), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1081), .A2(new_n1047), .ZN(new_n1082));
  NOR3_X1   g657(.A1(new_n1015), .A2(new_n1016), .A3(G286), .ZN(new_n1083));
  NAND2_X1  g658(.A1(new_n1046), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g659(.A(new_n1044), .B1(new_n1042), .B2(G8), .ZN(new_n1085));
  NOR3_X1   g660(.A1(new_n1084), .A2(new_n1061), .A3(new_n1085), .ZN(new_n1086));
  INV_X1    g661(.A(KEYINPUT63), .ZN(new_n1087));
  OAI211_X1 g662(.A(new_n1079), .B(new_n1082), .C1(new_n1086), .C2(new_n1087), .ZN(new_n1088));
  NAND2_X1  g663(.A1(new_n1023), .A2(KEYINPUT62), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT62), .ZN(new_n1090));
  NAND4_X1  g665(.A1(new_n1017), .A2(new_n1021), .A3(new_n1090), .A4(new_n1022), .ZN(new_n1091));
  NAND4_X1  g666(.A1(new_n1089), .A2(G171), .A3(new_n1091), .A4(new_n1031), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1083), .ZN(new_n1093));
  OAI21_X1  g668(.A(new_n1092), .B1(KEYINPUT63), .B2(new_n1093), .ZN(new_n1094));
  AND3_X1   g669(.A1(new_n1046), .A2(new_n1065), .A3(new_n1068), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n1088), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n1078), .A2(new_n1096), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n591), .B(G1986), .ZN(new_n1098));
  NOR2_X1   g673(.A1(new_n924), .A2(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n940), .A2(new_n1099), .ZN(new_n1100));
  AOI21_X1  g675(.A(new_n950), .B1(new_n1097), .B2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(new_n1100), .ZN(new_n1102));
  AOI211_X1 g677(.A(KEYINPUT124), .B(new_n1102), .C1(new_n1078), .C2(new_n1096), .ZN(new_n1103));
  OAI211_X1 g678(.A(new_n934), .B(new_n949), .C1(new_n1101), .C2(new_n1103), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g679(.A(new_n460), .B(G229), .C1(new_n914), .C2(new_n915), .ZN(new_n1106));
  NOR2_X1   g680(.A1(G401), .A2(G227), .ZN(new_n1107));
  NAND3_X1  g681(.A1(new_n1106), .A2(new_n865), .A3(new_n1107), .ZN(G225));
  INV_X1    g682(.A(G225), .ZN(G308));
endmodule


