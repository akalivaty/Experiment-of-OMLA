

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588;

  XNOR2_X1 U326 ( .A(n302), .B(n301), .ZN(n303) );
  NOR2_X1 U327 ( .A1(n536), .A2(n479), .ZN(n571) );
  XNOR2_X1 U328 ( .A(n473), .B(n472), .ZN(n552) );
  XNOR2_X1 U329 ( .A(n312), .B(n400), .ZN(n536) );
  XOR2_X1 U330 ( .A(n328), .B(n327), .Z(n294) );
  XOR2_X1 U331 ( .A(G15GAT), .B(G127GAT), .Z(n370) );
  INV_X1 U332 ( .A(KEYINPUT84), .ZN(n301) );
  XNOR2_X1 U333 ( .A(KEYINPUT48), .B(KEYINPUT122), .ZN(n472) );
  NAND2_X1 U334 ( .A1(n454), .A2(n453), .ZN(n488) );
  XNOR2_X1 U335 ( .A(n329), .B(n294), .ZN(n330) );
  NOR2_X1 U336 ( .A1(n586), .A2(n455), .ZN(n456) );
  XNOR2_X1 U337 ( .A(n304), .B(n303), .ZN(n307) );
  XNOR2_X1 U338 ( .A(n331), .B(n330), .ZN(n332) );
  INV_X1 U339 ( .A(G190GAT), .ZN(n480) );
  INV_X1 U340 ( .A(G43GAT), .ZN(n458) );
  XNOR2_X1 U341 ( .A(n457), .B(KEYINPUT38), .ZN(n508) );
  XNOR2_X1 U342 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U343 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U344 ( .A(n483), .B(n482), .ZN(G1351GAT) );
  XNOR2_X1 U345 ( .A(n461), .B(n460), .ZN(G1330GAT) );
  XOR2_X1 U346 ( .A(KEYINPUT20), .B(KEYINPUT83), .Z(n296) );
  XNOR2_X1 U347 ( .A(G113GAT), .B(G183GAT), .ZN(n295) );
  XNOR2_X1 U348 ( .A(n296), .B(n295), .ZN(n300) );
  XOR2_X1 U349 ( .A(KEYINPUT0), .B(n370), .Z(n298) );
  XOR2_X1 U350 ( .A(G190GAT), .B(G134GAT), .Z(n361) );
  XNOR2_X1 U351 ( .A(G43GAT), .B(n361), .ZN(n297) );
  XNOR2_X1 U352 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U353 ( .A(n300), .B(n299), .Z(n304) );
  NAND2_X1 U354 ( .A1(G227GAT), .A2(G233GAT), .ZN(n302) );
  XNOR2_X1 U355 ( .A(G99GAT), .B(G71GAT), .ZN(n305) );
  XNOR2_X1 U356 ( .A(n305), .B(G120GAT), .ZN(n315) );
  XNOR2_X1 U357 ( .A(n315), .B(KEYINPUT86), .ZN(n306) );
  XNOR2_X1 U358 ( .A(n307), .B(n306), .ZN(n312) );
  XOR2_X1 U359 ( .A(KEYINPUT19), .B(G176GAT), .Z(n309) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT18), .ZN(n308) );
  XNOR2_X1 U361 ( .A(n309), .B(n308), .ZN(n311) );
  XOR2_X1 U362 ( .A(KEYINPUT85), .B(KEYINPUT17), .Z(n310) );
  XNOR2_X1 U363 ( .A(n311), .B(n310), .ZN(n400) );
  XOR2_X1 U364 ( .A(G78GAT), .B(G148GAT), .Z(n314) );
  XNOR2_X1 U365 ( .A(G106GAT), .B(KEYINPUT71), .ZN(n313) );
  XNOR2_X1 U366 ( .A(n314), .B(n313), .ZN(n397) );
  XOR2_X1 U367 ( .A(n315), .B(n397), .Z(n333) );
  INV_X1 U368 ( .A(KEYINPUT70), .ZN(n316) );
  NAND2_X1 U369 ( .A1(G64GAT), .A2(n316), .ZN(n319) );
  INV_X1 U370 ( .A(G64GAT), .ZN(n317) );
  NAND2_X1 U371 ( .A1(n317), .A2(KEYINPUT70), .ZN(n318) );
  NAND2_X1 U372 ( .A1(n319), .A2(n318), .ZN(n321) );
  XNOR2_X1 U373 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n320) );
  XNOR2_X1 U374 ( .A(n321), .B(n320), .ZN(n368) );
  XOR2_X1 U375 ( .A(G85GAT), .B(G92GAT), .Z(n354) );
  XOR2_X1 U376 ( .A(n368), .B(n354), .Z(n323) );
  XNOR2_X1 U377 ( .A(G176GAT), .B(G204GAT), .ZN(n322) );
  XNOR2_X1 U378 ( .A(n323), .B(n322), .ZN(n331) );
  XOR2_X1 U379 ( .A(KEYINPUT72), .B(KEYINPUT33), .Z(n325) );
  XNOR2_X1 U380 ( .A(KEYINPUT73), .B(KEYINPUT74), .ZN(n324) );
  XNOR2_X1 U381 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n326), .B(KEYINPUT32), .ZN(n329) );
  XOR2_X1 U383 ( .A(KEYINPUT31), .B(KEYINPUT75), .Z(n328) );
  NAND2_X1 U384 ( .A1(G230GAT), .A2(G233GAT), .ZN(n327) );
  XNOR2_X1 U385 ( .A(n333), .B(n332), .ZN(n579) );
  XNOR2_X1 U386 ( .A(G36GAT), .B(KEYINPUT7), .ZN(n334) );
  XNOR2_X1 U387 ( .A(n334), .B(G29GAT), .ZN(n335) );
  XOR2_X1 U388 ( .A(n335), .B(KEYINPUT8), .Z(n337) );
  XNOR2_X1 U389 ( .A(G43GAT), .B(G50GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n337), .B(n336), .ZN(n353) );
  XOR2_X1 U391 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n339) );
  XNOR2_X1 U392 ( .A(G15GAT), .B(KEYINPUT68), .ZN(n338) );
  XNOR2_X1 U393 ( .A(n339), .B(n338), .ZN(n344) );
  XNOR2_X1 U394 ( .A(G141GAT), .B(G113GAT), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n340), .B(G1GAT), .ZN(n434) );
  XOR2_X1 U396 ( .A(n434), .B(KEYINPUT29), .Z(n342) );
  NAND2_X1 U397 ( .A1(G229GAT), .A2(G233GAT), .ZN(n341) );
  XNOR2_X1 U398 ( .A(n342), .B(n341), .ZN(n343) );
  XNOR2_X1 U399 ( .A(n344), .B(n343), .ZN(n347) );
  XNOR2_X1 U400 ( .A(G169GAT), .B(G22GAT), .ZN(n345) );
  XOR2_X1 U401 ( .A(G197GAT), .B(G8GAT), .Z(n404) );
  XOR2_X1 U402 ( .A(n345), .B(n404), .Z(n346) );
  XNOR2_X1 U403 ( .A(n347), .B(n346), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n353), .B(n348), .ZN(n575) );
  XNOR2_X1 U405 ( .A(n575), .B(KEYINPUT69), .ZN(n564) );
  NAND2_X1 U406 ( .A1(n579), .A2(n564), .ZN(n349) );
  XOR2_X1 U407 ( .A(KEYINPUT76), .B(n349), .Z(n491) );
  XOR2_X1 U408 ( .A(KEYINPUT78), .B(KEYINPUT9), .Z(n351) );
  XNOR2_X1 U409 ( .A(G106GAT), .B(KEYINPUT11), .ZN(n350) );
  XNOR2_X1 U410 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U411 ( .A(n353), .B(n352), .ZN(n365) );
  XOR2_X1 U412 ( .A(KEYINPUT10), .B(n354), .Z(n356) );
  XOR2_X1 U413 ( .A(KEYINPUT77), .B(G162GAT), .Z(n384) );
  XNOR2_X1 U414 ( .A(G218GAT), .B(n384), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U416 ( .A(KEYINPUT79), .B(KEYINPUT65), .Z(n358) );
  NAND2_X1 U417 ( .A1(G232GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U418 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U419 ( .A(n360), .B(n359), .Z(n363) );
  XNOR2_X1 U420 ( .A(G99GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n562) );
  XNOR2_X1 U423 ( .A(KEYINPUT36), .B(n562), .ZN(n586) );
  XOR2_X1 U424 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n367) );
  XNOR2_X1 U425 ( .A(G8GAT), .B(G1GAT), .ZN(n366) );
  XNOR2_X1 U426 ( .A(n367), .B(n366), .ZN(n369) );
  XOR2_X1 U427 ( .A(n369), .B(n368), .Z(n372) );
  XOR2_X1 U428 ( .A(G22GAT), .B(G155GAT), .Z(n383) );
  XNOR2_X1 U429 ( .A(n370), .B(n383), .ZN(n371) );
  XNOR2_X1 U430 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U431 ( .A(G183GAT), .B(G211GAT), .Z(n403) );
  XOR2_X1 U432 ( .A(n373), .B(n403), .Z(n375) );
  XNOR2_X1 U433 ( .A(G71GAT), .B(G78GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n377) );
  NAND2_X1 U436 ( .A1(G231GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U437 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U438 ( .A(KEYINPUT81), .B(n378), .Z(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n582) );
  XOR2_X1 U440 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n382) );
  XNOR2_X1 U441 ( .A(G197GAT), .B(G141GAT), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n388) );
  XOR2_X1 U443 ( .A(G211GAT), .B(n383), .Z(n386) );
  XNOR2_X1 U444 ( .A(G50GAT), .B(n384), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U446 ( .A(n388), .B(n387), .Z(n390) );
  NAND2_X1 U447 ( .A1(G228GAT), .A2(G233GAT), .ZN(n389) );
  XNOR2_X1 U448 ( .A(n390), .B(n389), .ZN(n391) );
  XOR2_X1 U449 ( .A(n391), .B(KEYINPUT23), .Z(n394) );
  XNOR2_X1 U450 ( .A(KEYINPUT2), .B(KEYINPUT3), .ZN(n392) );
  XNOR2_X1 U451 ( .A(n392), .B(KEYINPUT89), .ZN(n433) );
  XNOR2_X1 U452 ( .A(n433), .B(KEYINPUT90), .ZN(n393) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n399) );
  XOR2_X1 U454 ( .A(G204GAT), .B(KEYINPUT21), .Z(n396) );
  XNOR2_X1 U455 ( .A(G218GAT), .B(KEYINPUT88), .ZN(n395) );
  XNOR2_X1 U456 ( .A(n396), .B(n395), .ZN(n412) );
  XOR2_X1 U457 ( .A(n412), .B(n397), .Z(n398) );
  XNOR2_X1 U458 ( .A(n399), .B(n398), .ZN(n477) );
  INV_X1 U459 ( .A(n400), .ZN(n416) );
  XOR2_X1 U460 ( .A(KEYINPUT98), .B(KEYINPUT95), .Z(n402) );
  XNOR2_X1 U461 ( .A(G92GAT), .B(G64GAT), .ZN(n401) );
  XNOR2_X1 U462 ( .A(n402), .B(n401), .ZN(n408) );
  XOR2_X1 U463 ( .A(n403), .B(G190GAT), .Z(n406) );
  XNOR2_X1 U464 ( .A(G36GAT), .B(n404), .ZN(n405) );
  XNOR2_X1 U465 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U466 ( .A(n408), .B(n407), .Z(n410) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U468 ( .A(n410), .B(n409), .ZN(n411) );
  XOR2_X1 U469 ( .A(n411), .B(KEYINPUT96), .Z(n414) );
  XNOR2_X1 U470 ( .A(n412), .B(KEYINPUT97), .ZN(n413) );
  XNOR2_X1 U471 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U472 ( .A(n416), .B(n415), .ZN(n526) );
  NOR2_X1 U473 ( .A1(n536), .A2(n526), .ZN(n417) );
  XNOR2_X1 U474 ( .A(n417), .B(KEYINPUT102), .ZN(n418) );
  NOR2_X1 U475 ( .A1(n477), .A2(n418), .ZN(n419) );
  XNOR2_X1 U476 ( .A(KEYINPUT25), .B(n419), .ZN(n424) );
  NAND2_X1 U477 ( .A1(n477), .A2(n536), .ZN(n420) );
  XNOR2_X1 U478 ( .A(n420), .B(KEYINPUT26), .ZN(n573) );
  XNOR2_X1 U479 ( .A(KEYINPUT27), .B(KEYINPUT99), .ZN(n421) );
  XNOR2_X1 U480 ( .A(n421), .B(n526), .ZN(n449) );
  INV_X1 U481 ( .A(n449), .ZN(n422) );
  NOR2_X1 U482 ( .A1(n573), .A2(n422), .ZN(n554) );
  XNOR2_X1 U483 ( .A(n554), .B(KEYINPUT101), .ZN(n423) );
  NAND2_X1 U484 ( .A1(n424), .A2(n423), .ZN(n447) );
  XOR2_X1 U485 ( .A(KEYINPUT91), .B(KEYINPUT1), .Z(n426) );
  XNOR2_X1 U486 ( .A(KEYINPUT4), .B(KEYINPUT94), .ZN(n425) );
  XNOR2_X1 U487 ( .A(n426), .B(n425), .ZN(n438) );
  XOR2_X1 U488 ( .A(KEYINPUT92), .B(KEYINPUT0), .Z(n428) );
  XNOR2_X1 U489 ( .A(G120GAT), .B(G127GAT), .ZN(n427) );
  XNOR2_X1 U490 ( .A(n428), .B(n427), .ZN(n432) );
  XOR2_X1 U491 ( .A(G57GAT), .B(KEYINPUT5), .Z(n430) );
  XNOR2_X1 U492 ( .A(KEYINPUT93), .B(KEYINPUT6), .ZN(n429) );
  XNOR2_X1 U493 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U494 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U496 ( .A(n436), .B(n435), .ZN(n437) );
  XNOR2_X1 U497 ( .A(n438), .B(n437), .ZN(n446) );
  NAND2_X1 U498 ( .A1(G225GAT), .A2(G233GAT), .ZN(n444) );
  XOR2_X1 U499 ( .A(G85GAT), .B(G155GAT), .Z(n440) );
  XNOR2_X1 U500 ( .A(G148GAT), .B(G162GAT), .ZN(n439) );
  XNOR2_X1 U501 ( .A(n440), .B(n439), .ZN(n442) );
  XOR2_X1 U502 ( .A(G29GAT), .B(G134GAT), .Z(n441) );
  XNOR2_X1 U503 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U504 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(n551) );
  NAND2_X1 U506 ( .A1(n447), .A2(n551), .ZN(n454) );
  XOR2_X1 U507 ( .A(n536), .B(KEYINPUT87), .Z(n452) );
  XOR2_X1 U508 ( .A(KEYINPUT28), .B(KEYINPUT66), .Z(n448) );
  XNOR2_X1 U509 ( .A(n477), .B(n448), .ZN(n533) );
  NAND2_X1 U510 ( .A1(n533), .A2(n449), .ZN(n450) );
  NOR2_X1 U511 ( .A1(n551), .A2(n450), .ZN(n538) );
  XNOR2_X1 U512 ( .A(KEYINPUT100), .B(n538), .ZN(n451) );
  NAND2_X1 U513 ( .A1(n452), .A2(n451), .ZN(n453) );
  NAND2_X1 U514 ( .A1(n582), .A2(n488), .ZN(n455) );
  XOR2_X1 U515 ( .A(KEYINPUT37), .B(n456), .Z(n524) );
  NAND2_X1 U516 ( .A1(n491), .A2(n524), .ZN(n457) );
  NOR2_X1 U517 ( .A1(n536), .A2(n508), .ZN(n461) );
  XNOR2_X1 U518 ( .A(KEYINPUT40), .B(KEYINPUT112), .ZN(n459) );
  XNOR2_X1 U519 ( .A(n579), .B(KEYINPUT41), .ZN(n566) );
  INV_X1 U520 ( .A(n566), .ZN(n556) );
  NOR2_X1 U521 ( .A1(n556), .A2(n575), .ZN(n462) );
  XNOR2_X1 U522 ( .A(n462), .B(KEYINPUT46), .ZN(n465) );
  XNOR2_X1 U523 ( .A(KEYINPUT121), .B(n582), .ZN(n570) );
  INV_X1 U524 ( .A(n570), .ZN(n463) );
  NAND2_X1 U525 ( .A1(n562), .A2(n463), .ZN(n464) );
  OR2_X1 U526 ( .A1(n465), .A2(n464), .ZN(n466) );
  XNOR2_X1 U527 ( .A(n466), .B(KEYINPUT47), .ZN(n471) );
  NOR2_X1 U528 ( .A1(n586), .A2(n582), .ZN(n467) );
  XNOR2_X1 U529 ( .A(n467), .B(KEYINPUT45), .ZN(n468) );
  NAND2_X1 U530 ( .A1(n468), .A2(n579), .ZN(n469) );
  NOR2_X1 U531 ( .A1(n564), .A2(n469), .ZN(n470) );
  NOR2_X1 U532 ( .A1(n471), .A2(n470), .ZN(n473) );
  NOR2_X1 U533 ( .A1(n552), .A2(n526), .ZN(n474) );
  XNOR2_X1 U534 ( .A(n474), .B(KEYINPUT54), .ZN(n475) );
  NAND2_X1 U535 ( .A1(n475), .A2(n551), .ZN(n476) );
  XNOR2_X1 U536 ( .A(n476), .B(KEYINPUT64), .ZN(n574) );
  NOR2_X1 U537 ( .A1(n574), .A2(n477), .ZN(n478) );
  XNOR2_X1 U538 ( .A(n478), .B(KEYINPUT55), .ZN(n479) );
  INV_X1 U539 ( .A(n562), .ZN(n547) );
  NAND2_X1 U540 ( .A1(n571), .A2(n547), .ZN(n483) );
  XOR2_X1 U541 ( .A(KEYINPUT126), .B(KEYINPUT58), .Z(n481) );
  XOR2_X1 U542 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n485) );
  XNOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n484) );
  XNOR2_X1 U544 ( .A(n485), .B(n484), .ZN(n494) );
  NOR2_X1 U545 ( .A1(n547), .A2(n582), .ZN(n487) );
  XNOR2_X1 U546 ( .A(KEYINPUT16), .B(KEYINPUT82), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n487), .B(n486), .ZN(n489) );
  NAND2_X1 U548 ( .A1(n489), .A2(n488), .ZN(n490) );
  XNOR2_X1 U549 ( .A(KEYINPUT103), .B(n490), .ZN(n511) );
  NAND2_X1 U550 ( .A1(n511), .A2(n491), .ZN(n492) );
  XNOR2_X1 U551 ( .A(KEYINPUT104), .B(n492), .ZN(n501) );
  NOR2_X1 U552 ( .A1(n501), .A2(n551), .ZN(n493) );
  XOR2_X1 U553 ( .A(n494), .B(n493), .Z(G1324GAT) );
  NOR2_X1 U554 ( .A1(n501), .A2(n526), .ZN(n496) );
  XNOR2_X1 U555 ( .A(G8GAT), .B(KEYINPUT107), .ZN(n495) );
  XNOR2_X1 U556 ( .A(n496), .B(n495), .ZN(G1325GAT) );
  NOR2_X1 U557 ( .A1(n501), .A2(n536), .ZN(n500) );
  XOR2_X1 U558 ( .A(KEYINPUT108), .B(KEYINPUT109), .Z(n498) );
  XNOR2_X1 U559 ( .A(G15GAT), .B(KEYINPUT35), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(G1326GAT) );
  NOR2_X1 U562 ( .A1(n533), .A2(n501), .ZN(n502) );
  XOR2_X1 U563 ( .A(G22GAT), .B(n502), .Z(G1327GAT) );
  NOR2_X1 U564 ( .A1(n508), .A2(n551), .ZN(n504) );
  XNOR2_X1 U565 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1328GAT) );
  NOR2_X1 U567 ( .A1(n508), .A2(n526), .ZN(n506) );
  XNOR2_X1 U568 ( .A(KEYINPUT110), .B(KEYINPUT111), .ZN(n505) );
  XNOR2_X1 U569 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U570 ( .A(G36GAT), .B(n507), .ZN(G1329GAT) );
  XNOR2_X1 U571 ( .A(G50GAT), .B(KEYINPUT113), .ZN(n510) );
  NOR2_X1 U572 ( .A1(n533), .A2(n508), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n510), .B(n509), .ZN(G1331GAT) );
  AND2_X1 U574 ( .A1(n575), .A2(n566), .ZN(n523) );
  NAND2_X1 U575 ( .A1(n511), .A2(n523), .ZN(n519) );
  NOR2_X1 U576 ( .A1(n551), .A2(n519), .ZN(n512) );
  XOR2_X1 U577 ( .A(G57GAT), .B(n512), .Z(n513) );
  XNOR2_X1 U578 ( .A(KEYINPUT42), .B(n513), .ZN(G1332GAT) );
  NOR2_X1 U579 ( .A1(n526), .A2(n519), .ZN(n514) );
  XOR2_X1 U580 ( .A(G64GAT), .B(n514), .Z(G1333GAT) );
  NOR2_X1 U581 ( .A1(n536), .A2(n519), .ZN(n515) );
  XOR2_X1 U582 ( .A(KEYINPUT114), .B(n515), .Z(n516) );
  XNOR2_X1 U583 ( .A(G71GAT), .B(n516), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT117), .B(KEYINPUT116), .Z(n518) );
  XNOR2_X1 U585 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n521) );
  NOR2_X1 U587 ( .A1(n533), .A2(n519), .ZN(n520) );
  XOR2_X1 U588 ( .A(n521), .B(n520), .Z(n522) );
  XNOR2_X1 U589 ( .A(KEYINPUT115), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n523), .ZN(n532) );
  NOR2_X1 U591 ( .A1(n551), .A2(n532), .ZN(n525) );
  XOR2_X1 U592 ( .A(G85GAT), .B(n525), .Z(G1336GAT) );
  NOR2_X1 U593 ( .A1(n526), .A2(n532), .ZN(n528) );
  XNOR2_X1 U594 ( .A(KEYINPUT118), .B(KEYINPUT119), .ZN(n527) );
  XNOR2_X1 U595 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U596 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NOR2_X1 U597 ( .A1(n536), .A2(n532), .ZN(n530) );
  XOR2_X1 U598 ( .A(KEYINPUT120), .B(n530), .Z(n531) );
  XNOR2_X1 U599 ( .A(G99GAT), .B(n531), .ZN(G1338GAT) );
  NOR2_X1 U600 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT44), .B(n534), .Z(n535) );
  XNOR2_X1 U602 ( .A(G106GAT), .B(n535), .ZN(G1339GAT) );
  NOR2_X1 U603 ( .A1(n536), .A2(n552), .ZN(n537) );
  NAND2_X1 U604 ( .A1(n538), .A2(n537), .ZN(n539) );
  XNOR2_X1 U605 ( .A(KEYINPUT123), .B(n539), .ZN(n548) );
  NAND2_X1 U606 ( .A1(n564), .A2(n548), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n540), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U608 ( .A(KEYINPUT124), .B(KEYINPUT49), .Z(n542) );
  NAND2_X1 U609 ( .A1(n548), .A2(n566), .ZN(n541) );
  XNOR2_X1 U610 ( .A(n542), .B(n541), .ZN(n543) );
  XNOR2_X1 U611 ( .A(G120GAT), .B(n543), .ZN(G1341GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT50), .B(KEYINPUT125), .Z(n545) );
  NAND2_X1 U613 ( .A1(n548), .A2(n570), .ZN(n544) );
  XNOR2_X1 U614 ( .A(n545), .B(n544), .ZN(n546) );
  XNOR2_X1 U615 ( .A(G127GAT), .B(n546), .ZN(G1342GAT) );
  XOR2_X1 U616 ( .A(G134GAT), .B(KEYINPUT51), .Z(n550) );
  NAND2_X1 U617 ( .A1(n548), .A2(n547), .ZN(n549) );
  XNOR2_X1 U618 ( .A(n550), .B(n549), .ZN(G1343GAT) );
  NOR2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n554), .A2(n553), .ZN(n561) );
  NOR2_X1 U621 ( .A1(n575), .A2(n561), .ZN(n555) );
  XOR2_X1 U622 ( .A(G141GAT), .B(n555), .Z(G1344GAT) );
  NOR2_X1 U623 ( .A1(n556), .A2(n561), .ZN(n558) );
  XNOR2_X1 U624 ( .A(KEYINPUT53), .B(KEYINPUT52), .ZN(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(n559) );
  XNOR2_X1 U626 ( .A(G148GAT), .B(n559), .ZN(G1345GAT) );
  NOR2_X1 U627 ( .A1(n582), .A2(n561), .ZN(n560) );
  XOR2_X1 U628 ( .A(G155GAT), .B(n560), .Z(G1346GAT) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XOR2_X1 U630 ( .A(G162GAT), .B(n563), .Z(G1347GAT) );
  NAND2_X1 U631 ( .A1(n564), .A2(n571), .ZN(n565) );
  XNOR2_X1 U632 ( .A(n565), .B(G169GAT), .ZN(G1348GAT) );
  XOR2_X1 U633 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n568) );
  NAND2_X1 U634 ( .A1(n571), .A2(n566), .ZN(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(n569) );
  XNOR2_X1 U636 ( .A(G176GAT), .B(n569), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n571), .A2(n570), .ZN(n572) );
  XNOR2_X1 U638 ( .A(n572), .B(G183GAT), .ZN(G1350GAT) );
  OR2_X1 U639 ( .A1(n574), .A2(n573), .ZN(n585) );
  NOR2_X1 U640 ( .A1(n575), .A2(n585), .ZN(n577) );
  XNOR2_X1 U641 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n576) );
  XNOR2_X1 U642 ( .A(n577), .B(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(G197GAT), .B(n578), .ZN(G1352GAT) );
  NOR2_X1 U644 ( .A1(n579), .A2(n585), .ZN(n581) );
  XNOR2_X1 U645 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n580) );
  XNOR2_X1 U646 ( .A(n581), .B(n580), .ZN(G1353GAT) );
  NOR2_X1 U647 ( .A1(n582), .A2(n585), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G211GAT), .B(KEYINPUT127), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(G1354GAT) );
  NOR2_X1 U650 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT62), .B(n587), .Z(n588) );
  XNOR2_X1 U652 ( .A(G218GAT), .B(n588), .ZN(G1355GAT) );
endmodule

