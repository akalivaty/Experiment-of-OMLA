//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 0 0 0 0 1 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 1 1 0 0 1 1 0 1 1 1 0 0 1 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 0 1 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:52 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n767, new_n768, new_n769, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n801, new_n802, new_n803,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n811, new_n812,
    new_n813, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n823, new_n824, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n857, new_n858, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n956, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n987, new_n988, new_n989, new_n990, new_n991, new_n992,
    new_n993, new_n994, new_n995, new_n996, new_n997, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1012, new_n1013;
  XOR2_X1   g000(.A(G78gat), .B(G106gat), .Z(new_n202));
  XNOR2_X1  g001(.A(KEYINPUT31), .B(G50gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G22gat), .ZN(new_n205));
  INV_X1    g004(.A(G228gat), .ZN(new_n206));
  INV_X1    g005(.A(G233gat), .ZN(new_n207));
  NOR2_X1   g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  XNOR2_X1  g007(.A(G197gat), .B(G204gat), .ZN(new_n209));
  INV_X1    g008(.A(G211gat), .ZN(new_n210));
  INV_X1    g009(.A(G218gat), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT74), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n213), .A2(G218gat), .ZN(new_n214));
  AOI21_X1  g013(.A(new_n210), .B1(new_n212), .B2(new_n214), .ZN(new_n215));
  OAI21_X1  g014(.A(new_n209), .B1(new_n215), .B2(KEYINPUT22), .ZN(new_n216));
  XNOR2_X1  g015(.A(G211gat), .B(G218gat), .ZN(new_n217));
  AND3_X1   g016(.A1(new_n216), .A2(KEYINPUT75), .A3(new_n217), .ZN(new_n218));
  AOI21_X1  g017(.A(new_n217), .B1(new_n216), .B2(KEYINPUT75), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT29), .ZN(new_n221));
  AOI21_X1  g020(.A(KEYINPUT3), .B1(new_n220), .B2(new_n221), .ZN(new_n222));
  AND2_X1   g021(.A1(G155gat), .A2(G162gat), .ZN(new_n223));
  NOR2_X1   g022(.A1(G155gat), .A2(G162gat), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  XNOR2_X1  g024(.A(G141gat), .B(G148gat), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(G155gat), .ZN(new_n228));
  INV_X1    g027(.A(G162gat), .ZN(new_n229));
  OAI21_X1  g028(.A(KEYINPUT2), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  OR2_X1    g029(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n231));
  INV_X1    g030(.A(G141gat), .ZN(new_n232));
  INV_X1    g031(.A(G148gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  NAND2_X1  g033(.A1(G141gat), .A2(G148gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n231), .A2(new_n234), .A3(new_n235), .A4(new_n236), .ZN(new_n237));
  AOI22_X1  g036(.A1(new_n227), .A2(new_n230), .B1(new_n225), .B2(new_n237), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n208), .B1(new_n222), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n237), .A2(new_n225), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT3), .ZN(new_n241));
  AND2_X1   g040(.A1(G141gat), .A2(G148gat), .ZN(new_n242));
  NOR2_X1   g041(.A1(G141gat), .A2(G148gat), .ZN(new_n243));
  NOR2_X1   g042(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G155gat), .B(G162gat), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n244), .A2(new_n245), .A3(new_n230), .ZN(new_n246));
  NAND3_X1  g045(.A1(new_n240), .A2(new_n241), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n247), .A2(new_n221), .ZN(new_n248));
  OAI211_X1 g047(.A(new_n248), .B(KEYINPUT83), .C1(new_n218), .C2(new_n219), .ZN(new_n249));
  INV_X1    g048(.A(new_n249), .ZN(new_n250));
  INV_X1    g049(.A(new_n217), .ZN(new_n251));
  XOR2_X1   g050(.A(G197gat), .B(G204gat), .Z(new_n252));
  NOR2_X1   g051(.A1(new_n213), .A2(G218gat), .ZN(new_n253));
  NOR2_X1   g052(.A1(new_n211), .A2(KEYINPUT74), .ZN(new_n254));
  OAI21_X1  g053(.A(G211gat), .B1(new_n253), .B2(new_n254), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT22), .ZN(new_n256));
  AOI21_X1  g055(.A(new_n252), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT75), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n251), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n216), .A2(KEYINPUT75), .A3(new_n217), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(KEYINPUT83), .B1(new_n261), .B2(new_n248), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n250), .A2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT84), .B1(new_n239), .B2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(new_n262), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n265), .A2(new_n249), .ZN(new_n266));
  INV_X1    g065(.A(new_n208), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n241), .B1(new_n261), .B2(KEYINPUT29), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n240), .A2(new_n246), .ZN(new_n269));
  AOI21_X1  g068(.A(new_n267), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT84), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n266), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  NOR2_X1   g072(.A1(new_n257), .A2(new_n251), .ZN(new_n274));
  OAI21_X1  g073(.A(new_n221), .B1(new_n216), .B2(new_n217), .ZN(new_n275));
  OAI21_X1  g074(.A(new_n241), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n276), .A2(new_n269), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n248), .ZN(new_n278));
  AOI21_X1  g077(.A(new_n208), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n205), .B1(new_n273), .B2(new_n280), .ZN(new_n281));
  AOI211_X1 g080(.A(G22gat), .B(new_n279), .C1(new_n264), .C2(new_n272), .ZN(new_n282));
  OAI21_X1  g081(.A(new_n204), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(KEYINPUT85), .ZN(new_n284));
  INV_X1    g083(.A(KEYINPUT85), .ZN(new_n285));
  OAI211_X1 g084(.A(new_n285), .B(new_n204), .C1(new_n281), .C2(new_n282), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n281), .A2(new_n287), .ZN(new_n288));
  AOI21_X1  g087(.A(new_n279), .B1(new_n264), .B2(new_n272), .ZN(new_n289));
  OAI21_X1  g088(.A(KEYINPUT86), .B1(new_n289), .B2(new_n205), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n204), .B1(new_n289), .B2(new_n205), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n288), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  NAND3_X1  g091(.A1(new_n284), .A2(new_n286), .A3(new_n292), .ZN(new_n293));
  INV_X1    g092(.A(G127gat), .ZN(new_n294));
  INV_X1    g093(.A(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(G127gat), .A2(G134gat), .ZN(new_n297));
  XNOR2_X1  g096(.A(G113gat), .B(G120gat), .ZN(new_n298));
  OAI211_X1 g097(.A(new_n296), .B(new_n297), .C1(new_n298), .C2(KEYINPUT1), .ZN(new_n299));
  INV_X1    g098(.A(KEYINPUT67), .ZN(new_n300));
  AND2_X1   g099(.A1(G113gat), .A2(G120gat), .ZN(new_n301));
  NOR2_X1   g100(.A1(G113gat), .A2(G120gat), .ZN(new_n302));
  OAI21_X1  g101(.A(new_n300), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(G127gat), .A2(G134gat), .ZN(new_n304));
  NOR2_X1   g103(.A1(G127gat), .A2(G134gat), .ZN(new_n305));
  OAI21_X1  g104(.A(KEYINPUT68), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT68), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n296), .A2(new_n307), .A3(new_n297), .ZN(new_n308));
  NAND3_X1  g107(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  XNOR2_X1  g108(.A(KEYINPUT69), .B(KEYINPUT1), .ZN(new_n310));
  OAI21_X1  g109(.A(new_n310), .B1(new_n298), .B2(new_n300), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n299), .B1(new_n309), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(new_n312), .ZN(new_n313));
  NOR2_X1   g112(.A1(G169gat), .A2(G176gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(KEYINPUT23), .ZN(new_n315));
  NAND2_X1  g114(.A1(G169gat), .A2(G176gat), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT23), .ZN(new_n317));
  OAI21_X1  g116(.A(new_n317), .B1(G169gat), .B2(G176gat), .ZN(new_n318));
  AND4_X1   g117(.A1(KEYINPUT25), .A2(new_n315), .A3(new_n316), .A4(new_n318), .ZN(new_n319));
  NAND2_X1  g118(.A1(G183gat), .A2(G190gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT24), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G183gat), .ZN(new_n323));
  INV_X1    g122(.A(G190gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n322), .A2(new_n325), .A3(new_n326), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n319), .A2(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n326), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT64), .ZN(new_n331));
  AOI21_X1  g130(.A(new_n331), .B1(new_n320), .B2(new_n321), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  AOI21_X1  g132(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n334), .A2(new_n331), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n329), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n328), .B1(new_n336), .B2(KEYINPUT25), .ZN(new_n337));
  INV_X1    g136(.A(G169gat), .ZN(new_n338));
  INV_X1    g137(.A(G176gat), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT26), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT26), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n316), .A2(new_n341), .ZN(new_n342));
  OAI211_X1 g141(.A(new_n320), .B(new_n340), .C1(new_n342), .C2(new_n314), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT66), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  AOI22_X1  g144(.A1(new_n314), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(KEYINPUT66), .C1(new_n314), .C2(new_n342), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT65), .ZN(new_n348));
  INV_X1    g147(.A(KEYINPUT27), .ZN(new_n349));
  NOR2_X1   g148(.A1(new_n349), .A2(G183gat), .ZN(new_n350));
  NOR2_X1   g149(.A1(new_n323), .A2(KEYINPUT27), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n348), .B1(new_n350), .B2(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n323), .A2(KEYINPUT27), .ZN(new_n353));
  AOI21_X1  g152(.A(G190gat), .B1(new_n353), .B2(KEYINPUT65), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT28), .B1(new_n352), .B2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n324), .A2(KEYINPUT28), .ZN(new_n356));
  NOR3_X1   g155(.A1(new_n350), .A2(new_n351), .A3(new_n356), .ZN(new_n357));
  OAI211_X1 g156(.A(new_n345), .B(new_n347), .C1(new_n355), .C2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n313), .B1(new_n337), .B2(new_n358), .ZN(new_n359));
  INV_X1    g158(.A(new_n359), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n337), .A2(new_n358), .A3(new_n313), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(KEYINPUT70), .ZN(new_n362));
  NAND2_X1  g161(.A1(G227gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT70), .ZN(new_n364));
  NAND4_X1  g163(.A1(new_n337), .A2(new_n358), .A3(new_n313), .A4(new_n364), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n360), .A2(new_n362), .A3(new_n363), .A4(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(new_n366), .B(KEYINPUT34), .ZN(new_n367));
  INV_X1    g166(.A(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G71gat), .B(G99gat), .ZN(new_n370));
  XNOR2_X1  g169(.A(new_n369), .B(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n359), .B1(KEYINPUT70), .B2(new_n361), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n363), .B1(new_n373), .B2(new_n365), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT32), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n372), .B1(new_n374), .B2(new_n375), .ZN(new_n376));
  NOR2_X1   g175(.A1(new_n374), .A2(KEYINPUT33), .ZN(new_n377));
  OAI21_X1  g176(.A(KEYINPUT71), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n362), .A3(new_n365), .ZN(new_n379));
  INV_X1    g178(.A(new_n363), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n379), .A2(new_n380), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n371), .B1(new_n381), .B2(KEYINPUT32), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT71), .ZN(new_n383));
  INV_X1    g182(.A(KEYINPUT33), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n381), .A2(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n383), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n378), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n381), .A2(KEYINPUT32), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n371), .A2(new_n384), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(new_n390), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n368), .B1(new_n387), .B2(new_n391), .ZN(new_n392));
  AOI211_X1 g191(.A(new_n367), .B(new_n390), .C1(new_n378), .C2(new_n386), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G8gat), .B(G36gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(G64gat), .B(G92gat), .ZN(new_n396));
  XOR2_X1   g195(.A(new_n395), .B(new_n396), .Z(new_n397));
  INV_X1    g196(.A(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g198(.A1(G226gat), .A2(G233gat), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(KEYINPUT27), .B(G183gat), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n354), .B1(KEYINPUT65), .B2(new_n402), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT28), .ZN(new_n404));
  AOI21_X1  g203(.A(new_n357), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n345), .A2(new_n347), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n322), .A2(KEYINPUT64), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n407), .A2(new_n335), .A3(new_n325), .A4(new_n326), .ZN(new_n408));
  INV_X1    g207(.A(new_n329), .ZN(new_n409));
  AOI21_X1  g208(.A(KEYINPUT25), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n327), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT25), .ZN(new_n412));
  NOR3_X1   g211(.A1(new_n411), .A2(new_n329), .A3(new_n412), .ZN(new_n413));
  OAI22_X1  g212(.A1(new_n405), .A2(new_n406), .B1(new_n410), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n401), .B1(new_n414), .B2(new_n221), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n400), .B1(new_n337), .B2(new_n358), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n399), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(KEYINPUT29), .B1(new_n337), .B2(new_n358), .ZN(new_n418));
  OAI21_X1  g217(.A(KEYINPUT76), .B1(new_n418), .B2(new_n401), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n220), .B1(new_n417), .B2(new_n419), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n414), .A2(new_n401), .ZN(new_n421));
  OAI21_X1  g220(.A(new_n421), .B1(new_n418), .B2(new_n401), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(new_n261), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n398), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n422), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n425), .A2(new_n220), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n405), .A2(new_n406), .ZN(new_n427));
  AND2_X1   g226(.A1(new_n318), .A2(new_n316), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n325), .B(new_n326), .C1(new_n334), .C2(new_n331), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n322), .A2(KEYINPUT64), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n428), .B(new_n315), .C1(new_n429), .C2(new_n430), .ZN(new_n431));
  AOI22_X1  g230(.A1(new_n431), .A2(new_n412), .B1(new_n327), .B2(new_n319), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n221), .B1(new_n427), .B2(new_n432), .ZN(new_n433));
  AOI21_X1  g232(.A(new_n399), .B1(new_n433), .B2(new_n400), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(new_n399), .B2(new_n422), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n426), .B(new_n397), .C1(new_n435), .C2(new_n220), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n424), .A2(new_n436), .A3(KEYINPUT30), .ZN(new_n437));
  NOR2_X1   g236(.A1(new_n420), .A2(new_n423), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT30), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n438), .A2(new_n439), .A3(new_n397), .ZN(new_n440));
  AND2_X1   g239(.A1(new_n437), .A2(new_n440), .ZN(new_n441));
  AND2_X1   g240(.A1(new_n306), .A2(new_n308), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT1), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n443), .A2(KEYINPUT69), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT69), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(KEYINPUT1), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n301), .A2(new_n302), .ZN(new_n448));
  AOI21_X1  g247(.A(new_n447), .B1(KEYINPUT67), .B2(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n442), .A2(new_n449), .A3(new_n303), .ZN(new_n450));
  INV_X1    g249(.A(KEYINPUT4), .ZN(new_n451));
  NAND4_X1  g250(.A1(new_n450), .A2(new_n238), .A3(new_n451), .A4(new_n299), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT81), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT4), .B1(new_n312), .B2(new_n269), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n450), .A2(new_n238), .A3(new_n299), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n457), .A2(new_n453), .A3(KEYINPUT4), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g258(.A1(new_n244), .A2(new_n245), .A3(new_n230), .ZN(new_n460));
  AND2_X1   g259(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n461));
  NOR2_X1   g260(.A1(KEYINPUT77), .A2(KEYINPUT2), .ZN(new_n462));
  NOR2_X1   g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  AOI21_X1  g262(.A(new_n245), .B1(new_n244), .B2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(KEYINPUT3), .B1(new_n460), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n465), .A2(new_n312), .A3(new_n247), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n466), .A2(KEYINPUT78), .ZN(new_n467));
  INV_X1    g266(.A(KEYINPUT78), .ZN(new_n468));
  NAND4_X1  g267(.A1(new_n465), .A2(new_n312), .A3(new_n468), .A4(new_n247), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n467), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g269(.A1(G225gat), .A2(G233gat), .ZN(new_n471));
  INV_X1    g270(.A(new_n471), .ZN(new_n472));
  NOR2_X1   g271(.A1(new_n472), .A2(KEYINPUT5), .ZN(new_n473));
  AND3_X1   g272(.A1(new_n459), .A2(new_n470), .A3(new_n473), .ZN(new_n474));
  INV_X1    g273(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n312), .A2(new_n269), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n476), .A3(KEYINPUT79), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT79), .ZN(new_n478));
  NAND3_X1  g277(.A1(new_n312), .A2(new_n478), .A3(new_n269), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n477), .A2(new_n472), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT5), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n455), .A2(new_n452), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n470), .A2(new_n483), .A3(new_n471), .ZN(new_n484));
  AOI21_X1  g283(.A(KEYINPUT80), .B1(new_n482), .B2(new_n484), .ZN(new_n485));
  AOI221_X4 g284(.A(new_n472), .B1(new_n455), .B2(new_n452), .C1(new_n467), .C2(new_n469), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT80), .ZN(new_n487));
  NOR3_X1   g286(.A1(new_n486), .A2(new_n481), .A3(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(new_n475), .B1(new_n485), .B2(new_n488), .ZN(new_n489));
  XNOR2_X1  g288(.A(G1gat), .B(G29gat), .ZN(new_n490));
  XNOR2_X1  g289(.A(new_n490), .B(KEYINPUT0), .ZN(new_n491));
  XNOR2_X1  g290(.A(G57gat), .B(G85gat), .ZN(new_n492));
  XOR2_X1   g291(.A(new_n491), .B(new_n492), .Z(new_n493));
  INV_X1    g292(.A(new_n493), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n489), .A2(KEYINPUT82), .A3(new_n494), .ZN(new_n495));
  OAI21_X1  g294(.A(new_n487), .B1(new_n486), .B2(new_n481), .ZN(new_n496));
  NAND4_X1  g295(.A1(new_n484), .A2(KEYINPUT80), .A3(KEYINPUT5), .A4(new_n480), .ZN(new_n497));
  AOI21_X1  g296(.A(new_n474), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g297(.A(KEYINPUT6), .B1(new_n498), .B2(new_n493), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT82), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n500), .B1(new_n498), .B2(new_n493), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n499), .A3(new_n501), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n489), .A2(KEYINPUT6), .A3(new_n494), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n441), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n293), .A2(new_n394), .A3(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n505), .A2(KEYINPUT35), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT92), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND3_X1  g307(.A1(new_n505), .A2(KEYINPUT92), .A3(KEYINPUT35), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT35), .ZN(new_n510));
  AND2_X1   g309(.A1(new_n293), .A2(new_n510), .ZN(new_n511));
  NOR3_X1   g310(.A1(new_n376), .A2(new_n377), .A3(KEYINPUT71), .ZN(new_n512));
  AOI21_X1  g311(.A(new_n383), .B1(new_n382), .B2(new_n385), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n391), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(new_n367), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT73), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n390), .B1(new_n378), .B2(new_n386), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n517), .A2(new_n368), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  NOR3_X1   g318(.A1(new_n517), .A2(new_n516), .A3(new_n368), .ZN(new_n520));
  INV_X1    g319(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n437), .A2(new_n440), .ZN(new_n523));
  XNOR2_X1  g322(.A(new_n523), .B(KEYINPUT87), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n489), .A2(new_n494), .ZN(new_n525));
  AND3_X1   g324(.A1(new_n499), .A2(new_n525), .A3(KEYINPUT90), .ZN(new_n526));
  AOI21_X1  g325(.A(KEYINPUT90), .B1(new_n499), .B2(new_n525), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n503), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND4_X1  g327(.A1(new_n511), .A2(new_n522), .A3(new_n524), .A4(new_n528), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n508), .A2(new_n509), .A3(new_n529), .ZN(new_n530));
  INV_X1    g329(.A(KEYINPUT72), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n394), .A2(new_n531), .A3(KEYINPUT36), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n515), .A2(KEYINPUT36), .A3(new_n518), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(KEYINPUT72), .ZN(new_n534));
  OAI211_X1 g333(.A(new_n532), .B(new_n534), .C1(new_n522), .C2(KEYINPUT36), .ZN(new_n535));
  INV_X1    g334(.A(new_n293), .ZN(new_n536));
  NAND2_X1  g335(.A1(new_n499), .A2(new_n525), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT90), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n499), .A2(new_n525), .A3(KEYINPUT90), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  OAI21_X1  g340(.A(new_n426), .B1(new_n435), .B2(new_n220), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n398), .B1(new_n542), .B2(KEYINPUT37), .ZN(new_n543));
  INV_X1    g342(.A(KEYINPUT37), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n438), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g344(.A(KEYINPUT38), .B1(new_n543), .B2(new_n545), .ZN(new_n546));
  OR2_X1    g345(.A1(new_n435), .A2(new_n261), .ZN(new_n547));
  OAI21_X1  g346(.A(KEYINPUT37), .B1(new_n422), .B2(new_n220), .ZN(new_n548));
  INV_X1    g347(.A(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(KEYINPUT38), .B1(new_n547), .B2(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(new_n397), .B1(new_n438), .B2(new_n544), .ZN(new_n551));
  NAND3_X1  g350(.A1(new_n550), .A2(new_n551), .A3(KEYINPUT91), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n546), .A2(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  AOI21_X1  g353(.A(KEYINPUT91), .B1(new_n550), .B2(new_n551), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n503), .A2(new_n436), .ZN(new_n556));
  NOR2_X1   g355(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n541), .A2(new_n554), .A3(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(KEYINPUT87), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n523), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n459), .A2(new_n470), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n561), .A2(KEYINPUT88), .A3(new_n472), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT88), .ZN(new_n563));
  AOI22_X1  g362(.A1(new_n456), .A2(new_n458), .B1(new_n467), .B2(new_n469), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n563), .B1(new_n564), .B2(new_n471), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(KEYINPUT39), .ZN(new_n567));
  AOI21_X1  g366(.A(new_n494), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n477), .A2(new_n479), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n567), .B1(new_n569), .B2(new_n471), .ZN(new_n570));
  OR2_X1    g369(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n570), .A2(KEYINPUT89), .ZN(new_n572));
  NAND4_X1  g371(.A1(new_n571), .A2(new_n562), .A3(new_n565), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n568), .A2(KEYINPUT40), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n525), .ZN(new_n575));
  AOI21_X1  g374(.A(KEYINPUT40), .B1(new_n568), .B2(new_n573), .ZN(new_n576));
  NOR2_X1   g375(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n560), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g377(.A(new_n536), .B1(new_n558), .B2(new_n578), .ZN(new_n579));
  NAND2_X1  g378(.A1(new_n536), .A2(new_n504), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n535), .B1(new_n579), .B2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n530), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g382(.A1(G71gat), .A2(G78gat), .ZN(new_n584));
  NOR2_X1   g383(.A1(G71gat), .A2(G78gat), .ZN(new_n585));
  NOR2_X1   g384(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n586), .A2(KEYINPUT98), .ZN(new_n587));
  XNOR2_X1  g386(.A(G57gat), .B(G64gat), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT97), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT98), .ZN(new_n591));
  OAI21_X1  g390(.A(new_n591), .B1(new_n584), .B2(new_n585), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n587), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  OAI22_X1  g392(.A1(new_n588), .A2(new_n589), .B1(KEYINPUT9), .B2(new_n584), .ZN(new_n594));
  NOR2_X1   g393(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n595), .B(KEYINPUT99), .Z(new_n596));
  INV_X1    g395(.A(KEYINPUT9), .ZN(new_n597));
  OAI21_X1  g396(.A(new_n586), .B1(new_n588), .B2(new_n597), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n596), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT21), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(G231gat), .A2(G233gat), .ZN(new_n602));
  XNOR2_X1  g401(.A(new_n601), .B(new_n602), .ZN(new_n603));
  XNOR2_X1  g402(.A(new_n603), .B(G127gat), .ZN(new_n604));
  XNOR2_X1  g403(.A(G15gat), .B(G22gat), .ZN(new_n605));
  INV_X1    g404(.A(G1gat), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n606), .A2(KEYINPUT16), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n605), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n609));
  OAI211_X1 g408(.A(new_n608), .B(new_n609), .C1(G1gat), .C2(new_n605), .ZN(new_n610));
  NOR2_X1   g409(.A1(KEYINPUT94), .A2(G8gat), .ZN(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n612), .B1(new_n599), .B2(new_n600), .ZN(new_n613));
  OR2_X1    g412(.A1(new_n604), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n604), .A2(new_n613), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g415(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n228), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  XOR2_X1   g418(.A(new_n618), .B(new_n619), .Z(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g421(.A1(new_n614), .A2(new_n615), .A3(new_n620), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g423(.A(G43gat), .B(G50gat), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n625), .A2(KEYINPUT15), .ZN(new_n626));
  INV_X1    g425(.A(G50gat), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n627), .A2(KEYINPUT93), .A3(G43gat), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT15), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT93), .ZN(new_n631));
  AOI21_X1  g430(.A(new_n630), .B1(new_n625), .B2(new_n631), .ZN(new_n632));
  INV_X1    g431(.A(G29gat), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n633), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(KEYINPUT14), .B(G29gat), .ZN(new_n635));
  INV_X1    g434(.A(G36gat), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n626), .B1(new_n632), .B2(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(new_n638), .B1(new_n626), .B2(new_n637), .ZN(new_n639));
  OR2_X1    g438(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(KEYINPUT17), .ZN(new_n641));
  NAND2_X1  g440(.A1(G85gat), .A2(G92gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n642), .B(KEYINPUT7), .ZN(new_n643));
  INV_X1    g442(.A(G99gat), .ZN(new_n644));
  INV_X1    g443(.A(G106gat), .ZN(new_n645));
  OAI21_X1  g444(.A(KEYINPUT8), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n643), .B(new_n646), .C1(G85gat), .C2(G92gat), .ZN(new_n647));
  XNOR2_X1  g446(.A(G99gat), .B(G106gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n640), .A2(new_n641), .A3(new_n650), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT41), .ZN(new_n652));
  NAND2_X1  g451(.A1(G232gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(KEYINPUT100), .ZN(new_n654));
  OAI221_X1 g453(.A(new_n651), .B1(new_n652), .B2(new_n654), .C1(new_n639), .C2(new_n650), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(KEYINPUT101), .B1(new_n655), .B2(new_n656), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n654), .A2(new_n652), .ZN(new_n659));
  XOR2_X1   g458(.A(G134gat), .B(G162gat), .Z(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n657), .B(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n624), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n640), .A2(new_n612), .A3(new_n641), .ZN(new_n666));
  OR2_X1    g465(.A1(new_n612), .A2(new_n639), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(G229gat), .A2(G233gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(KEYINPUT18), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT95), .ZN(new_n673));
  OR2_X1    g472(.A1(new_n667), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n612), .A2(new_n639), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n667), .A2(new_n673), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n674), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g476(.A(new_n669), .B(KEYINPUT13), .Z(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  AND2_X1   g478(.A1(new_n672), .A2(new_n679), .ZN(new_n680));
  INV_X1    g479(.A(KEYINPUT96), .ZN(new_n681));
  XNOR2_X1  g480(.A(G113gat), .B(G141gat), .ZN(new_n682));
  XNOR2_X1  g481(.A(new_n682), .B(G197gat), .ZN(new_n683));
  XOR2_X1   g482(.A(KEYINPUT11), .B(G169gat), .Z(new_n684));
  XNOR2_X1  g483(.A(new_n683), .B(new_n684), .ZN(new_n685));
  XOR2_X1   g484(.A(new_n685), .B(KEYINPUT12), .Z(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n668), .A2(KEYINPUT18), .A3(new_n669), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n680), .A2(new_n681), .A3(new_n687), .A4(new_n688), .ZN(new_n689));
  NAND4_X1  g488(.A1(new_n672), .A2(new_n687), .A3(new_n688), .A4(new_n679), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(KEYINPUT96), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n689), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n680), .A2(new_n688), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n693), .A2(new_n686), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n695), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n599), .A2(new_n650), .ZN(new_n697));
  AOI21_X1  g496(.A(new_n649), .B1(new_n596), .B2(new_n598), .ZN(new_n698));
  OR3_X1    g497(.A1(new_n697), .A2(KEYINPUT10), .A3(new_n698), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n697), .A2(KEYINPUT10), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g500(.A1(G230gat), .A2(G233gat), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT102), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(G120gat), .B(G148gat), .ZN(new_n706));
  XNOR2_X1  g505(.A(G176gat), .B(G204gat), .ZN(new_n707));
  XOR2_X1   g506(.A(new_n706), .B(new_n707), .Z(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n697), .A2(new_n698), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n704), .ZN(new_n711));
  AOI21_X1  g510(.A(new_n709), .B1(new_n711), .B2(KEYINPUT103), .ZN(new_n712));
  OAI211_X1 g511(.A(new_n705), .B(new_n712), .C1(KEYINPUT103), .C2(new_n711), .ZN(new_n713));
  XOR2_X1   g512(.A(new_n708), .B(KEYINPUT104), .Z(new_n714));
  AOI21_X1  g513(.A(new_n703), .B1(new_n699), .B2(new_n700), .ZN(new_n715));
  OAI21_X1  g514(.A(new_n714), .B1(new_n715), .B2(new_n711), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n713), .A2(new_n716), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n665), .A2(new_n696), .A3(new_n717), .ZN(new_n718));
  AND3_X1   g517(.A1(new_n583), .A2(new_n718), .A3(KEYINPUT105), .ZN(new_n719));
  AOI21_X1  g518(.A(KEYINPUT105), .B1(new_n583), .B2(new_n718), .ZN(new_n720));
  NOR2_X1   g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n502), .A2(new_n503), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n723), .B(new_n606), .ZN(G1324gat));
  NOR2_X1   g523(.A1(new_n721), .A2(new_n524), .ZN(new_n725));
  INV_X1    g524(.A(G8gat), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  OR2_X1    g526(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n728));
  NAND2_X1  g527(.A1(new_n727), .A2(KEYINPUT106), .ZN(new_n729));
  XOR2_X1   g528(.A(KEYINPUT16), .B(G8gat), .Z(new_n730));
  NAND2_X1  g529(.A1(new_n725), .A2(new_n730), .ZN(new_n731));
  NOR2_X1   g530(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n732));
  AND2_X1   g531(.A1(new_n731), .A2(KEYINPUT42), .ZN(new_n733));
  OAI211_X1 g532(.A(new_n728), .B(new_n729), .C1(new_n732), .C2(new_n733), .ZN(G1325gat));
  AOI21_X1  g533(.A(new_n520), .B1(new_n394), .B2(new_n516), .ZN(new_n735));
  OR3_X1    g534(.A1(new_n721), .A2(G15gat), .A3(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(G15gat), .B1(new_n721), .B2(new_n535), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(G1326gat));
  NOR2_X1   g537(.A1(new_n721), .A2(new_n293), .ZN(new_n739));
  XOR2_X1   g538(.A(KEYINPUT43), .B(G22gat), .Z(new_n740));
  XNOR2_X1  g539(.A(new_n739), .B(new_n740), .ZN(G1327gat));
  INV_X1    g540(.A(KEYINPUT44), .ZN(new_n742));
  NAND4_X1  g541(.A1(new_n528), .A2(new_n524), .A3(new_n293), .A4(new_n510), .ZN(new_n743));
  NOR2_X1   g542(.A1(new_n743), .A2(new_n735), .ZN(new_n744));
  AOI21_X1  g543(.A(KEYINPUT92), .B1(new_n505), .B2(KEYINPUT35), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NOR3_X1   g545(.A1(new_n553), .A2(new_n555), .A3(new_n556), .ZN(new_n747));
  AOI22_X1  g546(.A1(new_n747), .A2(new_n541), .B1(new_n560), .B2(new_n577), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n580), .B1(new_n748), .B2(new_n536), .ZN(new_n749));
  AOI22_X1  g548(.A1(new_n746), .A2(new_n509), .B1(new_n749), .B2(new_n535), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n742), .B1(new_n750), .B2(new_n664), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n664), .B1(new_n530), .B2(new_n582), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(new_n754));
  NOR3_X1   g553(.A1(new_n624), .A2(new_n696), .A3(new_n717), .ZN(new_n755));
  INV_X1    g554(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  INV_X1    g556(.A(new_n722), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  AOI21_X1  g558(.A(new_n633), .B1(new_n759), .B2(KEYINPUT107), .ZN(new_n760));
  OAI21_X1  g559(.A(new_n760), .B1(KEYINPUT107), .B2(new_n759), .ZN(new_n761));
  INV_X1    g560(.A(new_n752), .ZN(new_n762));
  NOR2_X1   g561(.A1(new_n762), .A2(new_n756), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n763), .A2(new_n633), .A3(new_n758), .ZN(new_n764));
  XNOR2_X1  g563(.A(new_n764), .B(KEYINPUT45), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n761), .A2(new_n765), .ZN(G1328gat));
  NAND3_X1  g565(.A1(new_n763), .A2(new_n636), .A3(new_n560), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT46), .ZN(new_n768));
  AOI21_X1  g567(.A(new_n636), .B1(new_n757), .B2(new_n560), .ZN(new_n769));
  OR2_X1    g568(.A1(new_n768), .A2(new_n769), .ZN(G1329gat));
  INV_X1    g569(.A(KEYINPUT110), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT108), .ZN(new_n772));
  INV_X1    g571(.A(new_n535), .ZN(new_n773));
  NAND4_X1  g572(.A1(new_n751), .A2(new_n773), .A3(new_n753), .A4(new_n755), .ZN(new_n774));
  AOI21_X1  g573(.A(new_n772), .B1(new_n774), .B2(G43gat), .ZN(new_n775));
  INV_X1    g574(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n772), .A3(G43gat), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n735), .A2(G43gat), .ZN(new_n778));
  AOI21_X1  g577(.A(KEYINPUT47), .B1(new_n763), .B2(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n776), .A2(new_n777), .A3(new_n779), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n778), .ZN(new_n781));
  INV_X1    g580(.A(new_n781), .ZN(new_n782));
  INV_X1    g581(.A(G43gat), .ZN(new_n783));
  INV_X1    g582(.A(new_n774), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(KEYINPUT109), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n774), .A2(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n782), .B1(new_n785), .B2(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT47), .ZN(new_n789));
  OAI211_X1 g588(.A(new_n771), .B(new_n780), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  AOI21_X1  g589(.A(KEYINPUT44), .B1(new_n583), .B2(new_n663), .ZN(new_n791));
  AOI211_X1 g590(.A(new_n742), .B(new_n664), .C1(new_n530), .C2(new_n582), .ZN(new_n792));
  NOR2_X1   g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND4_X1  g592(.A1(new_n793), .A2(KEYINPUT109), .A3(new_n773), .A4(new_n755), .ZN(new_n794));
  NAND3_X1  g593(.A1(new_n787), .A2(new_n794), .A3(G43gat), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n789), .B1(new_n795), .B2(new_n781), .ZN(new_n796));
  NAND2_X1  g595(.A1(new_n777), .A2(new_n779), .ZN(new_n797));
  NOR2_X1   g596(.A1(new_n797), .A2(new_n775), .ZN(new_n798));
  OAI21_X1  g597(.A(KEYINPUT110), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n790), .A2(new_n799), .ZN(G1330gat));
  NAND3_X1  g599(.A1(new_n757), .A2(G50gat), .A3(new_n536), .ZN(new_n801));
  NOR3_X1   g600(.A1(new_n762), .A2(new_n293), .A3(new_n756), .ZN(new_n802));
  OAI21_X1  g601(.A(new_n801), .B1(G50gat), .B2(new_n802), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g603(.A(new_n717), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n665), .A2(new_n695), .A3(new_n805), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n583), .A2(new_n806), .ZN(new_n807));
  XOR2_X1   g606(.A(new_n807), .B(KEYINPUT111), .Z(new_n808));
  NAND2_X1  g607(.A1(new_n808), .A2(new_n758), .ZN(new_n809));
  XNOR2_X1  g608(.A(new_n809), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g609(.A1(new_n808), .A2(new_n560), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n811), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n812));
  XOR2_X1   g611(.A(KEYINPUT49), .B(G64gat), .Z(new_n813));
  OAI21_X1  g612(.A(new_n812), .B1(new_n811), .B2(new_n813), .ZN(G1333gat));
  INV_X1    g613(.A(G71gat), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n808), .A2(new_n815), .A3(new_n522), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n808), .A2(new_n773), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n816), .B1(new_n817), .B2(new_n815), .ZN(new_n818));
  INV_X1    g617(.A(KEYINPUT50), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OAI211_X1 g619(.A(KEYINPUT50), .B(new_n816), .C1(new_n817), .C2(new_n815), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(G1334gat));
  NAND2_X1  g621(.A1(new_n808), .A2(new_n536), .ZN(new_n823));
  XOR2_X1   g622(.A(KEYINPUT112), .B(G78gat), .Z(new_n824));
  XNOR2_X1  g623(.A(new_n823), .B(new_n824), .ZN(G1335gat));
  OR3_X1    g624(.A1(new_n624), .A2(KEYINPUT113), .A3(new_n695), .ZN(new_n826));
  OAI21_X1  g625(.A(KEYINPUT113), .B1(new_n624), .B2(new_n695), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n752), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT51), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n752), .A2(new_n828), .A3(KEYINPUT51), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n805), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(G85gat), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n833), .A2(new_n834), .A3(new_n758), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n717), .ZN(new_n836));
  OR3_X1    g635(.A1(new_n754), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n837));
  OAI21_X1  g636(.A(KEYINPUT114), .B1(new_n754), .B2(new_n836), .ZN(new_n838));
  AND3_X1   g637(.A1(new_n837), .A2(new_n758), .A3(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n835), .B1(new_n839), .B2(new_n834), .ZN(G1336gat));
  NOR2_X1   g639(.A1(new_n524), .A2(G92gat), .ZN(new_n841));
  INV_X1    g640(.A(new_n832), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT51), .B1(new_n752), .B2(new_n828), .ZN(new_n843));
  OAI211_X1 g642(.A(new_n717), .B(new_n841), .C1(new_n842), .C2(new_n843), .ZN(new_n844));
  XNOR2_X1  g643(.A(KEYINPUT116), .B(KEYINPUT52), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n754), .A2(new_n524), .A3(new_n836), .ZN(new_n846));
  INV_X1    g645(.A(G92gat), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n844), .B(new_n845), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n844), .A2(KEYINPUT115), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT115), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n833), .A2(new_n850), .A3(new_n841), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n837), .A2(new_n560), .A3(new_n838), .ZN(new_n853));
  AOI21_X1  g652(.A(new_n852), .B1(G92gat), .B2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n848), .B1(new_n854), .B2(new_n855), .ZN(G1337gat));
  NAND3_X1  g655(.A1(new_n833), .A2(new_n644), .A3(new_n522), .ZN(new_n857));
  AND3_X1   g656(.A1(new_n837), .A2(new_n773), .A3(new_n838), .ZN(new_n858));
  OAI21_X1  g657(.A(new_n857), .B1(new_n858), .B2(new_n644), .ZN(G1338gat));
  NOR2_X1   g658(.A1(new_n293), .A2(G106gat), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n833), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g660(.A(KEYINPUT117), .B(KEYINPUT53), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n754), .A2(new_n293), .A3(new_n836), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n861), .B(new_n862), .C1(new_n645), .C2(new_n863), .ZN(new_n864));
  NAND3_X1  g663(.A1(new_n837), .A2(new_n536), .A3(new_n838), .ZN(new_n865));
  AOI22_X1  g664(.A1(new_n865), .A2(G106gat), .B1(new_n833), .B2(new_n860), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n867));
  OAI21_X1  g666(.A(new_n864), .B1(new_n866), .B2(new_n867), .ZN(G1339gat));
  INV_X1    g667(.A(new_n624), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n699), .A2(new_n703), .A3(new_n700), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n705), .A2(KEYINPUT54), .A3(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872));
  AOI21_X1  g671(.A(new_n708), .B1(new_n715), .B2(new_n872), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n871), .A2(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT55), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g675(.A1(new_n871), .A2(KEYINPUT55), .A3(new_n873), .ZN(new_n877));
  NAND4_X1  g676(.A1(new_n876), .A2(new_n695), .A3(new_n713), .A4(new_n877), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n677), .A2(new_n678), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n668), .A2(new_n669), .ZN(new_n880));
  AOI21_X1  g679(.A(new_n879), .B1(KEYINPUT118), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(KEYINPUT118), .B2(new_n880), .ZN(new_n882));
  AOI22_X1  g681(.A1(new_n691), .A2(new_n689), .B1(new_n882), .B2(new_n685), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n883), .A2(new_n717), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n663), .B1(new_n878), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n876), .A2(new_n883), .A3(new_n663), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n877), .A2(new_n713), .ZN(new_n887));
  NOR2_X1   g686(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n869), .B1(new_n885), .B2(new_n888), .ZN(new_n889));
  NAND4_X1  g688(.A1(new_n624), .A2(new_n696), .A3(new_n664), .A4(new_n805), .ZN(new_n890));
  AOI211_X1 g689(.A(new_n735), .B(new_n536), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n560), .A2(new_n722), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  INV_X1    g692(.A(G113gat), .ZN(new_n894));
  NOR3_X1   g693(.A1(new_n893), .A2(new_n894), .A3(new_n696), .ZN(new_n895));
  AOI21_X1  g694(.A(new_n722), .B1(new_n889), .B2(new_n890), .ZN(new_n896));
  AND2_X1   g695(.A1(new_n293), .A2(new_n394), .ZN(new_n897));
  AND3_X1   g696(.A1(new_n896), .A2(new_n524), .A3(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G113gat), .B1(new_n898), .B2(new_n695), .ZN(new_n899));
  NOR2_X1   g698(.A1(new_n895), .A2(new_n899), .ZN(G1340gat));
  OAI21_X1  g699(.A(G120gat), .B1(new_n893), .B2(new_n805), .ZN(new_n901));
  XOR2_X1   g700(.A(new_n901), .B(KEYINPUT119), .Z(new_n902));
  INV_X1    g701(.A(G120gat), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n903), .A3(new_n717), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1341gat));
  OAI21_X1  g704(.A(G127gat), .B1(new_n893), .B2(new_n869), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n898), .A2(new_n294), .A3(new_n624), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n906), .A2(new_n907), .ZN(G1342gat));
  OAI21_X1  g707(.A(G134gat), .B1(new_n893), .B2(new_n664), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n664), .A2(new_n560), .ZN(new_n910));
  NAND4_X1  g709(.A1(new_n896), .A2(new_n295), .A3(new_n897), .A4(new_n910), .ZN(new_n911));
  OR2_X1    g710(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n911), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n909), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  AND2_X1   g713(.A1(new_n535), .A2(new_n892), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT57), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n293), .A2(new_n916), .ZN(new_n917));
  INV_X1    g716(.A(new_n917), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n696), .A2(new_n887), .ZN(new_n919));
  INV_X1    g718(.A(KEYINPUT120), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n876), .A2(new_n920), .ZN(new_n921));
  NAND3_X1  g720(.A1(new_n874), .A2(KEYINPUT120), .A3(new_n875), .ZN(new_n922));
  NAND3_X1  g721(.A1(new_n919), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n663), .B1(new_n923), .B2(new_n884), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n869), .B1(new_n924), .B2(new_n888), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n918), .B1(new_n925), .B2(new_n890), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n889), .A2(new_n890), .ZN(new_n927));
  AOI21_X1  g726(.A(KEYINPUT57), .B1(new_n927), .B2(new_n536), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n695), .B(new_n915), .C1(new_n926), .C2(new_n928), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n232), .B1(new_n929), .B2(KEYINPUT122), .ZN(new_n930));
  OAI21_X1  g729(.A(new_n930), .B1(KEYINPUT122), .B2(new_n929), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n773), .A2(new_n293), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n896), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n524), .ZN(new_n935));
  NOR3_X1   g734(.A1(new_n935), .A2(G141gat), .A3(new_n696), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(KEYINPUT58), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n931), .A2(new_n937), .ZN(new_n938));
  AND3_X1   g737(.A1(new_n929), .A2(KEYINPUT121), .A3(G141gat), .ZN(new_n939));
  AOI21_X1  g738(.A(KEYINPUT121), .B1(new_n929), .B2(G141gat), .ZN(new_n940));
  NOR3_X1   g739(.A1(new_n939), .A2(new_n940), .A3(new_n936), .ZN(new_n941));
  INV_X1    g740(.A(KEYINPUT58), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n938), .B1(new_n941), .B2(new_n942), .ZN(G1344gat));
  INV_X1    g742(.A(new_n935), .ZN(new_n944));
  NAND3_X1  g743(.A1(new_n944), .A2(new_n233), .A3(new_n717), .ZN(new_n945));
  OR2_X1    g744(.A1(new_n926), .A2(new_n928), .ZN(new_n946));
  AND2_X1   g745(.A1(new_n946), .A2(new_n915), .ZN(new_n947));
  AOI211_X1 g746(.A(KEYINPUT59), .B(new_n233), .C1(new_n947), .C2(new_n717), .ZN(new_n948));
  INV_X1    g747(.A(KEYINPUT59), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n927), .A2(new_n917), .ZN(new_n950));
  AOI21_X1  g749(.A(new_n293), .B1(new_n925), .B2(new_n890), .ZN(new_n951));
  OAI21_X1  g750(.A(new_n950), .B1(new_n951), .B2(KEYINPUT57), .ZN(new_n952));
  NAND3_X1  g751(.A1(new_n952), .A2(new_n717), .A3(new_n915), .ZN(new_n953));
  AOI21_X1  g752(.A(new_n949), .B1(new_n953), .B2(G148gat), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n945), .B1(new_n948), .B2(new_n954), .ZN(G1345gat));
  NAND3_X1  g754(.A1(new_n944), .A2(new_n228), .A3(new_n624), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n947), .A2(new_n624), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n956), .B1(new_n958), .B2(new_n228), .ZN(G1346gat));
  NAND3_X1  g758(.A1(new_n934), .A2(new_n229), .A3(new_n910), .ZN(new_n960));
  NAND2_X1  g759(.A1(new_n947), .A2(new_n663), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g761(.A(new_n960), .B1(new_n962), .B2(new_n229), .ZN(G1347gat));
  NOR2_X1   g762(.A1(new_n758), .A2(new_n524), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n891), .A2(new_n965), .ZN(new_n966));
  NOR3_X1   g765(.A1(new_n966), .A2(new_n338), .A3(new_n696), .ZN(new_n967));
  AOI21_X1  g766(.A(new_n758), .B1(new_n889), .B2(new_n890), .ZN(new_n968));
  AND3_X1   g767(.A1(new_n968), .A2(new_n560), .A3(new_n897), .ZN(new_n969));
  AOI21_X1  g768(.A(G169gat), .B1(new_n969), .B2(new_n695), .ZN(new_n970));
  NOR2_X1   g769(.A1(new_n967), .A2(new_n970), .ZN(G1348gat));
  OAI21_X1  g770(.A(G176gat), .B1(new_n966), .B2(new_n805), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n339), .A3(new_n717), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n972), .A2(new_n973), .ZN(G1349gat));
  OAI21_X1  g773(.A(G183gat), .B1(new_n966), .B2(new_n869), .ZN(new_n975));
  NAND3_X1  g774(.A1(new_n969), .A2(new_n402), .A3(new_n624), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  XNOR2_X1  g776(.A(new_n977), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g777(.A1(new_n969), .A2(new_n324), .A3(new_n663), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n891), .A2(new_n663), .A3(new_n965), .ZN(new_n980));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  NOR2_X1   g780(.A1(new_n981), .A2(KEYINPUT61), .ZN(new_n982));
  AOI21_X1  g781(.A(new_n324), .B1(new_n981), .B2(KEYINPUT61), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n980), .A2(new_n982), .A3(new_n983), .ZN(new_n984));
  AOI21_X1  g783(.A(new_n982), .B1(new_n980), .B2(new_n983), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n979), .B1(new_n984), .B2(new_n985), .ZN(G1351gat));
  NAND2_X1  g785(.A1(new_n932), .A2(new_n560), .ZN(new_n987));
  OR2_X1    g786(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n988));
  NAND2_X1  g787(.A1(new_n987), .A2(KEYINPUT125), .ZN(new_n989));
  NAND3_X1  g788(.A1(new_n988), .A2(new_n968), .A3(new_n989), .ZN(new_n990));
  INV_X1    g789(.A(new_n990), .ZN(new_n991));
  AOI21_X1  g790(.A(G197gat), .B1(new_n991), .B2(new_n695), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n965), .A2(new_n535), .ZN(new_n993));
  XNOR2_X1  g792(.A(new_n993), .B(KEYINPUT126), .ZN(new_n994));
  OR2_X1    g793(.A1(new_n951), .A2(KEYINPUT57), .ZN(new_n995));
  AOI21_X1  g794(.A(new_n994), .B1(new_n995), .B2(new_n950), .ZN(new_n996));
  AND2_X1   g795(.A1(new_n695), .A2(G197gat), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n992), .B1(new_n996), .B2(new_n997), .ZN(G1352gat));
  NAND2_X1  g797(.A1(new_n952), .A2(new_n717), .ZN(new_n999));
  OAI21_X1  g798(.A(G204gat), .B1(new_n999), .B2(new_n994), .ZN(new_n1000));
  OR2_X1    g799(.A1(new_n805), .A2(G204gat), .ZN(new_n1001));
  OR3_X1    g800(.A1(new_n990), .A2(KEYINPUT62), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g801(.A(KEYINPUT62), .B1(new_n990), .B2(new_n1001), .ZN(new_n1003));
  NAND3_X1  g802(.A1(new_n1000), .A2(new_n1002), .A3(new_n1003), .ZN(G1353gat));
  NOR2_X1   g803(.A1(new_n993), .A2(new_n869), .ZN(new_n1005));
  AOI21_X1  g804(.A(new_n210), .B1(new_n952), .B2(new_n1005), .ZN(new_n1006));
  OR3_X1    g805(.A1(new_n1006), .A2(KEYINPUT127), .A3(KEYINPUT63), .ZN(new_n1007));
  NAND3_X1  g806(.A1(new_n991), .A2(new_n210), .A3(new_n624), .ZN(new_n1008));
  AND2_X1   g807(.A1(new_n1006), .A2(KEYINPUT63), .ZN(new_n1009));
  OAI21_X1  g808(.A(KEYINPUT127), .B1(new_n1006), .B2(KEYINPUT63), .ZN(new_n1010));
  OAI211_X1 g809(.A(new_n1007), .B(new_n1008), .C1(new_n1009), .C2(new_n1010), .ZN(G1354gat));
  AOI21_X1  g810(.A(G218gat), .B1(new_n991), .B2(new_n663), .ZN(new_n1012));
  AOI21_X1  g811(.A(new_n664), .B1(new_n212), .B2(new_n214), .ZN(new_n1013));
  AOI21_X1  g812(.A(new_n1012), .B1(new_n996), .B2(new_n1013), .ZN(G1355gat));
endmodule


