//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 0 1 0 0 1 1 1 0 1 1 1 0 1 1 0 1 0 1 0 0 1 0 1 0 1 1 1 1 0 1 0 0 1 0 0 0 1 0 0 1 0 0 1 0 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:21 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n679,
    new_n680, new_n681, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n754, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n827,
    new_n828, new_n830, new_n831, new_n832, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n904, new_n905, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n915, new_n916, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n939, new_n940, new_n941, new_n942, new_n943, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n955, new_n956, new_n957;
  XNOR2_X1  g000(.A(G15gat), .B(G22gat), .ZN(new_n202));
  INV_X1    g001(.A(KEYINPUT16), .ZN(new_n203));
  AOI21_X1  g002(.A(G1gat), .B1(new_n202), .B2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G8gat), .ZN(new_n205));
  OR2_X1    g004(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n205), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g007(.A(new_n202), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT94), .ZN(new_n210));
  INV_X1    g009(.A(new_n210), .ZN(new_n211));
  NAND2_X1  g010(.A1(new_n208), .A2(new_n211), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n206), .A2(new_n210), .A3(new_n207), .ZN(new_n213));
  NAND2_X1  g012(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  NAND2_X1  g013(.A1(G29gat), .A2(G36gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G29gat), .A2(G36gat), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  NAND3_X1  g016(.A1(new_n216), .A2(KEYINPUT92), .A3(new_n217), .ZN(new_n218));
  XNOR2_X1  g017(.A(new_n216), .B(new_n217), .ZN(new_n219));
  OAI211_X1 g018(.A(new_n215), .B(new_n218), .C1(new_n219), .C2(KEYINPUT92), .ZN(new_n220));
  XNOR2_X1  g019(.A(G43gat), .B(G50gat), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n220), .A2(KEYINPUT15), .A3(new_n221), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT17), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224));
  OR3_X1    g023(.A1(new_n221), .A2(new_n224), .A3(KEYINPUT15), .ZN(new_n225));
  OAI21_X1  g024(.A(KEYINPUT15), .B1(new_n221), .B2(new_n224), .ZN(new_n226));
  NAND4_X1  g025(.A1(new_n225), .A2(new_n215), .A3(new_n226), .A4(new_n219), .ZN(new_n227));
  AND3_X1   g026(.A1(new_n222), .A2(new_n223), .A3(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n223), .B1(new_n222), .B2(new_n227), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n214), .B1(new_n228), .B2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(new_n222), .A2(new_n227), .ZN(new_n231));
  NAND3_X1  g030(.A1(new_n212), .A2(new_n231), .A3(new_n213), .ZN(new_n232));
  NAND2_X1  g031(.A1(G229gat), .A2(G233gat), .ZN(new_n233));
  XNOR2_X1  g032(.A(new_n233), .B(KEYINPUT95), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n230), .A2(new_n232), .A3(new_n234), .ZN(new_n235));
  INV_X1    g034(.A(KEYINPUT18), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n235), .A2(new_n236), .ZN(new_n237));
  AND2_X1   g036(.A1(new_n222), .A2(new_n227), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n214), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT96), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n240), .A3(new_n232), .ZN(new_n241));
  NAND4_X1  g040(.A1(new_n212), .A2(new_n231), .A3(KEYINPUT96), .A4(new_n213), .ZN(new_n242));
  XOR2_X1   g041(.A(new_n234), .B(KEYINPUT13), .Z(new_n243));
  NAND3_X1  g042(.A1(new_n241), .A2(new_n242), .A3(new_n243), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n230), .A2(KEYINPUT18), .A3(new_n232), .A4(new_n234), .ZN(new_n245));
  NAND3_X1  g044(.A1(new_n237), .A2(new_n244), .A3(new_n245), .ZN(new_n246));
  XNOR2_X1  g045(.A(KEYINPUT11), .B(G169gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n247), .B(G197gat), .ZN(new_n248));
  XOR2_X1   g047(.A(G113gat), .B(G141gat), .Z(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(KEYINPUT12), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n246), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g052(.A1(new_n237), .A2(new_n244), .A3(new_n251), .A4(new_n245), .ZN(new_n254));
  AND2_X1   g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  AND2_X1   g054(.A1(G71gat), .A2(G78gat), .ZN(new_n256));
  NOR2_X1   g055(.A1(G71gat), .A2(G78gat), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(KEYINPUT9), .B2(new_n257), .ZN(new_n258));
  INV_X1    g057(.A(G64gat), .ZN(new_n259));
  INV_X1    g058(.A(G57gat), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n259), .B1(new_n260), .B2(KEYINPUT97), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT97), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n262), .A2(G57gat), .A3(G64gat), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n261), .A2(new_n263), .ZN(new_n264));
  OAI21_X1  g063(.A(KEYINPUT98), .B1(new_n258), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G71gat), .A2(G78gat), .ZN(new_n266));
  INV_X1    g065(.A(G71gat), .ZN(new_n267));
  INV_X1    g066(.A(G78gat), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT9), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n266), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n271), .A2(new_n272), .A3(new_n261), .A4(new_n263), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n265), .A2(new_n273), .ZN(new_n274));
  OAI21_X1  g073(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n275), .B1(G57gat), .B2(G64gat), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n269), .A2(new_n266), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  INV_X1    g077(.A(new_n278), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n274), .A2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT99), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT7), .ZN(new_n282));
  OAI211_X1 g081(.A(G85gat), .B(G92gat), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n281), .A2(new_n282), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g084(.A1(new_n281), .A2(new_n282), .A3(G85gat), .A4(G92gat), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(KEYINPUT8), .ZN(new_n288));
  NOR2_X1   g087(.A1(G99gat), .A2(G106gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n288), .B1(new_n289), .B2(KEYINPUT100), .ZN(new_n290));
  NAND2_X1  g089(.A1(G99gat), .A2(G106gat), .ZN(new_n291));
  INV_X1    g090(.A(G85gat), .ZN(new_n292));
  INV_X1    g091(.A(G92gat), .ZN(new_n293));
  AOI22_X1  g092(.A1(new_n290), .A2(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n289), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(new_n291), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT100), .ZN(new_n298));
  INV_X1    g097(.A(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n295), .A2(new_n299), .ZN(new_n300));
  NAND3_X1  g099(.A1(new_n287), .A2(new_n294), .A3(new_n298), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n280), .A2(new_n300), .A3(new_n301), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n278), .B1(new_n265), .B2(new_n273), .ZN(new_n303));
  AND3_X1   g102(.A1(new_n287), .A2(new_n298), .A3(new_n294), .ZN(new_n304));
  AOI21_X1  g103(.A(new_n298), .B1(new_n287), .B2(new_n294), .ZN(new_n305));
  OAI21_X1  g104(.A(new_n303), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT101), .B(KEYINPUT10), .ZN(new_n307));
  NAND3_X1  g106(.A1(new_n302), .A2(new_n306), .A3(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT102), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n300), .A2(new_n301), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT10), .A3(new_n303), .ZN(new_n312));
  NAND4_X1  g111(.A1(new_n302), .A2(new_n306), .A3(KEYINPUT102), .A4(new_n307), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n310), .A2(new_n312), .A3(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(G230gat), .A2(G233gat), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n302), .A2(new_n306), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(G230gat), .A3(G233gat), .ZN(new_n318));
  AND2_X1   g117(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XNOR2_X1  g118(.A(G176gat), .B(G204gat), .ZN(new_n320));
  XNOR2_X1  g119(.A(new_n320), .B(G148gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(new_n321), .B(KEYINPUT104), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  XNOR2_X1  g122(.A(new_n322), .B(new_n323), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(KEYINPUT103), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n314), .A2(new_n326), .A3(new_n315), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n326), .B1(new_n314), .B2(new_n315), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n318), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n325), .A2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(KEYINPUT87), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT85), .ZN(new_n332));
  XOR2_X1   g131(.A(G141gat), .B(G148gat), .Z(new_n333));
  INV_X1    g132(.A(G155gat), .ZN(new_n334));
  INV_X1    g133(.A(G162gat), .ZN(new_n335));
  OAI21_X1  g134(.A(KEYINPUT2), .B1(new_n334), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G155gat), .B(G162gat), .ZN(new_n338));
  INV_X1    g137(.A(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n337), .A2(new_n339), .ZN(new_n340));
  NAND3_X1  g139(.A1(new_n333), .A2(new_n338), .A3(new_n336), .ZN(new_n341));
  NAND2_X1  g140(.A1(new_n340), .A2(new_n341), .ZN(new_n342));
  AND2_X1   g141(.A1(G197gat), .A2(G204gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(G197gat), .A2(G204gat), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT73), .ZN(new_n345));
  NOR3_X1   g144(.A1(new_n343), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  INV_X1    g145(.A(G197gat), .ZN(new_n347));
  INV_X1    g146(.A(G204gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  NAND2_X1  g148(.A1(G197gat), .A2(G204gat), .ZN(new_n350));
  AOI21_X1  g149(.A(KEYINPUT73), .B1(new_n349), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g150(.A(KEYINPUT22), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g151(.A1(G211gat), .A2(G218gat), .ZN(new_n353));
  NOR2_X1   g152(.A1(G211gat), .A2(G218gat), .ZN(new_n354));
  NOR2_X1   g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n355), .ZN(new_n357));
  OAI221_X1 g156(.A(new_n357), .B1(KEYINPUT22), .B2(new_n353), .C1(new_n346), .C2(new_n351), .ZN(new_n358));
  AOI21_X1  g157(.A(KEYINPUT29), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OAI211_X1 g158(.A(new_n332), .B(new_n342), .C1(new_n359), .C2(KEYINPUT3), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(G228gat), .A3(G233gat), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363));
  INV_X1    g162(.A(KEYINPUT3), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n340), .A2(new_n364), .A3(new_n341), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT29), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n356), .A2(new_n358), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT74), .ZN(new_n369));
  NOR2_X1   g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  AOI21_X1  g169(.A(KEYINPUT74), .B1(new_n356), .B2(new_n358), .ZN(new_n371));
  OAI21_X1  g170(.A(new_n367), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n342), .B1(new_n359), .B2(KEYINPUT3), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT85), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n362), .A2(new_n363), .A3(new_n372), .A4(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n372), .ZN(new_n376));
  OAI21_X1  g175(.A(KEYINPUT86), .B1(new_n376), .B2(new_n361), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n352), .A2(KEYINPUT82), .A3(new_n355), .ZN(new_n379));
  INV_X1    g178(.A(KEYINPUT82), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT22), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n345), .B1(new_n343), .B2(new_n344), .ZN(new_n382));
  NAND3_X1  g181(.A1(new_n349), .A2(KEYINPUT73), .A3(new_n350), .ZN(new_n383));
  AOI21_X1  g182(.A(new_n381), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  OAI21_X1  g183(.A(new_n380), .B1(new_n384), .B2(new_n357), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n379), .A2(new_n385), .A3(new_n358), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(new_n366), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(new_n364), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT77), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n342), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g189(.A1(new_n340), .A2(KEYINPUT77), .A3(new_n341), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(new_n392), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n388), .A2(KEYINPUT83), .A3(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT83), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT3), .B1(new_n386), .B2(new_n366), .ZN(new_n396));
  OAI21_X1  g195(.A(new_n395), .B1(new_n396), .B2(new_n392), .ZN(new_n397));
  NAND3_X1  g196(.A1(new_n394), .A2(new_n372), .A3(new_n397), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT84), .ZN(new_n399));
  NAND2_X1  g198(.A1(G228gat), .A2(G233gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n400), .B(KEYINPUT81), .Z(new_n401));
  AND3_X1   g200(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n399), .B1(new_n398), .B2(new_n401), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n378), .B1(new_n402), .B2(new_n403), .ZN(new_n404));
  XNOR2_X1  g203(.A(KEYINPUT31), .B(G50gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  XNOR2_X1  g205(.A(G78gat), .B(G106gat), .ZN(new_n407));
  XOR2_X1   g206(.A(new_n407), .B(G22gat), .Z(new_n408));
  INV_X1    g207(.A(new_n405), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n378), .B(new_n409), .C1(new_n402), .C2(new_n403), .ZN(new_n410));
  AND3_X1   g209(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n408), .B1(new_n406), .B2(new_n410), .ZN(new_n412));
  OAI21_X1  g211(.A(new_n331), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  XNOR2_X1  g212(.A(KEYINPUT0), .B(G57gat), .ZN(new_n414));
  XNOR2_X1  g213(.A(new_n414), .B(G85gat), .ZN(new_n415));
  XNOR2_X1  g214(.A(G1gat), .B(G29gat), .ZN(new_n416));
  XOR2_X1   g215(.A(new_n415), .B(new_n416), .Z(new_n417));
  INV_X1    g216(.A(new_n342), .ZN(new_n418));
  INV_X1    g217(.A(KEYINPUT1), .ZN(new_n419));
  INV_X1    g218(.A(G113gat), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n420), .A2(G120gat), .ZN(new_n421));
  NOR2_X1   g220(.A1(new_n323), .A2(G113gat), .ZN(new_n422));
  OAI21_X1  g221(.A(new_n419), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n423), .A2(KEYINPUT68), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT68), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n425), .B(new_n419), .C1(new_n421), .C2(new_n422), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n424), .A2(new_n426), .ZN(new_n427));
  XOR2_X1   g226(.A(G127gat), .B(G134gat), .Z(new_n428));
  NAND2_X1  g227(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  AOI21_X1  g228(.A(new_n428), .B1(new_n423), .B2(KEYINPUT68), .ZN(new_n430));
  INV_X1    g229(.A(new_n430), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n418), .A2(new_n429), .A3(new_n431), .ZN(new_n432));
  INV_X1    g231(.A(KEYINPUT79), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n432), .A2(new_n433), .A3(KEYINPUT4), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n429), .A2(new_n431), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n342), .A2(KEYINPUT3), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n436), .A3(new_n365), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT4), .ZN(new_n439));
  INV_X1    g238(.A(new_n428), .ZN(new_n440));
  AOI21_X1  g239(.A(new_n440), .B1(new_n424), .B2(new_n426), .ZN(new_n441));
  NOR2_X1   g240(.A1(new_n441), .A2(new_n430), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n392), .A2(new_n439), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n432), .A2(KEYINPUT4), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n443), .A2(new_n444), .A3(KEYINPUT79), .ZN(new_n445));
  NAND2_X1  g244(.A1(G225gat), .A2(G233gat), .ZN(new_n446));
  INV_X1    g245(.A(new_n446), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n447), .A2(KEYINPUT5), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n438), .A2(new_n445), .A3(new_n448), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n342), .B1(new_n441), .B2(new_n430), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n432), .A2(new_n450), .ZN(new_n451));
  AOI21_X1  g250(.A(KEYINPUT78), .B1(new_n451), .B2(new_n447), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT78), .ZN(new_n453));
  AOI211_X1 g252(.A(new_n453), .B(new_n446), .C1(new_n432), .C2(new_n450), .ZN(new_n454));
  OAI21_X1  g253(.A(KEYINPUT5), .B1(new_n452), .B2(new_n454), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n342), .A2(new_n441), .A3(new_n430), .ZN(new_n456));
  AOI21_X1  g255(.A(new_n456), .B1(new_n437), .B2(KEYINPUT4), .ZN(new_n457));
  AND3_X1   g256(.A1(new_n392), .A2(KEYINPUT4), .A3(new_n442), .ZN(new_n458));
  NOR3_X1   g257(.A1(new_n457), .A2(new_n458), .A3(new_n447), .ZN(new_n459));
  OAI211_X1 g258(.A(new_n417), .B(new_n449), .C1(new_n455), .C2(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT6), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  INV_X1    g261(.A(KEYINPUT80), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n449), .B1(new_n455), .B2(new_n459), .ZN(new_n465));
  INV_X1    g264(.A(new_n417), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n460), .A2(KEYINPUT80), .A3(new_n461), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n464), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n467), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n470), .A2(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n471), .ZN(new_n472));
  XNOR2_X1  g271(.A(G8gat), .B(G36gat), .ZN(new_n473));
  XNOR2_X1  g272(.A(new_n473), .B(new_n259), .ZN(new_n474));
  XNOR2_X1  g273(.A(new_n474), .B(new_n293), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g275(.A(KEYINPUT65), .B(G183gat), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT27), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT28), .ZN(new_n479));
  INV_X1    g278(.A(G183gat), .ZN(new_n480));
  NOR2_X1   g279(.A1(new_n480), .A2(KEYINPUT27), .ZN(new_n481));
  AOI21_X1  g280(.A(G190gat), .B1(new_n481), .B2(KEYINPUT66), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT66), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n480), .B2(KEYINPUT27), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n478), .A2(new_n479), .A3(new_n482), .A4(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(KEYINPUT27), .B(G183gat), .Z(new_n486));
  OAI21_X1  g285(.A(KEYINPUT28), .B1(new_n486), .B2(G190gat), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n485), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT67), .ZN(new_n489));
  NAND2_X1  g288(.A1(G183gat), .A2(G190gat), .ZN(new_n490));
  INV_X1    g289(.A(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(G169gat), .ZN(new_n492));
  INV_X1    g291(.A(G176gat), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g293(.A1(G169gat), .A2(G176gat), .ZN(new_n495));
  NOR3_X1   g294(.A1(new_n494), .A2(KEYINPUT26), .A3(new_n495), .ZN(new_n496));
  AOI211_X1 g295(.A(new_n491), .B(new_n496), .C1(KEYINPUT26), .C2(new_n495), .ZN(new_n497));
  INV_X1    g296(.A(KEYINPUT67), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n485), .A2(new_n498), .A3(new_n487), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n489), .A2(new_n497), .A3(new_n499), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT23), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n495), .A2(new_n501), .ZN(new_n502));
  OAI21_X1  g301(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n503));
  AOI21_X1  g302(.A(new_n494), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  XOR2_X1   g303(.A(new_n490), .B(KEYINPUT24), .Z(new_n505));
  NOR2_X1   g304(.A1(G183gat), .A2(G190gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT64), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n504), .B1(new_n505), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT25), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(new_n477), .ZN(new_n511));
  NOR2_X1   g310(.A1(new_n511), .A2(G190gat), .ZN(new_n512));
  OAI211_X1 g311(.A(KEYINPUT25), .B(new_n504), .C1(new_n512), .C2(new_n505), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n510), .A2(new_n513), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n500), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(KEYINPUT75), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT75), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n500), .A2(new_n517), .A3(new_n514), .ZN(new_n518));
  AND2_X1   g317(.A1(G226gat), .A2(G233gat), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n519), .A2(KEYINPUT29), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n516), .A2(new_n518), .A3(new_n520), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n370), .A2(new_n371), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n500), .A2(new_n514), .A3(new_n519), .ZN(new_n523));
  AND3_X1   g322(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n518), .ZN(new_n525));
  AOI21_X1  g324(.A(new_n517), .B1(new_n500), .B2(new_n514), .ZN(new_n526));
  OAI21_X1  g325(.A(new_n519), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  NAND2_X1  g326(.A1(new_n515), .A2(new_n520), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  OAI211_X1 g328(.A(KEYINPUT30), .B(new_n476), .C1(new_n524), .C2(new_n529), .ZN(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT76), .ZN(new_n531));
  INV_X1    g330(.A(new_n524), .ZN(new_n532));
  INV_X1    g331(.A(new_n529), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n532), .A2(new_n533), .A3(new_n475), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n534), .A2(KEYINPUT30), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n475), .B1(new_n532), .B2(new_n533), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g337(.A1(new_n472), .A2(new_n531), .A3(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(new_n408), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n398), .A2(new_n401), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n541), .A2(KEYINPUT84), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n398), .A2(new_n399), .A3(new_n401), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n409), .B1(new_n544), .B2(new_n378), .ZN(new_n545));
  INV_X1    g344(.A(new_n410), .ZN(new_n546));
  OAI21_X1  g345(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND3_X1  g346(.A1(new_n406), .A2(new_n408), .A3(new_n410), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n547), .A2(KEYINPUT87), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n413), .A2(new_n539), .A3(new_n549), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT36), .ZN(new_n551));
  OR3_X1    g350(.A1(new_n515), .A2(KEYINPUT69), .A3(new_n435), .ZN(new_n552));
  NAND2_X1  g351(.A1(G227gat), .A2(G233gat), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n515), .A2(new_n435), .ZN(new_n554));
  OAI21_X1  g353(.A(KEYINPUT69), .B1(new_n515), .B2(new_n435), .ZN(new_n555));
  NAND4_X1  g354(.A1(new_n552), .A2(new_n553), .A3(new_n554), .A4(new_n555), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n556), .B(KEYINPUT34), .ZN(new_n557));
  INV_X1    g356(.A(new_n557), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n552), .A2(new_n554), .A3(new_n555), .ZN(new_n559));
  INV_X1    g358(.A(new_n553), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT32), .ZN(new_n561));
  AOI22_X1  g360(.A1(new_n559), .A2(new_n560), .B1(new_n561), .B2(KEYINPUT33), .ZN(new_n562));
  XNOR2_X1  g361(.A(G15gat), .B(G43gat), .ZN(new_n563));
  XNOR2_X1  g362(.A(G71gat), .B(G99gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  XNOR2_X1  g364(.A(KEYINPUT70), .B(KEYINPUT71), .ZN(new_n566));
  XNOR2_X1  g365(.A(new_n565), .B(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(new_n567), .ZN(new_n568));
  NOR2_X1   g367(.A1(new_n562), .A2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(new_n561), .B1(new_n559), .B2(new_n560), .ZN(new_n571));
  OR2_X1    g370(.A1(new_n567), .A2(KEYINPUT72), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n572), .A2(KEYINPUT33), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n573), .B1(KEYINPUT72), .B2(new_n567), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n558), .B1(new_n570), .B2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n576), .ZN(new_n578));
  NOR3_X1   g377(.A1(new_n578), .A2(new_n569), .A3(new_n557), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n551), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(new_n558), .A3(new_n576), .ZN(new_n581));
  OAI21_X1  g380(.A(new_n557), .B1(new_n578), .B2(new_n569), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(KEYINPUT36), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g383(.A1(new_n550), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n585), .A2(KEYINPUT88), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n532), .A2(new_n533), .ZN(new_n587));
  NAND4_X1  g386(.A1(new_n587), .A2(KEYINPUT76), .A3(KEYINPUT30), .A4(new_n476), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT76), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n530), .A2(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  AOI21_X1  g390(.A(new_n536), .B1(new_n534), .B2(KEYINPUT30), .ZN(new_n592));
  OAI21_X1  g391(.A(KEYINPUT89), .B1(new_n591), .B2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT89), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n531), .A2(new_n594), .A3(new_n538), .ZN(new_n595));
  XOR2_X1   g394(.A(new_n417), .B(KEYINPUT90), .Z(new_n596));
  NAND2_X1  g395(.A1(new_n465), .A2(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT91), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n597), .B(new_n598), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n446), .B1(new_n438), .B2(new_n445), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT39), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n451), .A2(new_n447), .ZN(new_n602));
  NOR3_X1   g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  AOI211_X1 g402(.A(new_n596), .B(new_n603), .C1(new_n601), .C2(new_n600), .ZN(new_n604));
  AOI21_X1  g403(.A(new_n599), .B1(KEYINPUT40), .B2(new_n604), .ZN(new_n605));
  OR2_X1    g404(.A1(new_n604), .A2(KEYINPUT40), .ZN(new_n606));
  NAND4_X1  g405(.A1(new_n593), .A2(new_n595), .A3(new_n605), .A4(new_n606), .ZN(new_n607));
  INV_X1    g406(.A(KEYINPUT37), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n608), .ZN(new_n609));
  NAND3_X1  g408(.A1(new_n532), .A2(new_n533), .A3(KEYINPUT37), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(KEYINPUT38), .A3(new_n475), .A4(new_n610), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n527), .A2(new_n522), .A3(new_n528), .ZN(new_n612));
  AND2_X1   g411(.A1(new_n521), .A2(new_n523), .ZN(new_n613));
  OAI211_X1 g412(.A(new_n612), .B(KEYINPUT37), .C1(new_n522), .C2(new_n613), .ZN(new_n614));
  AND3_X1   g413(.A1(new_n609), .A2(new_n475), .A3(new_n614), .ZN(new_n615));
  OAI21_X1  g414(.A(new_n611), .B1(new_n615), .B2(KEYINPUT38), .ZN(new_n616));
  XNOR2_X1  g415(.A(new_n597), .B(KEYINPUT91), .ZN(new_n617));
  INV_X1    g416(.A(new_n462), .ZN(new_n618));
  AOI22_X1  g417(.A1(new_n617), .A2(new_n618), .B1(KEYINPUT6), .B2(new_n470), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n619), .A3(new_n537), .ZN(new_n620));
  NOR2_X1   g419(.A1(new_n411), .A2(new_n412), .ZN(new_n621));
  NAND3_X1  g420(.A1(new_n607), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT88), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n550), .A2(new_n623), .A3(new_n584), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n586), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n593), .A2(new_n595), .ZN(new_n626));
  INV_X1    g425(.A(new_n619), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n577), .A2(new_n579), .ZN(new_n628));
  NAND4_X1  g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .A4(new_n621), .ZN(new_n629));
  INV_X1    g428(.A(KEYINPUT35), .ZN(new_n630));
  AND3_X1   g429(.A1(new_n621), .A2(new_n628), .A3(KEYINPUT35), .ZN(new_n631));
  INV_X1    g430(.A(new_n539), .ZN(new_n632));
  AOI22_X1  g431(.A1(new_n629), .A2(new_n630), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  AOI211_X1 g432(.A(new_n255), .B(new_n330), .C1(new_n625), .C2(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n300), .B(new_n301), .C1(new_n228), .C2(new_n229), .ZN(new_n635));
  AND2_X1   g434(.A1(G232gat), .A2(G233gat), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n231), .A2(new_n311), .B1(KEYINPUT41), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n635), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(G134gat), .B(G162gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n638), .B(new_n640), .ZN(new_n641));
  NOR2_X1   g440(.A1(new_n636), .A2(KEYINPUT41), .ZN(new_n642));
  XNOR2_X1  g441(.A(G190gat), .B(G218gat), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n642), .B(new_n643), .ZN(new_n644));
  XOR2_X1   g443(.A(new_n641), .B(new_n644), .Z(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n303), .A2(KEYINPUT21), .ZN(new_n647));
  XNOR2_X1  g446(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n212), .A2(new_n213), .B1(KEYINPUT21), .B2(new_n303), .ZN(new_n651));
  XNOR2_X1  g450(.A(new_n651), .B(G183gat), .ZN(new_n652));
  NAND2_X1  g451(.A1(G231gat), .A2(G233gat), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g453(.A(G127gat), .B(G155gat), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n655), .B(G211gat), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n654), .A2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n657), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n654), .A2(new_n656), .ZN(new_n659));
  OAI21_X1  g458(.A(new_n650), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n659), .ZN(new_n661));
  NAND3_X1  g460(.A1(new_n661), .A2(new_n649), .A3(new_n657), .ZN(new_n662));
  AOI21_X1  g461(.A(new_n646), .B1(new_n660), .B2(new_n662), .ZN(new_n663));
  AND2_X1   g462(.A1(new_n634), .A2(new_n663), .ZN(new_n664));
  INV_X1    g463(.A(new_n472), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(G1gat), .ZN(G1324gat));
  INV_X1    g466(.A(new_n626), .ZN(new_n668));
  NAND2_X1  g467(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n203), .A2(new_n205), .ZN(new_n670));
  NAND4_X1  g469(.A1(new_n664), .A2(new_n668), .A3(new_n669), .A4(new_n670), .ZN(new_n671));
  INV_X1    g470(.A(KEYINPUT105), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  OR3_X1    g472(.A1(new_n671), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n205), .B1(new_n664), .B2(new_n668), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n675), .B1(new_n673), .B2(new_n671), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n672), .B1(new_n671), .B2(new_n673), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n674), .A2(new_n676), .A3(new_n677), .ZN(G1325gat));
  AOI21_X1  g477(.A(G15gat), .B1(new_n664), .B2(new_n628), .ZN(new_n679));
  INV_X1    g478(.A(new_n584), .ZN(new_n680));
  AND2_X1   g479(.A1(new_n664), .A2(G15gat), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n679), .B1(new_n680), .B2(new_n681), .ZN(G1326gat));
  NAND2_X1  g481(.A1(new_n413), .A2(new_n549), .ZN(new_n683));
  INV_X1    g482(.A(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n664), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(KEYINPUT43), .B(G22gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n685), .B(new_n686), .ZN(G1327gat));
  AOI21_X1  g486(.A(new_n645), .B1(new_n625), .B2(new_n633), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n660), .A2(new_n662), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n689), .A2(new_n255), .A3(new_n330), .ZN(new_n690));
  AND2_X1   g489(.A1(new_n688), .A2(new_n690), .ZN(new_n691));
  INV_X1    g490(.A(G29gat), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n665), .ZN(new_n693));
  XNOR2_X1  g492(.A(new_n693), .B(KEYINPUT45), .ZN(new_n694));
  NAND3_X1  g493(.A1(new_n622), .A2(new_n550), .A3(new_n584), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n695), .A2(new_n633), .ZN(new_n696));
  INV_X1    g495(.A(KEYINPUT44), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n696), .A2(new_n697), .A3(new_n646), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n698), .B1(new_n688), .B2(new_n697), .ZN(new_n699));
  XOR2_X1   g498(.A(new_n690), .B(KEYINPUT106), .Z(new_n700));
  AND2_X1   g499(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n701), .A2(new_n665), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n694), .B1(new_n692), .B2(new_n702), .ZN(G1328gat));
  INV_X1    g502(.A(G36gat), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n691), .A2(new_n704), .A3(new_n668), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT46), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n704), .B1(new_n701), .B2(new_n668), .ZN(new_n707));
  OR2_X1    g506(.A1(new_n706), .A2(new_n707), .ZN(G1329gat));
  INV_X1    g507(.A(KEYINPUT47), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n699), .A2(G43gat), .A3(new_n680), .A4(new_n700), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT107), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n688), .A2(new_n628), .A3(new_n690), .ZN(new_n712));
  INV_X1    g511(.A(G43gat), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(new_n711), .B1(new_n710), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n710), .A2(new_n714), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(KEYINPUT107), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n710), .A2(new_n711), .A3(new_n714), .ZN(new_n720));
  NAND3_X1  g519(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n720), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n717), .A2(new_n721), .ZN(G1330gat));
  INV_X1    g521(.A(G50gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n688), .A2(new_n723), .A3(new_n684), .A4(new_n690), .ZN(new_n724));
  INV_X1    g523(.A(new_n621), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n701), .A2(new_n725), .ZN(new_n726));
  OAI211_X1 g525(.A(KEYINPUT48), .B(new_n724), .C1(new_n726), .C2(new_n723), .ZN(new_n727));
  NAND3_X1  g526(.A1(new_n699), .A2(new_n684), .A3(new_n700), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT108), .ZN(new_n729));
  AND3_X1   g528(.A1(new_n728), .A2(new_n729), .A3(G50gat), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n729), .B1(new_n728), .B2(G50gat), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n724), .B(KEYINPUT109), .ZN(new_n732));
  NOR3_X1   g531(.A1(new_n730), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n727), .B1(new_n733), .B2(KEYINPUT48), .ZN(G1331gat));
  INV_X1    g533(.A(new_n330), .ZN(new_n735));
  AOI21_X1  g534(.A(new_n735), .B1(new_n695), .B2(new_n633), .ZN(new_n736));
  AND2_X1   g535(.A1(new_n663), .A2(new_n255), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n738), .A2(new_n472), .ZN(new_n739));
  XNOR2_X1  g538(.A(new_n739), .B(new_n260), .ZN(G1332gat));
  NOR2_X1   g539(.A1(new_n738), .A2(new_n626), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g544(.A(new_n628), .ZN(new_n746));
  OR3_X1    g545(.A1(new_n738), .A2(KEYINPUT111), .A3(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(KEYINPUT111), .B1(new_n738), .B2(new_n746), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n747), .A2(new_n267), .A3(new_n748), .ZN(new_n749));
  NAND4_X1  g548(.A1(new_n736), .A2(G71gat), .A3(new_n680), .A4(new_n737), .ZN(new_n750));
  XNOR2_X1  g549(.A(new_n750), .B(KEYINPUT110), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n752), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n683), .ZN(new_n754));
  XNOR2_X1  g553(.A(new_n754), .B(new_n268), .ZN(G1335gat));
  INV_X1    g554(.A(new_n255), .ZN(new_n756));
  NOR2_X1   g555(.A1(new_n689), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n699), .A2(new_n330), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n758), .A2(new_n292), .A3(new_n472), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n696), .A2(new_n646), .A3(new_n757), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT51), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n696), .A2(KEYINPUT51), .A3(new_n646), .A4(new_n757), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n735), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(G85gat), .B1(new_n764), .B2(new_n665), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n759), .A2(new_n765), .ZN(G1336gat));
  OAI21_X1  g565(.A(G92gat), .B1(new_n758), .B2(new_n626), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n762), .A2(new_n763), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n668), .A2(new_n293), .A3(new_n330), .ZN(new_n769));
  XNOR2_X1  g568(.A(new_n769), .B(KEYINPUT112), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n768), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT113), .B(KEYINPUT52), .Z(new_n773));
  XNOR2_X1  g572(.A(new_n772), .B(new_n773), .ZN(G1337gat));
  INV_X1    g573(.A(new_n758), .ZN(new_n775));
  AND3_X1   g574(.A1(new_n775), .A2(G99gat), .A3(new_n680), .ZN(new_n776));
  AOI21_X1  g575(.A(G99gat), .B1(new_n764), .B2(new_n628), .ZN(new_n777));
  NOR2_X1   g576(.A1(new_n776), .A2(new_n777), .ZN(G1338gat));
  AOI211_X1 g577(.A(G106gat), .B(new_n735), .C1(new_n762), .C2(new_n763), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n725), .ZN(new_n780));
  OAI21_X1  g579(.A(G106gat), .B1(new_n758), .B2(new_n621), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT53), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n775), .A2(new_n684), .ZN(new_n784));
  AOI22_X1  g583(.A1(new_n784), .A2(G106gat), .B1(new_n725), .B2(new_n779), .ZN(new_n785));
  OAI21_X1  g584(.A(new_n783), .B1(new_n785), .B2(new_n782), .ZN(G1339gat));
  NAND3_X1  g585(.A1(new_n663), .A2(new_n255), .A3(new_n735), .ZN(new_n787));
  INV_X1    g586(.A(new_n787), .ZN(new_n788));
  AOI21_X1  g587(.A(new_n243), .B1(new_n241), .B2(new_n242), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n234), .B1(new_n230), .B2(new_n232), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n250), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  AND2_X1   g590(.A1(new_n791), .A2(new_n254), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n330), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g592(.A1(new_n314), .A2(new_n315), .ZN(new_n794));
  OAI211_X1 g593(.A(KEYINPUT54), .B(new_n794), .C1(new_n327), .C2(new_n328), .ZN(new_n795));
  INV_X1    g594(.A(new_n316), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT54), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n324), .B1(new_n796), .B2(new_n797), .ZN(new_n798));
  NAND2_X1  g597(.A1(new_n795), .A2(new_n798), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT55), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n799), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n756), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n795), .A2(KEYINPUT55), .A3(new_n798), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n803), .A2(new_n329), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n793), .B1(new_n802), .B2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n805), .A2(new_n645), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n803), .A2(new_n329), .ZN(new_n807));
  NAND4_X1  g606(.A1(new_n807), .A2(new_n646), .A3(new_n792), .A4(new_n801), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n689), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n788), .B1(new_n809), .B2(new_n810), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n811), .A2(new_n472), .ZN(new_n812));
  NOR3_X1   g611(.A1(new_n668), .A2(new_n746), .A3(new_n725), .ZN(new_n813));
  NAND2_X1  g612(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n815), .A2(new_n420), .A3(new_n756), .ZN(new_n816));
  AOI22_X1  g615(.A1(new_n799), .A2(new_n800), .B1(new_n253), .B2(new_n254), .ZN(new_n817));
  NAND2_X1  g616(.A1(new_n807), .A2(new_n817), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n646), .B1(new_n818), .B2(new_n793), .ZN(new_n819));
  INV_X1    g618(.A(new_n808), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n810), .B1(new_n819), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n821), .A2(new_n787), .ZN(new_n822));
  NOR3_X1   g621(.A1(new_n684), .A2(new_n668), .A3(new_n472), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n628), .A3(new_n823), .ZN(new_n824));
  OAI21_X1  g623(.A(G113gat), .B1(new_n824), .B2(new_n255), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n816), .A2(new_n825), .ZN(G1340gat));
  NAND3_X1  g625(.A1(new_n815), .A2(new_n323), .A3(new_n330), .ZN(new_n827));
  OAI21_X1  g626(.A(G120gat), .B1(new_n824), .B2(new_n735), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(new_n828), .ZN(G1341gat));
  OAI21_X1  g628(.A(G127gat), .B1(new_n824), .B2(new_n810), .ZN(new_n830));
  OR2_X1    g629(.A1(new_n810), .A2(G127gat), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n830), .B1(new_n814), .B2(new_n831), .ZN(new_n832));
  XNOR2_X1  g631(.A(new_n832), .B(KEYINPUT114), .ZN(G1342gat));
  NOR3_X1   g632(.A1(new_n814), .A2(G134gat), .A3(new_n645), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT56), .ZN(new_n835));
  OAI21_X1  g634(.A(G134gat), .B1(new_n824), .B2(new_n645), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(G1343gat));
  AOI22_X1  g636(.A1(new_n807), .A2(new_n817), .B1(new_n330), .B2(new_n792), .ZN(new_n838));
  OAI21_X1  g637(.A(KEYINPUT115), .B1(new_n838), .B2(new_n646), .ZN(new_n839));
  INV_X1    g638(.A(KEYINPUT115), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n805), .A2(new_n840), .A3(new_n645), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n839), .A2(new_n841), .A3(new_n808), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n842), .A2(new_n810), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n843), .A2(new_n787), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n845));
  INV_X1    g644(.A(KEYINPUT57), .ZN(new_n846));
  NOR2_X1   g645(.A1(new_n683), .A2(new_n846), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n844), .A2(new_n845), .A3(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n621), .B1(new_n821), .B2(new_n787), .ZN(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n846), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n788), .B1(new_n842), .B2(new_n810), .ZN(new_n852));
  INV_X1    g651(.A(new_n847), .ZN(new_n853));
  OAI21_X1  g652(.A(KEYINPUT116), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND3_X1  g653(.A1(new_n848), .A2(new_n851), .A3(new_n854), .ZN(new_n855));
  NOR3_X1   g654(.A1(new_n680), .A2(new_n668), .A3(new_n472), .ZN(new_n856));
  NAND3_X1  g655(.A1(new_n855), .A2(new_n756), .A3(new_n856), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n857), .A2(G141gat), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n472), .B(new_n680), .C1(new_n821), .C2(new_n787), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n859), .A2(KEYINPUT117), .A3(new_n725), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n822), .A2(new_n665), .A3(new_n725), .A4(new_n584), .ZN(new_n861));
  INV_X1    g660(.A(KEYINPUT117), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n668), .B1(new_n860), .B2(new_n863), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n255), .A2(G141gat), .ZN(new_n865));
  AOI21_X1  g664(.A(KEYINPUT58), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n858), .A2(new_n866), .ZN(new_n867));
  NOR2_X1   g666(.A1(new_n861), .A2(new_n668), .ZN(new_n868));
  AOI22_X1  g667(.A1(new_n857), .A2(G141gat), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n867), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT118), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n867), .B(KEYINPUT118), .C1(new_n870), .C2(new_n869), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n873), .A2(new_n874), .ZN(G1344gat));
  NAND2_X1  g674(.A1(new_n860), .A2(new_n863), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n626), .ZN(new_n877));
  OR3_X1    g676(.A1(new_n877), .A2(G148gat), .A3(new_n735), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n855), .A2(new_n330), .A3(new_n856), .ZN(new_n879));
  INV_X1    g678(.A(KEYINPUT59), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n879), .A2(new_n880), .A3(G148gat), .ZN(new_n881));
  XNOR2_X1  g680(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n882));
  OAI21_X1  g681(.A(new_n846), .B1(new_n811), .B2(new_n683), .ZN(new_n883));
  AOI22_X1  g682(.A1(new_n883), .A2(KEYINPUT120), .B1(KEYINPUT57), .B2(new_n849), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n849), .A2(KEYINPUT120), .A3(KEYINPUT57), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  OAI211_X1 g685(.A(new_n330), .B(new_n856), .C1(new_n884), .C2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n882), .B1(new_n887), .B2(G148gat), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n878), .B1(new_n881), .B2(new_n888), .ZN(new_n889));
  INV_X1    g688(.A(KEYINPUT121), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g690(.A(new_n878), .B(KEYINPUT121), .C1(new_n881), .C2(new_n888), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(G1345gat));
  OAI21_X1  g692(.A(KEYINPUT122), .B1(new_n877), .B2(new_n810), .ZN(new_n894));
  INV_X1    g693(.A(KEYINPUT122), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n864), .A2(new_n895), .A3(new_n689), .ZN(new_n896));
  NAND3_X1  g695(.A1(new_n894), .A2(new_n896), .A3(new_n334), .ZN(new_n897));
  NAND4_X1  g696(.A1(new_n855), .A2(G155gat), .A3(new_n689), .A4(new_n856), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT123), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NAND3_X1  g700(.A1(new_n897), .A2(KEYINPUT123), .A3(new_n898), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n901), .A2(new_n902), .ZN(G1346gat));
  AOI21_X1  g702(.A(G162gat), .B1(new_n864), .B2(new_n646), .ZN(new_n904));
  AND3_X1   g703(.A1(new_n855), .A2(new_n646), .A3(new_n856), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n904), .B1(new_n905), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g705(.A1(new_n626), .A2(new_n665), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  NOR3_X1   g707(.A1(new_n811), .A2(new_n746), .A3(new_n908), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n909), .A2(new_n621), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n492), .A3(new_n756), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n909), .A2(new_n683), .ZN(new_n912));
  OAI21_X1  g711(.A(G169gat), .B1(new_n912), .B2(new_n255), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1348gat));
  AOI21_X1  g713(.A(G176gat), .B1(new_n910), .B2(new_n330), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n912), .A2(new_n493), .A3(new_n735), .ZN(new_n916));
  NOR2_X1   g715(.A1(new_n915), .A2(new_n916), .ZN(G1349gat));
  OAI21_X1  g716(.A(new_n511), .B1(new_n912), .B2(new_n810), .ZN(new_n918));
  INV_X1    g717(.A(new_n910), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n810), .A2(new_n486), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n918), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  XNOR2_X1  g720(.A(new_n921), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g721(.A(G190gat), .B1(new_n912), .B2(new_n645), .ZN(new_n923));
  XNOR2_X1  g722(.A(new_n923), .B(KEYINPUT61), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n645), .A2(G190gat), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n924), .B1(new_n919), .B2(new_n925), .ZN(G1351gat));
  AOI21_X1  g725(.A(KEYINPUT57), .B1(new_n822), .B2(new_n684), .ZN(new_n927));
  INV_X1    g726(.A(KEYINPUT120), .ZN(new_n928));
  OAI22_X1  g727(.A1(new_n927), .A2(new_n928), .B1(new_n850), .B2(new_n846), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n885), .ZN(new_n930));
  NOR2_X1   g729(.A1(new_n908), .A2(new_n680), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  OAI21_X1  g731(.A(G197gat), .B1(new_n932), .B2(new_n255), .ZN(new_n933));
  INV_X1    g732(.A(new_n931), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n850), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n347), .A3(new_n756), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n933), .A2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT124), .ZN(G1352gat));
  XNOR2_X1  g737(.A(KEYINPUT125), .B(G204gat), .ZN(new_n939));
  NOR4_X1   g738(.A1(new_n850), .A2(new_n934), .A3(new_n735), .A4(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT62), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n930), .A2(new_n330), .A3(new_n931), .ZN(new_n942));
  NAND2_X1  g741(.A1(new_n942), .A2(new_n939), .ZN(new_n943));
  NAND2_X1  g742(.A1(new_n941), .A2(new_n943), .ZN(G1353gat));
  INV_X1    g743(.A(KEYINPUT127), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n945), .B1(new_n932), .B2(new_n810), .ZN(new_n946));
  NAND4_X1  g745(.A1(new_n930), .A2(KEYINPUT127), .A3(new_n689), .A4(new_n931), .ZN(new_n947));
  NAND3_X1  g746(.A1(new_n946), .A2(G211gat), .A3(new_n947), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n948), .A2(KEYINPUT63), .ZN(new_n949));
  INV_X1    g748(.A(KEYINPUT63), .ZN(new_n950));
  NAND4_X1  g749(.A1(new_n946), .A2(new_n950), .A3(G211gat), .A4(new_n947), .ZN(new_n951));
  NOR4_X1   g750(.A1(new_n850), .A2(new_n934), .A3(G211gat), .A4(new_n810), .ZN(new_n952));
  XNOR2_X1  g751(.A(new_n952), .B(KEYINPUT126), .ZN(new_n953));
  NAND3_X1  g752(.A1(new_n949), .A2(new_n951), .A3(new_n953), .ZN(G1354gat));
  OAI21_X1  g753(.A(G218gat), .B1(new_n932), .B2(new_n645), .ZN(new_n955));
  INV_X1    g754(.A(G218gat), .ZN(new_n956));
  NAND3_X1  g755(.A1(new_n935), .A2(new_n956), .A3(new_n646), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(new_n957), .ZN(G1355gat));
endmodule


