

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583;

  XOR2_X1 U324 ( .A(n403), .B(n402), .Z(n551) );
  XNOR2_X1 U325 ( .A(n442), .B(n441), .ZN(n491) );
  XOR2_X1 U326 ( .A(n395), .B(n394), .Z(n292) );
  XOR2_X1 U327 ( .A(KEYINPUT62), .B(n583), .Z(n293) );
  NOR2_X1 U328 ( .A1(n523), .A2(n526), .ZN(n341) );
  XNOR2_X1 U329 ( .A(n342), .B(n320), .ZN(n321) );
  XNOR2_X1 U330 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U331 ( .A(n413), .B(n321), .ZN(n322) );
  XNOR2_X1 U332 ( .A(n396), .B(n292), .ZN(n397) );
  XNOR2_X1 U333 ( .A(n398), .B(n397), .ZN(n399) );
  NOR2_X1 U334 ( .A1(n507), .A2(n476), .ZN(n442) );
  NOR2_X1 U335 ( .A1(n568), .A2(n567), .ZN(n578) );
  NOR2_X1 U336 ( .A1(n528), .A2(n468), .ZN(n565) );
  XOR2_X1 U337 ( .A(n327), .B(n369), .Z(n513) );
  INV_X1 U338 ( .A(G29GAT), .ZN(n443) );
  XNOR2_X1 U339 ( .A(n469), .B(G190GAT), .ZN(n470) );
  XNOR2_X1 U340 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U341 ( .A(n471), .B(n470), .ZN(G1351GAT) );
  XNOR2_X1 U342 ( .A(n446), .B(n445), .ZN(G1328GAT) );
  INV_X1 U343 ( .A(KEYINPUT89), .ZN(n359) );
  XOR2_X1 U344 ( .A(KEYINPUT5), .B(G57GAT), .Z(n295) );
  XNOR2_X1 U345 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n294) );
  XNOR2_X1 U346 ( .A(n295), .B(n294), .ZN(n312) );
  XOR2_X1 U347 ( .A(G85GAT), .B(G148GAT), .Z(n297) );
  XNOR2_X1 U348 ( .A(G141GAT), .B(G120GAT), .ZN(n296) );
  XNOR2_X1 U349 ( .A(n297), .B(n296), .ZN(n299) );
  XOR2_X1 U350 ( .A(G29GAT), .B(G162GAT), .Z(n298) );
  XNOR2_X1 U351 ( .A(n299), .B(n298), .ZN(n308) );
  XNOR2_X1 U352 ( .A(KEYINPUT4), .B(KEYINPUT85), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n300), .B(KEYINPUT84), .ZN(n301) );
  XOR2_X1 U354 ( .A(n301), .B(KEYINPUT6), .Z(n306) );
  XOR2_X1 U355 ( .A(G127GAT), .B(KEYINPUT0), .Z(n303) );
  XNOR2_X1 U356 ( .A(G113GAT), .B(G134GAT), .ZN(n302) );
  XNOR2_X1 U357 ( .A(n303), .B(n302), .ZN(n346) );
  XNOR2_X1 U358 ( .A(G155GAT), .B(KEYINPUT2), .ZN(n304) );
  XNOR2_X1 U359 ( .A(n304), .B(KEYINPUT3), .ZN(n335) );
  XNOR2_X1 U360 ( .A(n346), .B(n335), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n307) );
  XNOR2_X1 U362 ( .A(n308), .B(n307), .ZN(n310) );
  NAND2_X1 U363 ( .A1(G225GAT), .A2(G233GAT), .ZN(n309) );
  XNOR2_X1 U364 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U365 ( .A(n312), .B(n311), .ZN(n510) );
  XOR2_X1 U366 ( .A(G211GAT), .B(KEYINPUT21), .Z(n314) );
  XNOR2_X1 U367 ( .A(G197GAT), .B(G218GAT), .ZN(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n334) );
  XOR2_X1 U369 ( .A(G36GAT), .B(G190GAT), .Z(n387) );
  XOR2_X1 U370 ( .A(G92GAT), .B(G64GAT), .Z(n316) );
  XNOR2_X1 U371 ( .A(G176GAT), .B(KEYINPUT72), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n317) );
  XOR2_X1 U373 ( .A(G204GAT), .B(n317), .Z(n413) );
  XOR2_X1 U374 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n319) );
  XNOR2_X1 U375 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n318) );
  XNOR2_X1 U376 ( .A(n319), .B(n318), .ZN(n342) );
  XOR2_X1 U377 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n320) );
  XOR2_X1 U378 ( .A(n387), .B(n322), .Z(n324) );
  NAND2_X1 U379 ( .A1(G226GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U380 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U381 ( .A(n334), .B(n325), .ZN(n327) );
  XNOR2_X1 U382 ( .A(G8GAT), .B(G183GAT), .ZN(n326) );
  XOR2_X1 U383 ( .A(n326), .B(KEYINPUT76), .Z(n369) );
  XNOR2_X1 U384 ( .A(KEYINPUT27), .B(n513), .ZN(n363) );
  NAND2_X1 U385 ( .A1(n510), .A2(n363), .ZN(n523) );
  XOR2_X1 U386 ( .A(G50GAT), .B(G162GAT), .Z(n393) );
  XOR2_X1 U387 ( .A(G78GAT), .B(G148GAT), .Z(n329) );
  XNOR2_X1 U388 ( .A(G106GAT), .B(KEYINPUT70), .ZN(n328) );
  XNOR2_X1 U389 ( .A(n329), .B(n328), .ZN(n416) );
  XNOR2_X1 U390 ( .A(n416), .B(KEYINPUT23), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n330), .B(G204GAT), .ZN(n333) );
  XOR2_X1 U392 ( .A(G141GAT), .B(G22GAT), .Z(n423) );
  XNOR2_X1 U393 ( .A(n423), .B(KEYINPUT24), .ZN(n331) );
  XNOR2_X1 U394 ( .A(n331), .B(KEYINPUT22), .ZN(n332) );
  XOR2_X1 U395 ( .A(n333), .B(n332), .Z(n337) );
  XNOR2_X1 U396 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U397 ( .A(n337), .B(n336), .ZN(n338) );
  XOR2_X1 U398 ( .A(n393), .B(n338), .Z(n340) );
  NAND2_X1 U399 ( .A1(G228GAT), .A2(G233GAT), .ZN(n339) );
  XNOR2_X1 U400 ( .A(n340), .B(n339), .ZN(n466) );
  XNOR2_X1 U401 ( .A(n466), .B(KEYINPUT28), .ZN(n526) );
  XNOR2_X1 U402 ( .A(n341), .B(KEYINPUT88), .ZN(n357) );
  XOR2_X1 U403 ( .A(G120GAT), .B(G71GAT), .Z(n417) );
  XOR2_X1 U404 ( .A(n417), .B(n342), .Z(n344) );
  NAND2_X1 U405 ( .A1(G227GAT), .A2(G233GAT), .ZN(n343) );
  XNOR2_X1 U406 ( .A(n344), .B(n343), .ZN(n345) );
  XOR2_X1 U407 ( .A(n345), .B(KEYINPUT83), .Z(n348) );
  XNOR2_X1 U408 ( .A(n346), .B(KEYINPUT82), .ZN(n347) );
  XNOR2_X1 U409 ( .A(n348), .B(n347), .ZN(n356) );
  XOR2_X1 U410 ( .A(G99GAT), .B(G190GAT), .Z(n350) );
  XNOR2_X1 U411 ( .A(G43GAT), .B(G15GAT), .ZN(n349) );
  XNOR2_X1 U412 ( .A(n350), .B(n349), .ZN(n354) );
  XOR2_X1 U413 ( .A(KEYINPUT81), .B(G183GAT), .Z(n352) );
  XNOR2_X1 U414 ( .A(G176GAT), .B(KEYINPUT20), .ZN(n351) );
  XNOR2_X1 U415 ( .A(n352), .B(n351), .ZN(n353) );
  XOR2_X1 U416 ( .A(n354), .B(n353), .Z(n355) );
  XOR2_X1 U417 ( .A(n356), .B(n355), .Z(n515) );
  INV_X1 U418 ( .A(n515), .ZN(n528) );
  NAND2_X1 U419 ( .A1(n357), .A2(n528), .ZN(n358) );
  XNOR2_X1 U420 ( .A(n359), .B(n358), .ZN(n368) );
  INV_X1 U421 ( .A(n510), .ZN(n464) );
  INV_X1 U422 ( .A(n513), .ZN(n460) );
  NOR2_X1 U423 ( .A1(n528), .A2(n460), .ZN(n360) );
  NOR2_X1 U424 ( .A1(n466), .A2(n360), .ZN(n361) );
  XNOR2_X1 U425 ( .A(n361), .B(KEYINPUT25), .ZN(n365) );
  NAND2_X1 U426 ( .A1(n528), .A2(n466), .ZN(n362) );
  XOR2_X1 U427 ( .A(n362), .B(KEYINPUT26), .Z(n542) );
  NAND2_X1 U428 ( .A1(n363), .A2(n542), .ZN(n364) );
  NAND2_X1 U429 ( .A1(n365), .A2(n364), .ZN(n366) );
  NAND2_X1 U430 ( .A1(n464), .A2(n366), .ZN(n367) );
  NAND2_X1 U431 ( .A1(n368), .A2(n367), .ZN(n474) );
  XOR2_X1 U432 ( .A(G57GAT), .B(KEYINPUT13), .Z(n411) );
  XNOR2_X1 U433 ( .A(n411), .B(n369), .ZN(n371) );
  NAND2_X1 U434 ( .A1(G231GAT), .A2(G233GAT), .ZN(n370) );
  XNOR2_X1 U435 ( .A(n371), .B(n370), .ZN(n386) );
  XOR2_X1 U436 ( .A(KEYINPUT77), .B(KEYINPUT78), .Z(n373) );
  XNOR2_X1 U437 ( .A(G64GAT), .B(KEYINPUT79), .ZN(n372) );
  XNOR2_X1 U438 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U439 ( .A(KEYINPUT80), .B(KEYINPUT12), .Z(n375) );
  XNOR2_X1 U440 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n374) );
  XNOR2_X1 U441 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U442 ( .A(n377), .B(n376), .ZN(n384) );
  XOR2_X1 U443 ( .A(G211GAT), .B(G155GAT), .Z(n379) );
  XNOR2_X1 U444 ( .A(G127GAT), .B(G71GAT), .ZN(n378) );
  XNOR2_X1 U445 ( .A(n379), .B(n378), .ZN(n380) );
  XOR2_X1 U446 ( .A(n380), .B(G78GAT), .Z(n382) );
  XOR2_X1 U447 ( .A(G15GAT), .B(G1GAT), .Z(n422) );
  XNOR2_X1 U448 ( .A(G22GAT), .B(n422), .ZN(n381) );
  XNOR2_X1 U449 ( .A(n382), .B(n381), .ZN(n383) );
  XNOR2_X1 U450 ( .A(n384), .B(n383), .ZN(n385) );
  XOR2_X1 U451 ( .A(n386), .B(n385), .Z(n472) );
  INV_X1 U452 ( .A(n472), .ZN(n579) );
  XOR2_X1 U453 ( .A(G99GAT), .B(G85GAT), .Z(n414) );
  XOR2_X1 U454 ( .A(n414), .B(n387), .Z(n389) );
  NAND2_X1 U455 ( .A1(G232GAT), .A2(G233GAT), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n398) );
  XOR2_X1 U457 ( .A(KEYINPUT73), .B(KEYINPUT74), .Z(n391) );
  XNOR2_X1 U458 ( .A(G218GAT), .B(KEYINPUT11), .ZN(n390) );
  XNOR2_X1 U459 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U460 ( .A(n393), .B(n392), .ZN(n396) );
  XOR2_X1 U461 ( .A(KEYINPUT10), .B(G92GAT), .Z(n395) );
  XNOR2_X1 U462 ( .A(G134GAT), .B(G106GAT), .ZN(n394) );
  XOR2_X1 U463 ( .A(n399), .B(KEYINPUT75), .Z(n403) );
  XOR2_X1 U464 ( .A(G29GAT), .B(G43GAT), .Z(n401) );
  XNOR2_X1 U465 ( .A(KEYINPUT8), .B(KEYINPUT7), .ZN(n400) );
  XNOR2_X1 U466 ( .A(n401), .B(n400), .ZN(n427) );
  XNOR2_X1 U467 ( .A(n427), .B(KEYINPUT9), .ZN(n402) );
  XNOR2_X1 U468 ( .A(n551), .B(KEYINPUT93), .ZN(n404) );
  XNOR2_X1 U469 ( .A(KEYINPUT36), .B(n404), .ZN(n582) );
  NOR2_X1 U470 ( .A1(n579), .A2(n582), .ZN(n405) );
  AND2_X1 U471 ( .A1(n474), .A2(n405), .ZN(n406) );
  XNOR2_X1 U472 ( .A(KEYINPUT37), .B(n406), .ZN(n507) );
  XOR2_X1 U473 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n408) );
  NAND2_X1 U474 ( .A1(G230GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U475 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U476 ( .A(KEYINPUT69), .B(n409), .ZN(n421) );
  XOR2_X1 U477 ( .A(KEYINPUT33), .B(KEYINPUT71), .Z(n410) );
  XNOR2_X1 U478 ( .A(n413), .B(n412), .ZN(n415) );
  XNOR2_X1 U479 ( .A(n415), .B(n414), .ZN(n419) );
  XOR2_X1 U480 ( .A(n417), .B(n416), .Z(n418) );
  XNOR2_X1 U481 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U482 ( .A(n421), .B(n420), .ZN(n573) );
  XOR2_X1 U483 ( .A(G36GAT), .B(G50GAT), .Z(n425) );
  XNOR2_X1 U484 ( .A(n423), .B(n422), .ZN(n424) );
  XNOR2_X1 U485 ( .A(n425), .B(n424), .ZN(n426) );
  XOR2_X1 U486 ( .A(n426), .B(G113GAT), .Z(n432) );
  XOR2_X1 U487 ( .A(n427), .B(KEYINPUT66), .Z(n429) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n428) );
  XNOR2_X1 U489 ( .A(n429), .B(n428), .ZN(n430) );
  XNOR2_X1 U490 ( .A(G169GAT), .B(n430), .ZN(n431) );
  XNOR2_X1 U491 ( .A(n432), .B(n431), .ZN(n440) );
  XOR2_X1 U492 ( .A(KEYINPUT65), .B(KEYINPUT30), .Z(n434) );
  XNOR2_X1 U493 ( .A(G197GAT), .B(G8GAT), .ZN(n433) );
  XNOR2_X1 U494 ( .A(n434), .B(n433), .ZN(n438) );
  XOR2_X1 U495 ( .A(KEYINPUT29), .B(KEYINPUT64), .Z(n436) );
  XNOR2_X1 U496 ( .A(KEYINPUT68), .B(KEYINPUT67), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U498 ( .A(n438), .B(n437), .Z(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n495) );
  INV_X1 U500 ( .A(n495), .ZN(n569) );
  NAND2_X1 U501 ( .A1(n573), .A2(n569), .ZN(n476) );
  XNOR2_X1 U502 ( .A(KEYINPUT94), .B(KEYINPUT38), .ZN(n441) );
  NAND2_X1 U503 ( .A1(n491), .A2(n510), .ZN(n446) );
  XOR2_X1 U504 ( .A(KEYINPUT95), .B(KEYINPUT39), .Z(n444) );
  XOR2_X1 U505 ( .A(KEYINPUT46), .B(KEYINPUT107), .Z(n448) );
  XNOR2_X1 U506 ( .A(n573), .B(KEYINPUT41), .ZN(n558) );
  NAND2_X1 U507 ( .A1(n569), .A2(n558), .ZN(n447) );
  XNOR2_X1 U508 ( .A(n448), .B(n447), .ZN(n449) );
  AND2_X1 U509 ( .A1(n472), .A2(n449), .ZN(n450) );
  XNOR2_X1 U510 ( .A(n450), .B(KEYINPUT108), .ZN(n452) );
  INV_X1 U511 ( .A(n551), .ZN(n451) );
  NAND2_X1 U512 ( .A1(n452), .A2(n451), .ZN(n453) );
  XNOR2_X1 U513 ( .A(n453), .B(KEYINPUT47), .ZN(n458) );
  NOR2_X1 U514 ( .A1(n472), .A2(n582), .ZN(n454) );
  XNOR2_X1 U515 ( .A(n454), .B(KEYINPUT45), .ZN(n455) );
  NAND2_X1 U516 ( .A1(n455), .A2(n573), .ZN(n456) );
  NOR2_X1 U517 ( .A1(n569), .A2(n456), .ZN(n457) );
  NOR2_X1 U518 ( .A1(n458), .A2(n457), .ZN(n459) );
  XNOR2_X1 U519 ( .A(KEYINPUT48), .B(n459), .ZN(n524) );
  NOR2_X1 U520 ( .A1(n524), .A2(n460), .ZN(n463) );
  XOR2_X1 U521 ( .A(KEYINPUT54), .B(KEYINPUT119), .Z(n461) );
  XNOR2_X1 U522 ( .A(KEYINPUT120), .B(n461), .ZN(n462) );
  XNOR2_X1 U523 ( .A(n463), .B(n462), .ZN(n465) );
  NAND2_X1 U524 ( .A1(n465), .A2(n464), .ZN(n567) );
  NOR2_X1 U525 ( .A1(n466), .A2(n567), .ZN(n467) );
  XNOR2_X1 U526 ( .A(n467), .B(KEYINPUT55), .ZN(n468) );
  NAND2_X1 U527 ( .A1(n565), .A2(n551), .ZN(n471) );
  XOR2_X1 U528 ( .A(KEYINPUT125), .B(KEYINPUT58), .Z(n469) );
  XOR2_X1 U529 ( .A(KEYINPUT34), .B(KEYINPUT90), .Z(n478) );
  NOR2_X1 U530 ( .A1(n472), .A2(n551), .ZN(n473) );
  XNOR2_X1 U531 ( .A(n473), .B(KEYINPUT16), .ZN(n475) );
  NAND2_X1 U532 ( .A1(n475), .A2(n474), .ZN(n496) );
  NOR2_X1 U533 ( .A1(n476), .A2(n496), .ZN(n485) );
  NAND2_X1 U534 ( .A1(n485), .A2(n510), .ZN(n477) );
  XNOR2_X1 U535 ( .A(n478), .B(n477), .ZN(n479) );
  XOR2_X1 U536 ( .A(G1GAT), .B(n479), .Z(G1324GAT) );
  XOR2_X1 U537 ( .A(KEYINPUT91), .B(KEYINPUT92), .Z(n481) );
  NAND2_X1 U538 ( .A1(n485), .A2(n513), .ZN(n480) );
  XNOR2_X1 U539 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U540 ( .A(G8GAT), .B(n482), .ZN(G1325GAT) );
  XOR2_X1 U541 ( .A(G15GAT), .B(KEYINPUT35), .Z(n484) );
  NAND2_X1 U542 ( .A1(n485), .A2(n515), .ZN(n483) );
  XNOR2_X1 U543 ( .A(n484), .B(n483), .ZN(G1326GAT) );
  NAND2_X1 U544 ( .A1(n526), .A2(n485), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n486), .B(G22GAT), .ZN(G1327GAT) );
  XNOR2_X1 U546 ( .A(G36GAT), .B(KEYINPUT96), .ZN(n488) );
  NAND2_X1 U547 ( .A1(n513), .A2(n491), .ZN(n487) );
  XNOR2_X1 U548 ( .A(n488), .B(n487), .ZN(G1329GAT) );
  NAND2_X1 U549 ( .A1(n491), .A2(n515), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n489), .B(KEYINPUT40), .ZN(n490) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n490), .ZN(G1330GAT) );
  XOR2_X1 U552 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n493) );
  NAND2_X1 U553 ( .A1(n491), .A2(n526), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U555 ( .A(G50GAT), .B(n494), .ZN(G1331GAT) );
  XOR2_X1 U556 ( .A(KEYINPUT99), .B(KEYINPUT42), .Z(n498) );
  NAND2_X1 U557 ( .A1(n495), .A2(n558), .ZN(n508) );
  NOR2_X1 U558 ( .A1(n508), .A2(n496), .ZN(n503) );
  NAND2_X1 U559 ( .A1(n503), .A2(n510), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U561 ( .A(G57GAT), .B(n499), .ZN(G1332GAT) );
  NAND2_X1 U562 ( .A1(n503), .A2(n513), .ZN(n500) );
  XNOR2_X1 U563 ( .A(n500), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U564 ( .A1(n503), .A2(n515), .ZN(n501) );
  XNOR2_X1 U565 ( .A(n501), .B(KEYINPUT100), .ZN(n502) );
  XNOR2_X1 U566 ( .A(G71GAT), .B(n502), .ZN(G1334GAT) );
  XOR2_X1 U567 ( .A(KEYINPUT101), .B(KEYINPUT43), .Z(n505) );
  NAND2_X1 U568 ( .A1(n503), .A2(n526), .ZN(n504) );
  XNOR2_X1 U569 ( .A(n505), .B(n504), .ZN(n506) );
  XOR2_X1 U570 ( .A(G78GAT), .B(n506), .Z(G1335GAT) );
  XOR2_X1 U571 ( .A(G85GAT), .B(KEYINPUT103), .Z(n512) );
  NOR2_X1 U572 ( .A1(n508), .A2(n507), .ZN(n509) );
  XNOR2_X1 U573 ( .A(n509), .B(KEYINPUT102), .ZN(n518) );
  NAND2_X1 U574 ( .A1(n518), .A2(n510), .ZN(n511) );
  XNOR2_X1 U575 ( .A(n512), .B(n511), .ZN(G1336GAT) );
  NAND2_X1 U576 ( .A1(n518), .A2(n513), .ZN(n514) );
  XNOR2_X1 U577 ( .A(n514), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U578 ( .A1(n518), .A2(n515), .ZN(n516) );
  XNOR2_X1 U579 ( .A(n516), .B(KEYINPUT104), .ZN(n517) );
  XNOR2_X1 U580 ( .A(G99GAT), .B(n517), .ZN(G1338GAT) );
  XNOR2_X1 U581 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n522) );
  XOR2_X1 U582 ( .A(KEYINPUT106), .B(KEYINPUT105), .Z(n520) );
  NAND2_X1 U583 ( .A1(n518), .A2(n526), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n520), .B(n519), .ZN(n521) );
  XNOR2_X1 U585 ( .A(n522), .B(n521), .ZN(G1339GAT) );
  XNOR2_X1 U586 ( .A(G113GAT), .B(KEYINPUT110), .ZN(n530) );
  NOR2_X1 U587 ( .A1(n524), .A2(n523), .ZN(n525) );
  XNOR2_X1 U588 ( .A(KEYINPUT109), .B(n525), .ZN(n543) );
  OR2_X1 U589 ( .A1(n543), .A2(n526), .ZN(n527) );
  NOR2_X1 U590 ( .A1(n528), .A2(n527), .ZN(n537) );
  NAND2_X1 U591 ( .A1(n537), .A2(n569), .ZN(n529) );
  XNOR2_X1 U592 ( .A(n530), .B(n529), .ZN(G1340GAT) );
  XOR2_X1 U593 ( .A(KEYINPUT111), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U594 ( .A1(n537), .A2(n558), .ZN(n531) );
  XNOR2_X1 U595 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U596 ( .A(G120GAT), .B(n533), .Z(G1341GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT112), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U598 ( .A1(n537), .A2(n579), .ZN(n534) );
  XNOR2_X1 U599 ( .A(n535), .B(n534), .ZN(n536) );
  XOR2_X1 U600 ( .A(G127GAT), .B(n536), .Z(G1342GAT) );
  XOR2_X1 U601 ( .A(KEYINPUT113), .B(KEYINPUT51), .Z(n539) );
  NAND2_X1 U602 ( .A1(n537), .A2(n551), .ZN(n538) );
  XNOR2_X1 U603 ( .A(n539), .B(n538), .ZN(n541) );
  XOR2_X1 U604 ( .A(G134GAT), .B(KEYINPUT114), .Z(n540) );
  XNOR2_X1 U605 ( .A(n541), .B(n540), .ZN(G1343GAT) );
  INV_X1 U606 ( .A(n542), .ZN(n568) );
  NOR2_X1 U607 ( .A1(n568), .A2(n543), .ZN(n552) );
  NAND2_X1 U608 ( .A1(n552), .A2(n569), .ZN(n544) );
  XNOR2_X1 U609 ( .A(G141GAT), .B(n544), .ZN(G1344GAT) );
  XOR2_X1 U610 ( .A(KEYINPUT115), .B(KEYINPUT52), .Z(n546) );
  NAND2_X1 U611 ( .A1(n552), .A2(n558), .ZN(n545) );
  XNOR2_X1 U612 ( .A(n546), .B(n545), .ZN(n548) );
  XOR2_X1 U613 ( .A(G148GAT), .B(KEYINPUT53), .Z(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(G1345GAT) );
  NAND2_X1 U615 ( .A1(n579), .A2(n552), .ZN(n549) );
  XNOR2_X1 U616 ( .A(n549), .B(KEYINPUT116), .ZN(n550) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(n550), .ZN(G1346GAT) );
  XOR2_X1 U618 ( .A(KEYINPUT117), .B(KEYINPUT118), .Z(n554) );
  NAND2_X1 U619 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U620 ( .A(n554), .B(n553), .ZN(n555) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT121), .Z(n557) );
  NAND2_X1 U623 ( .A1(n565), .A2(n569), .ZN(n556) );
  XNOR2_X1 U624 ( .A(n557), .B(n556), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n558), .A2(n565), .ZN(n564) );
  XOR2_X1 U626 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n560) );
  XNOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n559) );
  XNOR2_X1 U628 ( .A(n560), .B(n559), .ZN(n562) );
  XOR2_X1 U629 ( .A(G176GAT), .B(KEYINPUT122), .Z(n561) );
  XNOR2_X1 U630 ( .A(n562), .B(n561), .ZN(n563) );
  XNOR2_X1 U631 ( .A(n564), .B(n563), .ZN(G1349GAT) );
  NAND2_X1 U632 ( .A1(n579), .A2(n565), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n566), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n571) );
  NAND2_X1 U635 ( .A1(n578), .A2(n569), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(n572) );
  XNOR2_X1 U637 ( .A(G197GAT), .B(n572), .ZN(G1352GAT) );
  INV_X1 U638 ( .A(n578), .ZN(n581) );
  NOR2_X1 U639 ( .A1(n581), .A2(n573), .ZN(n577) );
  XOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .Z(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(KEYINPUT127), .ZN(n574) );
  XNOR2_X1 U642 ( .A(n575), .B(n574), .ZN(n576) );
  XNOR2_X1 U643 ( .A(n577), .B(n576), .ZN(G1353GAT) );
  NAND2_X1 U644 ( .A1(n579), .A2(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(n580), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(n293), .ZN(G1355GAT) );
endmodule

