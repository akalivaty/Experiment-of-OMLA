//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 0 0 1 0 0 1 0 0 0 1 1 0 0 1 1 1 1 1 0 1 0 1 1 1 1 1 0 0 0 0 1 0 1 0 1 1 0 1 1 1 1 1 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:12 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n208,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n602, new_n603, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n810, new_n811, new_n812, new_n813,
    new_n814, new_n815, new_n816, new_n817, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n824, new_n825, new_n826, new_n827,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR3_X1   g0006(.A1(new_n206), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0007(.A(G87), .B1(G97), .B2(G107), .ZN(new_n208));
  XNOR2_X1  g0008(.A(new_n208), .B(KEYINPUT65), .ZN(G355));
  NAND2_X1  g0009(.A1(G1), .A2(G20), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XNOR2_X1  g0012(.A(new_n212), .B(KEYINPUT0), .ZN(new_n213));
  NAND2_X1  g0013(.A1(new_n203), .A2(new_n205), .ZN(new_n214));
  INV_X1    g0014(.A(G50), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  INV_X1    g0017(.A(G20), .ZN(new_n218));
  NOR2_X1   g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  NAND2_X1  g0019(.A1(new_n216), .A2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(KEYINPUT66), .B(G238), .ZN(new_n221));
  NOR2_X1   g0021(.A1(new_n221), .A2(new_n202), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G77), .A2(G244), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G58), .A2(G232), .ZN(new_n226));
  NAND4_X1  g0026(.A1(new_n223), .A2(new_n224), .A3(new_n225), .A4(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n210), .B1(new_n222), .B2(new_n227), .ZN(new_n228));
  OAI211_X1 g0028(.A(new_n213), .B(new_n220), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  XNOR2_X1  g0031(.A(new_n231), .B(G232), .ZN(new_n232));
  XOR2_X1   g0032(.A(KEYINPUT2), .B(G226), .Z(new_n233));
  XNOR2_X1  g0033(.A(new_n232), .B(new_n233), .ZN(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(G264), .B(G270), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n234), .B(new_n237), .ZN(G358));
  XOR2_X1   g0038(.A(G87), .B(G97), .Z(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g0041(.A1(new_n215), .A2(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n202), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n241), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT77), .ZN(new_n248));
  INV_X1    g0048(.A(KEYINPUT69), .ZN(new_n249));
  NOR2_X1   g0049(.A1(new_n249), .A2(G58), .ZN(new_n250));
  NOR2_X1   g0050(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n251));
  OAI21_X1  g0051(.A(G68), .B1(new_n250), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g0052(.A(new_n218), .B1(new_n206), .B2(new_n252), .ZN(new_n253));
  NOR2_X1   g0053(.A1(G20), .A2(G33), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(G159), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n255), .A2(new_n256), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n253), .A2(new_n257), .ZN(new_n258));
  AND2_X1   g0058(.A1(KEYINPUT3), .A2(G33), .ZN(new_n259));
  NOR2_X1   g0059(.A1(KEYINPUT3), .A2(G33), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(new_n218), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT7), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n258), .B1(new_n263), .B2(new_n202), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT16), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  OAI21_X1  g0067(.A(new_n217), .B1(new_n210), .B2(new_n267), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  OAI21_X1  g0069(.A(KEYINPUT75), .B1(new_n253), .B2(new_n257), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n201), .A2(KEYINPUT69), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n249), .A2(G58), .ZN(new_n272));
  AOI21_X1  g0072(.A(new_n202), .B1(new_n271), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(G20), .B1(new_n273), .B2(new_n214), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT75), .ZN(new_n275));
  OAI211_X1 g0075(.A(new_n274), .B(new_n275), .C1(new_n256), .C2(new_n255), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n270), .A2(new_n276), .ZN(new_n277));
  OAI21_X1  g0077(.A(KEYINPUT73), .B1(new_n259), .B2(new_n260), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT3), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n267), .ZN(new_n280));
  INV_X1    g0080(.A(KEYINPUT73), .ZN(new_n281));
  NAND2_X1  g0081(.A1(KEYINPUT3), .A2(G33), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g0083(.A1(new_n278), .A2(new_n283), .A3(new_n218), .ZN(new_n284));
  INV_X1    g0084(.A(KEYINPUT7), .ZN(new_n285));
  AND2_X1   g0085(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  NAND4_X1  g0086(.A1(new_n280), .A2(KEYINPUT7), .A3(new_n218), .A4(new_n282), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(KEYINPUT74), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT74), .ZN(new_n289));
  NAND4_X1  g0089(.A1(new_n261), .A2(new_n289), .A3(KEYINPUT7), .A4(new_n218), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n288), .A2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(G68), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n277), .A2(KEYINPUT16), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(KEYINPUT76), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g0095(.A1(new_n277), .A2(new_n292), .A3(KEYINPUT76), .A4(KEYINPUT16), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n269), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G1), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n298), .A2(KEYINPUT67), .ZN(new_n299));
  INV_X1    g0099(.A(KEYINPUT67), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n300), .A2(G1), .ZN(new_n301));
  AND2_X1   g0101(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  AOI21_X1  g0102(.A(new_n268), .B1(new_n302), .B2(G20), .ZN(new_n303));
  INV_X1    g0103(.A(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(KEYINPUT8), .A2(G58), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n271), .A2(new_n272), .ZN(new_n306));
  AOI21_X1  g0106(.A(new_n305), .B1(new_n306), .B2(KEYINPUT8), .ZN(new_n307));
  NAND2_X1  g0107(.A1(new_n304), .A2(new_n307), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n302), .A2(G13), .A3(G20), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(new_n308), .B1(new_n307), .B2(new_n310), .ZN(new_n311));
  INV_X1    g0111(.A(new_n311), .ZN(new_n312));
  OAI21_X1  g0112(.A(new_n248), .B1(new_n297), .B2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n268), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n314), .B1(new_n264), .B2(new_n265), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n284), .A2(new_n285), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n316), .A2(new_n288), .A3(new_n290), .ZN(new_n317));
  AOI22_X1  g0117(.A1(new_n270), .A2(new_n276), .B1(new_n317), .B2(G68), .ZN(new_n318));
  AOI21_X1  g0118(.A(KEYINPUT76), .B1(new_n318), .B2(KEYINPUT16), .ZN(new_n319));
  AND4_X1   g0119(.A1(KEYINPUT76), .A2(new_n277), .A3(KEYINPUT16), .A4(new_n292), .ZN(new_n320));
  OAI21_X1  g0120(.A(new_n315), .B1(new_n319), .B2(new_n320), .ZN(new_n321));
  NAND3_X1  g0121(.A1(new_n321), .A2(KEYINPUT77), .A3(new_n311), .ZN(new_n322));
  INV_X1    g0122(.A(G226), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(G1698), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n324), .B1(G223), .B2(G1698), .ZN(new_n325));
  INV_X1    g0125(.A(G87), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n325), .A2(new_n261), .B1(new_n267), .B2(new_n326), .ZN(new_n327));
  AOI21_X1  g0127(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(G41), .ZN(new_n330));
  INV_X1    g0130(.A(G45), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g0132(.A1(new_n332), .A2(new_n298), .A3(G274), .ZN(new_n333));
  AOI21_X1  g0133(.A(new_n328), .B1(new_n302), .B2(new_n332), .ZN(new_n334));
  AOI21_X1  g0134(.A(new_n333), .B1(new_n334), .B2(G232), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n329), .A2(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G169), .ZN(new_n337));
  NOR2_X1   g0137(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AOI21_X1  g0138(.A(new_n338), .B1(G179), .B2(new_n336), .ZN(new_n339));
  INV_X1    g0139(.A(new_n339), .ZN(new_n340));
  NAND3_X1  g0140(.A1(new_n313), .A2(new_n322), .A3(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n341), .A2(KEYINPUT18), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n295), .A2(new_n296), .ZN(new_n343));
  AOI21_X1  g0143(.A(new_n312), .B1(new_n343), .B2(new_n315), .ZN(new_n344));
  NAND2_X1  g0144(.A1(new_n336), .A2(G190), .ZN(new_n345));
  INV_X1    g0145(.A(G200), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n345), .B1(new_n336), .B2(new_n346), .ZN(new_n347));
  INV_X1    g0147(.A(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(KEYINPUT17), .B1(new_n344), .B2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT17), .ZN(new_n350));
  NOR4_X1   g0150(.A1(new_n297), .A2(new_n350), .A3(new_n312), .A4(new_n347), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  INV_X1    g0152(.A(KEYINPUT18), .ZN(new_n353));
  NAND4_X1  g0153(.A1(new_n313), .A2(new_n322), .A3(new_n353), .A4(new_n340), .ZN(new_n354));
  NAND3_X1  g0154(.A1(new_n342), .A2(new_n352), .A3(new_n354), .ZN(new_n355));
  XOR2_X1   g0155(.A(new_n355), .B(KEYINPUT78), .Z(new_n356));
  NOR2_X1   g0156(.A1(new_n261), .A2(G1698), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G222), .ZN(new_n358));
  XNOR2_X1  g0158(.A(new_n358), .B(KEYINPUT68), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n280), .A2(new_n282), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G1698), .ZN(new_n361));
  INV_X1    g0161(.A(G223), .ZN(new_n362));
  INV_X1    g0162(.A(G77), .ZN(new_n363));
  OAI22_X1  g0163(.A1(new_n361), .A2(new_n362), .B1(new_n363), .B2(new_n360), .ZN(new_n364));
  OAI21_X1  g0164(.A(new_n328), .B1(new_n359), .B2(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n333), .B1(new_n334), .B2(G226), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  INV_X1    g0167(.A(G190), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n367), .A2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(G200), .B2(new_n367), .ZN(new_n370));
  NOR2_X1   g0170(.A1(new_n267), .A2(G20), .ZN(new_n371));
  AOI22_X1  g0171(.A1(new_n307), .A2(new_n371), .B1(G150), .B2(new_n254), .ZN(new_n372));
  OAI21_X1  g0172(.A(G20), .B1(new_n206), .B2(G50), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(new_n268), .ZN(new_n375));
  NOR2_X1   g0175(.A1(new_n309), .A2(G50), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n376), .B1(G50), .B2(new_n303), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  XNOR2_X1  g0178(.A(new_n378), .B(KEYINPUT9), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n370), .A2(new_n379), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n380), .A2(KEYINPUT10), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT10), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n370), .A2(new_n382), .A3(new_n379), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n381), .A2(new_n383), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n367), .A2(new_n337), .B1(new_n375), .B2(new_n377), .ZN(new_n385));
  INV_X1    g0185(.A(KEYINPUT70), .ZN(new_n386));
  OR2_X1    g0186(.A1(new_n385), .A2(new_n386), .ZN(new_n387));
  NOR2_X1   g0187(.A1(new_n367), .A2(G179), .ZN(new_n388));
  AOI21_X1  g0188(.A(new_n388), .B1(new_n385), .B2(new_n386), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  NAND2_X1  g0190(.A1(new_n384), .A2(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n255), .A2(new_n215), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n218), .A2(G33), .ZN(new_n393));
  OAI22_X1  g0193(.A1(new_n393), .A2(new_n363), .B1(new_n218), .B2(G68), .ZN(new_n394));
  OAI21_X1  g0194(.A(new_n268), .B1(new_n392), .B2(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT11), .ZN(new_n396));
  OAI21_X1  g0196(.A(new_n396), .B1(new_n202), .B2(new_n304), .ZN(new_n397));
  NOR2_X1   g0197(.A1(new_n309), .A2(G68), .ZN(new_n398));
  XNOR2_X1  g0198(.A(new_n398), .B(KEYINPUT12), .ZN(new_n399));
  NOR2_X1   g0199(.A1(new_n397), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(new_n400), .B(KEYINPUT71), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n360), .A2(G232), .A3(G1698), .ZN(new_n402));
  INV_X1    g0202(.A(G97), .ZN(new_n403));
  INV_X1    g0203(.A(G1698), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n360), .A2(new_n404), .ZN(new_n405));
  OAI221_X1 g0205(.A(new_n402), .B1(new_n267), .B2(new_n403), .C1(new_n405), .C2(new_n323), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n328), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n333), .B1(new_n334), .B2(G238), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g0209(.A(new_n409), .B(KEYINPUT13), .ZN(new_n410));
  INV_X1    g0210(.A(KEYINPUT14), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n410), .A2(new_n411), .A3(G169), .ZN(new_n412));
  INV_X1    g0212(.A(G179), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n412), .B1(new_n413), .B2(new_n410), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n411), .B1(new_n410), .B2(G169), .ZN(new_n415));
  OAI21_X1  g0215(.A(new_n401), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n410), .A2(G200), .ZN(new_n417));
  OAI211_X1 g0217(.A(new_n417), .B(new_n400), .C1(new_n368), .C2(new_n410), .ZN(new_n418));
  AND3_X1   g0218(.A1(new_n416), .A2(KEYINPUT72), .A3(new_n418), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT72), .B1(new_n416), .B2(new_n418), .ZN(new_n420));
  NAND3_X1  g0220(.A1(new_n360), .A2(G232), .A3(new_n404), .ZN(new_n421));
  INV_X1    g0221(.A(G107), .ZN(new_n422));
  OAI221_X1 g0222(.A(new_n421), .B1(new_n422), .B2(new_n360), .C1(new_n361), .C2(new_n221), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n423), .A2(new_n328), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n333), .B1(new_n334), .B2(G244), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n424), .A2(new_n425), .ZN(new_n426));
  INV_X1    g0226(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(new_n413), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n426), .A2(new_n337), .ZN(new_n429));
  XNOR2_X1  g0229(.A(KEYINPUT8), .B(G58), .ZN(new_n430));
  OAI22_X1  g0230(.A1(new_n430), .A2(new_n255), .B1(new_n218), .B2(new_n363), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT15), .B(G87), .ZN(new_n432));
  NOR2_X1   g0232(.A1(new_n432), .A2(new_n393), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n268), .B1(new_n431), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n303), .A2(G77), .ZN(new_n435));
  OAI211_X1 g0235(.A(new_n434), .B(new_n435), .C1(G77), .C2(new_n309), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n428), .A2(new_n429), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n436), .B1(new_n426), .B2(G200), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n438), .B1(new_n368), .B2(new_n426), .ZN(new_n439));
  NAND2_X1  g0239(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  NOR4_X1   g0240(.A1(new_n391), .A2(new_n419), .A3(new_n420), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n356), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g0243(.A1(new_n422), .A2(KEYINPUT6), .A3(G97), .ZN(new_n444));
  NOR2_X1   g0244(.A1(new_n403), .A2(new_n422), .ZN(new_n445));
  NOR2_X1   g0245(.A1(G97), .A2(G107), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g0247(.A(new_n444), .B1(new_n447), .B2(KEYINPUT6), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n448), .A2(G20), .B1(G77), .B2(new_n254), .ZN(new_n449));
  OAI21_X1  g0249(.A(new_n449), .B1(new_n263), .B2(new_n422), .ZN(new_n450));
  AOI22_X1  g0250(.A1(new_n450), .A2(new_n268), .B1(new_n403), .B2(new_n310), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n302), .A2(G33), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n309), .A2(new_n314), .A3(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(KEYINPUT79), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND4_X1  g0255(.A1(new_n309), .A2(new_n452), .A3(KEYINPUT79), .A4(new_n314), .ZN(new_n456));
  AND2_X1   g0256(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(G97), .ZN(new_n458));
  AND2_X1   g0258(.A1(new_n451), .A2(new_n458), .ZN(new_n459));
  AND3_X1   g0259(.A1(new_n299), .A2(new_n301), .A3(G45), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n460), .B1(KEYINPUT5), .B2(new_n330), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n461), .A2(KEYINPUT82), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT82), .ZN(new_n463));
  OAI211_X1 g0263(.A(new_n460), .B(new_n463), .C1(KEYINPUT5), .C2(new_n330), .ZN(new_n464));
  INV_X1    g0264(.A(G274), .ZN(new_n465));
  AND2_X1   g0265(.A1(new_n330), .A2(KEYINPUT5), .ZN(new_n466));
  NOR3_X1   g0266(.A1(new_n328), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n462), .A2(new_n464), .A3(new_n467), .ZN(new_n468));
  INV_X1    g0268(.A(new_n328), .ZN(new_n469));
  OAI211_X1 g0269(.A(G257), .B(new_n469), .C1(new_n461), .C2(new_n466), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(new_n471), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n357), .B(G244), .C1(KEYINPUT80), .C2(KEYINPUT4), .ZN(new_n473));
  NOR2_X1   g0273(.A1(KEYINPUT80), .A2(KEYINPUT4), .ZN(new_n474));
  INV_X1    g0274(.A(G244), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n474), .B1(new_n405), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(G33), .A2(G283), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n261), .A2(new_n404), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G250), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n473), .A2(new_n476), .A3(new_n477), .A4(new_n479), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(new_n328), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n472), .A2(G190), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n481), .A2(KEYINPUT81), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT81), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n480), .A2(new_n484), .A3(new_n328), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n471), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n459), .B(new_n482), .C1(new_n346), .C2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n472), .A2(new_n481), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n488), .A2(new_n337), .ZN(new_n489));
  AND3_X1   g0289(.A1(new_n480), .A2(new_n484), .A3(new_n328), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n484), .B1(new_n480), .B2(new_n328), .ZN(new_n491));
  OAI211_X1 g0291(.A(new_n413), .B(new_n472), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n451), .A2(new_n458), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n494));
  NAND3_X1  g0294(.A1(new_n360), .A2(new_n218), .A3(G87), .ZN(new_n495));
  XNOR2_X1  g0295(.A(new_n495), .B(KEYINPUT22), .ZN(new_n496));
  INV_X1    g0296(.A(KEYINPUT23), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n497), .B1(new_n218), .B2(G107), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n422), .A2(KEYINPUT23), .A3(G20), .ZN(new_n499));
  AOI22_X1  g0299(.A1(new_n498), .A2(new_n499), .B1(new_n371), .B2(G116), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n496), .A2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n501), .A2(KEYINPUT24), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT24), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n496), .A2(new_n503), .A3(new_n500), .ZN(new_n504));
  AOI21_X1  g0304(.A(new_n314), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(G33), .A2(G294), .ZN(new_n507));
  INV_X1    g0307(.A(G250), .ZN(new_n508));
  INV_X1    g0308(.A(G257), .ZN(new_n509));
  OAI221_X1 g0309(.A(new_n507), .B1(new_n405), .B2(new_n508), .C1(new_n509), .C2(new_n361), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n510), .A2(new_n328), .ZN(new_n511));
  OAI211_X1 g0311(.A(G264), .B(new_n469), .C1(new_n461), .C2(new_n466), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n511), .A2(new_n468), .A3(new_n512), .ZN(new_n513));
  OR2_X1    g0313(.A1(new_n513), .A2(new_n368), .ZN(new_n514));
  NOR2_X1   g0314(.A1(new_n309), .A2(G107), .ZN(new_n515));
  OR2_X1    g0315(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(KEYINPUT25), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n455), .A2(new_n456), .ZN(new_n519));
  OAI21_X1  g0319(.A(new_n518), .B1(new_n422), .B2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n513), .A2(G200), .ZN(new_n522));
  NAND4_X1  g0322(.A1(new_n506), .A2(new_n514), .A3(new_n521), .A4(new_n522), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n487), .A2(new_n494), .A3(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n478), .A2(G264), .ZN(new_n525));
  NAND2_X1  g0325(.A1(new_n357), .A2(G257), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n261), .A2(G303), .ZN(new_n527));
  NAND3_X1  g0327(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n528), .A2(new_n328), .ZN(new_n529));
  OAI211_X1 g0329(.A(G270), .B(new_n469), .C1(new_n461), .C2(new_n466), .ZN(new_n530));
  NAND3_X1  g0330(.A1(new_n529), .A2(new_n468), .A3(new_n530), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(KEYINPUT21), .A3(G169), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n529), .A2(new_n468), .A3(G179), .A4(new_n530), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  OAI211_X1 g0334(.A(new_n477), .B(new_n218), .C1(G33), .C2(new_n403), .ZN(new_n535));
  OAI211_X1 g0335(.A(new_n535), .B(new_n268), .C1(new_n218), .C2(G116), .ZN(new_n536));
  INV_X1    g0336(.A(KEYINPUT20), .ZN(new_n537));
  XNOR2_X1  g0337(.A(new_n536), .B(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G116), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n310), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n538), .B(new_n540), .C1(new_n539), .C2(new_n453), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n534), .A2(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n541), .B1(G200), .B2(new_n531), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n543), .B1(new_n368), .B2(new_n531), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n531), .A2(new_n541), .A3(G169), .ZN(new_n545));
  INV_X1    g0345(.A(KEYINPUT83), .ZN(new_n546));
  INV_X1    g0346(.A(KEYINPUT21), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  AOI21_X1  g0348(.A(new_n546), .B1(new_n545), .B2(new_n547), .ZN(new_n549));
  OAI211_X1 g0349(.A(new_n542), .B(new_n544), .C1(new_n548), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G116), .ZN(new_n551));
  INV_X1    g0351(.A(G238), .ZN(new_n552));
  OAI221_X1 g0352(.A(new_n551), .B1(new_n405), .B2(new_n552), .C1(new_n475), .C2(new_n361), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n460), .A2(new_n465), .ZN(new_n554));
  INV_X1    g0354(.A(new_n460), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n328), .B1(new_n555), .B2(new_n508), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n553), .A2(new_n328), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g0357(.A(new_n432), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n455), .A2(new_n558), .A3(new_n456), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n360), .A2(new_n218), .A3(G68), .ZN(new_n560));
  NOR2_X1   g0360(.A1(new_n393), .A2(new_n403), .ZN(new_n561));
  NOR2_X1   g0361(.A1(new_n267), .A2(new_n403), .ZN(new_n562));
  AOI21_X1  g0362(.A(G20), .B1(new_n562), .B2(KEYINPUT19), .ZN(new_n563));
  NOR3_X1   g0363(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n564));
  OAI221_X1 g0364(.A(new_n560), .B1(KEYINPUT19), .B2(new_n561), .C1(new_n563), .C2(new_n564), .ZN(new_n565));
  AOI22_X1  g0365(.A1(new_n565), .A2(new_n268), .B1(new_n310), .B2(new_n432), .ZN(new_n566));
  AOI22_X1  g0366(.A1(new_n413), .A2(new_n557), .B1(new_n559), .B2(new_n566), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n567), .B1(G169), .B2(new_n557), .ZN(new_n568));
  NAND3_X1  g0368(.A1(new_n455), .A2(G87), .A3(new_n456), .ZN(new_n569));
  AND2_X1   g0369(.A1(new_n569), .A2(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n557), .A2(G190), .ZN(new_n571));
  OAI211_X1 g0371(.A(new_n570), .B(new_n571), .C1(new_n346), .C2(new_n557), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n505), .A2(new_n520), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n513), .A2(new_n337), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n574), .B1(G179), .B2(new_n513), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n568), .B(new_n572), .C1(new_n573), .C2(new_n575), .ZN(new_n576));
  NOR3_X1   g0376(.A1(new_n524), .A2(new_n550), .A3(new_n576), .ZN(new_n577));
  AND2_X1   g0377(.A1(new_n443), .A2(new_n577), .ZN(G372));
  AND3_X1   g0378(.A1(new_n489), .A2(new_n492), .A3(new_n493), .ZN(new_n579));
  AND3_X1   g0379(.A1(new_n571), .A2(new_n566), .A3(new_n569), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n553), .A2(new_n328), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT84), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n556), .A2(new_n582), .A3(new_n554), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n582), .B1(new_n556), .B2(new_n554), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n585), .A2(G200), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n337), .ZN(new_n587));
  AOI22_X1  g0387(.A1(new_n580), .A2(new_n586), .B1(new_n587), .B2(new_n567), .ZN(new_n588));
  INV_X1    g0388(.A(KEYINPUT26), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n579), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n568), .A2(new_n572), .ZN(new_n591));
  OAI21_X1  g0391(.A(KEYINPUT26), .B1(new_n591), .B2(new_n494), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n587), .A2(new_n567), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n590), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n594), .A2(KEYINPUT85), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT85), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n590), .A2(new_n592), .A3(new_n596), .A4(new_n593), .ZN(new_n597));
  AND3_X1   g0397(.A1(new_n487), .A2(new_n494), .A3(new_n523), .ZN(new_n598));
  OAI221_X1 g0398(.A(new_n574), .B1(G179), .B2(new_n513), .C1(new_n505), .C2(new_n520), .ZN(new_n599));
  OAI211_X1 g0399(.A(new_n599), .B(new_n542), .C1(new_n549), .C2(new_n548), .ZN(new_n600));
  NAND3_X1  g0400(.A1(new_n598), .A2(new_n588), .A3(new_n600), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n595), .A2(new_n597), .A3(new_n601), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n443), .A2(new_n602), .ZN(new_n603));
  INV_X1    g0403(.A(new_n437), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n418), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n416), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g0406(.A1(new_n606), .A2(new_n352), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n321), .A2(new_n311), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n340), .ZN(new_n609));
  XNOR2_X1  g0409(.A(new_n609), .B(new_n353), .ZN(new_n610));
  AOI22_X1  g0410(.A1(new_n607), .A2(new_n610), .B1(new_n381), .B2(new_n383), .ZN(new_n611));
  INV_X1    g0411(.A(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT86), .ZN(new_n613));
  NAND3_X1  g0413(.A1(new_n612), .A2(new_n613), .A3(new_n390), .ZN(new_n614));
  INV_X1    g0414(.A(new_n390), .ZN(new_n615));
  OAI21_X1  g0415(.A(KEYINPUT86), .B1(new_n611), .B2(new_n615), .ZN(new_n616));
  NAND2_X1  g0416(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n603), .A2(new_n617), .ZN(G369));
  AND2_X1   g0418(.A1(new_n550), .A2(KEYINPUT87), .ZN(new_n619));
  AND2_X1   g0419(.A1(new_n218), .A2(G13), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n302), .A2(new_n620), .ZN(new_n621));
  OR2_X1    g0421(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n621), .A2(KEYINPUT27), .ZN(new_n623));
  NAND3_X1  g0423(.A1(new_n622), .A2(G213), .A3(new_n623), .ZN(new_n624));
  INV_X1    g0424(.A(G343), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n541), .A2(new_n626), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n627), .B1(new_n550), .B2(KEYINPUT87), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n545), .A2(new_n547), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n629), .A2(KEYINPUT83), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n630), .A2(new_n631), .B1(new_n534), .B2(new_n541), .ZN(new_n632));
  OAI22_X1  g0432(.A1(new_n619), .A2(new_n628), .B1(new_n632), .B2(new_n627), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G330), .ZN(new_n634));
  NOR2_X1   g0434(.A1(new_n573), .A2(new_n575), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n626), .B1(new_n505), .B2(new_n520), .ZN(new_n636));
  AOI21_X1  g0436(.A(new_n635), .B1(new_n523), .B2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n599), .A2(new_n626), .ZN(new_n638));
  NOR2_X1   g0438(.A1(new_n637), .A2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(new_n639), .ZN(new_n640));
  NOR2_X1   g0440(.A1(new_n634), .A2(new_n640), .ZN(new_n641));
  INV_X1    g0441(.A(new_n641), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n542), .B1(new_n548), .B2(new_n549), .ZN(new_n643));
  INV_X1    g0443(.A(new_n626), .ZN(new_n644));
  NAND2_X1  g0444(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  INV_X1    g0445(.A(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n523), .A2(new_n636), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n647), .A2(new_n599), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n638), .B1(new_n646), .B2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n642), .A2(new_n649), .ZN(G399));
  INV_X1    g0450(.A(new_n211), .ZN(new_n651));
  NOR2_X1   g0451(.A1(new_n651), .A2(G41), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n564), .A2(new_n539), .ZN(new_n653));
  NOR3_X1   g0453(.A1(new_n652), .A2(new_n653), .A3(new_n298), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n654), .B1(new_n216), .B2(new_n652), .ZN(new_n655));
  XOR2_X1   g0455(.A(new_n655), .B(KEYINPUT28), .Z(new_n656));
  INV_X1    g0456(.A(KEYINPUT89), .ZN(new_n657));
  AOI21_X1  g0457(.A(KEYINPUT29), .B1(new_n602), .B2(new_n644), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT29), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n600), .A2(KEYINPUT88), .ZN(new_n660));
  INV_X1    g0460(.A(KEYINPUT88), .ZN(new_n661));
  NAND3_X1  g0461(.A1(new_n632), .A2(new_n661), .A3(new_n599), .ZN(new_n662));
  NAND4_X1  g0462(.A1(new_n660), .A2(new_n662), .A3(new_n598), .A4(new_n588), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n589), .B1(new_n579), .B2(new_n588), .ZN(new_n664));
  NOR3_X1   g0464(.A1(new_n591), .A2(new_n494), .A3(KEYINPUT26), .ZN(new_n665));
  AND2_X1   g0465(.A1(new_n587), .A2(new_n567), .ZN(new_n666));
  NOR3_X1   g0466(.A1(new_n664), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  AOI211_X1 g0467(.A(new_n659), .B(new_n626), .C1(new_n663), .C2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n658), .A2(new_n668), .ZN(new_n669));
  INV_X1    g0469(.A(KEYINPUT31), .ZN(new_n670));
  INV_X1    g0470(.A(new_n550), .ZN(new_n671));
  INV_X1    g0471(.A(new_n576), .ZN(new_n672));
  NAND4_X1  g0472(.A1(new_n598), .A2(new_n671), .A3(new_n672), .A4(new_n644), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n557), .A2(new_n511), .A3(new_n512), .ZN(new_n674));
  NOR3_X1   g0474(.A1(new_n488), .A2(new_n674), .A3(new_n533), .ZN(new_n675));
  INV_X1    g0475(.A(new_n486), .ZN(new_n676));
  AND4_X1   g0476(.A1(new_n413), .A2(new_n585), .A3(new_n531), .A4(new_n513), .ZN(new_n677));
  AOI22_X1  g0477(.A1(KEYINPUT30), .A2(new_n675), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  OR2_X1    g0478(.A1(new_n675), .A2(KEYINPUT30), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n644), .B1(new_n678), .B2(new_n679), .ZN(new_n680));
  INV_X1    g0480(.A(new_n680), .ZN(new_n681));
  AOI21_X1  g0481(.A(new_n670), .B1(new_n673), .B2(new_n681), .ZN(new_n682));
  NOR2_X1   g0482(.A1(new_n680), .A2(KEYINPUT31), .ZN(new_n683));
  OAI21_X1  g0483(.A(G330), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g0484(.A(new_n684), .ZN(new_n685));
  OAI21_X1  g0485(.A(new_n657), .B1(new_n669), .B2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(KEYINPUT89), .B(new_n684), .C1(new_n658), .C2(new_n668), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n656), .B1(new_n688), .B2(G1), .ZN(G364));
  INV_X1    g0489(.A(new_n652), .ZN(new_n690));
  AOI21_X1  g0490(.A(new_n298), .B1(new_n620), .B2(G45), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n693), .B1(new_n633), .B2(G330), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n694), .B1(G330), .B2(new_n633), .ZN(new_n695));
  NOR2_X1   g0495(.A1(G13), .A2(G33), .ZN(new_n696));
  INV_X1    g0496(.A(new_n696), .ZN(new_n697));
  NOR2_X1   g0497(.A1(new_n697), .A2(G20), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n217), .B1(G20), .B2(new_n337), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  INV_X1    g0500(.A(new_n700), .ZN(new_n701));
  NOR2_X1   g0501(.A1(new_n246), .A2(new_n331), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n278), .A2(new_n283), .ZN(new_n703));
  NOR2_X1   g0503(.A1(new_n703), .A2(new_n651), .ZN(new_n704));
  INV_X1    g0504(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n705), .B1(new_n331), .B2(new_n216), .ZN(new_n706));
  INV_X1    g0506(.A(KEYINPUT90), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n702), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n707), .B2(new_n706), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n651), .A2(new_n261), .ZN(new_n710));
  AOI22_X1  g0510(.A1(new_n710), .A2(G355), .B1(new_n539), .B2(new_n651), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n701), .B1(new_n709), .B2(new_n711), .ZN(new_n712));
  NOR2_X1   g0512(.A1(new_n218), .A2(G179), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n713), .A2(G190), .A3(G200), .ZN(new_n714));
  INV_X1    g0514(.A(G303), .ZN(new_n715));
  NOR2_X1   g0515(.A1(G179), .A2(G200), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n218), .B1(new_n716), .B2(G190), .ZN(new_n717));
  INV_X1    g0517(.A(G294), .ZN(new_n718));
  OAI22_X1  g0518(.A1(new_n714), .A2(new_n715), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n218), .A2(new_n413), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n720), .A2(G200), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n721), .A2(new_n368), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  INV_X1    g0523(.A(G326), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n720), .ZN(new_n726));
  AOI21_X1  g0526(.A(G200), .B1(new_n726), .B2(KEYINPUT91), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(KEYINPUT91), .B2(new_n726), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n728), .A2(G190), .ZN(new_n729));
  AOI211_X1 g0529(.A(new_n719), .B(new_n725), .C1(new_n729), .C2(G311), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n716), .A2(G20), .A3(new_n368), .ZN(new_n731));
  OR2_X1    g0531(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n731), .A2(KEYINPUT92), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g0534(.A(new_n734), .ZN(new_n735));
  NAND2_X1  g0535(.A1(new_n735), .A2(G329), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n713), .A2(new_n368), .A3(G200), .ZN(new_n737));
  INV_X1    g0537(.A(G283), .ZN(new_n738));
  OAI21_X1  g0538(.A(new_n261), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g0539(.A(KEYINPUT33), .B(G317), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT93), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n721), .A2(G190), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n739), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n728), .A2(new_n368), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n744), .A2(G322), .ZN(new_n745));
  NAND4_X1  g0545(.A1(new_n730), .A2(new_n736), .A3(new_n743), .A4(new_n745), .ZN(new_n746));
  INV_X1    g0546(.A(new_n742), .ZN(new_n747));
  OAI22_X1  g0547(.A1(new_n747), .A2(new_n202), .B1(new_n717), .B2(new_n403), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n360), .B1(new_n723), .B2(new_n215), .ZN(new_n749));
  NOR2_X1   g0549(.A1(new_n714), .A2(new_n326), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n737), .A2(new_n422), .ZN(new_n751));
  NOR4_X1   g0551(.A1(new_n748), .A2(new_n749), .A3(new_n750), .A4(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n734), .A2(new_n256), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT32), .ZN(new_n754));
  AOI22_X1  g0554(.A1(G77), .A2(new_n729), .B1(new_n744), .B2(new_n306), .ZN(new_n755));
  NAND3_X1  g0555(.A1(new_n752), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n746), .A2(new_n756), .ZN(new_n757));
  AOI211_X1 g0557(.A(new_n692), .B(new_n712), .C1(new_n699), .C2(new_n757), .ZN(new_n758));
  INV_X1    g0558(.A(new_n698), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n758), .B1(new_n633), .B2(new_n759), .ZN(new_n760));
  AND2_X1   g0560(.A1(new_n695), .A2(new_n760), .ZN(new_n761));
  INV_X1    g0561(.A(new_n761), .ZN(G396));
  AND2_X1   g0562(.A1(new_n601), .A2(new_n597), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n626), .B1(new_n763), .B2(new_n595), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n626), .A2(new_n436), .ZN(new_n765));
  XNOR2_X1  g0565(.A(new_n765), .B(KEYINPUT95), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n440), .A2(new_n766), .ZN(new_n767));
  XNOR2_X1  g0567(.A(new_n767), .B(KEYINPUT96), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n604), .A2(new_n626), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n768), .A2(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n764), .A2(new_n770), .ZN(new_n771));
  INV_X1    g0571(.A(new_n768), .ZN(new_n772));
  AOI21_X1  g0572(.A(new_n771), .B1(new_n764), .B2(new_n772), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n693), .B1(new_n774), .B2(new_n684), .ZN(new_n775));
  OAI21_X1  g0575(.A(new_n775), .B1(new_n684), .B2(new_n774), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n699), .A2(new_n696), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n693), .B1(G77), .B2(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G137), .A2(new_n722), .B1(new_n742), .B2(G150), .ZN(new_n780));
  INV_X1    g0580(.A(new_n744), .ZN(new_n781));
  INV_X1    g0581(.A(G143), .ZN(new_n782));
  INV_X1    g0582(.A(new_n729), .ZN(new_n783));
  OAI221_X1 g0583(.A(new_n780), .B1(new_n781), .B2(new_n782), .C1(new_n256), .C2(new_n783), .ZN(new_n784));
  INV_X1    g0584(.A(KEYINPUT34), .ZN(new_n785));
  NAND2_X1  g0585(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  INV_X1    g0586(.A(new_n714), .ZN(new_n787));
  INV_X1    g0587(.A(new_n717), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n787), .A2(G50), .B1(new_n788), .B2(new_n306), .ZN(new_n789));
  INV_X1    g0589(.A(new_n737), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n790), .A2(G68), .ZN(new_n791));
  AND3_X1   g0591(.A1(new_n789), .A2(new_n703), .A3(new_n791), .ZN(new_n792));
  INV_X1    g0592(.A(G132), .ZN(new_n793));
  OAI211_X1 g0593(.A(new_n786), .B(new_n792), .C1(new_n793), .C2(new_n734), .ZN(new_n794));
  NOR2_X1   g0594(.A1(new_n784), .A2(new_n785), .ZN(new_n795));
  AOI22_X1  g0595(.A1(G283), .A2(new_n742), .B1(new_n722), .B2(G303), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n796), .B1(new_n783), .B2(new_n539), .ZN(new_n797));
  XOR2_X1   g0597(.A(new_n797), .B(KEYINPUT94), .Z(new_n798));
  NAND2_X1  g0598(.A1(new_n744), .A2(G294), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n735), .A2(G311), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n360), .B1(new_n788), .B2(G97), .ZN(new_n801));
  AOI22_X1  g0601(.A1(new_n787), .A2(G107), .B1(new_n790), .B2(G87), .ZN(new_n802));
  NAND4_X1  g0602(.A1(new_n799), .A2(new_n800), .A3(new_n801), .A4(new_n802), .ZN(new_n803));
  OAI22_X1  g0603(.A1(new_n794), .A2(new_n795), .B1(new_n798), .B2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n779), .B1(new_n804), .B2(new_n699), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n805), .B1(new_n770), .B2(new_n697), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n776), .A2(new_n806), .ZN(G384));
  OR2_X1    g0607(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n448), .A2(KEYINPUT35), .ZN(new_n809));
  NAND4_X1  g0609(.A1(new_n808), .A2(G116), .A3(new_n219), .A4(new_n809), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT36), .Z(new_n811));
  NAND3_X1  g0611(.A1(new_n216), .A2(G77), .A3(new_n252), .ZN(new_n812));
  AOI211_X1 g0612(.A(G13), .B(new_n302), .C1(new_n812), .C2(new_n242), .ZN(new_n813));
  NOR2_X1   g0613(.A1(new_n811), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(KEYINPUT39), .ZN(new_n815));
  XOR2_X1   g0615(.A(new_n624), .B(KEYINPUT98), .Z(new_n816));
  NAND3_X1  g0616(.A1(new_n313), .A2(new_n322), .A3(new_n816), .ZN(new_n817));
  AOI21_X1  g0617(.A(KEYINPUT37), .B1(new_n344), .B2(new_n348), .ZN(new_n818));
  NAND3_X1  g0618(.A1(new_n341), .A2(new_n817), .A3(new_n818), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT99), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  NAND4_X1  g0621(.A1(new_n341), .A2(new_n817), .A3(KEYINPUT99), .A4(new_n818), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NOR3_X1   g0623(.A1(new_n297), .A2(new_n312), .A3(new_n347), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NAND3_X1  g0625(.A1(new_n817), .A2(new_n825), .A3(new_n609), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n826), .A2(KEYINPUT37), .ZN(new_n827));
  NAND2_X1  g0627(.A1(new_n823), .A2(new_n827), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n817), .B1(new_n610), .B2(new_n352), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(KEYINPUT38), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n277), .A2(new_n292), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n314), .B1(new_n832), .B2(new_n265), .ZN(new_n833));
  AOI21_X1  g0633(.A(new_n312), .B1(new_n343), .B2(new_n833), .ZN(new_n834));
  OR3_X1    g0634(.A1(new_n834), .A2(KEYINPUT97), .A3(new_n624), .ZN(new_n835));
  OR2_X1    g0635(.A1(new_n834), .A2(new_n339), .ZN(new_n836));
  OAI21_X1  g0636(.A(KEYINPUT97), .B1(new_n834), .B2(new_n624), .ZN(new_n837));
  NAND4_X1  g0637(.A1(new_n835), .A2(new_n836), .A3(new_n825), .A4(new_n837), .ZN(new_n838));
  AOI22_X1  g0638(.A1(new_n821), .A2(new_n822), .B1(KEYINPUT37), .B2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n835), .A2(new_n837), .ZN(new_n840));
  AND2_X1   g0640(.A1(new_n355), .A2(new_n840), .ZN(new_n841));
  INV_X1    g0641(.A(KEYINPUT38), .ZN(new_n842));
  NOR3_X1   g0642(.A1(new_n839), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g0643(.A(new_n815), .B1(new_n831), .B2(new_n843), .ZN(new_n844));
  OR2_X1    g0644(.A1(new_n414), .A2(new_n415), .ZN(new_n845));
  NAND3_X1  g0645(.A1(new_n845), .A2(new_n401), .A3(new_n644), .ZN(new_n846));
  INV_X1    g0646(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n838), .A2(KEYINPUT37), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n823), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n355), .A2(new_n840), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n849), .A2(KEYINPUT38), .A3(new_n850), .ZN(new_n851));
  OAI21_X1  g0651(.A(new_n842), .B1(new_n839), .B2(new_n841), .ZN(new_n852));
  NAND3_X1  g0652(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT39), .ZN(new_n853));
  NAND3_X1  g0653(.A1(new_n844), .A2(new_n847), .A3(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n610), .A2(new_n816), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n851), .A2(new_n852), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n416), .A2(new_n418), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n401), .A2(new_n626), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n857), .A2(new_n859), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n416), .A2(new_n418), .A3(new_n858), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(new_n862), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n602), .A2(new_n644), .A3(new_n772), .ZN(new_n864));
  NOR2_X1   g0664(.A1(new_n437), .A2(new_n626), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n863), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  AOI21_X1  g0667(.A(new_n855), .B1(new_n856), .B2(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n854), .A2(new_n868), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n669), .A2(new_n356), .A3(new_n441), .ZN(new_n870));
  NAND2_X1  g0670(.A1(new_n870), .A2(new_n617), .ZN(new_n871));
  XNOR2_X1  g0671(.A(new_n869), .B(new_n871), .ZN(new_n872));
  INV_X1    g0672(.A(new_n856), .ZN(new_n873));
  INV_X1    g0673(.A(new_n683), .ZN(new_n874));
  AOI21_X1  g0674(.A(new_n680), .B1(new_n577), .B2(new_n644), .ZN(new_n875));
  OAI21_X1  g0675(.A(new_n874), .B1(new_n875), .B2(new_n670), .ZN(new_n876));
  INV_X1    g0676(.A(KEYINPUT40), .ZN(new_n877));
  NAND4_X1  g0677(.A1(new_n876), .A2(new_n877), .A3(new_n770), .A4(new_n862), .ZN(new_n878));
  OAI211_X1 g0678(.A(new_n862), .B(new_n770), .C1(new_n682), .C2(new_n683), .ZN(new_n879));
  AOI22_X1  g0679(.A1(new_n821), .A2(new_n822), .B1(KEYINPUT37), .B2(new_n826), .ZN(new_n880));
  OAI21_X1  g0680(.A(new_n842), .B1(new_n880), .B2(new_n829), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n879), .B1(new_n851), .B2(new_n881), .ZN(new_n882));
  OAI22_X1  g0682(.A1(new_n873), .A2(new_n878), .B1(new_n882), .B2(new_n877), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n883), .A2(new_n443), .A3(new_n876), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n878), .B1(new_n851), .B2(new_n852), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n851), .A2(new_n881), .ZN(new_n886));
  INV_X1    g0686(.A(new_n879), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  AOI21_X1  g0688(.A(new_n885), .B1(new_n888), .B2(KEYINPUT40), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n443), .A2(new_n876), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n884), .A2(new_n891), .A3(G330), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n872), .A2(new_n892), .ZN(new_n893));
  OAI21_X1  g0693(.A(new_n893), .B1(new_n302), .B2(new_n620), .ZN(new_n894));
  NOR2_X1   g0694(.A1(new_n872), .A2(new_n892), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n814), .B1(new_n894), .B2(new_n895), .ZN(G367));
  AOI22_X1  g0696(.A1(G50), .A2(new_n729), .B1(new_n744), .B2(G150), .ZN(new_n897));
  OAI22_X1  g0697(.A1(new_n723), .A2(new_n782), .B1(new_n363), .B2(new_n737), .ZN(new_n898));
  INV_X1    g0698(.A(new_n306), .ZN(new_n899));
  OAI22_X1  g0699(.A1(new_n747), .A2(new_n256), .B1(new_n714), .B2(new_n899), .ZN(new_n900));
  NOR2_X1   g0700(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n735), .A2(G137), .ZN(new_n902));
  AOI21_X1  g0702(.A(new_n261), .B1(new_n788), .B2(G68), .ZN(new_n903));
  NAND4_X1  g0703(.A1(new_n897), .A2(new_n901), .A3(new_n902), .A4(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n703), .ZN(new_n905));
  OAI21_X1  g0705(.A(new_n905), .B1(new_n422), .B2(new_n717), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n747), .A2(new_n718), .B1(new_n403), .B2(new_n737), .ZN(new_n907));
  AOI211_X1 g0707(.A(new_n906), .B(new_n907), .C1(G283), .C2(new_n729), .ZN(new_n908));
  AOI22_X1  g0708(.A1(new_n744), .A2(G303), .B1(G311), .B2(new_n722), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n910));
  AOI21_X1  g0710(.A(KEYINPUT46), .B1(new_n787), .B2(G116), .ZN(new_n911));
  AND3_X1   g0711(.A1(new_n787), .A2(KEYINPUT46), .A3(G116), .ZN(new_n912));
  XNOR2_X1  g0712(.A(KEYINPUT105), .B(G317), .ZN(new_n913));
  AOI211_X1 g0713(.A(new_n911), .B(new_n912), .C1(new_n735), .C2(new_n913), .ZN(new_n914));
  NAND3_X1  g0714(.A1(new_n908), .A2(new_n910), .A3(new_n914), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n909), .A2(KEYINPUT104), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n904), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  XNOR2_X1  g0717(.A(new_n917), .B(KEYINPUT47), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(new_n699), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n701), .B1(new_n651), .B2(new_n558), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n237), .A2(new_n704), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n692), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n588), .B1(new_n570), .B2(new_n644), .ZN(new_n923));
  OR3_X1    g0723(.A1(new_n593), .A2(new_n570), .A3(new_n644), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  OAI211_X1 g0725(.A(new_n919), .B(new_n922), .C1(new_n925), .C2(new_n759), .ZN(new_n926));
  XNOR2_X1  g0726(.A(new_n691), .B(KEYINPUT103), .ZN(new_n927));
  INV_X1    g0727(.A(new_n927), .ZN(new_n928));
  XNOR2_X1  g0728(.A(new_n639), .B(new_n646), .ZN(new_n929));
  XNOR2_X1  g0729(.A(new_n929), .B(new_n634), .ZN(new_n930));
  INV_X1    g0730(.A(new_n930), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n626), .B1(new_n663), .B2(new_n667), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n932), .A2(KEYINPUT29), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n933), .B1(new_n764), .B2(KEYINPUT29), .ZN(new_n934));
  AOI21_X1  g0734(.A(KEYINPUT89), .B1(new_n934), .B2(new_n684), .ZN(new_n935));
  INV_X1    g0735(.A(new_n687), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n931), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g0737(.A(KEYINPUT44), .ZN(new_n938));
  OAI211_X1 g0738(.A(new_n487), .B(new_n494), .C1(new_n459), .C2(new_n644), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n579), .A2(new_n626), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  OAI21_X1  g0741(.A(new_n938), .B1(new_n649), .B2(new_n941), .ZN(new_n942));
  OAI22_X1  g0742(.A1(new_n637), .A2(new_n645), .B1(new_n599), .B2(new_n626), .ZN(new_n943));
  INV_X1    g0743(.A(new_n941), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n943), .A2(new_n944), .A3(KEYINPUT44), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n942), .A2(new_n945), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT45), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n947), .B1(new_n943), .B2(new_n944), .ZN(new_n948));
  NAND3_X1  g0748(.A1(new_n649), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n946), .A2(new_n950), .ZN(new_n951));
  INV_X1    g0751(.A(KEYINPUT101), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n953), .A2(new_n642), .ZN(new_n954));
  AOI21_X1  g0754(.A(KEYINPUT101), .B1(new_n946), .B2(new_n950), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n641), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n954), .A2(new_n956), .ZN(new_n957));
  NOR3_X1   g0757(.A1(new_n937), .A2(new_n957), .A3(KEYINPUT102), .ZN(new_n958));
  INV_X1    g0758(.A(KEYINPUT102), .ZN(new_n959));
  AOI21_X1  g0759(.A(new_n930), .B1(new_n686), .B2(new_n687), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n955), .B(new_n642), .ZN(new_n961));
  AOI21_X1  g0761(.A(new_n959), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n688), .B1(new_n958), .B2(new_n962), .ZN(new_n963));
  XOR2_X1   g0763(.A(new_n652), .B(KEYINPUT41), .Z(new_n964));
  INV_X1    g0764(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g0765(.A(new_n928), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n641), .A2(new_n941), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n967), .B(KEYINPUT100), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n639), .A2(new_n646), .A3(new_n941), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n970));
  AND2_X1   g0770(.A1(new_n487), .A2(new_n635), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n644), .B1(new_n971), .B2(new_n579), .ZN(new_n972));
  NAND2_X1  g0772(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n969), .A2(KEYINPUT42), .ZN(new_n974));
  INV_X1    g0774(.A(KEYINPUT43), .ZN(new_n975));
  INV_X1    g0775(.A(new_n925), .ZN(new_n976));
  OAI22_X1  g0776(.A1(new_n973), .A2(new_n974), .B1(new_n975), .B2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n976), .A2(new_n975), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(new_n978), .ZN(new_n979));
  OR2_X1    g0779(.A1(new_n977), .A2(new_n978), .ZN(new_n980));
  AND3_X1   g0780(.A1(new_n968), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n968), .B1(new_n980), .B2(new_n979), .ZN(new_n982));
  NOR2_X1   g0782(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  INV_X1    g0783(.A(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n926), .B1(new_n966), .B2(new_n984), .ZN(G387));
  NAND3_X1  g0785(.A1(new_n686), .A2(new_n687), .A3(new_n930), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n937), .A2(new_n652), .A3(new_n986), .ZN(new_n987));
  NOR2_X1   g0787(.A1(new_n714), .A2(new_n363), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n788), .A2(new_n558), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n989), .B1(new_n723), .B2(new_n256), .ZN(new_n990));
  AOI211_X1 g0790(.A(new_n988), .B(new_n990), .C1(G50), .C2(new_n744), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n703), .B1(new_n403), .B2(new_n737), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n992), .B1(new_n307), .B2(new_n742), .ZN(new_n993));
  NAND2_X1  g0793(.A1(new_n735), .A2(G150), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n729), .A2(G68), .ZN(new_n995));
  NAND4_X1  g0795(.A1(new_n991), .A2(new_n993), .A3(new_n994), .A4(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n703), .B1(G116), .B2(new_n790), .ZN(new_n997));
  NAND2_X1  g0797(.A1(new_n744), .A2(new_n913), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G311), .A2(new_n742), .B1(new_n722), .B2(G322), .ZN(new_n999));
  OAI211_X1 g0799(.A(new_n998), .B(new_n999), .C1(new_n783), .C2(new_n715), .ZN(new_n1000));
  INV_X1    g0800(.A(KEYINPUT48), .ZN(new_n1001));
  OR2_X1    g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n787), .A2(G294), .B1(new_n788), .B2(G283), .ZN(new_n1004));
  NAND3_X1  g0804(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT49), .ZN(new_n1006));
  OAI221_X1 g0806(.A(new_n997), .B1(new_n724), .B2(new_n734), .C1(new_n1005), .C2(new_n1006), .ZN(new_n1007));
  AND2_X1   g0807(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n996), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1009), .A2(new_n699), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n639), .A2(new_n759), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n234), .A2(G45), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(KEYINPUT106), .ZN(new_n1013));
  AND2_X1   g0813(.A1(new_n653), .A2(KEYINPUT107), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n653), .A2(KEYINPUT107), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n331), .B1(new_n202), .B2(new_n363), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n1014), .A2(new_n1015), .A3(new_n1016), .ZN(new_n1017));
  INV_X1    g0817(.A(KEYINPUT108), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n1017), .A2(new_n1018), .ZN(new_n1019));
  NOR2_X1   g0819(.A1(new_n430), .A2(G50), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT50), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n1017), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n1021), .B1(new_n1022), .B2(KEYINPUT108), .ZN(new_n1023));
  OAI211_X1 g0823(.A(new_n1013), .B(new_n704), .C1(new_n1019), .C2(new_n1023), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n710), .A2(new_n653), .B1(new_n422), .B2(new_n651), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n701), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1026));
  NOR3_X1   g0826(.A1(new_n1011), .A2(new_n692), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g0827(.A1(new_n931), .A2(new_n928), .B1(new_n1010), .B2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n987), .A2(new_n1028), .ZN(G393));
  XNOR2_X1  g0829(.A(new_n951), .B(new_n642), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n652), .B1(new_n960), .B2(new_n1030), .ZN(new_n1031));
  OAI21_X1  g0831(.A(KEYINPUT102), .B1(new_n937), .B2(new_n957), .ZN(new_n1032));
  NAND3_X1  g0832(.A1(new_n960), .A2(new_n961), .A3(new_n959), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n1031), .B1(new_n1032), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n928), .ZN(new_n1035));
  OAI221_X1 g0835(.A(new_n700), .B1(new_n403), .B2(new_n211), .C1(new_n705), .C2(new_n241), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1036), .A2(new_n693), .ZN(new_n1037));
  XNOR2_X1  g0837(.A(new_n1037), .B(KEYINPUT109), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(new_n744), .A2(G159), .B1(G150), .B2(new_n722), .ZN(new_n1039));
  XOR2_X1   g0839(.A(new_n1039), .B(KEYINPUT51), .Z(new_n1040));
  OAI21_X1  g0840(.A(new_n703), .B1(new_n326), .B2(new_n737), .ZN(new_n1041));
  NAND2_X1  g0841(.A1(new_n788), .A2(G77), .ZN(new_n1042));
  OAI221_X1 g0842(.A(new_n1042), .B1(new_n202), .B2(new_n714), .C1(new_n747), .C2(new_n215), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(G143), .C2(new_n735), .ZN(new_n1044));
  OAI211_X1 g0844(.A(new_n1040), .B(new_n1044), .C1(new_n430), .C2(new_n783), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT110), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n1045), .A2(KEYINPUT110), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n744), .A2(G311), .B1(G317), .B2(new_n722), .ZN(new_n1048));
  XOR2_X1   g0848(.A(new_n1048), .B(KEYINPUT52), .Z(new_n1049));
  AND2_X1   g0849(.A1(new_n735), .A2(G322), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n742), .A2(G303), .B1(G116), .B2(new_n788), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n738), .B2(new_n714), .ZN(new_n1052));
  NOR4_X1   g0852(.A1(new_n1050), .A2(new_n1052), .A3(new_n360), .A4(new_n751), .ZN(new_n1053));
  OAI211_X1 g0853(.A(new_n1049), .B(new_n1053), .C1(new_n718), .C2(new_n783), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1046), .A2(new_n1047), .A3(new_n1054), .ZN(new_n1055));
  AOI21_X1  g0855(.A(new_n1038), .B1(new_n1055), .B2(new_n699), .ZN(new_n1056));
  OAI21_X1  g0856(.A(new_n1056), .B1(new_n941), .B2(new_n759), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1035), .A2(new_n1057), .ZN(new_n1058));
  NOR2_X1   g0858(.A1(new_n1034), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(G390));
  NAND4_X1  g0860(.A1(new_n876), .A2(G330), .A3(new_n770), .A4(new_n862), .ZN(new_n1061));
  INV_X1    g0861(.A(new_n1061), .ZN(new_n1062));
  NOR2_X1   g0862(.A1(new_n867), .A2(new_n847), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1063), .B1(new_n844), .B2(new_n853), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n865), .B1(new_n932), .B2(new_n772), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n846), .B1(new_n1065), .B2(new_n863), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n1066), .B1(new_n851), .B2(new_n881), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1062), .B1(new_n1064), .B2(new_n1067), .ZN(new_n1068));
  AND3_X1   g0868(.A1(new_n851), .A2(new_n852), .A3(KEYINPUT39), .ZN(new_n1069));
  AOI21_X1  g0869(.A(KEYINPUT39), .B1(new_n851), .B2(new_n881), .ZN(new_n1070));
  OAI22_X1  g0870(.A1(new_n1069), .A2(new_n1070), .B1(new_n847), .B2(new_n867), .ZN(new_n1071));
  OAI211_X1 g0871(.A(new_n886), .B(new_n846), .C1(new_n863), .C2(new_n1065), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1071), .A2(new_n1061), .A3(new_n1072), .ZN(new_n1073));
  OAI211_X1 g0873(.A(G330), .B(new_n770), .C1(new_n682), .C2(new_n683), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n863), .ZN(new_n1075));
  NAND3_X1  g0875(.A1(new_n1075), .A2(new_n1061), .A3(new_n1065), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  AOI22_X1  g0877(.A1(new_n1075), .A2(new_n1061), .B1(new_n864), .B2(new_n866), .ZN(new_n1078));
  NOR2_X1   g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n356), .A2(new_n685), .A3(new_n441), .ZN(new_n1080));
  NAND3_X1  g0880(.A1(new_n870), .A2(new_n617), .A3(new_n1080), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g0882(.A1(new_n1068), .A2(new_n1073), .A3(new_n1082), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n1083), .A2(KEYINPUT111), .ZN(new_n1084));
  INV_X1    g0884(.A(KEYINPUT111), .ZN(new_n1085));
  NAND4_X1  g0885(.A1(new_n1068), .A2(new_n1073), .A3(new_n1082), .A4(new_n1085), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1084), .A2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1088));
  AND3_X1   g0888(.A1(new_n870), .A2(new_n617), .A3(new_n1080), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1075), .A2(new_n1061), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n864), .A2(new_n866), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1090), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1092), .A2(new_n1076), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1094));
  AOI21_X1  g0894(.A(new_n690), .B1(new_n1088), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n1087), .A2(new_n1095), .ZN(new_n1096));
  OAI21_X1  g0896(.A(new_n696), .B1(new_n1069), .B2(new_n1070), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n693), .B1(new_n307), .B2(new_n778), .ZN(new_n1098));
  AOI22_X1  g0898(.A1(G107), .A2(new_n742), .B1(new_n722), .B2(G283), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n1099), .B1(new_n783), .B2(new_n403), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT112), .ZN(new_n1101));
  INV_X1    g0901(.A(new_n750), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1102), .A2(new_n791), .A3(new_n261), .A4(new_n1042), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1103), .B1(G294), .B2(new_n735), .ZN(new_n1104));
  OAI211_X1 g0904(.A(new_n1101), .B(new_n1104), .C1(new_n539), .C2(new_n781), .ZN(new_n1105));
  NOR2_X1   g0905(.A1(new_n1100), .A2(KEYINPUT112), .ZN(new_n1106));
  NAND2_X1  g0906(.A1(new_n735), .A2(G125), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n742), .A2(G137), .B1(G159), .B2(new_n788), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n722), .A2(G128), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n261), .B1(new_n790), .B2(G50), .ZN(new_n1110));
  NAND4_X1  g0910(.A1(new_n1107), .A2(new_n1108), .A3(new_n1109), .A4(new_n1110), .ZN(new_n1111));
  XOR2_X1   g0911(.A(KEYINPUT54), .B(G143), .Z(new_n1112));
  NAND2_X1  g0912(.A1(new_n729), .A2(new_n1112), .ZN(new_n1113));
  AOI21_X1  g0913(.A(KEYINPUT53), .B1(new_n787), .B2(G150), .ZN(new_n1114));
  AND3_X1   g0914(.A1(new_n787), .A2(KEYINPUT53), .A3(G150), .ZN(new_n1115));
  OAI221_X1 g0915(.A(new_n1113), .B1(new_n1114), .B2(new_n1115), .C1(new_n781), .C2(new_n793), .ZN(new_n1116));
  OAI22_X1  g0916(.A1(new_n1105), .A2(new_n1106), .B1(new_n1111), .B2(new_n1116), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1098), .B1(new_n1117), .B2(new_n699), .ZN(new_n1118));
  AND2_X1   g0918(.A1(new_n1097), .A2(new_n1118), .ZN(new_n1119));
  XNOR2_X1  g0919(.A(new_n1119), .B(KEYINPUT113), .ZN(new_n1120));
  NOR2_X1   g0920(.A1(new_n1088), .A2(new_n927), .ZN(new_n1121));
  NOR2_X1   g0921(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1096), .A2(new_n1122), .ZN(G378));
  INV_X1    g0923(.A(KEYINPUT57), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n624), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n378), .A2(new_n1126), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n1127), .B1(new_n384), .B2(new_n390), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n1128), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n384), .A2(new_n390), .A3(new_n1127), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1125), .B1(new_n1129), .B2(new_n1130), .ZN(new_n1131));
  INV_X1    g0931(.A(new_n1130), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1125), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1132), .A2(new_n1128), .A3(new_n1133), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n1131), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g0935(.A(G330), .ZN(new_n1136));
  OAI21_X1  g0936(.A(new_n1135), .B1(new_n889), .B2(new_n1136), .ZN(new_n1137));
  INV_X1    g0937(.A(KEYINPUT116), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n1138), .B1(new_n1131), .B2(new_n1134), .ZN(new_n1139));
  OAI21_X1  g0939(.A(new_n1133), .B1(new_n1132), .B2(new_n1128), .ZN(new_n1140));
  NAND3_X1  g0940(.A1(new_n1129), .A2(new_n1130), .A3(new_n1125), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1140), .A2(new_n1141), .A3(KEYINPUT116), .ZN(new_n1142));
  NAND2_X1  g0942(.A1(new_n1139), .A2(new_n1142), .ZN(new_n1143));
  AOI21_X1  g0943(.A(new_n877), .B1(new_n886), .B2(new_n887), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n1143), .C1(new_n1144), .C2(new_n885), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n869), .A2(KEYINPUT117), .ZN(new_n1147));
  INV_X1    g0947(.A(KEYINPUT117), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n854), .A2(new_n1148), .A3(new_n868), .ZN(new_n1149));
  NAND4_X1  g0949(.A1(new_n1146), .A2(KEYINPUT118), .A3(new_n1147), .A4(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1145), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1135), .ZN(new_n1152));
  AOI21_X1  g0952(.A(new_n1152), .B1(new_n883), .B2(G330), .ZN(new_n1153));
  NOR2_X1   g0953(.A1(new_n1151), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1147), .A2(new_n1149), .ZN(new_n1155));
  NOR2_X1   g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n869), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1137), .A2(new_n1157), .A3(new_n1145), .ZN(new_n1158));
  INV_X1    g0958(.A(KEYINPUT118), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  OAI21_X1  g0960(.A(new_n1150), .B1(new_n1156), .B2(new_n1160), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1081), .B1(new_n1084), .B2(new_n1086), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1124), .B1(new_n1161), .B2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1164));
  INV_X1    g0964(.A(KEYINPUT119), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1157), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n1166), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1124), .B1(new_n1167), .B2(new_n1158), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NOR3_X1   g0969(.A1(new_n1151), .A2(new_n1153), .A3(new_n869), .ZN(new_n1170));
  OAI21_X1  g0970(.A(KEYINPUT57), .B1(new_n1170), .B2(new_n1166), .ZN(new_n1171));
  OAI21_X1  g0971(.A(KEYINPUT119), .B1(new_n1162), .B2(new_n1171), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1163), .A2(new_n1169), .A3(new_n652), .A4(new_n1172), .ZN(new_n1173));
  NOR2_X1   g0973(.A1(new_n1161), .A2(new_n927), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n722), .A2(G125), .ZN(new_n1175));
  AOI22_X1  g0975(.A1(G128), .A2(new_n744), .B1(new_n729), .B2(G137), .ZN(new_n1176));
  AOI22_X1  g0976(.A1(new_n742), .A2(G132), .B1(G150), .B2(new_n788), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n787), .A2(new_n1112), .ZN(new_n1178));
  XOR2_X1   g0978(.A(new_n1178), .B(KEYINPUT115), .Z(new_n1179));
  AND4_X1   g0979(.A1(new_n1175), .A2(new_n1176), .A3(new_n1177), .A4(new_n1179), .ZN(new_n1180));
  INV_X1    g0980(.A(new_n1180), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n735), .A2(G124), .ZN(new_n1183));
  AOI211_X1 g0983(.A(G33), .B(G41), .C1(new_n790), .C2(G159), .ZN(new_n1184));
  AND3_X1   g0984(.A1(new_n1182), .A2(new_n1183), .A3(new_n1184), .ZN(new_n1185));
  OR2_X1    g0985(.A1(new_n1181), .A2(KEYINPUT59), .ZN(new_n1186));
  OAI22_X1  g0986(.A1(new_n723), .A2(new_n539), .B1(new_n737), .B2(new_n899), .ZN(new_n1187));
  AOI211_X1 g0987(.A(new_n988), .B(new_n1187), .C1(G68), .C2(new_n788), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n735), .A2(G283), .ZN(new_n1189));
  NOR2_X1   g0989(.A1(new_n703), .A2(G41), .ZN(new_n1190));
  NAND3_X1  g0990(.A1(new_n1188), .A2(new_n1189), .A3(new_n1190), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(new_n729), .A2(new_n558), .B1(G97), .B2(new_n742), .ZN(new_n1192));
  XNOR2_X1  g0992(.A(new_n1192), .B(KEYINPUT114), .ZN(new_n1193));
  AOI211_X1 g0993(.A(new_n1191), .B(new_n1193), .C1(G107), .C2(new_n744), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n1185), .A2(new_n1186), .B1(KEYINPUT58), .B2(new_n1194), .ZN(new_n1195));
  OAI21_X1  g0995(.A(new_n215), .B1(G33), .B2(G41), .ZN(new_n1196));
  OAI221_X1 g0996(.A(new_n1195), .B1(KEYINPUT58), .B2(new_n1194), .C1(new_n1190), .C2(new_n1196), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1197), .A2(new_n699), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n692), .B1(new_n215), .B2(new_n777), .ZN(new_n1199));
  OAI211_X1 g0999(.A(new_n1198), .B(new_n1199), .C1(new_n1143), .C2(new_n697), .ZN(new_n1200));
  INV_X1    g1000(.A(new_n1200), .ZN(new_n1201));
  NOR2_X1   g1001(.A1(new_n1174), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1173), .A2(new_n1202), .ZN(G375));
  NOR2_X1   g1003(.A1(new_n1089), .A2(new_n1093), .ZN(new_n1204));
  XOR2_X1   g1004(.A(new_n964), .B(KEYINPUT120), .Z(new_n1205));
  NOR3_X1   g1005(.A1(new_n1082), .A2(new_n1204), .A3(new_n1205), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n862), .A2(new_n697), .ZN(new_n1208));
  XNOR2_X1  g1008(.A(new_n1208), .B(KEYINPUT122), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n742), .A2(new_n1112), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1210), .B1(new_n723), .B2(new_n793), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n729), .A2(G150), .ZN(new_n1212));
  OAI22_X1  g1012(.A1(new_n714), .A2(new_n256), .B1(new_n717), .B2(new_n215), .ZN(new_n1213));
  AOI211_X1 g1013(.A(new_n1213), .B(new_n905), .C1(new_n306), .C2(new_n790), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n735), .A2(G128), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1212), .A2(new_n1214), .A3(new_n1215), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT123), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1211), .B(new_n1217), .C1(G137), .C2(new_n744), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n422), .A2(new_n783), .B1(new_n781), .B2(new_n738), .ZN(new_n1219));
  AOI22_X1  g1019(.A1(new_n722), .A2(G294), .B1(new_n787), .B2(G97), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1220), .B(new_n989), .C1(new_n539), .C2(new_n747), .ZN(new_n1221));
  OAI221_X1 g1021(.A(new_n261), .B1(new_n363), .B2(new_n737), .C1(new_n734), .C2(new_n715), .ZN(new_n1222));
  NOR3_X1   g1022(.A1(new_n1219), .A2(new_n1221), .A3(new_n1222), .ZN(new_n1223));
  OAI21_X1  g1023(.A(new_n699), .B1(new_n1218), .B2(new_n1223), .ZN(new_n1224));
  OAI211_X1 g1024(.A(new_n1224), .B(new_n693), .C1(G68), .C2(new_n778), .ZN(new_n1225));
  NOR2_X1   g1025(.A1(new_n1209), .A2(new_n1225), .ZN(new_n1226));
  AOI21_X1  g1026(.A(new_n1226), .B1(new_n1093), .B2(new_n928), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1207), .A2(new_n1227), .ZN(G381));
  INV_X1    g1028(.A(G378), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1173), .A2(new_n1229), .A3(new_n1202), .ZN(new_n1230));
  INV_X1    g1030(.A(new_n1230), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1032), .A2(new_n1033), .B1(new_n686), .B2(new_n687), .ZN(new_n1232));
  OAI21_X1  g1032(.A(new_n927), .B1(new_n1232), .B2(new_n964), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n983), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n987), .A2(new_n761), .A3(new_n1028), .ZN(new_n1235));
  NOR4_X1   g1035(.A1(G381), .A2(G384), .A3(G390), .A4(new_n1235), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1231), .A2(new_n1234), .A3(new_n926), .A4(new_n1236), .ZN(G407));
  OAI211_X1 g1037(.A(G407), .B(G213), .C1(G343), .C2(new_n1230), .ZN(G409));
  NAND2_X1  g1038(.A1(G393), .A2(G396), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1239), .A2(new_n1235), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1059), .A2(new_n1240), .ZN(new_n1241));
  OAI211_X1 g1041(.A(new_n1239), .B(new_n1235), .C1(new_n1034), .C2(new_n1058), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1241), .A2(new_n1242), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT126), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1244), .B1(new_n1234), .B2(new_n926), .ZN(new_n1245));
  INV_X1    g1045(.A(new_n926), .ZN(new_n1246));
  AOI211_X1 g1046(.A(KEYINPUT126), .B(new_n1246), .C1(new_n1233), .C2(new_n983), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1243), .B1(new_n1245), .B2(new_n1247), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(G387), .A2(KEYINPUT126), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1234), .A2(new_n1244), .A3(new_n926), .ZN(new_n1250));
  NAND4_X1  g1050(.A1(new_n1249), .A2(new_n1250), .A3(new_n1242), .A4(new_n1241), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1248), .A2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  INV_X1    g1053(.A(KEYINPUT124), .ZN(new_n1254));
  AOI21_X1  g1054(.A(new_n1204), .B1(KEYINPUT60), .B2(new_n1094), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1079), .A2(KEYINPUT60), .A3(new_n1081), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1256), .A2(new_n652), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1227), .B1(new_n1255), .B2(new_n1257), .ZN(new_n1258));
  INV_X1    g1058(.A(G384), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n1254), .B1(new_n1258), .B2(new_n1259), .ZN(new_n1260));
  AND2_X1   g1060(.A1(new_n1256), .A2(new_n652), .ZN(new_n1261));
  AND2_X1   g1061(.A1(new_n1094), .A2(KEYINPUT60), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1261), .B1(new_n1262), .B2(new_n1204), .ZN(new_n1263));
  NAND4_X1  g1063(.A1(new_n1263), .A2(KEYINPUT124), .A3(G384), .A4(new_n1227), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1258), .A2(new_n1259), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1260), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND3_X1  g1066(.A1(new_n625), .A2(G213), .A3(G2897), .ZN(new_n1267));
  INV_X1    g1067(.A(new_n1267), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n1266), .A2(new_n1268), .ZN(new_n1269));
  NAND4_X1  g1069(.A1(new_n1260), .A2(new_n1265), .A3(new_n1264), .A4(new_n1267), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  INV_X1    g1071(.A(new_n1271), .ZN(new_n1272));
  AOI21_X1  g1072(.A(new_n1229), .B1(new_n1173), .B2(new_n1202), .ZN(new_n1273));
  NAND2_X1  g1073(.A1(new_n625), .A2(G213), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1167), .A2(new_n1158), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1201), .B1(new_n1275), .B2(new_n928), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1276), .A2(new_n1096), .A3(new_n1122), .ZN(new_n1277));
  NOR3_X1   g1077(.A1(new_n1161), .A2(new_n1162), .A3(new_n1205), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1274), .B1(new_n1277), .B2(new_n1278), .ZN(new_n1279));
  OAI21_X1  g1079(.A(new_n1272), .B1(new_n1273), .B2(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1273), .A2(new_n1266), .A3(new_n1279), .ZN(new_n1281));
  INV_X1    g1081(.A(KEYINPUT62), .ZN(new_n1282));
  OAI211_X1 g1082(.A(new_n1253), .B(new_n1280), .C1(new_n1281), .C2(new_n1282), .ZN(new_n1283));
  NOR4_X1   g1083(.A1(new_n1273), .A2(KEYINPUT62), .A3(new_n1279), .A4(new_n1266), .ZN(new_n1284));
  OAI21_X1  g1084(.A(new_n1252), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1285));
  NOR2_X1   g1085(.A1(new_n1273), .A2(new_n1279), .ZN(new_n1286));
  NAND2_X1  g1086(.A1(new_n1271), .A2(KEYINPUT125), .ZN(new_n1287));
  INV_X1    g1087(.A(KEYINPUT125), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1269), .A2(new_n1288), .A3(new_n1270), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1287), .A2(new_n1289), .ZN(new_n1290));
  OAI21_X1  g1090(.A(KEYINPUT63), .B1(new_n1286), .B2(new_n1290), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1281), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1291), .A2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1248), .A2(new_n1251), .A3(new_n1253), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(KEYINPUT127), .ZN(new_n1295));
  INV_X1    g1095(.A(KEYINPUT127), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1248), .A2(new_n1251), .A3(new_n1296), .A4(new_n1253), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1295), .A2(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1298), .B1(KEYINPUT63), .B2(new_n1281), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(new_n1293), .A2(new_n1299), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1285), .A2(new_n1300), .ZN(G405));
  INV_X1    g1101(.A(new_n1266), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1302), .B1(new_n1231), .B2(new_n1273), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1273), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1304), .A2(new_n1230), .A3(new_n1266), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1303), .A2(new_n1305), .ZN(new_n1306));
  INV_X1    g1106(.A(new_n1252), .ZN(new_n1307));
  XNOR2_X1  g1107(.A(new_n1306), .B(new_n1307), .ZN(G402));
endmodule


