//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 1 0 0 0 1 0 0 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 0 0 0 1 0 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:07 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n715, new_n716, new_n718, new_n719, new_n720,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n755, new_n756, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n970, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1040, new_n1041, new_n1042,
    new_n1043, new_n1044, new_n1045, new_n1046, new_n1047, new_n1048,
    new_n1049, new_n1050, new_n1051, new_n1052, new_n1054, new_n1055,
    new_n1056, new_n1057, new_n1058, new_n1059, new_n1060, new_n1061,
    new_n1062, new_n1063, new_n1064;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT3), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(KEYINPUT73), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT73), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n191), .A2(KEYINPUT3), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(G107), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(G104), .ZN(new_n197));
  INV_X1    g011(.A(G104), .ZN(new_n198));
  NOR2_X1   g012(.A1(new_n198), .A2(G107), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n192), .B1(new_n197), .B2(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G101), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n196), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  XNOR2_X1  g016(.A(G143), .B(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  NOR2_X1   g018(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G143), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n207), .B(G146), .C1(new_n204), .C2(KEYINPUT1), .ZN(new_n208));
  INV_X1    g022(.A(G146), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n204), .A2(new_n209), .A3(G143), .ZN(new_n210));
  NAND3_X1  g024(.A1(new_n206), .A2(new_n208), .A3(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n198), .A2(G107), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(new_n195), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G101), .ZN(new_n214));
  NAND3_X1  g028(.A1(new_n202), .A2(new_n211), .A3(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(new_n214), .ZN(new_n216));
  AOI22_X1  g030(.A1(new_n195), .A2(new_n193), .B1(new_n213), .B2(new_n192), .ZN(new_n217));
  AOI21_X1  g031(.A(new_n216), .B1(new_n217), .B2(new_n201), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n208), .A2(new_n210), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(KEYINPUT65), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT65), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n208), .A2(new_n221), .A3(new_n210), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n220), .A2(new_n222), .A3(new_n206), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n215), .B1(new_n218), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(KEYINPUT64), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT64), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G134), .ZN(new_n228));
  INV_X1    g042(.A(G137), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT11), .ZN(new_n230));
  NAND3_X1  g044(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(G131), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n229), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  INV_X1    g047(.A(KEYINPUT11), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n234), .A2(G137), .ZN(new_n235));
  NAND4_X1  g049(.A1(new_n231), .A2(new_n232), .A3(new_n233), .A4(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(new_n236), .ZN(new_n237));
  AND2_X1   g051(.A1(new_n233), .A2(new_n235), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n232), .B1(new_n238), .B2(new_n231), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n237), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n240), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n224), .A2(KEYINPUT75), .A3(KEYINPUT12), .A4(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n202), .A2(new_n214), .ZN(new_n243));
  AND3_X1   g057(.A1(new_n208), .A2(new_n221), .A3(new_n210), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n221), .B1(new_n208), .B2(new_n210), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n209), .A2(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n207), .A2(G146), .ZN(new_n247));
  AND3_X1   g061(.A1(new_n205), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NOR3_X1   g062(.A1(new_n244), .A2(new_n245), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n243), .A2(new_n249), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n240), .B1(new_n250), .B2(new_n215), .ZN(new_n251));
  OAI21_X1  g065(.A(new_n242), .B1(KEYINPUT12), .B2(new_n251), .ZN(new_n252));
  AOI21_X1  g066(.A(KEYINPUT75), .B1(new_n251), .B2(KEYINPUT12), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n199), .B1(new_n190), .B2(new_n192), .ZN(new_n255));
  AOI22_X1  g069(.A1(new_n212), .A2(new_n195), .B1(new_n191), .B2(KEYINPUT3), .ZN(new_n256));
  OAI21_X1  g070(.A(G101), .B1(new_n255), .B2(new_n256), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n257), .A2(new_n202), .A3(KEYINPUT4), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n246), .A2(new_n247), .ZN(new_n259));
  INV_X1    g073(.A(KEYINPUT0), .ZN(new_n260));
  NOR2_X1   g074(.A1(new_n260), .A2(new_n204), .ZN(new_n261));
  NOR2_X1   g075(.A1(KEYINPUT0), .A2(G128), .ZN(new_n262));
  OAI21_X1  g076(.A(new_n259), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI211_X1 g077(.A(new_n246), .B(new_n247), .C1(new_n260), .C2(new_n204), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT4), .ZN(new_n266));
  OAI211_X1 g080(.A(new_n266), .B(G101), .C1(new_n255), .C2(new_n256), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n258), .A2(new_n265), .A3(new_n267), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT10), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n215), .A2(new_n269), .ZN(new_n270));
  AND2_X1   g084(.A1(new_n268), .A2(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n223), .A2(KEYINPUT10), .ZN(new_n272));
  OAI21_X1  g086(.A(KEYINPUT74), .B1(new_n272), .B2(new_n243), .ZN(new_n273));
  INV_X1    g087(.A(KEYINPUT74), .ZN(new_n274));
  NAND4_X1  g088(.A1(new_n218), .A2(new_n274), .A3(KEYINPUT10), .A4(new_n223), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n273), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g090(.A1(new_n271), .A2(new_n276), .A3(new_n240), .ZN(new_n277));
  INV_X1    g091(.A(G953), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(G227), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n279), .B(KEYINPUT71), .ZN(new_n280));
  XNOR2_X1  g094(.A(G110), .B(G140), .ZN(new_n281));
  XNOR2_X1  g095(.A(new_n280), .B(new_n281), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n277), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g097(.A1(new_n254), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n271), .A2(new_n276), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n285), .A2(new_n241), .ZN(new_n286));
  AOI21_X1  g100(.A(new_n282), .B1(new_n286), .B2(new_n277), .ZN(new_n287));
  OAI211_X1 g101(.A(new_n187), .B(new_n188), .C1(new_n284), .C2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(G469), .A2(G902), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n277), .B1(new_n252), .B2(new_n253), .ZN(new_n290));
  XOR2_X1   g104(.A(new_n282), .B(KEYINPUT72), .Z(new_n291));
  NAND2_X1  g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n286), .A2(new_n277), .A3(new_n282), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n292), .A2(G469), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n288), .A2(new_n289), .A3(new_n294), .ZN(new_n295));
  XNOR2_X1  g109(.A(KEYINPUT9), .B(G234), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  OAI21_X1  g112(.A(G214), .B1(G237), .B2(G902), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(G119), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n301), .A2(G116), .ZN(new_n302));
  INV_X1    g116(.A(G116), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n303), .A2(G119), .ZN(new_n304));
  INV_X1    g118(.A(G113), .ZN(new_n305));
  AND2_X1   g119(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n306));
  NOR2_X1   g120(.A1(new_n305), .A2(KEYINPUT2), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n302), .B(new_n304), .C1(new_n306), .C2(new_n307), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n302), .A2(new_n304), .ZN(new_n309));
  XNOR2_X1  g123(.A(KEYINPUT2), .B(G113), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g125(.A1(new_n308), .A2(new_n311), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n258), .A2(new_n312), .A3(new_n267), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n302), .A2(new_n304), .A3(KEYINPUT5), .ZN(new_n314));
  OR3_X1    g128(.A1(new_n303), .A2(KEYINPUT5), .A3(G119), .ZN(new_n315));
  NAND4_X1  g129(.A1(new_n314), .A2(new_n315), .A3(KEYINPUT76), .A4(G113), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n309), .A2(new_n310), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n314), .A2(new_n315), .A3(G113), .ZN(new_n318));
  INV_X1    g132(.A(KEYINPUT76), .ZN(new_n319));
  AOI21_X1  g133(.A(new_n317), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NAND3_X1  g134(.A1(new_n218), .A2(new_n316), .A3(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n313), .A2(new_n321), .ZN(new_n322));
  XNOR2_X1  g136(.A(G110), .B(G122), .ZN(new_n323));
  INV_X1    g137(.A(new_n323), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n322), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n313), .A2(new_n321), .A3(new_n323), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(KEYINPUT6), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n322), .A2(new_n328), .A3(new_n324), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n261), .A2(new_n262), .ZN(new_n330));
  OAI211_X1 g144(.A(new_n264), .B(G125), .C1(new_n330), .C2(new_n203), .ZN(new_n331));
  INV_X1    g145(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND4_X1  g147(.A1(new_n263), .A2(KEYINPUT77), .A3(G125), .A4(new_n264), .ZN(new_n334));
  AND2_X1   g148(.A1(new_n333), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G125), .ZN(new_n336));
  NAND4_X1  g150(.A1(new_n220), .A2(new_n336), .A3(new_n222), .A4(new_n206), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n278), .A2(G224), .ZN(new_n339));
  INV_X1    g153(.A(new_n339), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n335), .A2(new_n339), .A3(new_n337), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n327), .A2(new_n329), .A3(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n339), .A2(KEYINPUT7), .ZN(new_n345));
  NAND4_X1  g159(.A1(new_n333), .A2(new_n337), .A3(new_n334), .A4(new_n345), .ZN(new_n346));
  AND3_X1   g160(.A1(new_n243), .A2(new_n320), .A3(new_n316), .ZN(new_n347));
  XNOR2_X1  g161(.A(KEYINPUT78), .B(KEYINPUT8), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n323), .B(new_n348), .ZN(new_n349));
  AND2_X1   g163(.A1(new_n318), .A2(new_n308), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n349), .B1(new_n243), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n346), .B1(new_n347), .B2(new_n351), .ZN(new_n352));
  INV_X1    g166(.A(new_n331), .ZN(new_n353));
  AOI21_X1  g167(.A(new_n353), .B1(new_n337), .B2(KEYINPUT79), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT79), .ZN(new_n355));
  NAND3_X1  g169(.A1(new_n249), .A2(new_n355), .A3(new_n336), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n345), .B1(new_n354), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n352), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n358), .B2(new_n326), .ZN(new_n359));
  OAI21_X1  g173(.A(G210), .B1(G237), .B2(G902), .ZN(new_n360));
  AND3_X1   g174(.A1(new_n344), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(new_n360), .B1(new_n344), .B2(new_n359), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n298), .A2(new_n300), .A3(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G140), .ZN(new_n365));
  AOI21_X1  g179(.A(KEYINPUT16), .B1(new_n365), .B2(G125), .ZN(new_n366));
  OAI211_X1 g180(.A(KEYINPUT69), .B(G125), .C1(new_n365), .C2(KEYINPUT70), .ZN(new_n367));
  NAND2_X1  g181(.A1(KEYINPUT69), .A2(G125), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT70), .ZN(new_n369));
  NAND3_X1  g183(.A1(new_n368), .A2(new_n369), .A3(G140), .ZN(new_n370));
  OAI21_X1  g184(.A(KEYINPUT70), .B1(new_n365), .B2(G125), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  AOI21_X1  g186(.A(new_n366), .B1(new_n372), .B2(KEYINPUT16), .ZN(new_n373));
  NOR2_X1   g187(.A1(new_n373), .A2(new_n209), .ZN(new_n374));
  AOI211_X1 g188(.A(G146), .B(new_n366), .C1(new_n372), .C2(KEYINPUT16), .ZN(new_n375));
  NOR2_X1   g189(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  OR2_X1    g190(.A1(KEYINPUT80), .A2(G143), .ZN(new_n377));
  NOR2_X1   g191(.A1(G237), .A2(G953), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n377), .A2(G214), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g193(.A1(KEYINPUT80), .A2(G143), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n377), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G237), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n382), .A2(new_n278), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n379), .B1(new_n381), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g199(.A1(new_n385), .A2(KEYINPUT83), .A3(KEYINPUT17), .A4(G131), .ZN(new_n386));
  AOI22_X1  g200(.A1(new_n377), .A2(new_n380), .B1(new_n378), .B2(G214), .ZN(new_n387));
  NOR2_X1   g201(.A1(KEYINPUT80), .A2(G143), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n383), .A2(new_n388), .ZN(new_n389));
  OAI211_X1 g203(.A(KEYINPUT17), .B(G131), .C1(new_n387), .C2(new_n389), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT83), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n386), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n385), .A2(G131), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT17), .ZN(new_n395));
  OAI211_X1 g209(.A(new_n232), .B(new_n379), .C1(new_n381), .C2(new_n384), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n394), .A2(new_n395), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n376), .A2(new_n393), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(KEYINPUT18), .A2(G131), .ZN(new_n399));
  XNOR2_X1  g213(.A(new_n385), .B(new_n399), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT81), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n372), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n367), .A2(new_n370), .A3(new_n371), .A4(KEYINPUT81), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(G146), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n336), .A2(G140), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n365), .A2(G125), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n405), .A2(new_n406), .A3(new_n209), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n400), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g223(.A(G113), .B(G122), .ZN(new_n410));
  XNOR2_X1  g224(.A(new_n410), .B(new_n198), .ZN(new_n411));
  AND3_X1   g225(.A1(new_n398), .A2(new_n409), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n402), .A2(KEYINPUT19), .A3(new_n403), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT19), .ZN(new_n414));
  NAND3_X1  g228(.A1(new_n405), .A2(new_n406), .A3(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n209), .A3(new_n415), .ZN(new_n416));
  OR2_X1    g230(.A1(new_n373), .A2(new_n209), .ZN(new_n417));
  NAND3_X1  g231(.A1(new_n416), .A2(KEYINPUT82), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n394), .A2(new_n396), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g234(.A(KEYINPUT82), .B1(new_n416), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g235(.A(new_n409), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(new_n411), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n412), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(G475), .A2(G902), .ZN(new_n425));
  INV_X1    g239(.A(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(KEYINPUT20), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g241(.A(KEYINPUT20), .ZN(new_n428));
  NAND2_X1  g242(.A1(new_n416), .A2(new_n417), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT82), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n431), .A2(new_n418), .A3(new_n419), .ZN(new_n432));
  AOI21_X1  g246(.A(new_n411), .B1(new_n432), .B2(new_n409), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n428), .B(new_n425), .C1(new_n433), .C2(new_n412), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n427), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G475), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n398), .A2(new_n409), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(new_n423), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT84), .ZN(new_n439));
  NAND3_X1  g253(.A1(new_n398), .A2(new_n411), .A3(new_n409), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n438), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n411), .B1(new_n398), .B2(new_n409), .ZN(new_n442));
  AOI21_X1  g256(.A(G902), .B1(new_n442), .B2(KEYINPUT84), .ZN(new_n443));
  AOI21_X1  g257(.A(new_n436), .B1(new_n441), .B2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(new_n444), .ZN(new_n445));
  XNOR2_X1  g259(.A(KEYINPUT64), .B(G134), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n207), .A2(G128), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n204), .A2(G143), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n446), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(G122), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n450), .A2(G116), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n303), .A2(G122), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n453), .A2(G107), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n451), .A2(new_n452), .A3(new_n194), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  INV_X1    g270(.A(KEYINPUT13), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n448), .B1(new_n447), .B2(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT85), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n447), .A2(new_n459), .A3(new_n457), .ZN(new_n460));
  OAI21_X1  g274(.A(new_n457), .B1(new_n204), .B2(G143), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT85), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n458), .B1(new_n460), .B2(new_n462), .ZN(new_n463));
  OAI211_X1 g277(.A(new_n449), .B(new_n456), .C1(new_n463), .C2(new_n225), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n452), .A2(KEYINPUT14), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT14), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n303), .A3(G122), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n465), .A2(new_n467), .A3(new_n451), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(G107), .ZN(new_n469));
  INV_X1    g283(.A(new_n449), .ZN(new_n470));
  AOI21_X1  g284(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n471));
  OAI211_X1 g285(.A(new_n469), .B(new_n455), .C1(new_n470), .C2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n296), .ZN(new_n473));
  AND3_X1   g287(.A1(new_n473), .A2(G217), .A3(new_n278), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n464), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n474), .B1(new_n464), .B2(new_n472), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n188), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  INV_X1    g291(.A(G478), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT15), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  OAI221_X1 g294(.A(new_n188), .B1(KEYINPUT15), .B2(new_n478), .C1(new_n475), .C2(new_n476), .ZN(new_n481));
  AND2_X1   g295(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g296(.A1(G234), .A2(G237), .ZN(new_n483));
  AND3_X1   g297(.A1(new_n483), .A2(G902), .A3(G953), .ZN(new_n484));
  XNOR2_X1  g298(.A(KEYINPUT21), .B(G898), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n484), .A2(new_n485), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(G952), .A3(new_n278), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g302(.A(new_n488), .B(KEYINPUT86), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n482), .A2(new_n489), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n435), .A2(new_n445), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AOI21_X1  g307(.A(new_n444), .B1(new_n427), .B2(new_n434), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n494), .A2(KEYINPUT87), .A3(new_n490), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n493), .A2(new_n495), .ZN(new_n496));
  AND2_X1   g310(.A1(new_n364), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(G234), .ZN(new_n498));
  OAI21_X1  g312(.A(G217), .B1(new_n498), .B2(G902), .ZN(new_n499));
  XOR2_X1   g313(.A(new_n499), .B(KEYINPUT68), .Z(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n204), .A2(G119), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n301), .A2(G128), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT24), .B(G110), .ZN(new_n505));
  NOR2_X1   g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n507));
  NOR2_X1   g321(.A1(new_n301), .A2(G128), .ZN(new_n508));
  OAI211_X1 g322(.A(new_n503), .B(new_n507), .C1(new_n508), .C2(KEYINPUT23), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n506), .B1(G110), .B2(new_n509), .ZN(new_n510));
  OAI21_X1  g324(.A(new_n510), .B1(new_n374), .B2(new_n375), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n509), .A2(G110), .ZN(new_n512));
  AND2_X1   g326(.A1(new_n504), .A2(new_n505), .ZN(new_n513));
  OAI221_X1 g327(.A(new_n407), .B1(new_n512), .B2(new_n513), .C1(new_n373), .C2(new_n209), .ZN(new_n514));
  XNOR2_X1  g328(.A(KEYINPUT22), .B(G137), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n278), .A2(G221), .A3(G234), .ZN(new_n516));
  XNOR2_X1  g330(.A(new_n515), .B(new_n516), .ZN(new_n517));
  NAND3_X1  g331(.A1(new_n511), .A2(new_n514), .A3(new_n517), .ZN(new_n518));
  INV_X1    g332(.A(new_n518), .ZN(new_n519));
  AOI21_X1  g333(.A(new_n517), .B1(new_n511), .B2(new_n514), .ZN(new_n520));
  NOR2_X1   g334(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT25), .B1(new_n521), .B2(new_n188), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT25), .ZN(new_n523));
  NOR4_X1   g337(.A1(new_n519), .A2(new_n520), .A3(new_n523), .A4(G902), .ZN(new_n524));
  OAI21_X1  g338(.A(new_n501), .B1(new_n522), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n499), .A2(new_n188), .ZN(new_n526));
  INV_X1    g340(.A(new_n526), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n521), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n525), .A2(new_n528), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n378), .A2(G210), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n530), .B(KEYINPUT27), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT26), .B(G101), .ZN(new_n532));
  XNOR2_X1  g346(.A(new_n531), .B(new_n532), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n232), .B1(G134), .B2(G137), .ZN(new_n534));
  NAND2_X1  g348(.A1(new_n226), .A2(new_n228), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n534), .B1(new_n535), .B2(G137), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n236), .A2(new_n536), .ZN(new_n537));
  NOR2_X1   g351(.A1(new_n249), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n226), .A2(new_n228), .A3(new_n230), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n233), .A2(new_n235), .ZN(new_n540));
  OAI21_X1  g354(.A(G131), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n541), .A2(new_n236), .B1(new_n263), .B2(new_n264), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n538), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT28), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT66), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n312), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n308), .A2(new_n311), .A3(KEYINPUT66), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n543), .A2(new_n544), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g363(.A1(new_n223), .A2(new_n236), .A3(new_n536), .ZN(new_n550));
  OAI21_X1  g364(.A(new_n265), .B1(new_n237), .B2(new_n239), .ZN(new_n551));
  NAND3_X1  g365(.A1(new_n548), .A2(new_n550), .A3(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n550), .A2(new_n551), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n312), .ZN(new_n556));
  AOI21_X1  g370(.A(new_n533), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT30), .ZN(new_n558));
  AND3_X1   g372(.A1(new_n550), .A2(new_n551), .A3(new_n558), .ZN(new_n559));
  AOI21_X1  g373(.A(new_n558), .B1(new_n550), .B2(new_n551), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n312), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n561), .A2(new_n533), .A3(new_n552), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT31), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  INV_X1    g378(.A(new_n552), .ZN(new_n565));
  OAI21_X1  g379(.A(KEYINPUT30), .B1(new_n538), .B2(new_n542), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n550), .A2(new_n551), .A3(new_n558), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI21_X1  g382(.A(new_n565), .B1(new_n568), .B2(new_n312), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n569), .A2(KEYINPUT31), .A3(new_n533), .ZN(new_n570));
  AOI21_X1  g384(.A(new_n557), .B1(new_n564), .B2(new_n570), .ZN(new_n571));
  NOR2_X1   g385(.A1(G472), .A2(G902), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  OAI21_X1  g387(.A(KEYINPUT32), .B1(new_n571), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n554), .A2(new_n556), .ZN(new_n575));
  INV_X1    g389(.A(new_n533), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n575), .A2(new_n576), .ZN(new_n577));
  AOI21_X1  g391(.A(KEYINPUT31), .B1(new_n569), .B2(new_n533), .ZN(new_n578));
  AOI22_X1  g392(.A1(new_n566), .A2(new_n567), .B1(new_n311), .B2(new_n308), .ZN(new_n579));
  NOR4_X1   g393(.A1(new_n579), .A2(new_n563), .A3(new_n565), .A4(new_n576), .ZN(new_n580));
  OAI21_X1  g394(.A(new_n577), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT32), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n581), .A2(new_n582), .A3(new_n572), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n576), .B1(new_n579), .B2(new_n565), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n544), .B1(new_n543), .B2(new_n548), .ZN(new_n586));
  NOR2_X1   g400(.A1(new_n552), .A2(KEYINPUT28), .ZN(new_n587));
  OAI211_X1 g401(.A(new_n533), .B(new_n556), .C1(new_n586), .C2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT29), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n585), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT67), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NOR2_X1   g406(.A1(new_n543), .A2(new_n548), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n554), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n595), .ZN(new_n596));
  NOR2_X1   g410(.A1(new_n576), .A2(new_n589), .ZN(new_n597));
  AOI21_X1  g411(.A(G902), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n585), .A2(new_n588), .A3(KEYINPUT67), .A4(new_n589), .ZN(new_n599));
  NAND3_X1  g413(.A1(new_n592), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n600), .A2(G472), .ZN(new_n601));
  AOI21_X1  g415(.A(new_n529), .B1(new_n584), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n497), .A2(new_n602), .ZN(new_n603));
  XNOR2_X1  g417(.A(new_n603), .B(G101), .ZN(G3));
  NAND2_X1  g418(.A1(new_n435), .A2(new_n445), .ZN(new_n605));
  XNOR2_X1  g419(.A(KEYINPUT89), .B(KEYINPUT33), .ZN(new_n606));
  OAI21_X1  g420(.A(new_n606), .B1(new_n475), .B2(new_n476), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n478), .A2(G902), .ZN(new_n608));
  INV_X1    g422(.A(new_n475), .ZN(new_n609));
  INV_X1    g423(.A(KEYINPUT90), .ZN(new_n610));
  OAI211_X1 g424(.A(new_n609), .B(KEYINPUT33), .C1(new_n610), .C2(new_n476), .ZN(new_n611));
  AND2_X1   g425(.A1(new_n476), .A2(new_n610), .ZN(new_n612));
  OAI211_X1 g426(.A(new_n607), .B(new_n608), .C1(new_n611), .C2(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n477), .A2(new_n478), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n605), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n344), .A2(new_n359), .ZN(new_n617));
  INV_X1    g431(.A(new_n360), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT88), .ZN(new_n620));
  NAND3_X1  g434(.A1(new_n344), .A2(new_n359), .A3(new_n360), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  AOI21_X1  g436(.A(new_n300), .B1(new_n362), .B2(KEYINPUT88), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n622), .A2(new_n489), .A3(new_n623), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n616), .A2(new_n624), .ZN(new_n625));
  AND2_X1   g439(.A1(new_n295), .A2(new_n297), .ZN(new_n626));
  AND2_X1   g440(.A1(new_n525), .A2(new_n528), .ZN(new_n627));
  OAI21_X1  g441(.A(G472), .B1(new_n571), .B2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n581), .A2(new_n572), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n627), .A2(new_n628), .A3(new_n629), .ZN(new_n630));
  NAND3_X1  g444(.A1(new_n625), .A2(new_n626), .A3(new_n630), .ZN(new_n631));
  XOR2_X1   g445(.A(KEYINPUT34), .B(G104), .Z(new_n632));
  XNOR2_X1  g446(.A(new_n631), .B(new_n632), .ZN(G6));
  NAND3_X1  g447(.A1(new_n427), .A2(KEYINPUT91), .A3(new_n434), .ZN(new_n634));
  INV_X1    g448(.A(new_n424), .ZN(new_n635));
  INV_X1    g449(.A(KEYINPUT91), .ZN(new_n636));
  NAND4_X1  g450(.A1(new_n635), .A2(new_n636), .A3(new_n428), .A4(new_n425), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n444), .A2(new_n482), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n634), .A2(new_n637), .A3(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n624), .A2(new_n639), .ZN(new_n640));
  NAND3_X1  g454(.A1(new_n640), .A2(new_n626), .A3(new_n630), .ZN(new_n641));
  XOR2_X1   g455(.A(new_n641), .B(KEYINPUT92), .Z(new_n642));
  XOR2_X1   g456(.A(KEYINPUT35), .B(G107), .Z(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G9));
  AND2_X1   g458(.A1(new_n628), .A2(new_n629), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n511), .A2(new_n514), .ZN(new_n646));
  INV_X1    g460(.A(new_n517), .ZN(new_n647));
  NOR2_X1   g461(.A1(new_n647), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n646), .B(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n527), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n525), .A2(new_n650), .ZN(new_n651));
  AND2_X1   g465(.A1(new_n645), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n497), .A2(new_n652), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n653), .B(KEYINPUT93), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT37), .B(G110), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G12));
  AND4_X1   g470(.A1(new_n297), .A2(new_n295), .A3(new_n622), .A4(new_n623), .ZN(new_n657));
  INV_X1    g471(.A(new_n487), .ZN(new_n658));
  INV_X1    g472(.A(G900), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n658), .B1(new_n484), .B2(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n639), .A2(new_n660), .ZN(new_n661));
  INV_X1    g475(.A(new_n651), .ZN(new_n662));
  AOI21_X1  g476(.A(new_n662), .B1(new_n584), .B2(new_n601), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n657), .A2(new_n661), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(G128), .ZN(G30));
  XOR2_X1   g479(.A(new_n660), .B(KEYINPUT39), .Z(new_n666));
  XOR2_X1   g480(.A(KEYINPUT95), .B(KEYINPUT40), .Z(new_n667));
  NAND3_X1  g481(.A1(new_n626), .A2(new_n666), .A3(new_n667), .ZN(new_n668));
  INV_X1    g482(.A(G472), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n565), .A2(new_n533), .ZN(new_n670));
  AOI21_X1  g484(.A(G902), .B1(new_n594), .B2(new_n670), .ZN(new_n671));
  OAI21_X1  g485(.A(new_n533), .B1(new_n579), .B2(new_n565), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n669), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  AOI21_X1  g487(.A(new_n673), .B1(new_n574), .B2(new_n583), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n619), .A2(new_n621), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(KEYINPUT38), .ZN(new_n677));
  AND3_X1   g491(.A1(new_n668), .A2(new_n675), .A3(new_n677), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n626), .A2(new_n666), .ZN(new_n679));
  INV_X1    g493(.A(new_n667), .ZN(new_n680));
  NAND2_X1  g494(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(KEYINPUT96), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n482), .B1(new_n435), .B2(new_n445), .ZN(new_n684));
  NAND3_X1  g498(.A1(new_n684), .A2(new_n299), .A3(new_n662), .ZN(new_n685));
  XOR2_X1   g499(.A(new_n685), .B(KEYINPUT94), .Z(new_n686));
  OR3_X1    g500(.A1(new_n682), .A2(new_n683), .A3(new_n686), .ZN(new_n687));
  OAI21_X1  g501(.A(new_n683), .B1(new_n682), .B2(new_n686), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(new_n207), .ZN(G45));
  INV_X1    g504(.A(new_n615), .ZN(new_n691));
  NOR3_X1   g505(.A1(new_n494), .A2(new_n691), .A3(new_n660), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n657), .A2(new_n663), .A3(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G146), .ZN(G48));
  NAND2_X1  g508(.A1(new_n286), .A2(new_n277), .ZN(new_n695));
  INV_X1    g509(.A(new_n282), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n268), .A2(new_n270), .ZN(new_n697));
  AOI21_X1  g511(.A(new_n697), .B1(new_n275), .B2(new_n273), .ZN(new_n698));
  AOI21_X1  g512(.A(new_n696), .B1(new_n698), .B2(new_n240), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n224), .A2(KEYINPUT12), .A3(new_n241), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT75), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n224), .A2(new_n241), .ZN(new_n703));
  INV_X1    g517(.A(KEYINPUT12), .ZN(new_n704));
  NAND2_X1  g518(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  NAND3_X1  g519(.A1(new_n702), .A2(new_n705), .A3(new_n242), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n695), .A2(new_n696), .B1(new_n699), .B2(new_n706), .ZN(new_n707));
  OAI21_X1  g521(.A(G469), .B1(new_n707), .B2(G902), .ZN(new_n708));
  NAND3_X1  g522(.A1(new_n708), .A2(new_n297), .A3(new_n288), .ZN(new_n709));
  INV_X1    g523(.A(new_n709), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n625), .A2(new_n602), .A3(new_n710), .ZN(new_n711));
  XOR2_X1   g525(.A(KEYINPUT41), .B(G113), .Z(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(KEYINPUT97), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n711), .B(new_n713), .ZN(G15));
  NAND3_X1  g528(.A1(new_n602), .A2(new_n640), .A3(new_n710), .ZN(new_n715));
  XNOR2_X1  g529(.A(KEYINPUT98), .B(G116), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n715), .B(new_n716), .ZN(G18));
  NAND2_X1  g531(.A1(new_n622), .A2(new_n623), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n709), .A2(new_n718), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n496), .A2(new_n663), .A3(new_n719), .ZN(new_n720));
  XNOR2_X1  g534(.A(new_n720), .B(G119), .ZN(G21));
  AOI21_X1  g535(.A(new_n533), .B1(new_n554), .B2(new_n594), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n722), .B1(new_n564), .B2(new_n570), .ZN(new_n723));
  OAI21_X1  g537(.A(KEYINPUT99), .B1(new_n723), .B2(new_n573), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n595), .A2(new_n576), .ZN(new_n725));
  OAI21_X1  g539(.A(new_n725), .B1(new_n578), .B2(new_n580), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT99), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n726), .A2(new_n727), .A3(new_n572), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n724), .A2(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n581), .A2(new_n188), .ZN(new_n730));
  XOR2_X1   g544(.A(KEYINPUT100), .B(G472), .Z(new_n731));
  NAND2_X1  g545(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  AND3_X1   g546(.A1(new_n729), .A2(new_n627), .A3(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n709), .A2(new_n624), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n733), .A2(new_n734), .A3(new_n684), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AOI22_X1  g550(.A1(new_n724), .A2(new_n728), .B1(new_n730), .B2(new_n731), .ZN(new_n737));
  NAND4_X1  g551(.A1(new_n719), .A2(new_n692), .A3(new_n651), .A4(new_n737), .ZN(new_n738));
  XNOR2_X1  g552(.A(new_n738), .B(G125), .ZN(G27));
  INV_X1    g553(.A(KEYINPUT42), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n584), .A2(new_n601), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n741), .A2(new_n627), .ZN(new_n742));
  AOI21_X1  g556(.A(new_n691), .B1(new_n435), .B2(new_n445), .ZN(new_n743));
  INV_X1    g557(.A(new_n660), .ZN(new_n744));
  XNOR2_X1  g558(.A(new_n289), .B(KEYINPUT101), .ZN(new_n745));
  NAND3_X1  g559(.A1(new_n288), .A2(new_n294), .A3(new_n745), .ZN(new_n746));
  AND2_X1   g560(.A1(new_n297), .A2(new_n299), .ZN(new_n747));
  AND3_X1   g561(.A1(new_n619), .A2(new_n621), .A3(new_n747), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n743), .A2(new_n744), .A3(new_n746), .A4(new_n748), .ZN(new_n749));
  OAI21_X1  g563(.A(new_n740), .B1(new_n742), .B2(new_n749), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n743), .A2(new_n744), .A3(new_n746), .A4(new_n748), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n751), .A2(KEYINPUT42), .A3(new_n602), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n750), .A2(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(new_n753), .B(G131), .ZN(G33));
  AND2_X1   g568(.A1(new_n746), .A2(new_n748), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n602), .A2(new_n755), .A3(new_n661), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G134), .ZN(G36));
  NOR2_X1   g571(.A1(new_n645), .A2(new_n662), .ZN(new_n758));
  OR3_X1    g572(.A1(new_n605), .A2(KEYINPUT43), .A3(new_n691), .ZN(new_n759));
  OAI21_X1  g573(.A(KEYINPUT43), .B1(new_n605), .B2(new_n691), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT44), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n761), .A2(new_n762), .ZN(new_n763));
  NOR2_X1   g577(.A1(new_n761), .A2(new_n762), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n676), .A2(new_n300), .ZN(new_n765));
  INV_X1    g579(.A(new_n765), .ZN(new_n766));
  NOR3_X1   g580(.A1(new_n763), .A2(new_n764), .A3(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n292), .A2(new_n293), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n769));
  AOI21_X1  g583(.A(new_n187), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n292), .A2(KEYINPUT45), .A3(new_n293), .ZN(new_n771));
  AOI21_X1  g585(.A(KEYINPUT102), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(new_n291), .ZN(new_n773));
  AOI21_X1  g587(.A(new_n773), .B1(new_n706), .B2(new_n277), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n240), .B1(new_n271), .B2(new_n276), .ZN(new_n775));
  NOR2_X1   g589(.A1(new_n283), .A2(new_n775), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n769), .B1(new_n774), .B2(new_n776), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n777), .A2(new_n771), .A3(KEYINPUT102), .A4(G469), .ZN(new_n778));
  INV_X1    g592(.A(new_n778), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n745), .B1(new_n772), .B2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(KEYINPUT46), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g596(.A(new_n745), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n777), .A2(new_n771), .A3(G469), .ZN(new_n784));
  INV_X1    g598(.A(KEYINPUT102), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n784), .A2(new_n785), .ZN(new_n786));
  AOI21_X1  g600(.A(new_n783), .B1(new_n786), .B2(new_n778), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(KEYINPUT46), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n782), .A2(new_n288), .A3(new_n788), .ZN(new_n789));
  AND2_X1   g603(.A1(new_n666), .A2(new_n297), .ZN(new_n790));
  AOI21_X1  g604(.A(KEYINPUT103), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  OAI21_X1  g605(.A(new_n288), .B1(new_n787), .B2(KEYINPUT46), .ZN(new_n792));
  AOI211_X1 g606(.A(new_n781), .B(new_n783), .C1(new_n786), .C2(new_n778), .ZN(new_n793));
  OAI211_X1 g607(.A(KEYINPUT103), .B(new_n790), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  INV_X1    g608(.A(new_n794), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n767), .B1(new_n791), .B2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G137), .ZN(G39));
  OAI21_X1  g611(.A(new_n297), .B1(new_n792), .B2(new_n793), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n798), .A2(KEYINPUT47), .ZN(new_n799));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  NAND3_X1  g614(.A1(new_n789), .A2(new_n800), .A3(new_n297), .ZN(new_n801));
  AOI22_X1  g615(.A1(new_n574), .A2(new_n583), .B1(new_n600), .B2(G472), .ZN(new_n802));
  AND4_X1   g616(.A1(new_n802), .A2(new_n692), .A3(new_n529), .A4(new_n765), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(G140), .ZN(G42));
  INV_X1    g619(.A(new_n277), .ZN(new_n806));
  OAI21_X1  g620(.A(new_n696), .B1(new_n806), .B2(new_n775), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n706), .A2(new_n277), .A3(new_n282), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  AOI21_X1  g623(.A(new_n187), .B1(new_n809), .B2(new_n188), .ZN(new_n810));
  AOI211_X1 g624(.A(G469), .B(G902), .C1(new_n807), .C2(new_n808), .ZN(new_n811));
  NOR2_X1   g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  INV_X1    g626(.A(KEYINPUT49), .ZN(new_n813));
  OAI211_X1 g627(.A(new_n627), .B(new_n747), .C1(new_n812), .C2(new_n813), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n814), .B1(new_n813), .B2(new_n812), .ZN(new_n815));
  NOR2_X1   g629(.A1(new_n675), .A2(new_n677), .ZN(new_n816));
  NAND4_X1  g630(.A1(new_n815), .A2(new_n494), .A3(new_n615), .A4(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n710), .A2(new_n765), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n674), .A2(new_n627), .A3(new_n658), .ZN(new_n819));
  NOR2_X1   g633(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(KEYINPUT111), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(new_n743), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n823), .A2(G952), .A3(new_n278), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n759), .A2(new_n658), .A3(new_n760), .ZN(new_n825));
  INV_X1    g639(.A(KEYINPUT107), .ZN(new_n826));
  XNOR2_X1  g640(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n827), .A2(new_n733), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n824), .B1(new_n719), .B2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(new_n818), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n825), .A2(new_n826), .ZN(new_n831));
  NOR2_X1   g645(.A1(new_n825), .A2(new_n826), .ZN(new_n832));
  OAI21_X1  g646(.A(new_n830), .B1(new_n831), .B2(new_n832), .ZN(new_n833));
  INV_X1    g647(.A(KEYINPUT110), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(new_n834), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n827), .A2(KEYINPUT110), .A3(new_n830), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(KEYINPUT48), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n838), .A3(new_n602), .ZN(new_n839));
  INV_X1    g653(.A(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n838), .B1(new_n837), .B2(new_n602), .ZN(new_n841));
  OAI21_X1  g655(.A(new_n829), .B1(new_n840), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n605), .A2(new_n615), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n821), .A2(new_n822), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT112), .ZN(new_n845));
  NAND2_X1  g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR3_X1   g660(.A1(new_n677), .A2(new_n299), .A3(new_n709), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n733), .B(new_n847), .C1(new_n831), .C2(new_n832), .ZN(new_n848));
  XOR2_X1   g662(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NOR2_X1   g664(.A1(KEYINPUT109), .A2(KEYINPUT50), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n827), .A2(new_n733), .A3(new_n847), .A4(new_n851), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n821), .A2(KEYINPUT112), .A3(new_n822), .A4(new_n843), .ZN(new_n853));
  NAND4_X1  g667(.A1(new_n846), .A2(new_n850), .A3(new_n852), .A4(new_n853), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n729), .A2(new_n651), .A3(new_n732), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n855), .B1(new_n835), .B2(new_n836), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n854), .A2(new_n856), .ZN(new_n857));
  NAND2_X1  g671(.A1(new_n828), .A2(new_n765), .ZN(new_n858));
  INV_X1    g672(.A(new_n812), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n859), .A2(new_n297), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n799), .B2(new_n801), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT51), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n842), .B1(new_n857), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n861), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT108), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n867), .A3(new_n765), .A4(new_n828), .ZN(new_n868));
  OAI21_X1  g682(.A(KEYINPUT108), .B1(new_n858), .B2(new_n861), .ZN(new_n869));
  NAND3_X1  g683(.A1(new_n857), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(KEYINPUT113), .ZN(new_n871));
  AND3_X1   g685(.A1(new_n870), .A2(new_n871), .A3(new_n863), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n871), .B1(new_n870), .B2(new_n863), .ZN(new_n873));
  OAI21_X1  g687(.A(new_n865), .B1(new_n872), .B2(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT52), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n812), .A2(new_n297), .A3(new_n622), .A4(new_n623), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n876), .A2(new_n855), .ZN(new_n877));
  NOR3_X1   g691(.A1(new_n718), .A2(new_n494), .A3(new_n482), .ZN(new_n878));
  AND2_X1   g692(.A1(new_n744), .A2(new_n297), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n746), .A2(new_n662), .A3(new_n879), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n880), .A2(new_n674), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n877), .A2(new_n692), .B1(new_n878), .B2(new_n881), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n657), .B(new_n663), .C1(new_n661), .C2(new_n692), .ZN(new_n883));
  AOI21_X1  g697(.A(KEYINPUT105), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n878), .ZN(new_n885));
  AND4_X1   g699(.A1(KEYINPUT105), .A2(new_n883), .A3(new_n738), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n875), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  AND2_X1   g701(.A1(new_n720), .A2(new_n715), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n802), .A2(new_n529), .A3(new_n709), .ZN(new_n889));
  AND4_X1   g703(.A1(new_n627), .A2(new_n729), .A3(new_n684), .A4(new_n732), .ZN(new_n890));
  AOI22_X1  g704(.A1(new_n625), .A2(new_n889), .B1(new_n890), .B2(new_n734), .ZN(new_n891));
  AND3_X1   g705(.A1(new_n480), .A2(KEYINPUT104), .A3(new_n481), .ZN(new_n892));
  AOI21_X1  g706(.A(KEYINPUT104), .B1(new_n480), .B2(new_n481), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n494), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n616), .A2(new_n895), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n676), .A2(new_n489), .A3(new_n299), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n896), .A2(new_n626), .A3(new_n630), .A4(new_n898), .ZN(new_n899));
  OAI211_X1 g713(.A(new_n364), .B(new_n496), .C1(new_n652), .C2(new_n602), .ZN(new_n900));
  NAND4_X1  g714(.A1(new_n888), .A2(new_n891), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n744), .B1(new_n892), .B2(new_n893), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n902), .A2(new_n444), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n903), .A2(new_n363), .A3(new_n299), .A4(new_n651), .ZN(new_n904));
  NOR3_X1   g718(.A1(new_n802), .A2(new_n298), .A3(new_n904), .ZN(new_n905));
  AND2_X1   g719(.A1(new_n634), .A2(new_n637), .ZN(new_n906));
  INV_X1    g720(.A(new_n855), .ZN(new_n907));
  AOI22_X1  g721(.A1(new_n905), .A2(new_n906), .B1(new_n907), .B2(new_n751), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n753), .A2(new_n908), .A3(new_n756), .ZN(new_n909));
  NOR2_X1   g723(.A1(new_n901), .A2(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT105), .ZN(new_n911));
  INV_X1    g725(.A(new_n883), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n885), .A2(new_n738), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n911), .B1(new_n912), .B2(new_n913), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n882), .A2(KEYINPUT105), .A3(new_n883), .ZN(new_n915));
  NAND3_X1  g729(.A1(new_n914), .A2(new_n915), .A3(KEYINPUT52), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n887), .A2(new_n910), .A3(new_n916), .ZN(new_n917));
  INV_X1    g731(.A(KEYINPUT53), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  INV_X1    g733(.A(KEYINPUT54), .ZN(new_n920));
  OAI21_X1  g734(.A(KEYINPUT52), .B1(new_n912), .B2(new_n913), .ZN(new_n921));
  NAND4_X1  g735(.A1(new_n887), .A2(new_n910), .A3(KEYINPUT53), .A4(new_n921), .ZN(new_n922));
  AND3_X1   g736(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n923));
  NAND3_X1  g737(.A1(new_n887), .A2(new_n910), .A3(new_n921), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n924), .A2(new_n918), .ZN(new_n925));
  NAND4_X1  g739(.A1(new_n887), .A2(new_n910), .A3(new_n916), .A4(KEYINPUT53), .ZN(new_n926));
  AOI21_X1  g740(.A(new_n920), .B1(new_n925), .B2(new_n926), .ZN(new_n927));
  OAI21_X1  g741(.A(KEYINPUT106), .B1(new_n923), .B2(new_n927), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT52), .B1(new_n914), .B2(new_n915), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n735), .A2(new_n711), .A3(new_n899), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n720), .A2(new_n715), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n756), .ZN(new_n933));
  AOI21_X1  g747(.A(new_n933), .B1(new_n750), .B2(new_n752), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n932), .A2(new_n900), .A3(new_n934), .A4(new_n908), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n929), .A2(new_n935), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT53), .B1(new_n936), .B2(new_n921), .ZN(new_n937));
  INV_X1    g751(.A(new_n926), .ZN(new_n938));
  OAI21_X1  g752(.A(KEYINPUT54), .B1(new_n937), .B2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(KEYINPUT106), .ZN(new_n940));
  NAND3_X1  g754(.A1(new_n919), .A2(new_n920), .A3(new_n922), .ZN(new_n941));
  NAND3_X1  g755(.A1(new_n939), .A2(new_n940), .A3(new_n941), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n874), .B1(new_n928), .B2(new_n942), .ZN(new_n943));
  NOR2_X1   g757(.A1(G952), .A2(G953), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n817), .B1(new_n943), .B2(new_n944), .ZN(G75));
  AOI21_X1  g759(.A(new_n188), .B1(new_n919), .B2(new_n922), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n946), .A2(G210), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT56), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n327), .A2(new_n329), .ZN(new_n949));
  XNOR2_X1  g763(.A(new_n949), .B(new_n343), .ZN(new_n950));
  XNOR2_X1  g764(.A(KEYINPUT114), .B(KEYINPUT55), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n950), .B(new_n951), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n947), .A2(new_n948), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n952), .B1(new_n947), .B2(new_n948), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n278), .A2(G952), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n954), .A3(new_n955), .ZN(G51));
  NAND2_X1  g770(.A1(new_n919), .A2(new_n922), .ZN(new_n957));
  NAND4_X1  g771(.A1(new_n957), .A2(G902), .A3(new_n786), .A4(new_n778), .ZN(new_n958));
  INV_X1    g772(.A(KEYINPUT117), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n957), .A2(KEYINPUT54), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n941), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n745), .B(KEYINPUT57), .Z(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  XNOR2_X1  g778(.A(new_n707), .B(KEYINPUT115), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n964), .A2(new_n965), .ZN(new_n966));
  AOI21_X1  g780(.A(new_n960), .B1(new_n966), .B2(KEYINPUT116), .ZN(new_n967));
  OR2_X1    g781(.A1(new_n966), .A2(KEYINPUT116), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n955), .B1(new_n967), .B2(new_n968), .ZN(G54));
  NAND3_X1  g783(.A1(new_n946), .A2(KEYINPUT58), .A3(G475), .ZN(new_n970));
  AND2_X1   g784(.A1(new_n970), .A2(new_n424), .ZN(new_n971));
  NOR2_X1   g785(.A1(new_n970), .A2(new_n424), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n971), .A2(new_n972), .A3(new_n955), .ZN(G60));
  XNOR2_X1  g787(.A(KEYINPUT119), .B(KEYINPUT59), .ZN(new_n974));
  NOR2_X1   g788(.A1(new_n478), .A2(new_n188), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n974), .B(new_n975), .Z(new_n976));
  INV_X1    g790(.A(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n928), .A2(new_n942), .A3(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n607), .B1(new_n611), .B2(new_n612), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT118), .ZN(new_n980));
  NAND2_X1  g794(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n980), .A2(new_n976), .ZN(new_n982));
  AOI21_X1  g796(.A(new_n955), .B1(new_n962), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n981), .A2(new_n983), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n984), .A2(KEYINPUT120), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT120), .ZN(new_n986));
  NAND3_X1  g800(.A1(new_n981), .A2(new_n986), .A3(new_n983), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n985), .A2(new_n987), .ZN(G63));
  NAND2_X1  g802(.A1(G217), .A2(G902), .ZN(new_n989));
  XNOR2_X1  g803(.A(new_n989), .B(KEYINPUT121), .ZN(new_n990));
  XNOR2_X1  g804(.A(new_n990), .B(KEYINPUT60), .ZN(new_n991));
  NAND2_X1  g805(.A1(new_n957), .A2(new_n991), .ZN(new_n992));
  INV_X1    g806(.A(new_n521), .ZN(new_n993));
  AOI21_X1  g807(.A(new_n955), .B1(new_n992), .B2(new_n993), .ZN(new_n994));
  INV_X1    g808(.A(new_n992), .ZN(new_n995));
  AND3_X1   g809(.A1(new_n995), .A2(KEYINPUT122), .A3(new_n649), .ZN(new_n996));
  AOI21_X1  g810(.A(KEYINPUT122), .B1(new_n995), .B2(new_n649), .ZN(new_n997));
  OAI21_X1  g811(.A(new_n994), .B1(new_n996), .B2(new_n997), .ZN(new_n998));
  INV_X1    g812(.A(KEYINPUT123), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n999), .B1(new_n996), .B2(new_n997), .ZN(new_n1000));
  INV_X1    g814(.A(KEYINPUT61), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n998), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  OAI221_X1 g816(.A(new_n994), .B1(new_n999), .B2(KEYINPUT61), .C1(new_n996), .C2(new_n997), .ZN(new_n1003));
  NAND2_X1  g817(.A1(new_n1002), .A2(new_n1003), .ZN(G66));
  NAND2_X1  g818(.A1(G224), .A2(G953), .ZN(new_n1005));
  OAI22_X1  g819(.A1(new_n901), .A2(G953), .B1(new_n485), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g820(.A(G898), .ZN(new_n1007));
  AOI21_X1  g821(.A(new_n949), .B1(new_n1007), .B2(G953), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1006), .B(new_n1008), .ZN(G69));
  AOI21_X1  g823(.A(new_n278), .B1(G227), .B2(G900), .ZN(new_n1010));
  AND2_X1   g824(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1011));
  NOR2_X1   g825(.A1(new_n1010), .A2(KEYINPUT126), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n883), .A2(new_n738), .ZN(new_n1013));
  NAND2_X1  g827(.A1(new_n934), .A2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n790), .B1(new_n792), .B2(new_n793), .ZN(new_n1015));
  INV_X1    g829(.A(KEYINPUT103), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  NAND2_X1  g831(.A1(new_n1017), .A2(new_n794), .ZN(new_n1018));
  AOI21_X1  g832(.A(new_n1014), .B1(new_n1018), .B2(new_n767), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n878), .A2(new_n602), .ZN(new_n1020));
  INV_X1    g834(.A(new_n1020), .ZN(new_n1021));
  OAI21_X1  g835(.A(new_n1021), .B1(new_n791), .B2(new_n795), .ZN(new_n1022));
  NAND4_X1  g836(.A1(new_n1019), .A2(KEYINPUT124), .A3(new_n804), .A4(new_n1022), .ZN(new_n1023));
  INV_X1    g837(.A(new_n1023), .ZN(new_n1024));
  AND3_X1   g838(.A1(new_n799), .A2(new_n801), .A3(new_n803), .ZN(new_n1025));
  AOI21_X1  g839(.A(new_n1020), .B1(new_n1017), .B2(new_n794), .ZN(new_n1026));
  NOR2_X1   g840(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1027));
  AOI21_X1  g841(.A(KEYINPUT124), .B1(new_n1027), .B2(new_n1019), .ZN(new_n1028));
  OAI21_X1  g842(.A(new_n278), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  NOR2_X1   g843(.A1(new_n278), .A2(G900), .ZN(new_n1030));
  INV_X1    g844(.A(new_n1030), .ZN(new_n1031));
  NAND3_X1  g845(.A1(new_n1029), .A2(KEYINPUT125), .A3(new_n1031), .ZN(new_n1032));
  INV_X1    g846(.A(KEYINPUT125), .ZN(new_n1033));
  INV_X1    g847(.A(new_n1014), .ZN(new_n1034));
  NAND4_X1  g848(.A1(new_n796), .A2(new_n1022), .A3(new_n804), .A4(new_n1034), .ZN(new_n1035));
  INV_X1    g849(.A(KEYINPUT124), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AOI21_X1  g851(.A(G953), .B1(new_n1037), .B2(new_n1023), .ZN(new_n1038));
  OAI21_X1  g852(.A(new_n1033), .B1(new_n1038), .B2(new_n1030), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n413), .A2(new_n415), .ZN(new_n1040));
  XNOR2_X1  g854(.A(new_n568), .B(new_n1040), .ZN(new_n1041));
  NAND3_X1  g855(.A1(new_n1032), .A2(new_n1039), .A3(new_n1041), .ZN(new_n1042));
  INV_X1    g856(.A(new_n1041), .ZN(new_n1043));
  NAND3_X1  g857(.A1(new_n687), .A2(new_n688), .A3(new_n1013), .ZN(new_n1044));
  XNOR2_X1  g858(.A(new_n1044), .B(KEYINPUT62), .ZN(new_n1045));
  NOR3_X1   g859(.A1(new_n679), .A2(new_n742), .A3(new_n766), .ZN(new_n1046));
  NAND2_X1  g860(.A1(new_n1046), .A2(new_n896), .ZN(new_n1047));
  NAND3_X1  g861(.A1(new_n796), .A2(new_n804), .A3(new_n1047), .ZN(new_n1048));
  NOR2_X1   g862(.A1(new_n1045), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1043), .B1(new_n1049), .B2(G953), .ZN(new_n1050));
  AOI211_X1 g864(.A(new_n1011), .B(new_n1012), .C1(new_n1042), .C2(new_n1050), .ZN(new_n1051));
  AND4_X1   g865(.A1(KEYINPUT126), .A2(new_n1042), .A3(new_n1010), .A4(new_n1050), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n1051), .A2(new_n1052), .ZN(G72));
  INV_X1    g867(.A(new_n901), .ZN(new_n1054));
  NAND2_X1  g868(.A1(new_n1049), .A2(new_n1054), .ZN(new_n1055));
  NAND2_X1  g869(.A1(G472), .A2(G902), .ZN(new_n1056));
  XNOR2_X1  g870(.A(new_n1056), .B(KEYINPUT63), .ZN(new_n1057));
  XNOR2_X1  g871(.A(new_n1057), .B(KEYINPUT127), .ZN(new_n1058));
  AOI21_X1  g872(.A(new_n672), .B1(new_n1055), .B2(new_n1058), .ZN(new_n1059));
  NOR2_X1   g873(.A1(new_n937), .A2(new_n938), .ZN(new_n1060));
  AOI211_X1 g874(.A(new_n1057), .B(new_n1060), .C1(new_n585), .C2(new_n562), .ZN(new_n1061));
  NAND2_X1  g875(.A1(new_n670), .A2(new_n561), .ZN(new_n1062));
  NAND3_X1  g876(.A1(new_n1037), .A2(new_n1054), .A3(new_n1023), .ZN(new_n1063));
  AOI21_X1  g877(.A(new_n1062), .B1(new_n1063), .B2(new_n1058), .ZN(new_n1064));
  NOR4_X1   g878(.A1(new_n1059), .A2(new_n1061), .A3(new_n955), .A4(new_n1064), .ZN(G57));
endmodule


