//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 0 0 0 1 1 0 0 0 0 1 1 0 1 1 0 0 0 1 1 1 1 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 1 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0 1 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:56 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n434, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n555, new_n557, new_n558, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n565, new_n566, new_n569,
    new_n570, new_n571, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n591, new_n592,
    new_n593, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n609,
    new_n612, new_n614, new_n615, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1126, new_n1127;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XNOR2_X1  g002(.A(KEYINPUT64), .B(G452), .ZN(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XOR2_X1   g008(.A(KEYINPUT66), .B(G44), .Z(new_n434));
  INV_X1    g009(.A(new_n434), .ZN(G218));
  INV_X1    g010(.A(G132), .ZN(G219));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  XNOR2_X1  g014(.A(KEYINPUT67), .B(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT68), .Z(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G218), .A2(G221), .A3(G219), .A4(G220), .ZN(new_n452));
  XOR2_X1   g027(.A(new_n452), .B(KEYINPUT2), .Z(new_n453));
  NOR4_X1   g028(.A1(G236), .A2(G237), .A3(G235), .A4(G238), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT69), .Z(new_n455));
  OR2_X1    g030(.A1(new_n453), .A2(new_n455), .ZN(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  AOI21_X1  g032(.A(KEYINPUT70), .B1(new_n455), .B2(G567), .ZN(new_n458));
  AOI21_X1  g033(.A(new_n458), .B1(G2106), .B2(new_n453), .ZN(new_n459));
  NAND3_X1  g034(.A1(new_n455), .A2(KEYINPUT70), .A3(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  AND2_X1   g043(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n469));
  NOR2_X1   g044(.A1(KEYINPUT71), .A2(G2105), .ZN(new_n470));
  OAI211_X1 g045(.A(new_n466), .B(new_n468), .C1(new_n469), .C2(new_n470), .ZN(new_n471));
  INV_X1    g046(.A(G137), .ZN(new_n472));
  OAI21_X1  g047(.A(new_n465), .B1(new_n471), .B2(new_n472), .ZN(new_n473));
  XNOR2_X1  g048(.A(KEYINPUT71), .B(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n466), .A2(new_n468), .A3(G125), .ZN(new_n475));
  NAND2_X1  g050(.A1(G113), .A2(G2104), .ZN(new_n476));
  AOI21_X1  g051(.A(new_n474), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g052(.A1(new_n473), .A2(new_n477), .ZN(G160));
  XNOR2_X1  g053(.A(KEYINPUT3), .B(G2104), .ZN(new_n479));
  INV_X1    g054(.A(new_n479), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(new_n474), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n480), .A2(G2105), .ZN(new_n482));
  AOI22_X1  g057(.A1(G124), .A2(new_n481), .B1(new_n482), .B2(G136), .ZN(new_n483));
  OAI221_X1 g058(.A(G2104), .B1(G100), .B2(G2105), .C1(new_n474), .C2(G112), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  XNOR2_X1  g060(.A(new_n485), .B(KEYINPUT72), .ZN(G162));
  INV_X1    g061(.A(G138), .ZN(new_n487));
  OAI21_X1  g062(.A(KEYINPUT75), .B1(new_n471), .B2(new_n487), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT75), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n474), .A2(new_n479), .A3(new_n489), .A4(G138), .ZN(new_n490));
  NAND3_X1  g065(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n491));
  OAI21_X1  g066(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n492));
  INV_X1    g067(.A(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(G114), .ZN(new_n494));
  AND3_X1   g069(.A1(new_n494), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n495));
  AOI21_X1  g070(.A(KEYINPUT73), .B1(new_n494), .B2(G2105), .ZN(new_n496));
  OAI21_X1  g071(.A(new_n493), .B1(new_n495), .B2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT74), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  INV_X1    g075(.A(G2105), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n500), .B1(new_n501), .B2(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n494), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n503));
  AOI21_X1  g078(.A(new_n492), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  NAND2_X1  g079(.A1(new_n504), .A2(KEYINPUT74), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n499), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT4), .ZN(new_n507));
  OAI211_X1 g082(.A(KEYINPUT75), .B(new_n507), .C1(new_n471), .C2(new_n487), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n479), .A2(G126), .A3(G2105), .ZN(new_n509));
  NAND4_X1  g084(.A1(new_n491), .A2(new_n506), .A3(new_n508), .A4(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(new_n510), .ZN(G164));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n512), .A2(KEYINPUT5), .ZN(new_n513));
  INV_X1    g088(.A(KEYINPUT5), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n514), .A2(G543), .ZN(new_n515));
  AND2_X1   g090(.A1(new_n513), .A2(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  XNOR2_X1  g094(.A(KEYINPUT6), .B(G651), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n516), .A2(new_n520), .ZN(new_n521));
  INV_X1    g096(.A(G88), .ZN(new_n522));
  INV_X1    g097(.A(G50), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n520), .A2(G543), .ZN(new_n524));
  OAI22_X1  g099(.A1(new_n521), .A2(new_n522), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  OR2_X1    g100(.A1(new_n519), .A2(new_n525), .ZN(G303));
  INV_X1    g101(.A(G303), .ZN(G166));
  NAND3_X1  g102(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n528));
  XNOR2_X1  g103(.A(new_n528), .B(KEYINPUT76), .ZN(new_n529));
  XOR2_X1   g104(.A(new_n529), .B(KEYINPUT7), .Z(new_n530));
  AND2_X1   g105(.A1(new_n520), .A2(G543), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G51), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n518), .A2(KEYINPUT6), .ZN(new_n533));
  INV_X1    g108(.A(KEYINPUT6), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(G651), .ZN(new_n535));
  AND4_X1   g110(.A1(new_n513), .A2(new_n515), .A3(new_n533), .A4(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(G89), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n538));
  NAND3_X1  g113(.A1(new_n532), .A2(new_n537), .A3(new_n538), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n530), .A2(new_n539), .ZN(G168));
  AOI22_X1  g115(.A1(new_n531), .A2(G52), .B1(new_n536), .B2(G90), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n542));
  INV_X1    g117(.A(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT77), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(KEYINPUT77), .ZN(new_n545));
  OAI21_X1  g120(.A(new_n541), .B1(new_n544), .B2(new_n545), .ZN(G301));
  INV_X1    g121(.A(G301), .ZN(G171));
  AOI22_X1  g122(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n548), .A2(new_n518), .ZN(new_n549));
  INV_X1    g124(.A(G81), .ZN(new_n550));
  INV_X1    g125(.A(G43), .ZN(new_n551));
  OAI22_X1  g126(.A1(new_n521), .A2(new_n550), .B1(new_n551), .B2(new_n524), .ZN(new_n552));
  NOR2_X1   g127(.A1(new_n549), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G860), .ZN(G153));
  AND3_X1   g129(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G36), .ZN(G176));
  NAND2_X1  g131(.A1(G1), .A2(G3), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT8), .ZN(new_n558));
  NAND2_X1  g133(.A1(new_n555), .A2(new_n558), .ZN(G188));
  NAND2_X1  g134(.A1(new_n531), .A2(G53), .ZN(new_n560));
  INV_X1    g135(.A(KEYINPUT9), .ZN(new_n561));
  XNOR2_X1  g136(.A(new_n560), .B(new_n561), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n536), .A2(G91), .ZN(new_n563));
  AOI22_X1  g138(.A1(new_n516), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n564));
  OAI21_X1  g139(.A(new_n563), .B1(new_n564), .B2(new_n518), .ZN(new_n565));
  NOR2_X1   g140(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  INV_X1    g141(.A(new_n566), .ZN(G299));
  INV_X1    g142(.A(G168), .ZN(G286));
  NAND2_X1  g143(.A1(new_n531), .A2(G49), .ZN(new_n569));
  OAI21_X1  g144(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n536), .A2(G87), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n569), .A2(new_n570), .A3(new_n571), .ZN(G288));
  INV_X1    g147(.A(KEYINPUT79), .ZN(new_n573));
  INV_X1    g148(.A(G86), .ZN(new_n574));
  OAI21_X1  g149(.A(new_n573), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  NAND4_X1  g150(.A1(new_n533), .A2(new_n535), .A3(G48), .A4(G543), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT80), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g153(.A1(new_n520), .A2(KEYINPUT80), .A3(G48), .A4(G543), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n536), .A2(KEYINPUT79), .A3(G86), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n575), .A2(new_n580), .A3(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n513), .A2(new_n515), .A3(G61), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT78), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND4_X1  g160(.A1(new_n513), .A2(new_n515), .A3(KEYINPUT78), .A4(G61), .ZN(new_n586));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n585), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n588), .A2(G651), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n582), .A2(new_n589), .ZN(G305));
  XOR2_X1   g165(.A(KEYINPUT81), .B(G85), .Z(new_n591));
  AOI22_X1  g166(.A1(new_n531), .A2(G47), .B1(new_n536), .B2(new_n591), .ZN(new_n592));
  AOI22_X1  g167(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  OAI21_X1  g168(.A(new_n592), .B1(new_n518), .B2(new_n593), .ZN(G290));
  NAND2_X1  g169(.A1(G301), .A2(G868), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n536), .A2(G92), .ZN(new_n596));
  XOR2_X1   g171(.A(new_n596), .B(KEYINPUT82), .Z(new_n597));
  NAND2_X1  g172(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n516), .A2(G66), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  XNOR2_X1  g175(.A(new_n600), .B(KEYINPUT83), .ZN(new_n601));
  AOI21_X1  g176(.A(new_n518), .B1(new_n599), .B2(new_n601), .ZN(new_n602));
  AOI21_X1  g177(.A(new_n602), .B1(G54), .B2(new_n531), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n598), .A2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n597), .A2(KEYINPUT10), .ZN(new_n605));
  NOR2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G284));
  OAI21_X1  g182(.A(new_n595), .B1(new_n606), .B2(G868), .ZN(G321));
  NAND2_X1  g183(.A1(G286), .A2(G868), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n609), .B1(G868), .B2(new_n566), .ZN(G297));
  OAI21_X1  g185(.A(new_n609), .B1(G868), .B2(new_n566), .ZN(G280));
  INV_X1    g186(.A(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n606), .B1(new_n612), .B2(G860), .ZN(G148));
  OR2_X1    g188(.A1(new_n604), .A2(new_n605), .ZN(new_n614));
  OAI21_X1  g189(.A(G868), .B1(new_n614), .B2(G559), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n615), .B1(G868), .B2(new_n553), .ZN(G323));
  XNOR2_X1  g191(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g192(.A1(new_n481), .A2(G123), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n618), .B(KEYINPUT84), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n482), .A2(G135), .ZN(new_n620));
  NOR2_X1   g195(.A1(new_n474), .A2(G111), .ZN(new_n621));
  OAI21_X1  g196(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n622));
  OAI211_X1 g197(.A(new_n619), .B(new_n620), .C1(new_n621), .C2(new_n622), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2096), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n479), .A2(new_n464), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(KEYINPUT12), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT13), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2100), .ZN(new_n628));
  NAND2_X1  g203(.A1(new_n624), .A2(new_n628), .ZN(G156));
  INV_X1    g204(.A(KEYINPUT14), .ZN(new_n630));
  XNOR2_X1  g205(.A(KEYINPUT15), .B(G2430), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n631), .B(G2435), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2427), .B(G2438), .ZN(new_n633));
  AOI21_X1  g208(.A(new_n630), .B1(new_n632), .B2(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n634), .B1(new_n633), .B2(new_n632), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2451), .B(G2454), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT16), .B(G1341), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(G2443), .B(G2446), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n638), .B(new_n640), .ZN(new_n641));
  OAI21_X1  g216(.A(G14), .B1(new_n635), .B2(new_n641), .ZN(new_n642));
  AOI21_X1  g217(.A(new_n642), .B1(new_n635), .B2(new_n641), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(new_n644), .B(KEYINPUT17), .Z(new_n645));
  XOR2_X1   g220(.A(G2084), .B(G2090), .Z(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  NOR2_X1   g223(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g224(.A1(new_n647), .A2(new_n648), .ZN(new_n650));
  INV_X1    g225(.A(new_n650), .ZN(new_n651));
  OR3_X1    g226(.A1(new_n645), .A2(new_n649), .A3(new_n651), .ZN(new_n652));
  NOR3_X1   g227(.A1(new_n647), .A2(new_n644), .A3(new_n648), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT18), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n644), .A2(KEYINPUT85), .ZN(new_n655));
  OR2_X1    g230(.A1(new_n644), .A2(KEYINPUT85), .ZN(new_n656));
  NAND3_X1  g231(.A1(new_n651), .A2(new_n655), .A3(new_n656), .ZN(new_n657));
  NAND3_X1  g232(.A1(new_n652), .A2(new_n654), .A3(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(G2096), .B(G2100), .Z(new_n659));
  XNOR2_X1  g234(.A(new_n658), .B(new_n659), .ZN(G227));
  XNOR2_X1  g235(.A(G1971), .B(G1976), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT19), .ZN(new_n662));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  OR2_X1    g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n663), .A2(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n662), .A2(new_n665), .A3(new_n666), .ZN(new_n667));
  NOR2_X1   g242(.A1(new_n662), .A2(new_n666), .ZN(new_n668));
  INV_X1    g243(.A(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(KEYINPUT20), .ZN(new_n670));
  OAI221_X1 g245(.A(new_n667), .B1(new_n662), .B2(new_n665), .C1(new_n669), .C2(new_n670), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n671), .B1(new_n670), .B2(new_n669), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G1991), .ZN(new_n673));
  INV_X1    g248(.A(G1996), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1981), .B(G1986), .ZN(new_n676));
  XNOR2_X1  g251(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n678));
  NAND2_X1  g253(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  INV_X1    g254(.A(new_n676), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n675), .B(new_n680), .ZN(new_n681));
  INV_X1    g256(.A(new_n678), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n679), .A2(new_n683), .ZN(G229));
  INV_X1    g259(.A(G22), .ZN(new_n685));
  NOR2_X1   g260(.A1(new_n685), .A2(G16), .ZN(new_n686));
  AOI21_X1  g261(.A(new_n686), .B1(G303), .B2(G16), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(G1971), .ZN(new_n688));
  NOR2_X1   g263(.A1(G16), .A2(G23), .ZN(new_n689));
  INV_X1    g264(.A(G288), .ZN(new_n690));
  AOI21_X1  g265(.A(new_n689), .B1(new_n690), .B2(G16), .ZN(new_n691));
  XNOR2_X1  g266(.A(KEYINPUT33), .B(G1976), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n691), .B(new_n692), .ZN(new_n693));
  MUX2_X1   g268(.A(G6), .B(G305), .S(G16), .Z(new_n694));
  XNOR2_X1  g269(.A(KEYINPUT32), .B(G1981), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n695), .B(KEYINPUT87), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n688), .B(new_n693), .C1(new_n694), .C2(new_n696), .ZN(new_n697));
  AOI21_X1  g272(.A(new_n697), .B1(new_n694), .B2(new_n696), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT34), .ZN(new_n699));
  NOR2_X1   g274(.A1(G25), .A2(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n481), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n482), .A2(G131), .ZN(new_n702));
  OAI221_X1 g277(.A(G2104), .B1(G95), .B2(G2105), .C1(new_n474), .C2(G107), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n701), .A2(new_n702), .A3(new_n703), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n700), .B1(new_n705), .B2(G29), .ZN(new_n706));
  XOR2_X1   g281(.A(new_n706), .B(KEYINPUT86), .Z(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT35), .B(G1991), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  MUX2_X1   g285(.A(G24), .B(G290), .S(G16), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(G1986), .ZN(new_n712));
  NOR2_X1   g287(.A1(new_n707), .A2(new_n709), .ZN(new_n713));
  AOI211_X1 g288(.A(new_n712), .B(new_n713), .C1(KEYINPUT89), .C2(KEYINPUT36), .ZN(new_n714));
  NAND3_X1  g289(.A1(new_n699), .A2(new_n710), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g290(.A(KEYINPUT89), .B1(KEYINPUT88), .B2(KEYINPUT36), .ZN(new_n716));
  XOR2_X1   g291(.A(new_n715), .B(new_n716), .Z(new_n717));
  NAND2_X1  g292(.A1(new_n481), .A2(G129), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n482), .A2(G141), .ZN(new_n719));
  NAND3_X1  g294(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n720));
  INV_X1    g295(.A(KEYINPUT26), .ZN(new_n721));
  OR2_X1    g296(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n720), .A2(new_n721), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n722), .A2(new_n723), .B1(G105), .B2(new_n464), .ZN(new_n724));
  AND3_X1   g299(.A1(new_n718), .A2(new_n719), .A3(new_n724), .ZN(new_n725));
  NAND2_X1  g300(.A1(new_n725), .A2(G29), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n726), .B(KEYINPUT92), .ZN(new_n727));
  INV_X1    g302(.A(G29), .ZN(new_n728));
  INV_X1    g303(.A(G32), .ZN(new_n729));
  AOI21_X1  g304(.A(new_n727), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  XOR2_X1   g305(.A(KEYINPUT27), .B(G1996), .Z(new_n731));
  NAND2_X1  g306(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NOR2_X1   g307(.A1(G5), .A2(G16), .ZN(new_n733));
  AOI21_X1  g308(.A(new_n733), .B1(G171), .B2(G16), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT24), .ZN(new_n735));
  INV_X1    g310(.A(G34), .ZN(new_n736));
  AOI21_X1  g311(.A(G29), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(new_n735), .B2(new_n736), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(G160), .B2(new_n728), .ZN(new_n739));
  OAI221_X1 g314(.A(new_n732), .B1(G1961), .B2(new_n734), .C1(G2084), .C2(new_n739), .ZN(new_n740));
  AND2_X1   g315(.A1(new_n740), .A2(KEYINPUT94), .ZN(new_n741));
  OR2_X1    g316(.A1(G29), .A2(G33), .ZN(new_n742));
  NAND3_X1  g317(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n743));
  AOI22_X1  g318(.A1(new_n482), .A2(G139), .B1(KEYINPUT25), .B2(new_n743), .ZN(new_n744));
  AOI22_X1  g319(.A1(new_n479), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n745));
  OAI221_X1 g320(.A(new_n744), .B1(KEYINPUT25), .B2(new_n743), .C1(new_n474), .C2(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT90), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n742), .B1(new_n747), .B2(new_n728), .ZN(new_n748));
  INV_X1    g323(.A(G2072), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(KEYINPUT91), .Z(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G35), .ZN(new_n752));
  AOI21_X1  g327(.A(new_n752), .B1(G162), .B2(G29), .ZN(new_n753));
  XOR2_X1   g328(.A(KEYINPUT95), .B(KEYINPUT29), .Z(new_n754));
  XNOR2_X1  g329(.A(new_n753), .B(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2090), .ZN(new_n756));
  NOR2_X1   g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n751), .B1(KEYINPUT97), .B2(new_n757), .ZN(new_n758));
  AOI211_X1 g333(.A(new_n741), .B(new_n758), .C1(KEYINPUT97), .C2(new_n757), .ZN(new_n759));
  XNOR2_X1  g334(.A(KEYINPUT31), .B(G11), .ZN(new_n760));
  INV_X1    g335(.A(G28), .ZN(new_n761));
  AOI21_X1  g336(.A(G29), .B1(new_n761), .B2(KEYINPUT30), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n762), .A2(KEYINPUT93), .ZN(new_n763));
  INV_X1    g338(.A(new_n763), .ZN(new_n764));
  OAI22_X1  g339(.A1(new_n762), .A2(KEYINPUT93), .B1(KEYINPUT30), .B2(new_n761), .ZN(new_n765));
  OAI221_X1 g340(.A(new_n760), .B1(new_n764), .B2(new_n765), .C1(new_n623), .C2(new_n728), .ZN(new_n766));
  INV_X1    g341(.A(new_n553), .ZN(new_n767));
  MUX2_X1   g342(.A(G19), .B(new_n767), .S(G16), .Z(new_n768));
  XNOR2_X1  g343(.A(new_n768), .B(G1341), .ZN(new_n769));
  AOI211_X1 g344(.A(new_n766), .B(new_n769), .C1(G2084), .C2(new_n739), .ZN(new_n770));
  MUX2_X1   g345(.A(G21), .B(G286), .S(G16), .Z(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1966), .Z(new_n772));
  MUX2_X1   g347(.A(G4), .B(new_n614), .S(G16), .Z(new_n773));
  OAI211_X1 g348(.A(new_n770), .B(new_n772), .C1(G1348), .C2(new_n773), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n728), .A2(G27), .ZN(new_n775));
  OAI21_X1  g350(.A(new_n775), .B1(G164), .B2(new_n728), .ZN(new_n776));
  XNOR2_X1  g351(.A(new_n776), .B(G2078), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n734), .A2(G1961), .ZN(new_n778));
  INV_X1    g353(.A(KEYINPUT28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n481), .A2(G128), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n482), .A2(G140), .ZN(new_n781));
  OAI221_X1 g356(.A(G2104), .B1(G104), .B2(G2105), .C1(new_n474), .C2(G116), .ZN(new_n782));
  NAND3_X1  g357(.A1(new_n780), .A2(new_n781), .A3(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n783), .A2(G29), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n728), .A2(G26), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n779), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI21_X1  g361(.A(new_n786), .B1(new_n779), .B2(new_n785), .ZN(new_n787));
  INV_X1    g362(.A(G2067), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n778), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n787), .A2(new_n788), .ZN(new_n790));
  OAI21_X1  g365(.A(new_n790), .B1(new_n730), .B2(new_n731), .ZN(new_n791));
  NOR4_X1   g366(.A1(new_n774), .A2(new_n777), .A3(new_n789), .A4(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n755), .A2(new_n756), .ZN(new_n793));
  OAI22_X1  g368(.A1(new_n740), .A2(KEYINPUT94), .B1(KEYINPUT96), .B2(new_n793), .ZN(new_n794));
  INV_X1    g369(.A(KEYINPUT23), .ZN(new_n795));
  INV_X1    g370(.A(G20), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G16), .ZN(new_n797));
  AOI211_X1 g372(.A(new_n795), .B(new_n797), .C1(G299), .C2(G16), .ZN(new_n798));
  AOI21_X1  g373(.A(new_n798), .B1(new_n795), .B2(new_n797), .ZN(new_n799));
  XOR2_X1   g374(.A(new_n799), .B(G1956), .Z(new_n800));
  NAND2_X1  g375(.A1(new_n773), .A2(G1348), .ZN(new_n801));
  OAI211_X1 g376(.A(new_n800), .B(new_n801), .C1(new_n749), .C2(new_n748), .ZN(new_n802));
  AOI211_X1 g377(.A(new_n794), .B(new_n802), .C1(KEYINPUT96), .C2(new_n793), .ZN(new_n803));
  NAND4_X1  g378(.A1(new_n717), .A2(new_n759), .A3(new_n792), .A4(new_n803), .ZN(G150));
  INV_X1    g379(.A(G150), .ZN(G311));
  NAND2_X1  g380(.A1(new_n606), .A2(G559), .ZN(new_n806));
  INV_X1    g381(.A(G93), .ZN(new_n807));
  INV_X1    g382(.A(G55), .ZN(new_n808));
  OAI22_X1  g383(.A1(new_n521), .A2(new_n807), .B1(new_n808), .B2(new_n524), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n516), .A2(G67), .ZN(new_n810));
  NAND2_X1  g385(.A1(G80), .A2(G543), .ZN(new_n811));
  AOI21_X1  g386(.A(new_n518), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n809), .A2(new_n812), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n813), .B(KEYINPUT98), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n814), .B(new_n553), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n806), .B(new_n815), .ZN(new_n816));
  INV_X1    g391(.A(new_n816), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n818));
  AOI21_X1  g393(.A(G860), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  OAI21_X1  g394(.A(new_n819), .B1(new_n818), .B2(new_n817), .ZN(new_n820));
  OAI21_X1  g395(.A(G860), .B1(new_n809), .B2(new_n812), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n821), .B(KEYINPUT37), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n820), .A2(new_n822), .ZN(G145));
  XNOR2_X1  g398(.A(G162), .B(new_n725), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n623), .B(G160), .ZN(new_n825));
  XOR2_X1   g400(.A(new_n824), .B(new_n825), .Z(new_n826));
  XNOR2_X1  g401(.A(new_n783), .B(new_n704), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n827), .B(new_n510), .ZN(new_n828));
  OAI21_X1  g403(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n474), .A2(G118), .ZN(new_n830));
  AOI21_X1  g405(.A(new_n829), .B1(new_n830), .B2(KEYINPUT99), .ZN(new_n831));
  OAI21_X1  g406(.A(new_n831), .B1(KEYINPUT99), .B2(new_n830), .ZN(new_n832));
  AOI22_X1  g407(.A1(G130), .A2(new_n481), .B1(new_n482), .B2(G142), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n832), .A2(new_n833), .ZN(new_n834));
  OR2_X1    g409(.A1(new_n828), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n828), .A2(new_n834), .ZN(new_n836));
  AND2_X1   g411(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n826), .A2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n824), .B(new_n825), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n835), .A2(new_n836), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n838), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n747), .B(new_n626), .ZN(new_n843));
  INV_X1    g418(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g419(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G37), .ZN(new_n846));
  NAND3_X1  g421(.A1(new_n838), .A2(new_n843), .A3(new_n841), .ZN(new_n847));
  NAND3_X1  g422(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g423(.A1(new_n848), .A2(KEYINPUT100), .ZN(new_n849));
  INV_X1    g424(.A(KEYINPUT100), .ZN(new_n850));
  NAND4_X1  g425(.A1(new_n845), .A2(new_n850), .A3(new_n846), .A4(new_n847), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n849), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n852), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g428(.A(G305), .B(G288), .ZN(new_n854));
  XOR2_X1   g429(.A(G303), .B(G290), .Z(new_n855));
  XNOR2_X1  g430(.A(new_n854), .B(new_n855), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n858), .B(KEYINPUT42), .Z(new_n859));
  NAND2_X1  g434(.A1(new_n606), .A2(new_n612), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n815), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n614), .A2(new_n566), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n606), .A2(G299), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g439(.A1(new_n861), .A2(new_n864), .ZN(new_n865));
  AND3_X1   g440(.A1(new_n862), .A2(KEYINPUT41), .A3(new_n863), .ZN(new_n866));
  AOI21_X1  g441(.A(KEYINPUT41), .B1(new_n862), .B2(new_n863), .ZN(new_n867));
  OAI21_X1  g442(.A(KEYINPUT101), .B1(new_n866), .B2(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  INV_X1    g444(.A(KEYINPUT101), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n868), .A2(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n861), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n872), .A2(new_n873), .ZN(new_n874));
  AND3_X1   g449(.A1(new_n859), .A2(new_n865), .A3(new_n874), .ZN(new_n875));
  AOI21_X1  g450(.A(new_n859), .B1(new_n874), .B2(new_n865), .ZN(new_n876));
  OAI21_X1  g451(.A(G868), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  OAI21_X1  g452(.A(new_n877), .B1(G868), .B2(new_n813), .ZN(G295));
  OAI21_X1  g453(.A(new_n877), .B1(G868), .B2(new_n813), .ZN(G331));
  INV_X1    g454(.A(new_n864), .ZN(new_n880));
  XNOR2_X1  g455(.A(G286), .B(G301), .ZN(new_n881));
  OR2_X1    g456(.A1(new_n815), .A2(new_n881), .ZN(new_n882));
  INV_X1    g457(.A(KEYINPUT104), .ZN(new_n883));
  NAND2_X1  g458(.A1(new_n815), .A2(new_n881), .ZN(new_n884));
  NAND3_X1  g459(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND3_X1  g460(.A1(new_n815), .A2(KEYINPUT104), .A3(new_n881), .ZN(new_n886));
  AOI21_X1  g461(.A(new_n880), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n882), .A2(KEYINPUT103), .A3(new_n884), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT103), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n815), .A2(new_n889), .A3(new_n881), .ZN(new_n890));
  AND2_X1   g465(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  AOI21_X1  g466(.A(new_n887), .B1(new_n872), .B2(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(G37), .B1(new_n892), .B2(new_n857), .ZN(new_n893));
  AOI21_X1  g468(.A(new_n880), .B1(new_n888), .B2(new_n890), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT105), .ZN(new_n895));
  AND2_X1   g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OAI211_X1 g471(.A(new_n885), .B(new_n886), .C1(new_n866), .C2(new_n867), .ZN(new_n897));
  OAI21_X1  g472(.A(new_n897), .B1(new_n894), .B2(new_n895), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n856), .B1(new_n896), .B2(new_n898), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n893), .A2(new_n899), .A3(KEYINPUT43), .ZN(new_n900));
  OR2_X1    g475(.A1(new_n892), .A2(new_n857), .ZN(new_n901));
  AOI21_X1  g476(.A(KEYINPUT43), .B1(new_n901), .B2(new_n893), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT44), .B1(new_n900), .B2(new_n902), .ZN(new_n903));
  INV_X1    g478(.A(KEYINPUT44), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT43), .ZN(new_n905));
  AND3_X1   g480(.A1(new_n893), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  AOI21_X1  g481(.A(new_n905), .B1(new_n901), .B2(new_n893), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n903), .A2(new_n908), .ZN(G397));
  XNOR2_X1  g484(.A(new_n725), .B(G1996), .ZN(new_n910));
  XNOR2_X1  g485(.A(new_n783), .B(new_n788), .ZN(new_n911));
  XNOR2_X1  g486(.A(new_n704), .B(new_n709), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n910), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  NOR2_X1   g488(.A1(G290), .A2(G1986), .ZN(new_n914));
  AND2_X1   g489(.A1(G290), .A2(G1986), .ZN(new_n915));
  OR3_X1    g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(G1384), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n504), .A2(KEYINPUT74), .ZN(new_n918));
  AOI211_X1 g493(.A(new_n498), .B(new_n492), .C1(new_n502), .C2(new_n503), .ZN(new_n919));
  OAI211_X1 g494(.A(new_n508), .B(new_n509), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n488), .A2(KEYINPUT4), .A3(new_n490), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n917), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(KEYINPUT45), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  XOR2_X1   g499(.A(KEYINPUT106), .B(G40), .Z(new_n925));
  NOR3_X1   g500(.A1(new_n473), .A2(new_n477), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n926), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n924), .A2(new_n927), .ZN(new_n928));
  AND2_X1   g503(.A1(new_n916), .A2(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n930), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n931));
  INV_X1    g506(.A(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n930), .B1(new_n510), .B2(new_n917), .ZN(new_n933));
  NOR3_X1   g508(.A1(new_n932), .A2(new_n933), .A3(new_n927), .ZN(new_n934));
  OAI211_X1 g509(.A(KEYINPUT45), .B(new_n917), .C1(new_n920), .C2(new_n921), .ZN(new_n935));
  NAND3_X1  g510(.A1(new_n924), .A2(new_n926), .A3(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(G1971), .ZN(new_n937));
  AOI22_X1  g512(.A1(new_n934), .A2(new_n756), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT107), .ZN(new_n939));
  INV_X1    g514(.A(new_n935), .ZN(new_n940));
  AOI21_X1  g515(.A(KEYINPUT45), .B1(new_n510), .B2(new_n917), .ZN(new_n941));
  NOR3_X1   g516(.A1(new_n940), .A2(new_n941), .A3(new_n927), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n922), .A2(KEYINPUT50), .ZN(new_n943));
  NAND3_X1  g518(.A1(new_n943), .A2(new_n926), .A3(new_n931), .ZN(new_n944));
  OAI22_X1  g519(.A1(new_n942), .A2(G1971), .B1(new_n944), .B2(G2090), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT107), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(G303), .A2(G8), .ZN(new_n948));
  XNOR2_X1  g523(.A(new_n948), .B(KEYINPUT55), .ZN(new_n949));
  INV_X1    g524(.A(new_n949), .ZN(new_n950));
  AND4_X1   g525(.A1(G8), .A2(new_n939), .A3(new_n947), .A4(new_n950), .ZN(new_n951));
  OAI211_X1 g526(.A(new_n917), .B(new_n926), .C1(new_n920), .C2(new_n921), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n690), .A2(G1976), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n952), .A2(G8), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n954), .A2(KEYINPUT52), .ZN(new_n955));
  INV_X1    g530(.A(G1976), .ZN(new_n956));
  AOI21_X1  g531(.A(KEYINPUT52), .B1(G288), .B2(new_n956), .ZN(new_n957));
  NAND4_X1  g532(.A1(new_n952), .A2(new_n957), .A3(G8), .A4(new_n953), .ZN(new_n958));
  AND2_X1   g533(.A1(new_n955), .A2(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n952), .ZN(new_n960));
  INV_X1    g535(.A(G8), .ZN(new_n961));
  NOR2_X1   g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  AOI22_X1  g537(.A1(new_n578), .A2(new_n579), .B1(new_n536), .B2(G86), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT108), .ZN(new_n964));
  OAI21_X1  g539(.A(new_n589), .B1(new_n963), .B2(new_n964), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n536), .A2(G86), .ZN(new_n966));
  AND3_X1   g541(.A1(new_n580), .A2(new_n964), .A3(new_n966), .ZN(new_n967));
  OAI21_X1  g542(.A(G1981), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  INV_X1    g543(.A(G1981), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n582), .A2(new_n969), .A3(new_n589), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(KEYINPUT49), .A3(new_n970), .ZN(new_n971));
  AOI21_X1  g546(.A(KEYINPUT49), .B1(new_n968), .B2(new_n970), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT109), .ZN(new_n973));
  OAI211_X1 g548(.A(new_n962), .B(new_n971), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  AOI211_X1 g549(.A(KEYINPUT109), .B(KEYINPUT49), .C1(new_n968), .C2(new_n970), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n959), .B1(new_n974), .B2(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(new_n976), .ZN(new_n977));
  OAI211_X1 g552(.A(new_n956), .B(new_n690), .C1(new_n974), .C2(new_n975), .ZN(new_n978));
  XNOR2_X1  g553(.A(new_n970), .B(KEYINPUT110), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n978), .A2(new_n979), .ZN(new_n980));
  AOI22_X1  g555(.A1(new_n951), .A2(new_n977), .B1(new_n980), .B2(new_n962), .ZN(new_n981));
  AOI21_X1  g556(.A(new_n927), .B1(new_n922), .B2(KEYINPUT50), .ZN(new_n982));
  INV_X1    g557(.A(G2084), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n982), .A2(new_n983), .A3(new_n931), .ZN(new_n984));
  OAI211_X1 g559(.A(G168), .B(new_n984), .C1(new_n942), .C2(G1966), .ZN(new_n985));
  INV_X1    g560(.A(KEYINPUT51), .ZN(new_n986));
  AND2_X1   g561(.A1(KEYINPUT119), .A2(G8), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n985), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  OAI21_X1  g563(.A(new_n984), .B1(new_n942), .B2(G1966), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n989), .A2(G8), .A3(G286), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(new_n990), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n986), .B1(new_n985), .B2(new_n987), .ZN(new_n992));
  OAI21_X1  g567(.A(KEYINPUT62), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g568(.A1(new_n985), .A2(new_n987), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(KEYINPUT51), .ZN(new_n995));
  INV_X1    g570(.A(KEYINPUT62), .ZN(new_n996));
  NAND4_X1  g571(.A1(new_n995), .A2(new_n996), .A3(new_n990), .A4(new_n988), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n993), .A2(new_n997), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n976), .A2(KEYINPUT111), .ZN(new_n999));
  INV_X1    g574(.A(KEYINPUT111), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n959), .B(new_n1000), .C1(new_n974), .C2(new_n975), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n999), .A2(new_n1001), .ZN(new_n1002));
  NAND4_X1  g577(.A1(new_n939), .A2(new_n947), .A3(G8), .A4(new_n950), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n949), .B1(new_n938), .B2(new_n961), .ZN(new_n1004));
  INV_X1    g579(.A(G2078), .ZN(new_n1005));
  NAND4_X1  g580(.A1(new_n924), .A2(new_n1005), .A3(new_n926), .A4(new_n935), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT121), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n941), .A2(new_n927), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1011));
  NAND4_X1  g586(.A1(new_n1009), .A2(new_n1005), .A3(new_n935), .A4(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n1008), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g588(.A(KEYINPUT122), .B(G1961), .Z(new_n1014));
  AOI22_X1  g589(.A1(new_n1010), .A2(new_n1006), .B1(new_n944), .B2(new_n1014), .ZN(new_n1015));
  AOI21_X1  g590(.A(G301), .B1(new_n1013), .B2(new_n1015), .ZN(new_n1016));
  NAND4_X1  g591(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(new_n981), .B1(new_n998), .B2(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1348), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n944), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(KEYINPUT115), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n952), .A2(G2067), .ZN(new_n1022));
  INV_X1    g597(.A(new_n1022), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1020), .A2(new_n1021), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1348), .B1(new_n982), .B2(new_n931), .ZN(new_n1025));
  OAI21_X1  g600(.A(KEYINPUT115), .B1(new_n1025), .B2(new_n1022), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1024), .A2(new_n1026), .A3(new_n606), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n566), .A2(KEYINPUT57), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT57), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1029), .B1(new_n562), .B2(new_n565), .ZN(new_n1030));
  AND2_X1   g605(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1031));
  XOR2_X1   g606(.A(KEYINPUT56), .B(G2072), .Z(new_n1032));
  XNOR2_X1  g607(.A(new_n1032), .B(KEYINPUT114), .ZN(new_n1033));
  NAND4_X1  g608(.A1(new_n924), .A2(new_n926), .A3(new_n935), .A4(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1034), .ZN(new_n1035));
  XNOR2_X1  g610(.A(KEYINPUT113), .B(G1956), .ZN(new_n1036));
  AOI21_X1  g611(.A(new_n1036), .B1(new_n982), .B2(new_n931), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1031), .B1(new_n1035), .B2(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1027), .A2(new_n1038), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1028), .A2(new_n1030), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1040), .B(new_n1034), .C1(new_n934), .C2(new_n1036), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1039), .A2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND3_X1  g619(.A1(new_n1039), .A2(KEYINPUT116), .A3(new_n1041), .ZN(new_n1045));
  NAND3_X1  g620(.A1(new_n1038), .A2(new_n1041), .A3(KEYINPUT61), .ZN(new_n1046));
  XOR2_X1   g621(.A(KEYINPUT58), .B(G1341), .Z(new_n1047));
  NAND2_X1  g622(.A1(new_n952), .A2(new_n1047), .ZN(new_n1048));
  OAI21_X1  g623(.A(new_n1048), .B1(new_n936), .B2(G1996), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1049), .A2(new_n553), .ZN(new_n1050));
  XNOR2_X1  g625(.A(new_n1050), .B(KEYINPUT59), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1038), .A2(new_n1041), .ZN(new_n1052));
  XNOR2_X1  g627(.A(KEYINPUT117), .B(KEYINPUT61), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT118), .B1(new_n1052), .B2(new_n1054), .ZN(new_n1055));
  INV_X1    g630(.A(KEYINPUT118), .ZN(new_n1056));
  AOI211_X1 g631(.A(new_n1056), .B(new_n1053), .C1(new_n1038), .C2(new_n1041), .ZN(new_n1057));
  OAI211_X1 g632(.A(new_n1046), .B(new_n1051), .C1(new_n1055), .C2(new_n1057), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1021), .B1(new_n1020), .B2(new_n1023), .ZN(new_n1059));
  AOI211_X1 g634(.A(KEYINPUT115), .B(new_n1022), .C1(new_n944), .C2(new_n1019), .ZN(new_n1060));
  NOR3_X1   g635(.A1(new_n1059), .A2(new_n1060), .A3(KEYINPUT60), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT60), .B1(new_n1059), .B2(new_n1060), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(new_n606), .ZN(new_n1063));
  OAI211_X1 g638(.A(KEYINPUT60), .B(new_n614), .C1(new_n1059), .C2(new_n1060), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1061), .B1(new_n1063), .B2(new_n1064), .ZN(new_n1065));
  OAI211_X1 g640(.A(new_n1044), .B(new_n1045), .C1(new_n1058), .C2(new_n1065), .ZN(new_n1066));
  XNOR2_X1  g641(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n1067));
  NOR3_X1   g642(.A1(new_n940), .A2(new_n1010), .A3(G2078), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT124), .ZN(new_n1069));
  OR2_X1    g644(.A1(new_n473), .A2(KEYINPUT123), .ZN(new_n1070));
  INV_X1    g645(.A(new_n477), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n473), .A2(KEYINPUT123), .ZN(new_n1072));
  NAND4_X1  g647(.A1(new_n1070), .A2(G40), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1073), .ZN(new_n1074));
  NAND3_X1  g649(.A1(new_n924), .A2(new_n1069), .A3(new_n1074), .ZN(new_n1075));
  OAI21_X1  g650(.A(KEYINPUT124), .B1(new_n941), .B2(new_n1073), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1068), .A2(new_n1075), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1015), .A2(G301), .A3(new_n1077), .ZN(new_n1078));
  OAI21_X1  g653(.A(new_n1067), .B1(new_n1016), .B2(new_n1078), .ZN(new_n1079));
  NAND3_X1  g654(.A1(new_n1013), .A2(G301), .A3(new_n1015), .ZN(new_n1080));
  AND2_X1   g655(.A1(new_n1015), .A2(new_n1077), .ZN(new_n1081));
  OAI211_X1 g656(.A(new_n1080), .B(KEYINPUT54), .C1(G301), .C2(new_n1081), .ZN(new_n1082));
  NAND3_X1  g657(.A1(new_n995), .A2(new_n990), .A3(new_n988), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n1079), .A2(new_n1082), .A3(new_n1083), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1084), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1018), .B1(new_n1066), .B2(new_n1086), .ZN(new_n1087));
  XOR2_X1   g662(.A(KEYINPUT112), .B(KEYINPUT63), .Z(new_n1088));
  NAND3_X1  g663(.A1(new_n989), .A2(G8), .A3(G168), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1088), .B1(new_n1085), .B2(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n939), .A2(new_n947), .A3(G8), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(new_n949), .ZN(new_n1092));
  INV_X1    g667(.A(new_n1089), .ZN(new_n1093));
  NAND4_X1  g668(.A1(new_n1092), .A2(KEYINPUT63), .A3(new_n977), .A4(new_n1093), .ZN(new_n1094));
  NAND2_X1  g669(.A1(new_n1090), .A2(new_n1094), .ZN(new_n1095));
  AOI21_X1  g670(.A(new_n929), .B1(new_n1087), .B2(new_n1095), .ZN(new_n1096));
  NAND2_X1  g671(.A1(new_n928), .A2(new_n674), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT126), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT46), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1100));
  XNOR2_X1  g675(.A(new_n1097), .B(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n911), .A2(new_n725), .ZN(new_n1102));
  AOI22_X1  g677(.A1(new_n1102), .A2(new_n928), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n1104), .B(KEYINPUT47), .ZN(new_n1105));
  AOI21_X1  g680(.A(KEYINPUT48), .B1(new_n928), .B2(new_n914), .ZN(new_n1106));
  AOI21_X1  g681(.A(new_n1106), .B1(new_n928), .B2(new_n913), .ZN(new_n1107));
  NAND3_X1  g682(.A1(new_n928), .A2(KEYINPUT48), .A3(new_n914), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n705), .A2(new_n709), .ZN(new_n1109));
  XNOR2_X1  g684(.A(new_n1109), .B(KEYINPUT125), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n910), .A2(new_n911), .ZN(new_n1111));
  OAI22_X1  g686(.A1(new_n1110), .A2(new_n1111), .B1(G2067), .B2(new_n783), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1107), .A2(new_n1108), .B1(new_n928), .B2(new_n1112), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1105), .A2(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(KEYINPUT127), .B1(new_n1096), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1066), .A2(new_n1086), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1018), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1116), .A2(new_n1095), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g693(.A(new_n929), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT127), .ZN(new_n1121));
  INV_X1    g696(.A(new_n1114), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1120), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1115), .A2(new_n1123), .ZN(G329));
  assign    G231 = 1'b0;
  OR3_X1    g699(.A1(G227), .A2(new_n461), .A3(G401), .ZN(new_n1126));
  NOR2_X1   g700(.A1(G229), .A2(new_n1126), .ZN(new_n1127));
  OAI211_X1 g701(.A(new_n1127), .B(new_n852), .C1(new_n906), .C2(new_n907), .ZN(G225));
  INV_X1    g702(.A(G225), .ZN(G308));
endmodule


