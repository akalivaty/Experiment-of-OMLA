//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 0 0 0 0 0 1 1 1 1 1 1 1 1 1 1 1 1 1 1 0 1 1 1 0 1 1 0 1 1 0 1 0 0 1 1 0 1 0 0 1 0 1 0 0 1 0 1 1 0 0 1 0 1 0 1 1 1 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:06 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n734, new_n735, new_n736,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n813, new_n814, new_n815, new_n816, new_n818, new_n819, new_n820,
    new_n821, new_n822, new_n823, new_n825, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n903,
    new_n904, new_n905, new_n907, new_n908, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n958, new_n959,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n972, new_n973, new_n974, new_n976,
    new_n977, new_n978, new_n979, new_n980, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n995, new_n996, new_n997, new_n998, new_n999,
    new_n1000, new_n1001, new_n1002, new_n1003, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1017, new_n1018;
  AOI21_X1  g000(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n202));
  OR2_X1    g001(.A1(new_n202), .A2(KEYINPUT96), .ZN(new_n203));
  XOR2_X1   g002(.A(G57gat), .B(G64gat), .Z(new_n204));
  NAND2_X1  g003(.A1(new_n202), .A2(KEYINPUT96), .ZN(new_n205));
  NAND3_X1  g004(.A1(new_n203), .A2(new_n204), .A3(new_n205), .ZN(new_n206));
  XNOR2_X1  g005(.A(G71gat), .B(G78gat), .ZN(new_n207));
  INV_X1    g006(.A(new_n207), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND4_X1  g008(.A1(new_n203), .A2(new_n204), .A3(new_n207), .A4(new_n205), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT21), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  NAND2_X1  g012(.A1(G231gat), .A2(G233gat), .ZN(new_n214));
  XNOR2_X1  g013(.A(new_n213), .B(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(G127gat), .ZN(new_n216));
  XNOR2_X1  g015(.A(new_n215), .B(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G15gat), .B(G22gat), .ZN(new_n218));
  INV_X1    g017(.A(G1gat), .ZN(new_n219));
  NAND2_X1  g018(.A1(new_n219), .A2(KEYINPUT16), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n218), .A2(new_n220), .ZN(new_n221));
  OAI21_X1  g020(.A(new_n221), .B1(G1gat), .B2(new_n218), .ZN(new_n222));
  OR2_X1    g021(.A1(new_n222), .A2(G8gat), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n222), .A2(G8gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  NOR2_X1   g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  INV_X1    g026(.A(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(KEYINPUT92), .B1(new_n223), .B2(new_n224), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  OAI211_X1 g029(.A(new_n228), .B(new_n230), .C1(new_n212), .C2(new_n211), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n217), .B(new_n231), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n233));
  INV_X1    g032(.A(G155gat), .ZN(new_n234));
  XNOR2_X1  g033(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g034(.A(G183gat), .B(G211gat), .ZN(new_n236));
  XOR2_X1   g035(.A(new_n235), .B(new_n236), .Z(new_n237));
  NAND2_X1  g036(.A1(new_n232), .A2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(new_n231), .ZN(new_n239));
  XNOR2_X1  g038(.A(new_n217), .B(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(new_n237), .ZN(new_n241));
  NAND2_X1  g040(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n238), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(new_n243), .ZN(new_n244));
  XNOR2_X1  g043(.A(G190gat), .B(G218gat), .ZN(new_n245));
  INV_X1    g044(.A(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT17), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT15), .ZN(new_n248));
  INV_X1    g047(.A(G50gat), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n249), .A2(KEYINPUT88), .A3(G43gat), .ZN(new_n250));
  XOR2_X1   g049(.A(G43gat), .B(G50gat), .Z(new_n251));
  OAI211_X1 g050(.A(new_n248), .B(new_n250), .C1(new_n251), .C2(KEYINPUT88), .ZN(new_n252));
  XNOR2_X1  g051(.A(G43gat), .B(G50gat), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n253), .A2(KEYINPUT15), .ZN(new_n254));
  INV_X1    g053(.A(G29gat), .ZN(new_n255));
  INV_X1    g054(.A(G36gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(KEYINPUT14), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT14), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(G29gat), .B2(G36gat), .ZN(new_n259));
  NAND2_X1  g058(.A1(G29gat), .A2(G36gat), .ZN(new_n260));
  AND3_X1   g059(.A1(new_n257), .A2(new_n259), .A3(new_n260), .ZN(new_n261));
  AND3_X1   g060(.A1(new_n252), .A2(new_n254), .A3(new_n261), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n261), .A2(new_n254), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT89), .ZN(new_n264));
  NOR2_X1   g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NOR2_X1   g064(.A1(new_n262), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n252), .A2(new_n254), .A3(new_n261), .ZN(new_n267));
  NOR2_X1   g066(.A1(new_n267), .A2(new_n264), .ZN(new_n268));
  OAI21_X1  g067(.A(new_n247), .B1(new_n266), .B2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n262), .A2(KEYINPUT89), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n267), .B1(new_n264), .B2(new_n263), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n270), .A2(new_n271), .A3(KEYINPUT17), .ZN(new_n272));
  NAND2_X1  g071(.A1(G99gat), .A2(G106gat), .ZN(new_n273));
  INV_X1    g072(.A(G85gat), .ZN(new_n274));
  INV_X1    g073(.A(G92gat), .ZN(new_n275));
  AOI22_X1  g074(.A1(KEYINPUT8), .A2(new_n273), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT7), .ZN(new_n277));
  OAI21_X1  g076(.A(new_n277), .B1(new_n274), .B2(new_n275), .ZN(new_n278));
  NAND3_X1  g077(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n276), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(G99gat), .B(G106gat), .Z(new_n281));
  OR2_X1    g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n281), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n282), .A2(KEYINPUT99), .A3(new_n283), .ZN(new_n284));
  OR2_X1    g083(.A1(new_n283), .A2(KEYINPUT99), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n284), .A2(new_n285), .ZN(new_n286));
  INV_X1    g085(.A(KEYINPUT100), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n284), .A2(KEYINPUT100), .A3(new_n285), .ZN(new_n289));
  NAND4_X1  g088(.A1(new_n269), .A2(new_n272), .A3(new_n288), .A4(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n270), .A2(new_n271), .ZN(new_n291));
  NAND2_X1  g090(.A1(G232gat), .A2(G233gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT97), .ZN(new_n293));
  INV_X1    g092(.A(new_n293), .ZN(new_n294));
  AOI22_X1  g093(.A1(new_n291), .A2(new_n286), .B1(KEYINPUT41), .B2(new_n294), .ZN(new_n295));
  AOI21_X1  g094(.A(new_n246), .B1(new_n290), .B2(new_n295), .ZN(new_n296));
  INV_X1    g095(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n290), .A2(new_n246), .A3(new_n295), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  XOR2_X1   g098(.A(G134gat), .B(G162gat), .Z(new_n300));
  XNOR2_X1  g099(.A(new_n300), .B(KEYINPUT98), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n294), .A2(KEYINPUT41), .ZN(new_n302));
  XOR2_X1   g101(.A(new_n301), .B(new_n302), .Z(new_n303));
  INV_X1    g102(.A(KEYINPUT101), .ZN(new_n304));
  OAI21_X1  g103(.A(new_n303), .B1(new_n296), .B2(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n299), .A2(new_n305), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n297), .A2(new_n304), .A3(new_n298), .A4(new_n303), .ZN(new_n307));
  AND2_X1   g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n244), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT10), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n209), .A2(new_n210), .ZN(new_n311));
  AOI21_X1  g110(.A(new_n311), .B1(new_n285), .B2(new_n284), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n282), .A2(new_n283), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  INV_X1    g113(.A(new_n314), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n310), .B1(new_n312), .B2(new_n315), .ZN(new_n316));
  NAND3_X1  g115(.A1(new_n286), .A2(KEYINPUT10), .A3(new_n311), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT102), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n318), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G230gat), .A2(G233gat), .ZN(new_n321));
  NAND3_X1  g120(.A1(new_n316), .A2(KEYINPUT102), .A3(new_n317), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n320), .A2(new_n321), .A3(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n312), .A2(new_n315), .ZN(new_n324));
  INV_X1    g123(.A(new_n321), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(new_n326), .ZN(new_n327));
  XNOR2_X1  g126(.A(G120gat), .B(G148gat), .ZN(new_n328));
  XNOR2_X1  g127(.A(G176gat), .B(G204gat), .ZN(new_n329));
  XOR2_X1   g128(.A(new_n328), .B(new_n329), .Z(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NOR2_X1   g130(.A1(new_n327), .A2(new_n331), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n323), .A2(new_n332), .ZN(new_n333));
  XOR2_X1   g132(.A(new_n321), .B(KEYINPUT103), .Z(new_n334));
  AOI21_X1  g133(.A(new_n334), .B1(new_n316), .B2(new_n317), .ZN(new_n335));
  OAI21_X1  g134(.A(new_n331), .B1(new_n335), .B2(new_n327), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n333), .A2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n309), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G113gat), .B(G120gat), .ZN(new_n340));
  NOR2_X1   g139(.A1(new_n216), .A2(G134gat), .ZN(new_n341));
  INV_X1    g140(.A(G134gat), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n342), .A2(G127gat), .ZN(new_n343));
  OAI22_X1  g142(.A1(new_n340), .A2(KEYINPUT1), .B1(new_n341), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(G120gat), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n345), .A2(G113gat), .ZN(new_n346));
  INV_X1    g145(.A(G113gat), .ZN(new_n347));
  NAND2_X1  g146(.A1(new_n347), .A2(G120gat), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n346), .A2(new_n348), .ZN(new_n349));
  XNOR2_X1  g148(.A(G127gat), .B(G134gat), .ZN(new_n350));
  INV_X1    g149(.A(KEYINPUT1), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n349), .A2(new_n350), .A3(new_n351), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n344), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  INV_X1    g153(.A(G169gat), .ZN(new_n355));
  INV_X1    g154(.A(G176gat), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n355), .A2(new_n356), .A3(KEYINPUT26), .ZN(new_n357));
  NAND2_X1  g156(.A1(G169gat), .A2(G176gat), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT26), .ZN(new_n359));
  NAND2_X1  g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NOR2_X1   g159(.A1(G169gat), .A2(G176gat), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n354), .B(new_n357), .C1(new_n360), .C2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  AND2_X1   g162(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n365));
  NOR2_X1   g164(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  XNOR2_X1  g165(.A(KEYINPUT27), .B(G183gat), .ZN(new_n367));
  AND3_X1   g166(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT28), .ZN(new_n368));
  AOI21_X1  g167(.A(KEYINPUT28), .B1(new_n366), .B2(new_n367), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n363), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT68), .ZN(new_n371));
  OR2_X1    g170(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n372));
  INV_X1    g171(.A(G183gat), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n373), .A2(KEYINPUT27), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT27), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(G183gat), .ZN(new_n376));
  NAND2_X1  g175(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n372), .A2(new_n374), .A3(new_n376), .A4(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT28), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n366), .A2(new_n367), .A3(KEYINPUT28), .ZN(new_n381));
  AOI21_X1  g180(.A(new_n362), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  INV_X1    g181(.A(KEYINPUT68), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n371), .A2(new_n384), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n361), .A2(KEYINPUT23), .ZN(new_n386));
  INV_X1    g185(.A(KEYINPUT23), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n387), .B1(G169gat), .B2(G176gat), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n386), .A2(KEYINPUT25), .A3(new_n388), .A4(new_n358), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  NAND2_X1  g189(.A1(new_n354), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g190(.A1(KEYINPUT64), .A2(G183gat), .A3(G190gat), .ZN(new_n392));
  INV_X1    g191(.A(KEYINPUT24), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n393), .A2(KEYINPUT65), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT65), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(KEYINPUT24), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n391), .A2(new_n392), .A3(new_n394), .A4(new_n396), .ZN(new_n397));
  NAND3_X1  g196(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n398));
  NAND3_X1  g197(.A1(new_n372), .A2(new_n373), .A3(new_n377), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n397), .A2(new_n398), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g199(.A(new_n389), .B1(new_n400), .B2(KEYINPUT67), .ZN(new_n401));
  INV_X1    g200(.A(KEYINPUT67), .ZN(new_n402));
  NAND4_X1  g201(.A1(new_n397), .A2(new_n402), .A3(new_n398), .A4(new_n399), .ZN(new_n403));
  INV_X1    g202(.A(KEYINPUT25), .ZN(new_n404));
  OAI21_X1  g203(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(new_n354), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n406), .A2(new_n398), .ZN(new_n407));
  NAND4_X1  g206(.A1(new_n407), .A2(new_n386), .A3(new_n358), .A4(new_n388), .ZN(new_n408));
  AOI22_X1  g207(.A1(new_n401), .A2(new_n403), .B1(new_n404), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n353), .B1(new_n385), .B2(new_n409), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n380), .A2(new_n381), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n383), .B1(new_n411), .B2(new_n363), .ZN(new_n412));
  AOI211_X1 g211(.A(KEYINPUT68), .B(new_n362), .C1(new_n380), .C2(new_n381), .ZN(new_n413));
  NOR2_X1   g212(.A1(new_n412), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n400), .A2(KEYINPUT67), .ZN(new_n415));
  INV_X1    g214(.A(new_n389), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n415), .A2(new_n403), .A3(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n408), .A2(new_n404), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  AND2_X1   g218(.A1(new_n344), .A2(new_n352), .ZN(new_n420));
  NAND3_X1  g219(.A1(new_n414), .A2(new_n419), .A3(new_n420), .ZN(new_n421));
  NAND2_X1  g220(.A1(G227gat), .A2(G233gat), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n410), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  XNOR2_X1  g222(.A(new_n423), .B(KEYINPUT34), .ZN(new_n424));
  XNOR2_X1  g223(.A(KEYINPUT69), .B(G71gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(G99gat), .ZN(new_n426));
  XNOR2_X1  g225(.A(G15gat), .B(G43gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  AOI21_X1  g227(.A(new_n422), .B1(new_n410), .B2(new_n421), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(new_n429), .B2(KEYINPUT33), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT32), .ZN(new_n431));
  NOR2_X1   g230(.A1(new_n429), .A2(new_n431), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n410), .A2(new_n421), .ZN(new_n434));
  INV_X1    g233(.A(new_n422), .ZN(new_n435));
  AOI221_X4 g234(.A(new_n431), .B1(KEYINPUT33), .B2(new_n428), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  OAI21_X1  g235(.A(new_n424), .B1(new_n433), .B2(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT70), .ZN(new_n438));
  NOR3_X1   g237(.A1(new_n385), .A2(new_n409), .A3(new_n353), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n420), .B1(new_n414), .B2(new_n419), .ZN(new_n440));
  OAI21_X1  g239(.A(new_n435), .B1(new_n439), .B2(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n441), .A2(KEYINPUT32), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT33), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n442), .A2(new_n444), .A3(new_n428), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT34), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n423), .B(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n445), .A2(new_n447), .A3(new_n448), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n437), .A2(new_n438), .A3(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n448), .ZN(new_n451));
  NAND3_X1  g250(.A1(new_n451), .A2(KEYINPUT70), .A3(new_n424), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(G155gat), .A2(G162gat), .ZN(new_n454));
  INV_X1    g253(.A(G162gat), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n234), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g255(.A(G141gat), .B(G148gat), .ZN(new_n457));
  OAI211_X1 g256(.A(new_n454), .B(new_n456), .C1(new_n457), .C2(KEYINPUT2), .ZN(new_n458));
  INV_X1    g257(.A(G141gat), .ZN(new_n459));
  NAND2_X1  g258(.A1(new_n459), .A2(G148gat), .ZN(new_n460));
  INV_X1    g259(.A(G148gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n461), .A2(G141gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n456), .A2(new_n454), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n454), .A2(KEYINPUT2), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n458), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(KEYINPUT3), .ZN(new_n468));
  XOR2_X1   g267(.A(KEYINPUT77), .B(KEYINPUT3), .Z(new_n469));
  NAND3_X1  g268(.A1(new_n458), .A2(new_n466), .A3(new_n469), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n353), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(G225gat), .A2(G233gat), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT4), .ZN(new_n473));
  AND2_X1   g272(.A1(new_n458), .A2(new_n466), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n473), .B1(new_n474), .B2(new_n420), .ZN(new_n475));
  NOR3_X1   g274(.A1(new_n467), .A2(new_n353), .A3(KEYINPUT4), .ZN(new_n476));
  OAI211_X1 g275(.A(new_n471), .B(new_n472), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  INV_X1    g276(.A(new_n472), .ZN(new_n478));
  NOR2_X1   g277(.A1(new_n467), .A2(new_n353), .ZN(new_n479));
  AOI22_X1  g278(.A1(new_n458), .A2(new_n466), .B1(new_n344), .B2(new_n352), .ZN(new_n480));
  OAI21_X1  g279(.A(new_n478), .B1(new_n479), .B2(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(KEYINPUT78), .ZN(new_n482));
  NAND2_X1  g281(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  OAI211_X1 g282(.A(KEYINPUT78), .B(new_n478), .C1(new_n479), .C2(new_n480), .ZN(new_n484));
  NAND4_X1  g283(.A1(new_n477), .A2(new_n483), .A3(KEYINPUT5), .A4(new_n484), .ZN(new_n485));
  XOR2_X1   g284(.A(G1gat), .B(G29gat), .Z(new_n486));
  XNOR2_X1  g285(.A(new_n486), .B(KEYINPUT0), .ZN(new_n487));
  XNOR2_X1  g286(.A(G57gat), .B(G85gat), .ZN(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n479), .A2(new_n473), .ZN(new_n490));
  OAI21_X1  g289(.A(KEYINPUT4), .B1(new_n467), .B2(new_n353), .ZN(new_n491));
  NAND3_X1  g290(.A1(new_n490), .A2(KEYINPUT79), .A3(new_n491), .ZN(new_n492));
  OR2_X1    g291(.A1(new_n491), .A2(KEYINPUT79), .ZN(new_n493));
  NOR2_X1   g292(.A1(new_n478), .A2(KEYINPUT5), .ZN(new_n494));
  NAND4_X1  g293(.A1(new_n492), .A2(new_n493), .A3(new_n471), .A4(new_n494), .ZN(new_n495));
  NAND3_X1  g294(.A1(new_n485), .A2(new_n489), .A3(new_n495), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT80), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n496), .A2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n485), .A2(new_n495), .ZN(new_n499));
  INV_X1    g298(.A(new_n489), .ZN(new_n500));
  NAND2_X1  g299(.A1(new_n499), .A2(new_n500), .ZN(new_n501));
  INV_X1    g300(.A(KEYINPUT6), .ZN(new_n502));
  NAND4_X1  g301(.A1(new_n485), .A2(KEYINPUT80), .A3(new_n489), .A4(new_n495), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n498), .A2(new_n501), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n499), .A2(KEYINPUT6), .A3(new_n500), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(KEYINPUT75), .B(KEYINPUT29), .Z(new_n507));
  NAND2_X1  g306(.A1(G226gat), .A2(G233gat), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n414), .B2(new_n419), .ZN(new_n510));
  NOR3_X1   g309(.A1(new_n409), .A2(new_n382), .A3(new_n508), .ZN(new_n511));
  XNOR2_X1  g310(.A(KEYINPUT72), .B(KEYINPUT22), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT73), .B(G218gat), .ZN(new_n513));
  INV_X1    g312(.A(G211gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n512), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  XNOR2_X1  g314(.A(G197gat), .B(G204gat), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(G211gat), .B(G218gat), .ZN(new_n518));
  INV_X1    g317(.A(new_n518), .ZN(new_n519));
  AND2_X1   g318(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n517), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n519), .A2(KEYINPUT74), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n522), .A2(new_n515), .A3(new_n516), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NOR3_X1   g323(.A1(new_n510), .A2(new_n511), .A3(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT29), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n527), .B(new_n508), .C1(new_n409), .C2(new_n382), .ZN(new_n528));
  INV_X1    g327(.A(new_n508), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n414), .A2(new_n419), .A3(new_n529), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n526), .B1(new_n528), .B2(new_n530), .ZN(new_n531));
  XOR2_X1   g330(.A(G64gat), .B(G92gat), .Z(new_n532));
  XNOR2_X1  g331(.A(G8gat), .B(G36gat), .ZN(new_n533));
  XNOR2_X1  g332(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(new_n534), .ZN(new_n535));
  NOR3_X1   g334(.A1(new_n525), .A2(new_n531), .A3(new_n535), .ZN(new_n536));
  XNOR2_X1  g335(.A(new_n534), .B(KEYINPUT76), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n528), .A2(new_n530), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n538), .A2(new_n524), .ZN(new_n539));
  NAND3_X1  g338(.A1(new_n419), .A2(new_n370), .A3(new_n529), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n385), .A2(new_n409), .ZN(new_n541));
  OAI211_X1 g340(.A(new_n526), .B(new_n540), .C1(new_n541), .C2(new_n509), .ZN(new_n542));
  AOI21_X1  g341(.A(new_n537), .B1(new_n539), .B2(new_n542), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT30), .B1(new_n536), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n539), .A2(new_n534), .A3(new_n542), .ZN(new_n545));
  INV_X1    g344(.A(KEYINPUT30), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n545), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n544), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n506), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G78gat), .B(G106gat), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n550), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(G228gat), .A2(G233gat), .ZN(new_n553));
  INV_X1    g352(.A(KEYINPUT81), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n470), .A2(new_n507), .ZN(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  OAI21_X1  g355(.A(new_n554), .B1(new_n556), .B2(new_n524), .ZN(new_n557));
  NAND4_X1  g356(.A1(new_n555), .A2(KEYINPUT81), .A3(new_n523), .A4(new_n521), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n517), .A2(new_n518), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n515), .A2(new_n519), .A3(new_n516), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n560), .A2(new_n507), .A3(new_n561), .ZN(new_n562));
  AOI21_X1  g361(.A(new_n474), .B1(new_n562), .B2(new_n469), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n553), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  OAI21_X1  g363(.A(KEYINPUT83), .B1(new_n556), .B2(new_n524), .ZN(new_n565));
  INV_X1    g364(.A(KEYINPUT83), .ZN(new_n566));
  NAND4_X1  g365(.A1(new_n555), .A2(new_n566), .A3(new_n523), .A4(new_n521), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n467), .A2(new_n527), .ZN(new_n569));
  AOI21_X1  g368(.A(new_n569), .B1(new_n523), .B2(new_n521), .ZN(new_n570));
  INV_X1    g369(.A(new_n468), .ZN(new_n571));
  OAI21_X1  g370(.A(KEYINPUT82), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n553), .ZN(new_n573));
  INV_X1    g372(.A(KEYINPUT82), .ZN(new_n574));
  OAI211_X1 g373(.A(new_n574), .B(new_n468), .C1(new_n526), .C2(new_n569), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n568), .A2(new_n572), .A3(new_n573), .A4(new_n575), .ZN(new_n576));
  XOR2_X1   g375(.A(KEYINPUT31), .B(G50gat), .Z(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AND3_X1   g377(.A1(new_n564), .A2(new_n576), .A3(new_n578), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n578), .B1(new_n564), .B2(new_n576), .ZN(new_n580));
  OAI21_X1  g379(.A(new_n552), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n564), .A2(new_n576), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(new_n577), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n564), .A2(new_n576), .A3(new_n578), .ZN(new_n584));
  NAND3_X1  g383(.A1(new_n583), .A2(new_n551), .A3(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n581), .A2(new_n585), .ZN(new_n586));
  INV_X1    g385(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n453), .A2(new_n549), .A3(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT71), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n437), .A2(new_n589), .A3(new_n449), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n451), .A2(KEYINPUT71), .A3(new_n424), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n505), .ZN(new_n593));
  AND3_X1   g392(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n594));
  INV_X1    g393(.A(KEYINPUT85), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n489), .B1(new_n499), .B2(new_n595), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n596), .B1(new_n595), .B2(new_n499), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n593), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT35), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n581), .A2(new_n585), .A3(new_n599), .ZN(new_n600));
  NOR3_X1   g399(.A1(new_n598), .A2(new_n600), .A3(new_n548), .ZN(new_n601));
  AOI22_X1  g400(.A1(new_n588), .A2(KEYINPUT35), .B1(new_n592), .B2(new_n601), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT87), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n525), .A2(new_n531), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT37), .ZN(new_n605));
  OAI21_X1  g404(.A(new_n535), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n539), .A2(new_n605), .A3(new_n542), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n607), .A2(KEYINPUT86), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT86), .ZN(new_n609));
  NAND4_X1  g408(.A1(new_n539), .A2(new_n609), .A3(new_n605), .A4(new_n542), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n606), .B1(new_n608), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT38), .ZN(new_n612));
  OAI21_X1  g411(.A(new_n603), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n608), .A2(new_n610), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n539), .A2(new_n542), .ZN(new_n615));
  AOI21_X1  g414(.A(new_n534), .B1(new_n615), .B2(KEYINPUT37), .ZN(new_n616));
  AOI21_X1  g415(.A(new_n612), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n617), .A2(KEYINPUT87), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n510), .A2(new_n511), .ZN(new_n619));
  AOI21_X1  g418(.A(new_n605), .B1(new_n619), .B2(new_n524), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n538), .A2(new_n526), .ZN(new_n621));
  AOI211_X1 g420(.A(KEYINPUT38), .B(new_n537), .C1(new_n620), .C2(new_n621), .ZN(new_n622));
  AOI21_X1  g421(.A(new_n536), .B1(new_n614), .B2(new_n622), .ZN(new_n623));
  NAND4_X1  g422(.A1(new_n613), .A2(new_n618), .A3(new_n598), .A4(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT40), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n492), .A2(new_n493), .A3(new_n471), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n626), .A2(new_n478), .ZN(new_n627));
  INV_X1    g426(.A(new_n479), .ZN(new_n628));
  INV_X1    g427(.A(new_n480), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n472), .A3(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(KEYINPUT84), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n630), .A2(new_n631), .ZN(new_n633));
  NAND4_X1  g432(.A1(new_n627), .A2(KEYINPUT39), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g434(.A(new_n489), .B1(new_n627), .B2(KEYINPUT39), .ZN(new_n636));
  OAI21_X1  g435(.A(new_n625), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  OR2_X1    g436(.A1(new_n627), .A2(KEYINPUT39), .ZN(new_n638));
  NAND4_X1  g437(.A1(new_n638), .A2(new_n634), .A3(KEYINPUT40), .A4(new_n489), .ZN(new_n639));
  AND3_X1   g438(.A1(new_n637), .A2(new_n639), .A3(new_n597), .ZN(new_n640));
  AOI21_X1  g439(.A(new_n586), .B1(new_n640), .B2(new_n548), .ZN(new_n641));
  NAND2_X1  g440(.A1(new_n453), .A2(KEYINPUT36), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT36), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n590), .A2(new_n591), .A3(new_n643), .ZN(new_n644));
  AOI22_X1  g443(.A1(new_n624), .A2(new_n641), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n537), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(new_n525), .B2(new_n531), .ZN(new_n647));
  AOI21_X1  g446(.A(new_n546), .B1(new_n647), .B2(new_n545), .ZN(new_n648));
  AOI21_X1  g447(.A(KEYINPUT30), .B1(new_n604), .B2(new_n534), .ZN(new_n649));
  NOR2_X1   g448(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n504), .A2(new_n505), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n652), .A2(new_n586), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n602), .B1(new_n645), .B2(new_n653), .ZN(new_n654));
  OR2_X1    g453(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n225), .A2(KEYINPUT90), .ZN(new_n656));
  NAND4_X1  g455(.A1(new_n655), .A2(new_n269), .A3(new_n272), .A4(new_n656), .ZN(new_n657));
  OAI21_X1  g456(.A(new_n291), .B1(new_n227), .B2(new_n229), .ZN(new_n658));
  NAND2_X1  g457(.A1(G229gat), .A2(G233gat), .ZN(new_n659));
  XNOR2_X1  g458(.A(new_n659), .B(KEYINPUT91), .ZN(new_n660));
  NAND3_X1  g459(.A1(new_n657), .A2(new_n658), .A3(new_n660), .ZN(new_n661));
  INV_X1    g460(.A(KEYINPUT93), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  INV_X1    g462(.A(KEYINPUT18), .ZN(new_n664));
  NAND4_X1  g463(.A1(new_n657), .A2(KEYINPUT93), .A3(new_n658), .A4(new_n660), .ZN(new_n665));
  NAND3_X1  g464(.A1(new_n663), .A2(new_n664), .A3(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT94), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  NAND4_X1  g467(.A1(new_n663), .A2(KEYINPUT94), .A3(new_n664), .A4(new_n665), .ZN(new_n669));
  XOR2_X1   g468(.A(new_n660), .B(KEYINPUT13), .Z(new_n670));
  NAND2_X1  g469(.A1(new_n228), .A2(new_n230), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n671), .A2(new_n291), .ZN(new_n672));
  INV_X1    g471(.A(new_n658), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n670), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND4_X1  g473(.A1(new_n657), .A2(KEYINPUT18), .A3(new_n658), .A4(new_n660), .ZN(new_n675));
  XNOR2_X1  g474(.A(G113gat), .B(G141gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n676), .B(G197gat), .ZN(new_n677));
  XOR2_X1   g476(.A(KEYINPUT11), .B(G169gat), .Z(new_n678));
  XNOR2_X1  g477(.A(new_n677), .B(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n679), .B(KEYINPUT12), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n674), .A2(new_n675), .A3(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n668), .A2(new_n669), .A3(new_n681), .ZN(new_n682));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n674), .A3(new_n675), .ZN(new_n683));
  INV_X1    g482(.A(new_n680), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  INV_X1    g485(.A(new_n686), .ZN(new_n687));
  OAI21_X1  g486(.A(KEYINPUT95), .B1(new_n654), .B2(new_n687), .ZN(new_n688));
  OAI211_X1 g487(.A(new_n623), .B(new_n598), .C1(new_n617), .C2(KEYINPUT87), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n611), .A2(new_n603), .A3(new_n612), .ZN(new_n690));
  OAI21_X1  g489(.A(new_n641), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n642), .A2(new_n644), .ZN(new_n692));
  NAND3_X1  g491(.A1(new_n691), .A2(new_n692), .A3(new_n653), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n588), .A2(KEYINPUT35), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n601), .A2(new_n592), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(new_n696), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT95), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n697), .A2(new_n698), .A3(new_n686), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n339), .B1(new_n688), .B2(new_n699), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n506), .ZN(new_n701));
  XOR2_X1   g500(.A(KEYINPUT104), .B(G1gat), .Z(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1324gat));
  INV_X1    g502(.A(G8gat), .ZN(new_n704));
  AOI21_X1  g503(.A(new_n704), .B1(new_n700), .B2(new_n548), .ZN(new_n705));
  INV_X1    g504(.A(new_n339), .ZN(new_n706));
  AOI21_X1  g505(.A(new_n698), .B1(new_n697), .B2(new_n686), .ZN(new_n707));
  AOI211_X1 g506(.A(KEYINPUT95), .B(new_n687), .C1(new_n693), .C2(new_n696), .ZN(new_n708));
  OAI211_X1 g507(.A(new_n548), .B(new_n706), .C1(new_n707), .C2(new_n708), .ZN(new_n709));
  XNOR2_X1  g508(.A(KEYINPUT16), .B(G8gat), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  OAI21_X1  g510(.A(KEYINPUT42), .B1(new_n705), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT105), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n688), .A2(new_n699), .ZN(new_n714));
  INV_X1    g513(.A(new_n710), .ZN(new_n715));
  NAND4_X1  g514(.A1(new_n714), .A2(new_n548), .A3(new_n706), .A4(new_n715), .ZN(new_n716));
  INV_X1    g515(.A(KEYINPUT42), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND3_X1  g517(.A1(new_n712), .A2(new_n713), .A3(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n709), .A2(G8gat), .ZN(new_n720));
  AOI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(new_n716), .ZN(new_n721));
  AND2_X1   g520(.A1(new_n716), .A2(new_n717), .ZN(new_n722));
  OAI21_X1  g521(.A(KEYINPUT105), .B1(new_n721), .B2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n719), .A2(new_n723), .ZN(G1325gat));
  INV_X1    g523(.A(new_n700), .ZN(new_n725));
  OR2_X1    g524(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n692), .A2(KEYINPUT106), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(new_n728), .ZN(new_n729));
  OAI21_X1  g528(.A(G15gat), .B1(new_n725), .B2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n592), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n731), .A2(G15gat), .ZN(new_n732));
  OAI21_X1  g531(.A(new_n730), .B1(new_n725), .B2(new_n732), .ZN(G1326gat));
  OAI21_X1  g532(.A(KEYINPUT107), .B1(new_n725), .B2(new_n587), .ZN(new_n734));
  INV_X1    g533(.A(KEYINPUT107), .ZN(new_n735));
  NAND3_X1  g534(.A1(new_n700), .A2(new_n735), .A3(new_n586), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n734), .A2(new_n736), .ZN(new_n737));
  XNOR2_X1  g536(.A(KEYINPUT43), .B(G22gat), .ZN(new_n738));
  INV_X1    g537(.A(new_n738), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  NAND3_X1  g539(.A1(new_n734), .A2(new_n736), .A3(new_n738), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n740), .A2(new_n741), .ZN(G1327gat));
  NOR2_X1   g541(.A1(new_n243), .A2(new_n337), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  INV_X1    g543(.A(new_n308), .ZN(new_n745));
  NOR2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n714), .A2(new_n746), .ZN(new_n747));
  INV_X1    g546(.A(KEYINPUT45), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n506), .A2(new_n255), .ZN(new_n749));
  OR3_X1    g548(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT108), .ZN(new_n751));
  AOI221_X4 g550(.A(new_n751), .B1(new_n581), .B2(new_n585), .C1(new_n650), .C2(new_n651), .ZN(new_n752));
  AOI21_X1  g551(.A(KEYINPUT108), .B1(new_n652), .B2(new_n586), .ZN(new_n753));
  NOR2_X1   g552(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND3_X1  g553(.A1(new_n754), .A2(new_n691), .A3(new_n692), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n755), .A2(new_n696), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n756), .A2(KEYINPUT109), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT109), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n755), .A2(new_n758), .A3(new_n696), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n745), .A2(KEYINPUT44), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n757), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT44), .ZN(new_n762));
  AOI21_X1  g561(.A(new_n762), .B1(new_n697), .B2(new_n308), .ZN(new_n763));
  INV_X1    g562(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n761), .A2(new_n764), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n744), .A2(new_n687), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(G29gat), .B1(new_n767), .B2(new_n651), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n748), .B1(new_n747), .B2(new_n749), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n750), .A2(new_n768), .A3(new_n769), .ZN(G1328gat));
  NAND4_X1  g569(.A1(new_n714), .A2(new_n256), .A3(new_n548), .A4(new_n746), .ZN(new_n771));
  XOR2_X1   g570(.A(new_n771), .B(KEYINPUT46), .Z(new_n772));
  INV_X1    g571(.A(KEYINPUT110), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n767), .B2(new_n650), .ZN(new_n774));
  INV_X1    g573(.A(new_n766), .ZN(new_n775));
  AOI21_X1  g574(.A(new_n775), .B1(new_n761), .B2(new_n764), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(KEYINPUT110), .A3(new_n548), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n774), .A2(G36gat), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n772), .A2(new_n778), .ZN(G1329gat));
  OAI21_X1  g578(.A(G43gat), .B1(new_n767), .B2(new_n692), .ZN(new_n780));
  INV_X1    g579(.A(G43gat), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n592), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n747), .A2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(new_n783), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n780), .A2(new_n784), .A3(KEYINPUT47), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n781), .B1(new_n776), .B2(new_n728), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n783), .ZN(new_n787));
  OAI21_X1  g586(.A(new_n785), .B1(KEYINPUT47), .B2(new_n787), .ZN(G1330gat));
  INV_X1    g587(.A(KEYINPUT48), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n249), .B1(new_n776), .B2(new_n586), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n586), .A2(new_n249), .ZN(new_n791));
  XOR2_X1   g590(.A(new_n791), .B(KEYINPUT111), .Z(new_n792));
  NOR2_X1   g591(.A1(new_n747), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n789), .B1(new_n790), .B2(new_n793), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n755), .A2(new_n758), .A3(new_n696), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n758), .B1(new_n755), .B2(new_n696), .ZN(new_n796));
  INV_X1    g595(.A(new_n760), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n795), .A2(new_n796), .A3(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n586), .B(new_n766), .C1(new_n798), .C2(new_n763), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT112), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT112), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n776), .A2(new_n801), .A3(new_n586), .ZN(new_n802));
  AND3_X1   g601(.A1(new_n800), .A2(G50gat), .A3(new_n802), .ZN(new_n803));
  OAI21_X1  g602(.A(KEYINPUT48), .B1(new_n747), .B2(new_n792), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n794), .B1(new_n803), .B2(new_n804), .ZN(G1331gat));
  NOR2_X1   g604(.A1(new_n795), .A2(new_n796), .ZN(new_n806));
  NOR2_X1   g605(.A1(new_n686), .A2(new_n338), .ZN(new_n807));
  AND2_X1   g606(.A1(new_n309), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g607(.A1(new_n806), .A2(new_n808), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  NAND2_X1  g609(.A1(new_n810), .A2(new_n506), .ZN(new_n811));
  XNOR2_X1  g610(.A(new_n811), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g611(.A1(new_n809), .A2(new_n650), .ZN(new_n813));
  NOR2_X1   g612(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n814));
  AND2_X1   g613(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n815));
  OAI21_X1  g614(.A(new_n813), .B1(new_n814), .B2(new_n815), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n816), .B1(new_n813), .B2(new_n814), .ZN(G1333gat));
  OR3_X1    g616(.A1(new_n809), .A2(G71gat), .A3(new_n731), .ZN(new_n818));
  OAI21_X1  g617(.A(G71gat), .B1(new_n809), .B2(new_n729), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT50), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n818), .A2(new_n819), .A3(KEYINPUT50), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(G1334gat));
  NAND2_X1  g623(.A1(new_n810), .A2(new_n586), .ZN(new_n825));
  XNOR2_X1  g624(.A(new_n825), .B(G78gat), .ZN(G1335gat));
  NAND2_X1  g625(.A1(new_n807), .A2(new_n244), .ZN(new_n827));
  XOR2_X1   g626(.A(new_n827), .B(KEYINPUT113), .Z(new_n828));
  INV_X1    g627(.A(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n829), .B1(new_n761), .B2(new_n764), .ZN(new_n830));
  INV_X1    g629(.A(new_n830), .ZN(new_n831));
  OAI21_X1  g630(.A(G85gat), .B1(new_n831), .B2(new_n651), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n686), .A2(new_n745), .A3(new_n243), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n756), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g633(.A(new_n834), .B(KEYINPUT51), .ZN(new_n835));
  NAND3_X1  g634(.A1(new_n506), .A2(new_n274), .A3(new_n337), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n832), .B1(new_n835), .B2(new_n836), .ZN(G1336gat));
  AOI21_X1  g636(.A(new_n275), .B1(new_n830), .B2(new_n548), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n337), .A2(new_n548), .A3(new_n275), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n835), .A2(new_n839), .ZN(new_n840));
  OR3_X1    g639(.A1(new_n838), .A2(KEYINPUT52), .A3(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(KEYINPUT52), .B1(new_n838), .B2(new_n840), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(new_n842), .ZN(G1337gat));
  OAI21_X1  g642(.A(G99gat), .B1(new_n831), .B2(new_n729), .ZN(new_n844));
  OR3_X1    g643(.A1(new_n731), .A2(G99gat), .A3(new_n338), .ZN(new_n845));
  OAI21_X1  g644(.A(new_n844), .B1(new_n835), .B2(new_n845), .ZN(G1338gat));
  INV_X1    g645(.A(G106gat), .ZN(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n830), .B2(new_n586), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT51), .ZN(new_n849));
  XNOR2_X1  g648(.A(new_n834), .B(new_n849), .ZN(new_n850));
  NOR3_X1   g649(.A1(new_n338), .A2(new_n587), .A3(G106gat), .ZN(new_n851));
  AND2_X1   g650(.A1(new_n850), .A2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(KEYINPUT53), .B1(new_n848), .B2(new_n852), .ZN(new_n853));
  OAI211_X1 g652(.A(new_n586), .B(new_n828), .C1(new_n798), .C2(new_n763), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(G106gat), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT115), .ZN(new_n856));
  XOR2_X1   g655(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n857));
  AOI21_X1  g656(.A(new_n857), .B1(new_n850), .B2(new_n851), .ZN(new_n858));
  AND3_X1   g657(.A1(new_n855), .A2(new_n856), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g658(.A(new_n856), .B1(new_n855), .B2(new_n858), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n853), .B1(new_n859), .B2(new_n860), .ZN(G1339gat));
  INV_X1    g660(.A(KEYINPUT54), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n316), .A2(new_n317), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n862), .B1(new_n863), .B2(new_n334), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n323), .A2(new_n864), .ZN(new_n865));
  INV_X1    g664(.A(new_n334), .ZN(new_n866));
  NAND3_X1  g665(.A1(new_n318), .A2(new_n862), .A3(new_n866), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n867), .A2(new_n331), .ZN(new_n868));
  INV_X1    g667(.A(new_n868), .ZN(new_n869));
  NAND3_X1  g668(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT55), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n870), .A2(KEYINPUT116), .ZN(new_n871));
  AOI21_X1  g670(.A(new_n868), .B1(new_n323), .B2(new_n864), .ZN(new_n872));
  INV_X1    g671(.A(KEYINPUT116), .ZN(new_n873));
  NAND3_X1  g672(.A1(new_n872), .A2(new_n873), .A3(KEYINPUT55), .ZN(new_n874));
  NAND2_X1  g673(.A1(new_n871), .A2(new_n874), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n865), .A2(new_n869), .ZN(new_n876));
  INV_X1    g675(.A(KEYINPUT55), .ZN(new_n877));
  AOI22_X1  g676(.A1(new_n876), .A2(new_n877), .B1(new_n323), .B2(new_n332), .ZN(new_n878));
  NAND3_X1  g677(.A1(new_n875), .A2(new_n686), .A3(new_n878), .ZN(new_n879));
  OR2_X1    g678(.A1(new_n672), .A2(new_n673), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT117), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n660), .B1(new_n657), .B2(new_n658), .ZN(new_n882));
  OAI22_X1  g681(.A1(new_n880), .A2(new_n670), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  AND2_X1   g682(.A1(new_n882), .A2(new_n881), .ZN(new_n884));
  OAI21_X1  g683(.A(new_n679), .B1(new_n883), .B2(new_n884), .ZN(new_n885));
  NAND3_X1  g684(.A1(new_n682), .A2(new_n885), .A3(new_n337), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n308), .B1(new_n879), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n873), .B1(new_n872), .B2(KEYINPUT55), .ZN(new_n888));
  AND4_X1   g687(.A1(new_n873), .A2(new_n865), .A3(KEYINPUT55), .A4(new_n869), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n878), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n682), .A2(new_n885), .A3(new_n308), .ZN(new_n891));
  NOR2_X1   g690(.A1(new_n890), .A2(new_n891), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n244), .B1(new_n887), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n706), .A2(new_n687), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n651), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n453), .A2(new_n587), .ZN(new_n896));
  NOR2_X1   g695(.A1(new_n896), .A2(new_n548), .ZN(new_n897));
  AND2_X1   g696(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(G113gat), .B1(new_n898), .B2(new_n686), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n586), .B1(new_n893), .B2(new_n894), .ZN(new_n900));
  INV_X1    g699(.A(new_n900), .ZN(new_n901));
  NOR2_X1   g700(.A1(new_n548), .A2(new_n651), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n592), .A2(new_n902), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n901), .A2(new_n903), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n687), .A2(new_n347), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n899), .B1(new_n904), .B2(new_n905), .ZN(G1340gat));
  AOI21_X1  g705(.A(G120gat), .B1(new_n898), .B2(new_n337), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n338), .A2(new_n345), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n907), .B1(new_n904), .B2(new_n908), .ZN(G1341gat));
  NAND3_X1  g708(.A1(new_n898), .A2(new_n216), .A3(new_n243), .ZN(new_n910));
  NOR3_X1   g709(.A1(new_n901), .A2(new_n244), .A3(new_n903), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n910), .B1(new_n216), .B2(new_n911), .ZN(G1342gat));
  NAND3_X1  g711(.A1(new_n898), .A2(new_n342), .A3(new_n308), .ZN(new_n913));
  OR2_X1    g712(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(KEYINPUT56), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n901), .A2(new_n745), .A3(new_n903), .ZN(new_n916));
  OAI211_X1 g715(.A(new_n914), .B(new_n915), .C1(new_n342), .C2(new_n916), .ZN(G1343gat));
  INV_X1    g716(.A(KEYINPUT119), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n918), .A2(KEYINPUT58), .ZN(new_n919));
  INV_X1    g718(.A(new_n919), .ZN(new_n920));
  NAND2_X1  g719(.A1(new_n692), .A2(new_n902), .ZN(new_n921));
  INV_X1    g720(.A(new_n921), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n893), .A2(new_n894), .ZN(new_n923));
  AOI21_X1  g722(.A(KEYINPUT57), .B1(new_n923), .B2(new_n586), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT57), .ZN(new_n925));
  AOI211_X1 g724(.A(new_n925), .B(new_n587), .C1(new_n893), .C2(new_n894), .ZN(new_n926));
  OAI211_X1 g725(.A(new_n686), .B(new_n922), .C1(new_n924), .C2(new_n926), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(G141gat), .ZN(new_n928));
  AND4_X1   g727(.A1(new_n650), .A2(new_n726), .A3(new_n586), .A4(new_n727), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n686), .A2(new_n459), .ZN(new_n930));
  XNOR2_X1  g729(.A(new_n930), .B(KEYINPUT118), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n895), .A2(new_n929), .A3(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n918), .A2(KEYINPUT58), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  INV_X1    g733(.A(new_n934), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n920), .B1(new_n928), .B2(new_n935), .ZN(new_n936));
  AOI211_X1 g735(.A(new_n919), .B(new_n934), .C1(new_n927), .C2(G141gat), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n936), .A2(new_n937), .ZN(G1344gat));
  INV_X1    g737(.A(KEYINPUT120), .ZN(new_n939));
  AOI21_X1  g738(.A(new_n338), .B1(new_n921), .B2(new_n939), .ZN(new_n940));
  OAI221_X1 g739(.A(new_n940), .B1(new_n939), .B2(new_n921), .C1(new_n924), .C2(new_n926), .ZN(new_n941));
  AND2_X1   g740(.A1(KEYINPUT59), .A2(G148gat), .ZN(new_n942));
  AND2_X1   g741(.A1(new_n895), .A2(new_n929), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n338), .A2(G148gat), .ZN(new_n944));
  AOI22_X1  g743(.A1(new_n941), .A2(new_n942), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  INV_X1    g744(.A(new_n924), .ZN(new_n946));
  INV_X1    g745(.A(new_n926), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n921), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g747(.A(new_n461), .B1(new_n948), .B2(new_n337), .ZN(new_n949));
  OAI21_X1  g748(.A(new_n945), .B1(new_n949), .B2(KEYINPUT59), .ZN(G1345gat));
  NAND2_X1  g749(.A1(new_n943), .A2(new_n243), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT121), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n953), .A2(G155gat), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n951), .A2(new_n952), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n244), .A2(new_n234), .ZN(new_n956));
  AOI22_X1  g755(.A1(new_n954), .A2(new_n955), .B1(new_n948), .B2(new_n956), .ZN(G1346gat));
  AOI21_X1  g756(.A(G162gat), .B1(new_n943), .B2(new_n308), .ZN(new_n958));
  NOR2_X1   g757(.A1(new_n745), .A2(new_n455), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n958), .B1(new_n948), .B2(new_n959), .ZN(G1347gat));
  AOI21_X1  g759(.A(new_n506), .B1(new_n893), .B2(new_n894), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n896), .A2(new_n650), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  INV_X1    g762(.A(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(G169gat), .B1(new_n964), .B2(new_n686), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n506), .A2(new_n650), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  NOR2_X1   g766(.A1(new_n731), .A2(new_n967), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n900), .A2(new_n968), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n687), .A2(new_n355), .ZN(new_n970));
  AOI21_X1  g769(.A(new_n965), .B1(new_n969), .B2(new_n970), .ZN(G1348gat));
  NOR2_X1   g770(.A1(new_n338), .A2(G176gat), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n900), .A2(new_n337), .A3(new_n968), .ZN(new_n973));
  AOI22_X1  g772(.A1(new_n964), .A2(new_n972), .B1(new_n973), .B2(G176gat), .ZN(new_n974));
  XNOR2_X1  g773(.A(new_n974), .B(KEYINPUT122), .ZN(G1349gat));
  NAND4_X1  g774(.A1(new_n923), .A2(new_n587), .A3(new_n243), .A4(new_n968), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT123), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NAND4_X1  g777(.A1(new_n900), .A2(KEYINPUT123), .A3(new_n243), .A4(new_n968), .ZN(new_n979));
  NAND3_X1  g778(.A1(new_n978), .A2(G183gat), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g779(.A1(new_n243), .A2(new_n367), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n980), .B1(new_n963), .B2(new_n981), .ZN(new_n982));
  INV_X1    g781(.A(KEYINPUT124), .ZN(new_n983));
  INV_X1    g782(.A(KEYINPUT60), .ZN(new_n984));
  NOR2_X1   g783(.A1(new_n983), .A2(new_n984), .ZN(new_n985));
  NAND2_X1  g784(.A1(new_n982), .A2(new_n985), .ZN(new_n986));
  OAI221_X1 g785(.A(new_n980), .B1(new_n983), .B2(new_n984), .C1(new_n963), .C2(new_n981), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n986), .A2(new_n987), .ZN(G1350gat));
  NAND3_X1  g787(.A1(new_n964), .A2(new_n366), .A3(new_n308), .ZN(new_n989));
  NAND2_X1  g788(.A1(new_n969), .A2(new_n308), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT61), .ZN(new_n991));
  AND3_X1   g790(.A1(new_n990), .A2(new_n991), .A3(G190gat), .ZN(new_n992));
  AOI21_X1  g791(.A(new_n991), .B1(new_n990), .B2(G190gat), .ZN(new_n993));
  OAI21_X1  g792(.A(new_n989), .B1(new_n992), .B2(new_n993), .ZN(G1351gat));
  NOR3_X1   g793(.A1(new_n728), .A2(new_n650), .A3(new_n587), .ZN(new_n995));
  AND2_X1   g794(.A1(new_n995), .A2(new_n961), .ZN(new_n996));
  XOR2_X1   g795(.A(KEYINPUT125), .B(G197gat), .Z(new_n997));
  NAND3_X1  g796(.A1(new_n996), .A2(new_n686), .A3(new_n997), .ZN(new_n998));
  AND2_X1   g797(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n999));
  NOR2_X1   g798(.A1(new_n998), .A2(KEYINPUT126), .ZN(new_n1000));
  NOR2_X1   g799(.A1(new_n728), .A2(new_n967), .ZN(new_n1001));
  OAI21_X1  g800(.A(new_n1001), .B1(new_n924), .B2(new_n926), .ZN(new_n1002));
  NOR2_X1   g801(.A1(new_n1002), .A2(new_n687), .ZN(new_n1003));
  OAI22_X1  g802(.A1(new_n999), .A2(new_n1000), .B1(new_n1003), .B2(new_n997), .ZN(G1352gat));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n1005));
  AOI21_X1  g804(.A(G204gat), .B1(new_n1005), .B2(KEYINPUT62), .ZN(new_n1006));
  NAND3_X1  g805(.A1(new_n996), .A2(new_n337), .A3(new_n1006), .ZN(new_n1007));
  NOR2_X1   g806(.A1(new_n1005), .A2(KEYINPUT62), .ZN(new_n1008));
  XNOR2_X1  g807(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  OAI21_X1  g808(.A(G204gat), .B1(new_n1002), .B2(new_n338), .ZN(new_n1010));
  NAND2_X1  g809(.A1(new_n1009), .A2(new_n1010), .ZN(G1353gat));
  NAND3_X1  g810(.A1(new_n996), .A2(new_n514), .A3(new_n243), .ZN(new_n1012));
  OAI211_X1 g811(.A(new_n243), .B(new_n1001), .C1(new_n924), .C2(new_n926), .ZN(new_n1013));
  AND3_X1   g812(.A1(new_n1013), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n1014));
  AOI21_X1  g813(.A(KEYINPUT63), .B1(new_n1013), .B2(G211gat), .ZN(new_n1015));
  OAI21_X1  g814(.A(new_n1012), .B1(new_n1014), .B2(new_n1015), .ZN(G1354gat));
  NOR3_X1   g815(.A1(new_n1002), .A2(new_n513), .A3(new_n745), .ZN(new_n1017));
  AOI21_X1  g816(.A(G218gat), .B1(new_n996), .B2(new_n308), .ZN(new_n1018));
  NOR2_X1   g817(.A1(new_n1017), .A2(new_n1018), .ZN(G1355gat));
endmodule


