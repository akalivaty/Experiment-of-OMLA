

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593;

  NAND2_X1 U324 ( .A1(n397), .A2(n396), .ZN(n398) );
  NOR2_X1 U325 ( .A1(n531), .A2(n530), .ZN(n532) );
  XNOR2_X1 U326 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U327 ( .A(n328), .B(n327), .ZN(n392) );
  NOR2_X1 U328 ( .A1(n368), .A2(n583), .ZN(n369) );
  XNOR2_X1 U329 ( .A(KEYINPUT75), .B(G85GAT), .ZN(n308) );
  INV_X1 U330 ( .A(KEYINPUT120), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n312), .B(n311), .ZN(n352) );
  XNOR2_X1 U332 ( .A(n453), .B(n452), .ZN(n454) );
  XOR2_X1 U333 ( .A(KEYINPUT36), .B(n457), .Z(n591) );
  XNOR2_X1 U334 ( .A(n455), .B(n454), .ZN(n456) );
  NOR2_X1 U335 ( .A1(n535), .A2(n534), .ZN(n545) );
  XOR2_X1 U336 ( .A(n413), .B(n412), .Z(n518) );
  XNOR2_X1 U337 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n458) );
  XNOR2_X1 U338 ( .A(n459), .B(n458), .ZN(G1351GAT) );
  XOR2_X1 U339 ( .A(KEYINPUT89), .B(KEYINPUT88), .Z(n293) );
  XNOR2_X1 U340 ( .A(G43GAT), .B(KEYINPUT20), .ZN(n292) );
  XNOR2_X1 U341 ( .A(n293), .B(n292), .ZN(n306) );
  XOR2_X1 U342 ( .A(G15GAT), .B(G127GAT), .Z(n341) );
  XOR2_X1 U343 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n295) );
  XNOR2_X1 U344 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n294) );
  XNOR2_X1 U345 ( .A(n295), .B(n294), .ZN(n403) );
  XOR2_X1 U346 ( .A(n341), .B(n403), .Z(n297) );
  NAND2_X1 U347 ( .A1(G227GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U348 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U349 ( .A(n298), .B(G176GAT), .Z(n301) );
  XNOR2_X1 U350 ( .A(G113GAT), .B(G134GAT), .ZN(n299) );
  XNOR2_X1 U351 ( .A(n299), .B(KEYINPUT0), .ZN(n442) );
  XNOR2_X1 U352 ( .A(n442), .B(G183GAT), .ZN(n300) );
  XNOR2_X1 U353 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U354 ( .A(G120GAT), .B(G71GAT), .Z(n363) );
  XOR2_X1 U355 ( .A(n302), .B(n363), .Z(n304) );
  XNOR2_X1 U356 ( .A(G99GAT), .B(G190GAT), .ZN(n303) );
  XNOR2_X1 U357 ( .A(n304), .B(n303), .ZN(n305) );
  XOR2_X2 U358 ( .A(n306), .B(n305), .Z(n520) );
  INV_X1 U359 ( .A(n520), .ZN(n535) );
  XNOR2_X1 U360 ( .A(G36GAT), .B(G190GAT), .ZN(n307) );
  XNOR2_X1 U361 ( .A(n307), .B(G92GAT), .ZN(n399) );
  INV_X1 U362 ( .A(G99GAT), .ZN(n312) );
  INV_X1 U363 ( .A(n308), .ZN(n310) );
  XNOR2_X1 U364 ( .A(G106GAT), .B(KEYINPUT74), .ZN(n309) );
  XNOR2_X1 U365 ( .A(n310), .B(n309), .ZN(n311) );
  XNOR2_X1 U366 ( .A(n399), .B(n352), .ZN(n314) );
  XOR2_X1 U367 ( .A(KEYINPUT10), .B(KEYINPUT65), .Z(n313) );
  XNOR2_X1 U368 ( .A(n314), .B(n313), .ZN(n328) );
  NAND2_X1 U369 ( .A1(G232GAT), .A2(G233GAT), .ZN(n320) );
  XOR2_X1 U370 ( .A(KEYINPUT11), .B(KEYINPUT82), .Z(n316) );
  XNOR2_X1 U371 ( .A(KEYINPUT66), .B(KEYINPUT9), .ZN(n315) );
  XNOR2_X1 U372 ( .A(n316), .B(n315), .ZN(n318) );
  XOR2_X1 U373 ( .A(G134GAT), .B(KEYINPUT83), .Z(n317) );
  XNOR2_X1 U374 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U375 ( .A(n320), .B(n319), .ZN(n326) );
  XOR2_X1 U376 ( .A(G29GAT), .B(G43GAT), .Z(n322) );
  XNOR2_X1 U377 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n321) );
  XNOR2_X1 U378 ( .A(n322), .B(n321), .ZN(n373) );
  XOR2_X1 U379 ( .A(G162GAT), .B(KEYINPUT81), .Z(n324) );
  XNOR2_X1 U380 ( .A(G50GAT), .B(G218GAT), .ZN(n323) );
  XNOR2_X1 U381 ( .A(n324), .B(n323), .ZN(n430) );
  XNOR2_X1 U382 ( .A(n373), .B(n430), .ZN(n325) );
  INV_X1 U383 ( .A(KEYINPUT84), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n392), .B(n329), .ZN(n457) );
  XOR2_X1 U385 ( .A(KEYINPUT13), .B(G57GAT), .Z(n359) );
  XOR2_X1 U386 ( .A(G8GAT), .B(G183GAT), .Z(n409) );
  XOR2_X1 U387 ( .A(n359), .B(n409), .Z(n331) );
  XOR2_X1 U388 ( .A(KEYINPUT70), .B(G1GAT), .Z(n372) );
  XOR2_X1 U389 ( .A(G22GAT), .B(G155GAT), .Z(n421) );
  XNOR2_X1 U390 ( .A(n372), .B(n421), .ZN(n330) );
  XNOR2_X1 U391 ( .A(n331), .B(n330), .ZN(n345) );
  XOR2_X1 U392 ( .A(KEYINPUT86), .B(KEYINPUT87), .Z(n333) );
  NAND2_X1 U393 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U394 ( .A(n333), .B(n332), .ZN(n337) );
  XOR2_X1 U395 ( .A(KEYINPUT12), .B(KEYINPUT14), .Z(n335) );
  XNOR2_X1 U396 ( .A(KEYINPUT15), .B(KEYINPUT85), .ZN(n334) );
  XNOR2_X1 U397 ( .A(n335), .B(n334), .ZN(n336) );
  XOR2_X1 U398 ( .A(n337), .B(n336), .Z(n343) );
  XOR2_X1 U399 ( .A(G64GAT), .B(G78GAT), .Z(n339) );
  XNOR2_X1 U400 ( .A(G71GAT), .B(G211GAT), .ZN(n338) );
  XNOR2_X1 U401 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U402 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U403 ( .A(n343), .B(n342), .ZN(n344) );
  XOR2_X1 U404 ( .A(n345), .B(n344), .Z(n587) );
  INV_X1 U405 ( .A(n587), .ZN(n486) );
  NOR2_X1 U406 ( .A1(n591), .A2(n486), .ZN(n346) );
  XOR2_X1 U407 ( .A(n346), .B(KEYINPUT45), .Z(n368) );
  XOR2_X1 U408 ( .A(G64GAT), .B(KEYINPUT78), .Z(n348) );
  XNOR2_X1 U409 ( .A(G176GAT), .B(G204GAT), .ZN(n347) );
  XNOR2_X1 U410 ( .A(n348), .B(n347), .ZN(n400) );
  XOR2_X1 U411 ( .A(KEYINPUT76), .B(n400), .Z(n350) );
  NAND2_X1 U412 ( .A1(G230GAT), .A2(G233GAT), .ZN(n349) );
  XNOR2_X1 U413 ( .A(n350), .B(n349), .ZN(n351) );
  XNOR2_X1 U414 ( .A(n352), .B(n351), .ZN(n367) );
  XOR2_X1 U415 ( .A(KEYINPUT31), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U416 ( .A(KEYINPUT71), .B(KEYINPUT80), .ZN(n353) );
  XNOR2_X1 U417 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U418 ( .A(KEYINPUT33), .B(KEYINPUT73), .Z(n356) );
  XNOR2_X1 U419 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n355) );
  XNOR2_X1 U420 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U421 ( .A(n358), .B(n357), .Z(n365) );
  XOR2_X1 U422 ( .A(KEYINPUT72), .B(n359), .Z(n361) );
  XOR2_X1 U423 ( .A(G148GAT), .B(G78GAT), .Z(n418) );
  XNOR2_X1 U424 ( .A(n418), .B(G92GAT), .ZN(n360) );
  XNOR2_X1 U425 ( .A(n361), .B(n360), .ZN(n362) );
  XNOR2_X1 U426 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U427 ( .A(n365), .B(n364), .ZN(n366) );
  XNOR2_X1 U428 ( .A(n367), .B(n366), .ZN(n583) );
  XNOR2_X1 U429 ( .A(n369), .B(KEYINPUT109), .ZN(n387) );
  XOR2_X1 U430 ( .A(G197GAT), .B(G15GAT), .Z(n371) );
  XNOR2_X1 U431 ( .A(G169GAT), .B(G113GAT), .ZN(n370) );
  XNOR2_X1 U432 ( .A(n371), .B(n370), .ZN(n386) );
  XOR2_X1 U433 ( .A(n372), .B(G50GAT), .Z(n375) );
  XNOR2_X1 U434 ( .A(G36GAT), .B(n373), .ZN(n374) );
  XNOR2_X1 U435 ( .A(n375), .B(n374), .ZN(n379) );
  XOR2_X1 U436 ( .A(KEYINPUT29), .B(KEYINPUT69), .Z(n377) );
  NAND2_X1 U437 ( .A1(G229GAT), .A2(G233GAT), .ZN(n376) );
  XNOR2_X1 U438 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U439 ( .A(n379), .B(n378), .Z(n384) );
  XOR2_X1 U440 ( .A(KEYINPUT68), .B(G8GAT), .Z(n381) );
  XNOR2_X1 U441 ( .A(G141GAT), .B(G22GAT), .ZN(n380) );
  XNOR2_X1 U442 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U443 ( .A(n382), .B(KEYINPUT30), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U445 ( .A(n386), .B(n385), .ZN(n503) );
  INV_X1 U446 ( .A(n503), .ZN(n580) );
  NOR2_X1 U447 ( .A1(n387), .A2(n580), .ZN(n389) );
  INV_X1 U448 ( .A(KEYINPUT110), .ZN(n388) );
  XNOR2_X1 U449 ( .A(n389), .B(n388), .ZN(n397) );
  XOR2_X1 U450 ( .A(KEYINPUT41), .B(KEYINPUT64), .Z(n390) );
  XNOR2_X1 U451 ( .A(n583), .B(n390), .ZN(n563) );
  NAND2_X1 U452 ( .A1(n580), .A2(n563), .ZN(n391) );
  XNOR2_X1 U453 ( .A(KEYINPUT46), .B(n391), .ZN(n393) );
  NAND2_X1 U454 ( .A1(n393), .A2(n392), .ZN(n394) );
  NOR2_X1 U455 ( .A1(n587), .A2(n394), .ZN(n395) );
  XNOR2_X1 U456 ( .A(KEYINPUT47), .B(n395), .ZN(n396) );
  XNOR2_X1 U457 ( .A(n398), .B(KEYINPUT48), .ZN(n529) );
  XOR2_X1 U458 ( .A(n400), .B(n399), .Z(n405) );
  XOR2_X1 U459 ( .A(G211GAT), .B(KEYINPUT91), .Z(n402) );
  XNOR2_X1 U460 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n401) );
  XNOR2_X1 U461 ( .A(n402), .B(n401), .ZN(n429) );
  XNOR2_X1 U462 ( .A(n403), .B(n429), .ZN(n404) );
  XNOR2_X1 U463 ( .A(n405), .B(n404), .ZN(n413) );
  XOR2_X1 U464 ( .A(KEYINPUT95), .B(KEYINPUT96), .Z(n407) );
  XNOR2_X1 U465 ( .A(G218GAT), .B(KEYINPUT94), .ZN(n406) );
  XNOR2_X1 U466 ( .A(n407), .B(n406), .ZN(n408) );
  XOR2_X1 U467 ( .A(n409), .B(n408), .Z(n411) );
  NAND2_X1 U468 ( .A1(G226GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U469 ( .A(n411), .B(n410), .ZN(n412) );
  NAND2_X1 U470 ( .A1(n529), .A2(n518), .ZN(n415) );
  XNOR2_X1 U471 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n414) );
  XNOR2_X1 U472 ( .A(n415), .B(n414), .ZN(n575) );
  XOR2_X1 U473 ( .A(KEYINPUT3), .B(KEYINPUT92), .Z(n417) );
  XNOR2_X1 U474 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n416) );
  XNOR2_X1 U475 ( .A(n417), .B(n416), .ZN(n441) );
  XOR2_X1 U476 ( .A(n418), .B(n441), .Z(n420) );
  NAND2_X1 U477 ( .A1(G228GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U478 ( .A(n420), .B(n419), .ZN(n422) );
  XOR2_X1 U479 ( .A(n422), .B(n421), .Z(n424) );
  XNOR2_X1 U480 ( .A(G106GAT), .B(G204GAT), .ZN(n423) );
  XNOR2_X1 U481 ( .A(n424), .B(n423), .ZN(n428) );
  XOR2_X1 U482 ( .A(KEYINPUT23), .B(KEYINPUT90), .Z(n426) );
  XNOR2_X1 U483 ( .A(KEYINPUT22), .B(KEYINPUT24), .ZN(n425) );
  XNOR2_X1 U484 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U485 ( .A(n428), .B(n427), .Z(n432) );
  XNOR2_X1 U486 ( .A(n430), .B(n429), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n465) );
  XOR2_X1 U488 ( .A(KEYINPUT4), .B(G57GAT), .Z(n434) );
  XNOR2_X1 U489 ( .A(G1GAT), .B(G155GAT), .ZN(n433) );
  XNOR2_X1 U490 ( .A(n434), .B(n433), .ZN(n450) );
  XOR2_X1 U491 ( .A(G148GAT), .B(G162GAT), .Z(n436) );
  XNOR2_X1 U492 ( .A(G120GAT), .B(G127GAT), .ZN(n435) );
  XNOR2_X1 U493 ( .A(n436), .B(n435), .ZN(n438) );
  XOR2_X1 U494 ( .A(G29GAT), .B(G85GAT), .Z(n437) );
  XNOR2_X1 U495 ( .A(n438), .B(n437), .ZN(n446) );
  XNOR2_X1 U496 ( .A(KEYINPUT1), .B(KEYINPUT93), .ZN(n439) );
  XNOR2_X1 U497 ( .A(n439), .B(KEYINPUT6), .ZN(n440) );
  XOR2_X1 U498 ( .A(n440), .B(KEYINPUT5), .Z(n444) );
  XNOR2_X1 U499 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n448) );
  NAND2_X1 U502 ( .A1(G225GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n450), .B(n449), .ZN(n528) );
  INV_X1 U505 ( .A(n528), .ZN(n574) );
  AND2_X1 U506 ( .A1(n465), .A2(n574), .ZN(n451) );
  NAND2_X1 U507 ( .A1(n575), .A2(n451), .ZN(n455) );
  XOR2_X1 U508 ( .A(KEYINPUT121), .B(KEYINPUT55), .Z(n453) );
  NOR2_X1 U509 ( .A1(n535), .A2(n456), .ZN(n570) );
  BUF_X1 U510 ( .A(n457), .Z(n544) );
  NAND2_X1 U511 ( .A1(n570), .A2(n544), .ZN(n459) );
  XOR2_X1 U512 ( .A(KEYINPUT34), .B(KEYINPUT98), .Z(n476) );
  NOR2_X1 U513 ( .A1(n583), .A2(n503), .ZN(n490) );
  XOR2_X1 U514 ( .A(n465), .B(KEYINPUT67), .Z(n460) );
  XOR2_X1 U515 ( .A(KEYINPUT28), .B(n460), .Z(n522) );
  INV_X1 U516 ( .A(n522), .ZN(n533) );
  XOR2_X1 U517 ( .A(n518), .B(KEYINPUT27), .Z(n531) );
  NOR2_X1 U518 ( .A1(n531), .A2(n520), .ZN(n461) );
  NAND2_X1 U519 ( .A1(n533), .A2(n461), .ZN(n462) );
  NAND2_X1 U520 ( .A1(n528), .A2(n462), .ZN(n471) );
  NAND2_X1 U521 ( .A1(n520), .A2(n518), .ZN(n463) );
  NAND2_X1 U522 ( .A1(n465), .A2(n463), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT25), .B(n464), .Z(n469) );
  NOR2_X1 U524 ( .A1(n465), .A2(n520), .ZN(n466) );
  XOR2_X1 U525 ( .A(n466), .B(KEYINPUT26), .Z(n548) );
  NOR2_X1 U526 ( .A1(n548), .A2(n531), .ZN(n467) );
  NOR2_X1 U527 ( .A1(n467), .A2(n528), .ZN(n468) );
  NAND2_X1 U528 ( .A1(n469), .A2(n468), .ZN(n470) );
  NAND2_X1 U529 ( .A1(n471), .A2(n470), .ZN(n485) );
  NOR2_X1 U530 ( .A1(n544), .A2(n486), .ZN(n472) );
  XOR2_X1 U531 ( .A(KEYINPUT16), .B(n472), .Z(n473) );
  NOR2_X1 U532 ( .A1(n485), .A2(n473), .ZN(n502) );
  NAND2_X1 U533 ( .A1(n490), .A2(n502), .ZN(n474) );
  XNOR2_X1 U534 ( .A(KEYINPUT97), .B(n474), .ZN(n483) );
  NAND2_X1 U535 ( .A1(n483), .A2(n528), .ZN(n475) );
  XNOR2_X1 U536 ( .A(n476), .B(n475), .ZN(n477) );
  XOR2_X1 U537 ( .A(G1GAT), .B(n477), .Z(G1324GAT) );
  NAND2_X1 U538 ( .A1(n483), .A2(n518), .ZN(n478) );
  XNOR2_X1 U539 ( .A(n478), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U540 ( .A(KEYINPUT100), .B(KEYINPUT35), .Z(n480) );
  NAND2_X1 U541 ( .A1(n483), .A2(n520), .ZN(n479) );
  XNOR2_X1 U542 ( .A(n480), .B(n479), .ZN(n482) );
  XOR2_X1 U543 ( .A(G15GAT), .B(KEYINPUT99), .Z(n481) );
  XNOR2_X1 U544 ( .A(n482), .B(n481), .ZN(G1326GAT) );
  NAND2_X1 U545 ( .A1(n483), .A2(n522), .ZN(n484) );
  XNOR2_X1 U546 ( .A(n484), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U547 ( .A(KEYINPUT102), .B(KEYINPUT38), .Z(n492) );
  NOR2_X1 U548 ( .A1(n591), .A2(n485), .ZN(n487) );
  NAND2_X1 U549 ( .A1(n487), .A2(n486), .ZN(n488) );
  XOR2_X1 U550 ( .A(KEYINPUT37), .B(n488), .Z(n516) );
  INV_X1 U551 ( .A(n516), .ZN(n489) );
  NAND2_X1 U552 ( .A1(n490), .A2(n489), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n492), .B(n491), .ZN(n500) );
  NAND2_X1 U554 ( .A1(n528), .A2(n500), .ZN(n496) );
  XOR2_X1 U555 ( .A(KEYINPUT101), .B(KEYINPUT39), .Z(n494) );
  XNOR2_X1 U556 ( .A(G29GAT), .B(KEYINPUT103), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n494), .B(n493), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1328GAT) );
  NAND2_X1 U559 ( .A1(n500), .A2(n518), .ZN(n497) );
  XNOR2_X1 U560 ( .A(n497), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U561 ( .A1(n500), .A2(n520), .ZN(n498) );
  XNOR2_X1 U562 ( .A(n498), .B(KEYINPUT40), .ZN(n499) );
  XNOR2_X1 U563 ( .A(G43GAT), .B(n499), .ZN(G1330GAT) );
  NAND2_X1 U564 ( .A1(n522), .A2(n500), .ZN(n501) );
  XNOR2_X1 U565 ( .A(G50GAT), .B(n501), .ZN(G1331GAT) );
  INV_X1 U566 ( .A(n502), .ZN(n504) );
  NAND2_X1 U567 ( .A1(n503), .A2(n563), .ZN(n515) );
  NOR2_X1 U568 ( .A1(n504), .A2(n515), .ZN(n512) );
  NAND2_X1 U569 ( .A1(n528), .A2(n512), .ZN(n508) );
  XOR2_X1 U570 ( .A(KEYINPUT105), .B(KEYINPUT106), .Z(n506) );
  XNOR2_X1 U571 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n505) );
  XNOR2_X1 U572 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U573 ( .A(n508), .B(n507), .ZN(n509) );
  XNOR2_X1 U574 ( .A(KEYINPUT104), .B(n509), .ZN(G1332GAT) );
  NAND2_X1 U575 ( .A1(n512), .A2(n518), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n510), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U577 ( .A1(n512), .A2(n520), .ZN(n511) );
  XNOR2_X1 U578 ( .A(n511), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U579 ( .A(G78GAT), .B(KEYINPUT43), .Z(n514) );
  NAND2_X1 U580 ( .A1(n512), .A2(n522), .ZN(n513) );
  XNOR2_X1 U581 ( .A(n514), .B(n513), .ZN(G1335GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n515), .ZN(n523) );
  NAND2_X1 U583 ( .A1(n523), .A2(n528), .ZN(n517) );
  XNOR2_X1 U584 ( .A(G85GAT), .B(n517), .ZN(G1336GAT) );
  NAND2_X1 U585 ( .A1(n523), .A2(n518), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U587 ( .A1(n523), .A2(n520), .ZN(n521) );
  XNOR2_X1 U588 ( .A(n521), .B(G99GAT), .ZN(G1338GAT) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(KEYINPUT107), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT44), .B(KEYINPUT108), .Z(n525) );
  NAND2_X1 U591 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U592 ( .A(n525), .B(n524), .ZN(n526) );
  XNOR2_X1 U593 ( .A(n527), .B(n526), .ZN(G1339GAT) );
  XOR2_X1 U594 ( .A(KEYINPUT112), .B(KEYINPUT113), .Z(n537) );
  NAND2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n530) );
  XOR2_X1 U596 ( .A(KEYINPUT111), .B(n532), .Z(n549) );
  NAND2_X1 U597 ( .A1(n549), .A2(n533), .ZN(n534) );
  NAND2_X1 U598 ( .A1(n545), .A2(n580), .ZN(n536) );
  XNOR2_X1 U599 ( .A(n537), .B(n536), .ZN(n538) );
  XNOR2_X1 U600 ( .A(G113GAT), .B(n538), .ZN(G1340GAT) );
  XOR2_X1 U601 ( .A(G120GAT), .B(KEYINPUT49), .Z(n540) );
  NAND2_X1 U602 ( .A1(n545), .A2(n563), .ZN(n539) );
  XNOR2_X1 U603 ( .A(n540), .B(n539), .ZN(G1341GAT) );
  XOR2_X1 U604 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n542) );
  NAND2_X1 U605 ( .A1(n545), .A2(n587), .ZN(n541) );
  XNOR2_X1 U606 ( .A(n542), .B(n541), .ZN(n543) );
  XOR2_X1 U607 ( .A(G127GAT), .B(n543), .Z(G1342GAT) );
  XOR2_X1 U608 ( .A(G134GAT), .B(KEYINPUT51), .Z(n547) );
  NAND2_X1 U609 ( .A1(n545), .A2(n544), .ZN(n546) );
  XNOR2_X1 U610 ( .A(n547), .B(n546), .ZN(G1343GAT) );
  INV_X1 U611 ( .A(n548), .ZN(n577) );
  NAND2_X1 U612 ( .A1(n549), .A2(n577), .ZN(n559) );
  INV_X1 U613 ( .A(n559), .ZN(n556) );
  NAND2_X1 U614 ( .A1(n580), .A2(n556), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT115), .B(n550), .Z(n551) );
  XNOR2_X1 U616 ( .A(G141GAT), .B(n551), .ZN(G1344GAT) );
  XNOR2_X1 U617 ( .A(G148GAT), .B(KEYINPUT116), .ZN(n555) );
  XOR2_X1 U618 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n553) );
  NAND2_X1 U619 ( .A1(n556), .A2(n563), .ZN(n552) );
  XNOR2_X1 U620 ( .A(n553), .B(n552), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(G1345GAT) );
  XOR2_X1 U622 ( .A(G155GAT), .B(KEYINPUT117), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n587), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1346GAT) );
  NOR2_X1 U625 ( .A1(n392), .A2(n559), .ZN(n560) );
  XOR2_X1 U626 ( .A(KEYINPUT118), .B(n560), .Z(n561) );
  XNOR2_X1 U627 ( .A(G162GAT), .B(n561), .ZN(G1347GAT) );
  NAND2_X1 U628 ( .A1(n570), .A2(n580), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U630 ( .A1(n563), .A2(n570), .ZN(n569) );
  XOR2_X1 U631 ( .A(KEYINPUT124), .B(KEYINPUT123), .Z(n565) );
  XNOR2_X1 U632 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n564) );
  XNOR2_X1 U633 ( .A(n565), .B(n564), .ZN(n567) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT122), .Z(n566) );
  XNOR2_X1 U635 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(G1349GAT) );
  NAND2_X1 U637 ( .A1(n570), .A2(n587), .ZN(n571) );
  XNOR2_X1 U638 ( .A(n571), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT126), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n572), .B(KEYINPUT60), .ZN(n573) );
  XOR2_X1 U641 ( .A(KEYINPUT59), .B(n573), .Z(n582) );
  AND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n576) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n579) );
  INV_X1 U644 ( .A(KEYINPUT125), .ZN(n578) );
  XNOR2_X1 U645 ( .A(n579), .B(n578), .ZN(n590) );
  INV_X1 U646 ( .A(n590), .ZN(n588) );
  NAND2_X1 U647 ( .A1(n588), .A2(n580), .ZN(n581) );
  XNOR2_X1 U648 ( .A(n582), .B(n581), .ZN(G1352GAT) );
  XOR2_X1 U649 ( .A(KEYINPUT127), .B(KEYINPUT61), .Z(n585) );
  NAND2_X1 U650 ( .A1(n588), .A2(n583), .ZN(n584) );
  XNOR2_X1 U651 ( .A(n585), .B(n584), .ZN(n586) );
  XOR2_X1 U652 ( .A(G204GAT), .B(n586), .Z(G1353GAT) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n589), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  XOR2_X1 U656 ( .A(KEYINPUT62), .B(n592), .Z(n593) );
  XNOR2_X1 U657 ( .A(G218GAT), .B(n593), .ZN(G1355GAT) );
endmodule

