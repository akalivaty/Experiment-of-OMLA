

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  INV_X1 U546 ( .A(n623), .ZN(n654) );
  NOR2_X1 U547 ( .A1(n612), .A2(n924), .ZN(n615) );
  AND2_X2 U548 ( .A1(n589), .A2(n697), .ZN(n623) );
  INV_X1 U549 ( .A(KEYINPUT99), .ZN(n682) );
  AND2_X1 U550 ( .A1(n676), .A2(n675), .ZN(n677) );
  NOR2_X1 U551 ( .A1(G2105), .A2(n529), .ZN(n581) );
  XNOR2_X1 U552 ( .A(n532), .B(KEYINPUT17), .ZN(n698) );
  NAND2_X1 U553 ( .A1(n695), .A2(n514), .ZN(n732) );
  BUF_X1 U554 ( .A(n698), .Z(n864) );
  NOR2_X1 U555 ( .A1(n663), .A2(n642), .ZN(n510) );
  XOR2_X1 U556 ( .A(KEYINPUT31), .B(n650), .Z(n511) );
  XOR2_X1 U557 ( .A(KEYINPUT14), .B(n603), .Z(n512) );
  OR2_X1 U558 ( .A1(n693), .A2(n692), .ZN(n513) );
  AND2_X1 U559 ( .A1(n694), .A2(n513), .ZN(n514) );
  AND2_X1 U560 ( .A1(n914), .A2(n744), .ZN(n515) );
  INV_X1 U561 ( .A(G8), .ZN(n642) );
  XNOR2_X1 U562 ( .A(KEYINPUT30), .B(KEYINPUT94), .ZN(n644) );
  XNOR2_X1 U563 ( .A(n645), .B(n644), .ZN(n646) );
  INV_X1 U564 ( .A(KEYINPUT29), .ZN(n635) );
  INV_X1 U565 ( .A(KEYINPUT95), .ZN(n652) );
  INV_X1 U566 ( .A(n921), .ZN(n674) );
  NAND2_X1 U567 ( .A1(G8), .A2(n654), .ZN(n693) );
  INV_X1 U568 ( .A(G2105), .ZN(n531) );
  NAND2_X1 U569 ( .A1(n749), .A2(n588), .ZN(n696) );
  XNOR2_X1 U570 ( .A(KEYINPUT23), .B(KEYINPUT65), .ZN(n582) );
  NOR2_X1 U571 ( .A1(n730), .A2(n515), .ZN(n731) );
  XNOR2_X1 U572 ( .A(n583), .B(n582), .ZN(n584) );
  XOR2_X1 U573 ( .A(KEYINPUT1), .B(n521), .Z(n780) );
  NOR2_X1 U574 ( .A1(G651), .A2(n541), .ZN(n781) );
  AND2_X1 U575 ( .A1(n585), .A2(n584), .ZN(n749) );
  NOR2_X2 U576 ( .A1(G651), .A2(G543), .ZN(n776) );
  NAND2_X1 U577 ( .A1(n776), .A2(G89), .ZN(n516) );
  XNOR2_X1 U578 ( .A(n516), .B(KEYINPUT4), .ZN(n518) );
  XOR2_X1 U579 ( .A(KEYINPUT0), .B(G543), .Z(n541) );
  INV_X1 U580 ( .A(G651), .ZN(n520) );
  NOR2_X1 U581 ( .A1(n541), .A2(n520), .ZN(n777) );
  NAND2_X1 U582 ( .A1(G76), .A2(n777), .ZN(n517) );
  NAND2_X1 U583 ( .A1(n518), .A2(n517), .ZN(n519) );
  XNOR2_X1 U584 ( .A(n519), .B(KEYINPUT5), .ZN(n527) );
  XNOR2_X1 U585 ( .A(KEYINPUT6), .B(KEYINPUT71), .ZN(n525) );
  NOR2_X1 U586 ( .A1(G543), .A2(n520), .ZN(n521) );
  NAND2_X1 U587 ( .A1(G63), .A2(n780), .ZN(n523) );
  NAND2_X1 U588 ( .A1(G51), .A2(n781), .ZN(n522) );
  NAND2_X1 U589 ( .A1(n523), .A2(n522), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(n526) );
  NAND2_X1 U591 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U592 ( .A(KEYINPUT7), .B(n528), .ZN(G168) );
  XOR2_X1 U593 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  INV_X1 U594 ( .A(G2104), .ZN(n529) );
  BUF_X1 U595 ( .A(n581), .Z(n530) );
  NAND2_X1 U596 ( .A1(G102), .A2(n530), .ZN(n534) );
  NAND2_X1 U597 ( .A1(n529), .A2(n531), .ZN(n532) );
  NAND2_X1 U598 ( .A1(G138), .A2(n698), .ZN(n533) );
  NAND2_X1 U599 ( .A1(n534), .A2(n533), .ZN(n539) );
  INV_X1 U600 ( .A(G2104), .ZN(n535) );
  AND2_X1 U601 ( .A1(n535), .A2(G2105), .ZN(n860) );
  NAND2_X1 U602 ( .A1(G126), .A2(n860), .ZN(n537) );
  AND2_X1 U603 ( .A1(G2104), .A2(G2105), .ZN(n861) );
  NAND2_X1 U604 ( .A1(G114), .A2(n861), .ZN(n536) );
  NAND2_X1 U605 ( .A1(n537), .A2(n536), .ZN(n538) );
  NOR2_X1 U606 ( .A1(n539), .A2(n538), .ZN(G164) );
  NAND2_X1 U607 ( .A1(G49), .A2(n781), .ZN(n540) );
  XNOR2_X1 U608 ( .A(n540), .B(KEYINPUT76), .ZN(n546) );
  NAND2_X1 U609 ( .A1(G87), .A2(n541), .ZN(n543) );
  NAND2_X1 U610 ( .A1(G74), .A2(G651), .ZN(n542) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  NOR2_X1 U612 ( .A1(n780), .A2(n544), .ZN(n545) );
  NAND2_X1 U613 ( .A1(n546), .A2(n545), .ZN(G288) );
  NAND2_X1 U614 ( .A1(G78), .A2(n777), .ZN(n548) );
  NAND2_X1 U615 ( .A1(G65), .A2(n780), .ZN(n547) );
  NAND2_X1 U616 ( .A1(n548), .A2(n547), .ZN(n551) );
  NAND2_X1 U617 ( .A1(G91), .A2(n776), .ZN(n549) );
  XNOR2_X1 U618 ( .A(KEYINPUT67), .B(n549), .ZN(n550) );
  NOR2_X1 U619 ( .A1(n551), .A2(n550), .ZN(n553) );
  NAND2_X1 U620 ( .A1(n781), .A2(G53), .ZN(n552) );
  NAND2_X1 U621 ( .A1(n553), .A2(n552), .ZN(G299) );
  NAND2_X1 U622 ( .A1(G64), .A2(n780), .ZN(n555) );
  NAND2_X1 U623 ( .A1(G52), .A2(n781), .ZN(n554) );
  NAND2_X1 U624 ( .A1(n555), .A2(n554), .ZN(n560) );
  NAND2_X1 U625 ( .A1(G90), .A2(n776), .ZN(n557) );
  NAND2_X1 U626 ( .A1(G77), .A2(n777), .ZN(n556) );
  NAND2_X1 U627 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U628 ( .A(KEYINPUT9), .B(n558), .Z(n559) );
  NOR2_X1 U629 ( .A1(n560), .A2(n559), .ZN(G171) );
  NAND2_X1 U630 ( .A1(G88), .A2(n776), .ZN(n562) );
  NAND2_X1 U631 ( .A1(G75), .A2(n777), .ZN(n561) );
  NAND2_X1 U632 ( .A1(n562), .A2(n561), .ZN(n566) );
  NAND2_X1 U633 ( .A1(G62), .A2(n780), .ZN(n564) );
  NAND2_X1 U634 ( .A1(G50), .A2(n781), .ZN(n563) );
  NAND2_X1 U635 ( .A1(n564), .A2(n563), .ZN(n565) );
  NOR2_X1 U636 ( .A1(n566), .A2(n565), .ZN(G166) );
  INV_X1 U637 ( .A(G166), .ZN(G303) );
  NAND2_X1 U638 ( .A1(G86), .A2(n776), .ZN(n568) );
  NAND2_X1 U639 ( .A1(G61), .A2(n780), .ZN(n567) );
  NAND2_X1 U640 ( .A1(n568), .A2(n567), .ZN(n571) );
  NAND2_X1 U641 ( .A1(n777), .A2(G73), .ZN(n569) );
  XOR2_X1 U642 ( .A(KEYINPUT2), .B(n569), .Z(n570) );
  NOR2_X1 U643 ( .A1(n571), .A2(n570), .ZN(n573) );
  NAND2_X1 U644 ( .A1(n781), .A2(G48), .ZN(n572) );
  NAND2_X1 U645 ( .A1(n573), .A2(n572), .ZN(G305) );
  NAND2_X1 U646 ( .A1(G85), .A2(n776), .ZN(n575) );
  NAND2_X1 U647 ( .A1(G72), .A2(n777), .ZN(n574) );
  NAND2_X1 U648 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U649 ( .A1(G47), .A2(n781), .ZN(n576) );
  XOR2_X1 U650 ( .A(KEYINPUT66), .B(n576), .Z(n577) );
  NOR2_X1 U651 ( .A1(n578), .A2(n577), .ZN(n580) );
  NAND2_X1 U652 ( .A1(n780), .A2(G60), .ZN(n579) );
  NAND2_X1 U653 ( .A1(n580), .A2(n579), .ZN(G290) );
  NAND2_X1 U654 ( .A1(G137), .A2(n698), .ZN(n585) );
  NAND2_X1 U655 ( .A1(G101), .A2(n581), .ZN(n583) );
  NAND2_X1 U656 ( .A1(G125), .A2(n860), .ZN(n587) );
  NAND2_X1 U657 ( .A1(G113), .A2(n861), .ZN(n586) );
  AND2_X1 U658 ( .A1(n587), .A2(n586), .ZN(n750) );
  AND2_X1 U659 ( .A1(G40), .A2(n750), .ZN(n588) );
  XNOR2_X1 U660 ( .A(KEYINPUT87), .B(n696), .ZN(n589) );
  NOR2_X1 U661 ( .A1(G164), .A2(G1384), .ZN(n697) );
  NOR2_X1 U662 ( .A1(G1976), .A2(G288), .ZN(n919) );
  NAND2_X1 U663 ( .A1(n919), .A2(KEYINPUT33), .ZN(n590) );
  NOR2_X1 U664 ( .A1(n693), .A2(n590), .ZN(n681) );
  NAND2_X1 U665 ( .A1(G92), .A2(n776), .ZN(n592) );
  NAND2_X1 U666 ( .A1(G66), .A2(n780), .ZN(n591) );
  NAND2_X1 U667 ( .A1(n592), .A2(n591), .ZN(n596) );
  NAND2_X1 U668 ( .A1(G79), .A2(n777), .ZN(n594) );
  NAND2_X1 U669 ( .A1(G54), .A2(n781), .ZN(n593) );
  NAND2_X1 U670 ( .A1(n594), .A2(n593), .ZN(n595) );
  NOR2_X1 U671 ( .A1(n596), .A2(n595), .ZN(n597) );
  XOR2_X1 U672 ( .A(KEYINPUT15), .B(n597), .Z(n888) );
  INV_X1 U673 ( .A(n888), .ZN(n614) );
  NAND2_X1 U674 ( .A1(n623), .A2(G1996), .ZN(n598) );
  XNOR2_X1 U675 ( .A(n598), .B(KEYINPUT26), .ZN(n600) );
  NAND2_X1 U676 ( .A1(G1341), .A2(n654), .ZN(n599) );
  NAND2_X1 U677 ( .A1(n600), .A2(n599), .ZN(n602) );
  INV_X1 U678 ( .A(KEYINPUT91), .ZN(n601) );
  XNOR2_X1 U679 ( .A(n602), .B(n601), .ZN(n612) );
  NAND2_X1 U680 ( .A1(G56), .A2(n780), .ZN(n603) );
  NAND2_X1 U681 ( .A1(G81), .A2(n776), .ZN(n604) );
  XNOR2_X1 U682 ( .A(n604), .B(KEYINPUT12), .ZN(n605) );
  XNOR2_X1 U683 ( .A(n605), .B(KEYINPUT68), .ZN(n607) );
  NAND2_X1 U684 ( .A1(G68), .A2(n777), .ZN(n606) );
  NAND2_X1 U685 ( .A1(n607), .A2(n606), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT13), .B(n608), .Z(n609) );
  NOR2_X1 U687 ( .A1(n512), .A2(n609), .ZN(n611) );
  NAND2_X1 U688 ( .A1(n781), .A2(G43), .ZN(n610) );
  NAND2_X1 U689 ( .A1(n611), .A2(n610), .ZN(n924) );
  INV_X1 U690 ( .A(n615), .ZN(n613) );
  NAND2_X1 U691 ( .A1(n614), .A2(n613), .ZN(n622) );
  NAND2_X1 U692 ( .A1(n615), .A2(n888), .ZN(n620) );
  NAND2_X1 U693 ( .A1(G1348), .A2(n654), .ZN(n617) );
  NAND2_X1 U694 ( .A1(G2067), .A2(n623), .ZN(n616) );
  NAND2_X1 U695 ( .A1(n617), .A2(n616), .ZN(n618) );
  XNOR2_X1 U696 ( .A(KEYINPUT92), .B(n618), .ZN(n619) );
  NAND2_X1 U697 ( .A1(n620), .A2(n619), .ZN(n621) );
  NAND2_X1 U698 ( .A1(n622), .A2(n621), .ZN(n629) );
  NAND2_X1 U699 ( .A1(n623), .A2(G2072), .ZN(n624) );
  XOR2_X1 U700 ( .A(KEYINPUT27), .B(n624), .Z(n626) );
  NAND2_X1 U701 ( .A1(G1956), .A2(n654), .ZN(n625) );
  NAND2_X1 U702 ( .A1(n626), .A2(n625), .ZN(n630) );
  NOR2_X1 U703 ( .A1(G299), .A2(n630), .ZN(n627) );
  XNOR2_X1 U704 ( .A(n627), .B(KEYINPUT93), .ZN(n628) );
  NAND2_X1 U705 ( .A1(n629), .A2(n628), .ZN(n634) );
  NAND2_X1 U706 ( .A1(n630), .A2(G299), .ZN(n631) );
  XNOR2_X1 U707 ( .A(n631), .B(KEYINPUT28), .ZN(n632) );
  XNOR2_X1 U708 ( .A(n632), .B(KEYINPUT90), .ZN(n633) );
  NAND2_X1 U709 ( .A1(n634), .A2(n633), .ZN(n636) );
  XNOR2_X1 U710 ( .A(n636), .B(n635), .ZN(n641) );
  XOR2_X1 U711 ( .A(G1961), .B(KEYINPUT88), .Z(n959) );
  NAND2_X1 U712 ( .A1(n959), .A2(n654), .ZN(n638) );
  XNOR2_X1 U713 ( .A(KEYINPUT25), .B(G2078), .ZN(n945) );
  NAND2_X1 U714 ( .A1(n623), .A2(n945), .ZN(n637) );
  NAND2_X1 U715 ( .A1(n638), .A2(n637), .ZN(n647) );
  AND2_X1 U716 ( .A1(n647), .A2(G171), .ZN(n639) );
  XNOR2_X1 U717 ( .A(n639), .B(KEYINPUT89), .ZN(n640) );
  NAND2_X1 U718 ( .A1(n641), .A2(n640), .ZN(n651) );
  NOR2_X1 U719 ( .A1(G1966), .A2(n693), .ZN(n666) );
  INV_X1 U720 ( .A(n666), .ZN(n643) );
  NOR2_X1 U721 ( .A1(G2084), .A2(n654), .ZN(n663) );
  NAND2_X1 U722 ( .A1(n643), .A2(n510), .ZN(n645) );
  NOR2_X1 U723 ( .A1(G168), .A2(n646), .ZN(n649) );
  NOR2_X1 U724 ( .A1(G171), .A2(n647), .ZN(n648) );
  NOR2_X1 U725 ( .A1(n649), .A2(n648), .ZN(n650) );
  NAND2_X1 U726 ( .A1(n651), .A2(n511), .ZN(n664) );
  NAND2_X1 U727 ( .A1(n664), .A2(G286), .ZN(n653) );
  XNOR2_X1 U728 ( .A(n653), .B(n652), .ZN(n660) );
  NOR2_X1 U729 ( .A1(G1971), .A2(n693), .ZN(n656) );
  NOR2_X1 U730 ( .A1(G2090), .A2(n654), .ZN(n655) );
  NOR2_X1 U731 ( .A1(n656), .A2(n655), .ZN(n657) );
  NAND2_X1 U732 ( .A1(n657), .A2(G303), .ZN(n658) );
  XNOR2_X1 U733 ( .A(KEYINPUT96), .B(n658), .ZN(n659) );
  NAND2_X1 U734 ( .A1(n660), .A2(n659), .ZN(n661) );
  NAND2_X1 U735 ( .A1(n661), .A2(G8), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n662), .B(KEYINPUT32), .ZN(n670) );
  NAND2_X1 U737 ( .A1(G8), .A2(n663), .ZN(n668) );
  INV_X1 U738 ( .A(n664), .ZN(n665) );
  NOR2_X1 U739 ( .A1(n666), .A2(n665), .ZN(n667) );
  NAND2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  NAND2_X1 U741 ( .A1(n670), .A2(n669), .ZN(n686) );
  NOR2_X1 U742 ( .A1(G1971), .A2(G303), .ZN(n671) );
  NOR2_X1 U743 ( .A1(n919), .A2(n671), .ZN(n672) );
  NAND2_X1 U744 ( .A1(n686), .A2(n672), .ZN(n676) );
  NAND2_X1 U745 ( .A1(G288), .A2(G1976), .ZN(n673) );
  XOR2_X1 U746 ( .A(KEYINPUT97), .B(n673), .Z(n921) );
  NOR2_X1 U747 ( .A1(n674), .A2(n693), .ZN(n675) );
  XNOR2_X1 U748 ( .A(n677), .B(KEYINPUT64), .ZN(n678) );
  NOR2_X1 U749 ( .A1(n678), .A2(KEYINPUT33), .ZN(n679) );
  XNOR2_X1 U750 ( .A(n679), .B(KEYINPUT98), .ZN(n680) );
  NOR2_X1 U751 ( .A1(n681), .A2(n680), .ZN(n683) );
  XNOR2_X1 U752 ( .A(n683), .B(n682), .ZN(n685) );
  XOR2_X1 U753 ( .A(G1981), .B(KEYINPUT100), .Z(n684) );
  XNOR2_X1 U754 ( .A(G305), .B(n684), .ZN(n910) );
  NAND2_X1 U755 ( .A1(n685), .A2(n910), .ZN(n695) );
  NOR2_X1 U756 ( .A1(G2090), .A2(G303), .ZN(n687) );
  NAND2_X1 U757 ( .A1(G8), .A2(n687), .ZN(n688) );
  NAND2_X1 U758 ( .A1(n686), .A2(n688), .ZN(n689) );
  XOR2_X1 U759 ( .A(KEYINPUT101), .B(n689), .Z(n690) );
  NAND2_X1 U760 ( .A1(n690), .A2(n693), .ZN(n694) );
  NOR2_X1 U761 ( .A1(G1981), .A2(G305), .ZN(n691) );
  XOR2_X1 U762 ( .A(n691), .B(KEYINPUT24), .Z(n692) );
  NOR2_X1 U763 ( .A1(n697), .A2(n696), .ZN(n744) );
  NAND2_X1 U764 ( .A1(G104), .A2(n530), .ZN(n700) );
  NAND2_X1 U765 ( .A1(G140), .A2(n864), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n700), .A2(n699), .ZN(n701) );
  XNOR2_X1 U767 ( .A(KEYINPUT34), .B(n701), .ZN(n706) );
  NAND2_X1 U768 ( .A1(G128), .A2(n860), .ZN(n703) );
  NAND2_X1 U769 ( .A1(G116), .A2(n861), .ZN(n702) );
  NAND2_X1 U770 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U771 ( .A(KEYINPUT35), .B(n704), .Z(n705) );
  NOR2_X1 U772 ( .A1(n706), .A2(n705), .ZN(n707) );
  XNOR2_X1 U773 ( .A(KEYINPUT36), .B(n707), .ZN(n883) );
  XNOR2_X1 U774 ( .A(G2067), .B(KEYINPUT37), .ZN(n742) );
  NOR2_X1 U775 ( .A1(n883), .A2(n742), .ZN(n988) );
  NAND2_X1 U776 ( .A1(n744), .A2(n988), .ZN(n708) );
  XOR2_X1 U777 ( .A(KEYINPUT81), .B(n708), .Z(n739) );
  NAND2_X1 U778 ( .A1(n860), .A2(G129), .ZN(n709) );
  XNOR2_X1 U779 ( .A(n709), .B(KEYINPUT82), .ZN(n711) );
  NAND2_X1 U780 ( .A1(G117), .A2(n861), .ZN(n710) );
  NAND2_X1 U781 ( .A1(n711), .A2(n710), .ZN(n715) );
  NAND2_X1 U782 ( .A1(G105), .A2(n530), .ZN(n712) );
  XNOR2_X1 U783 ( .A(n712), .B(KEYINPUT83), .ZN(n713) );
  XNOR2_X1 U784 ( .A(n713), .B(KEYINPUT38), .ZN(n714) );
  NOR2_X1 U785 ( .A1(n715), .A2(n714), .ZN(n716) );
  XNOR2_X1 U786 ( .A(n716), .B(KEYINPUT84), .ZN(n718) );
  NAND2_X1 U787 ( .A1(G141), .A2(n864), .ZN(n717) );
  NAND2_X1 U788 ( .A1(n718), .A2(n717), .ZN(n872) );
  NAND2_X1 U789 ( .A1(G1996), .A2(n872), .ZN(n719) );
  XOR2_X1 U790 ( .A(KEYINPUT85), .B(n719), .Z(n727) );
  NAND2_X1 U791 ( .A1(G95), .A2(n530), .ZN(n721) );
  NAND2_X1 U792 ( .A1(G131), .A2(n864), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n725) );
  NAND2_X1 U794 ( .A1(G119), .A2(n860), .ZN(n723) );
  NAND2_X1 U795 ( .A1(G107), .A2(n861), .ZN(n722) );
  NAND2_X1 U796 ( .A1(n723), .A2(n722), .ZN(n724) );
  OR2_X1 U797 ( .A1(n725), .A2(n724), .ZN(n859) );
  NAND2_X1 U798 ( .A1(G1991), .A2(n859), .ZN(n726) );
  NAND2_X1 U799 ( .A1(n727), .A2(n726), .ZN(n1003) );
  NAND2_X1 U800 ( .A1(n744), .A2(n1003), .ZN(n728) );
  NAND2_X1 U801 ( .A1(n739), .A2(n728), .ZN(n729) );
  XNOR2_X1 U802 ( .A(n729), .B(KEYINPUT86), .ZN(n730) );
  XNOR2_X1 U803 ( .A(G1986), .B(G290), .ZN(n914) );
  NAND2_X1 U804 ( .A1(n732), .A2(n731), .ZN(n747) );
  NOR2_X1 U805 ( .A1(G1996), .A2(n872), .ZN(n996) );
  NOR2_X1 U806 ( .A1(G1986), .A2(G290), .ZN(n733) );
  NOR2_X1 U807 ( .A1(G1991), .A2(n859), .ZN(n992) );
  NOR2_X1 U808 ( .A1(n733), .A2(n992), .ZN(n734) );
  XNOR2_X1 U809 ( .A(n734), .B(KEYINPUT102), .ZN(n735) );
  NOR2_X1 U810 ( .A1(n1003), .A2(n735), .ZN(n736) );
  NOR2_X1 U811 ( .A1(n996), .A2(n736), .ZN(n737) );
  XOR2_X1 U812 ( .A(KEYINPUT39), .B(n737), .Z(n738) );
  XNOR2_X1 U813 ( .A(KEYINPUT103), .B(n738), .ZN(n740) );
  NAND2_X1 U814 ( .A1(n740), .A2(n739), .ZN(n741) );
  XNOR2_X1 U815 ( .A(n741), .B(KEYINPUT104), .ZN(n743) );
  NAND2_X1 U816 ( .A1(n883), .A2(n742), .ZN(n993) );
  NAND2_X1 U817 ( .A1(n743), .A2(n993), .ZN(n745) );
  NAND2_X1 U818 ( .A1(n745), .A2(n744), .ZN(n746) );
  NAND2_X1 U819 ( .A1(n747), .A2(n746), .ZN(n748) );
  XNOR2_X1 U820 ( .A(n748), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U821 ( .A1(n749), .A2(n750), .ZN(G160) );
  AND2_X1 U822 ( .A1(G452), .A2(G94), .ZN(G173) );
  NAND2_X1 U823 ( .A1(G99), .A2(n530), .ZN(n751) );
  XNOR2_X1 U824 ( .A(n751), .B(KEYINPUT74), .ZN(n760) );
  NAND2_X1 U825 ( .A1(G123), .A2(n860), .ZN(n752) );
  XNOR2_X1 U826 ( .A(n752), .B(KEYINPUT18), .ZN(n753) );
  XNOR2_X1 U827 ( .A(n753), .B(KEYINPUT72), .ZN(n755) );
  NAND2_X1 U828 ( .A1(G135), .A2(n864), .ZN(n754) );
  NAND2_X1 U829 ( .A1(n755), .A2(n754), .ZN(n758) );
  NAND2_X1 U830 ( .A1(G111), .A2(n861), .ZN(n756) );
  XNOR2_X1 U831 ( .A(KEYINPUT73), .B(n756), .ZN(n757) );
  NOR2_X1 U832 ( .A1(n758), .A2(n757), .ZN(n759) );
  NAND2_X1 U833 ( .A1(n760), .A2(n759), .ZN(n989) );
  XNOR2_X1 U834 ( .A(G2096), .B(n989), .ZN(n761) );
  OR2_X1 U835 ( .A1(G2100), .A2(n761), .ZN(G156) );
  INV_X1 U836 ( .A(G57), .ZN(G237) );
  INV_X1 U837 ( .A(G132), .ZN(G219) );
  INV_X1 U838 ( .A(G82), .ZN(G220) );
  NAND2_X1 U839 ( .A1(G7), .A2(G661), .ZN(n762) );
  XNOR2_X1 U840 ( .A(n762), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U841 ( .A(G223), .ZN(n816) );
  NAND2_X1 U842 ( .A1(n816), .A2(G567), .ZN(n763) );
  XOR2_X1 U843 ( .A(KEYINPUT11), .B(n763), .Z(G234) );
  XNOR2_X1 U844 ( .A(G860), .B(KEYINPUT69), .ZN(n769) );
  OR2_X1 U845 ( .A1(n924), .A2(n769), .ZN(G153) );
  INV_X1 U846 ( .A(G171), .ZN(G301) );
  NAND2_X1 U847 ( .A1(G301), .A2(G868), .ZN(n764) );
  XNOR2_X1 U848 ( .A(n764), .B(KEYINPUT70), .ZN(n766) );
  INV_X1 U849 ( .A(G868), .ZN(n797) );
  NAND2_X1 U850 ( .A1(n797), .A2(n614), .ZN(n765) );
  NAND2_X1 U851 ( .A1(n766), .A2(n765), .ZN(G284) );
  NOR2_X1 U852 ( .A1(G286), .A2(n797), .ZN(n768) );
  NOR2_X1 U853 ( .A1(G868), .A2(G299), .ZN(n767) );
  NOR2_X1 U854 ( .A1(n768), .A2(n767), .ZN(G297) );
  NAND2_X1 U855 ( .A1(n769), .A2(G559), .ZN(n770) );
  NAND2_X1 U856 ( .A1(n770), .A2(n888), .ZN(n771) );
  XNOR2_X1 U857 ( .A(n771), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U858 ( .A1(G868), .A2(n924), .ZN(n774) );
  NAND2_X1 U859 ( .A1(G868), .A2(n888), .ZN(n772) );
  NOR2_X1 U860 ( .A1(G559), .A2(n772), .ZN(n773) );
  NOR2_X1 U861 ( .A1(n774), .A2(n773), .ZN(G282) );
  NAND2_X1 U862 ( .A1(n888), .A2(G559), .ZN(n794) );
  XNOR2_X1 U863 ( .A(n924), .B(n794), .ZN(n775) );
  NOR2_X1 U864 ( .A1(n775), .A2(G860), .ZN(n787) );
  NAND2_X1 U865 ( .A1(G93), .A2(n776), .ZN(n779) );
  NAND2_X1 U866 ( .A1(G80), .A2(n777), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n786) );
  NAND2_X1 U868 ( .A1(G67), .A2(n780), .ZN(n783) );
  NAND2_X1 U869 ( .A1(G55), .A2(n781), .ZN(n782) );
  NAND2_X1 U870 ( .A1(n783), .A2(n782), .ZN(n784) );
  XOR2_X1 U871 ( .A(KEYINPUT75), .B(n784), .Z(n785) );
  OR2_X1 U872 ( .A1(n786), .A2(n785), .ZN(n796) );
  XOR2_X1 U873 ( .A(n787), .B(n796), .Z(G145) );
  XNOR2_X1 U874 ( .A(G299), .B(G288), .ZN(n793) );
  XOR2_X1 U875 ( .A(n796), .B(KEYINPUT19), .Z(n789) );
  XNOR2_X1 U876 ( .A(n924), .B(G166), .ZN(n788) );
  XNOR2_X1 U877 ( .A(n789), .B(n788), .ZN(n790) );
  XOR2_X1 U878 ( .A(n790), .B(G290), .Z(n791) );
  XNOR2_X1 U879 ( .A(G305), .B(n791), .ZN(n792) );
  XNOR2_X1 U880 ( .A(n793), .B(n792), .ZN(n886) );
  XNOR2_X1 U881 ( .A(n794), .B(n886), .ZN(n795) );
  NAND2_X1 U882 ( .A1(n795), .A2(G868), .ZN(n799) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n798) );
  NAND2_X1 U884 ( .A1(n799), .A2(n798), .ZN(G295) );
  NAND2_X1 U885 ( .A1(G2078), .A2(G2084), .ZN(n800) );
  XNOR2_X1 U886 ( .A(n800), .B(KEYINPUT20), .ZN(n801) );
  XNOR2_X1 U887 ( .A(n801), .B(KEYINPUT77), .ZN(n802) );
  NAND2_X1 U888 ( .A1(n802), .A2(G2090), .ZN(n803) );
  XNOR2_X1 U889 ( .A(KEYINPUT21), .B(n803), .ZN(n804) );
  NAND2_X1 U890 ( .A1(n804), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U891 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U892 ( .A1(G220), .A2(G219), .ZN(n805) );
  XOR2_X1 U893 ( .A(KEYINPUT22), .B(n805), .Z(n806) );
  NOR2_X1 U894 ( .A1(G218), .A2(n806), .ZN(n807) );
  NAND2_X1 U895 ( .A1(G96), .A2(n807), .ZN(n821) );
  NAND2_X1 U896 ( .A1(G2106), .A2(n821), .ZN(n808) );
  XNOR2_X1 U897 ( .A(n808), .B(KEYINPUT78), .ZN(n812) );
  NAND2_X1 U898 ( .A1(G120), .A2(G69), .ZN(n809) );
  NOR2_X1 U899 ( .A1(G237), .A2(n809), .ZN(n810) );
  NAND2_X1 U900 ( .A1(G108), .A2(n810), .ZN(n822) );
  NAND2_X1 U901 ( .A1(G567), .A2(n822), .ZN(n811) );
  NAND2_X1 U902 ( .A1(n812), .A2(n811), .ZN(n823) );
  NAND2_X1 U903 ( .A1(G661), .A2(G483), .ZN(n813) );
  XOR2_X1 U904 ( .A(KEYINPUT79), .B(n813), .Z(n814) );
  NOR2_X1 U905 ( .A1(n823), .A2(n814), .ZN(n815) );
  XNOR2_X1 U906 ( .A(KEYINPUT80), .B(n815), .ZN(n819) );
  NAND2_X1 U907 ( .A1(G36), .A2(n819), .ZN(G176) );
  NAND2_X1 U908 ( .A1(G2106), .A2(n816), .ZN(G217) );
  AND2_X1 U909 ( .A1(G15), .A2(G2), .ZN(n817) );
  NAND2_X1 U910 ( .A1(G661), .A2(n817), .ZN(G259) );
  NAND2_X1 U911 ( .A1(G3), .A2(G1), .ZN(n818) );
  XNOR2_X1 U912 ( .A(n818), .B(KEYINPUT108), .ZN(n820) );
  NAND2_X1 U913 ( .A1(n820), .A2(n819), .ZN(G188) );
  XNOR2_X1 U914 ( .A(G69), .B(KEYINPUT109), .ZN(G235) );
  INV_X1 U916 ( .A(G120), .ZN(G236) );
  INV_X1 U917 ( .A(G96), .ZN(G221) );
  NOR2_X1 U918 ( .A1(n822), .A2(n821), .ZN(G325) );
  INV_X1 U919 ( .A(G325), .ZN(G261) );
  XOR2_X1 U920 ( .A(KEYINPUT110), .B(n823), .Z(G319) );
  XOR2_X1 U921 ( .A(G2100), .B(G2096), .Z(n825) );
  XNOR2_X1 U922 ( .A(KEYINPUT42), .B(G2678), .ZN(n824) );
  XNOR2_X1 U923 ( .A(n825), .B(n824), .ZN(n829) );
  XOR2_X1 U924 ( .A(KEYINPUT43), .B(G2090), .Z(n827) );
  XNOR2_X1 U925 ( .A(G2067), .B(G2072), .ZN(n826) );
  XNOR2_X1 U926 ( .A(n827), .B(n826), .ZN(n828) );
  XOR2_X1 U927 ( .A(n829), .B(n828), .Z(n831) );
  XNOR2_X1 U928 ( .A(G2078), .B(G2084), .ZN(n830) );
  XNOR2_X1 U929 ( .A(n831), .B(n830), .ZN(G227) );
  XOR2_X1 U930 ( .A(G1961), .B(G1956), .Z(n833) );
  XNOR2_X1 U931 ( .A(G1996), .B(G1986), .ZN(n832) );
  XNOR2_X1 U932 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U933 ( .A(G1976), .B(G1981), .Z(n835) );
  XNOR2_X1 U934 ( .A(G1966), .B(G1971), .ZN(n834) );
  XNOR2_X1 U935 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U936 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U937 ( .A(KEYINPUT111), .B(G2474), .ZN(n838) );
  XNOR2_X1 U938 ( .A(n839), .B(n838), .ZN(n841) );
  XOR2_X1 U939 ( .A(G1991), .B(KEYINPUT41), .Z(n840) );
  XNOR2_X1 U940 ( .A(n841), .B(n840), .ZN(G229) );
  NAND2_X1 U941 ( .A1(G112), .A2(n861), .ZN(n842) );
  XNOR2_X1 U942 ( .A(n842), .B(KEYINPUT112), .ZN(n845) );
  NAND2_X1 U943 ( .A1(G100), .A2(n530), .ZN(n843) );
  XOR2_X1 U944 ( .A(KEYINPUT113), .B(n843), .Z(n844) );
  NAND2_X1 U945 ( .A1(n845), .A2(n844), .ZN(n850) );
  NAND2_X1 U946 ( .A1(G124), .A2(n860), .ZN(n846) );
  XNOR2_X1 U947 ( .A(n846), .B(KEYINPUT44), .ZN(n848) );
  NAND2_X1 U948 ( .A1(n864), .A2(G136), .ZN(n847) );
  NAND2_X1 U949 ( .A1(n848), .A2(n847), .ZN(n849) );
  NOR2_X1 U950 ( .A1(n850), .A2(n849), .ZN(G162) );
  NAND2_X1 U951 ( .A1(G103), .A2(n530), .ZN(n852) );
  NAND2_X1 U952 ( .A1(G139), .A2(n864), .ZN(n851) );
  NAND2_X1 U953 ( .A1(n852), .A2(n851), .ZN(n857) );
  NAND2_X1 U954 ( .A1(G127), .A2(n860), .ZN(n854) );
  NAND2_X1 U955 ( .A1(G115), .A2(n861), .ZN(n853) );
  NAND2_X1 U956 ( .A1(n854), .A2(n853), .ZN(n855) );
  XOR2_X1 U957 ( .A(KEYINPUT47), .B(n855), .Z(n856) );
  NOR2_X1 U958 ( .A1(n857), .A2(n856), .ZN(n983) );
  XOR2_X1 U959 ( .A(G164), .B(n983), .Z(n858) );
  XNOR2_X1 U960 ( .A(n859), .B(n858), .ZN(n871) );
  NAND2_X1 U961 ( .A1(G130), .A2(n860), .ZN(n863) );
  NAND2_X1 U962 ( .A1(G118), .A2(n861), .ZN(n862) );
  NAND2_X1 U963 ( .A1(n863), .A2(n862), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G106), .A2(n530), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G142), .A2(n864), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(n867), .B(KEYINPUT45), .Z(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U969 ( .A(n871), .B(n870), .Z(n873) );
  XNOR2_X1 U970 ( .A(n873), .B(n872), .ZN(n882) );
  XOR2_X1 U971 ( .A(KEYINPUT115), .B(KEYINPUT46), .Z(n875) );
  XNOR2_X1 U972 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n874) );
  XNOR2_X1 U973 ( .A(n875), .B(n874), .ZN(n876) );
  XNOR2_X1 U974 ( .A(KEYINPUT114), .B(n876), .ZN(n878) );
  XNOR2_X1 U975 ( .A(n989), .B(KEYINPUT48), .ZN(n877) );
  XNOR2_X1 U976 ( .A(n878), .B(n877), .ZN(n880) );
  XOR2_X1 U977 ( .A(G160), .B(G162), .Z(n879) );
  XNOR2_X1 U978 ( .A(n880), .B(n879), .ZN(n881) );
  XNOR2_X1 U979 ( .A(n882), .B(n881), .ZN(n884) );
  XOR2_X1 U980 ( .A(n884), .B(n883), .Z(n885) );
  NOR2_X1 U981 ( .A1(G37), .A2(n885), .ZN(G395) );
  XNOR2_X1 U982 ( .A(G286), .B(G301), .ZN(n887) );
  XNOR2_X1 U983 ( .A(n887), .B(n886), .ZN(n889) );
  XNOR2_X1 U984 ( .A(n889), .B(n888), .ZN(n890) );
  NOR2_X1 U985 ( .A1(G37), .A2(n890), .ZN(G397) );
  XOR2_X1 U986 ( .A(G2443), .B(G2451), .Z(n892) );
  XNOR2_X1 U987 ( .A(KEYINPUT106), .B(G2427), .ZN(n891) );
  XNOR2_X1 U988 ( .A(n892), .B(n891), .ZN(n893) );
  XOR2_X1 U989 ( .A(n893), .B(G2430), .Z(n895) );
  XNOR2_X1 U990 ( .A(G1341), .B(G1348), .ZN(n894) );
  XNOR2_X1 U991 ( .A(n895), .B(n894), .ZN(n899) );
  XOR2_X1 U992 ( .A(G2438), .B(G2435), .Z(n897) );
  XNOR2_X1 U993 ( .A(KEYINPUT107), .B(G2454), .ZN(n896) );
  XNOR2_X1 U994 ( .A(n897), .B(n896), .ZN(n898) );
  XOR2_X1 U995 ( .A(n899), .B(n898), .Z(n901) );
  XNOR2_X1 U996 ( .A(G2446), .B(KEYINPUT105), .ZN(n900) );
  XNOR2_X1 U997 ( .A(n901), .B(n900), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n902), .A2(G14), .ZN(n908) );
  NAND2_X1 U999 ( .A1(n908), .A2(G319), .ZN(n905) );
  NOR2_X1 U1000 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U1001 ( .A(KEYINPUT49), .B(n903), .ZN(n904) );
  NOR2_X1 U1002 ( .A1(n905), .A2(n904), .ZN(n907) );
  NOR2_X1 U1003 ( .A1(G395), .A2(G397), .ZN(n906) );
  NAND2_X1 U1004 ( .A1(n907), .A2(n906), .ZN(G225) );
  INV_X1 U1005 ( .A(G225), .ZN(G308) );
  INV_X1 U1006 ( .A(G108), .ZN(G238) );
  INV_X1 U1007 ( .A(n908), .ZN(G401) );
  XNOR2_X1 U1008 ( .A(G16), .B(KEYINPUT56), .ZN(n937) );
  XNOR2_X1 U1009 ( .A(G1966), .B(G168), .ZN(n909) );
  XNOR2_X1 U1010 ( .A(n909), .B(KEYINPUT120), .ZN(n911) );
  NAND2_X1 U1011 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1012 ( .A(KEYINPUT57), .B(n912), .ZN(n935) );
  XNOR2_X1 U1013 ( .A(G1956), .B(G299), .ZN(n913) );
  NOR2_X1 U1014 ( .A1(n914), .A2(n913), .ZN(n932) );
  XNOR2_X1 U1015 ( .A(G171), .B(G1961), .ZN(n917) );
  XNOR2_X1 U1016 ( .A(G1348), .B(KEYINPUT121), .ZN(n915) );
  XNOR2_X1 U1017 ( .A(n915), .B(n614), .ZN(n916) );
  NAND2_X1 U1018 ( .A1(n917), .A2(n916), .ZN(n918) );
  XNOR2_X1 U1019 ( .A(n918), .B(KEYINPUT122), .ZN(n930) );
  INV_X1 U1020 ( .A(n919), .ZN(n920) );
  NAND2_X1 U1021 ( .A1(n921), .A2(n920), .ZN(n922) );
  XNOR2_X1 U1022 ( .A(n922), .B(KEYINPUT123), .ZN(n928) );
  XNOR2_X1 U1023 ( .A(G1971), .B(KEYINPUT124), .ZN(n923) );
  XNOR2_X1 U1024 ( .A(n923), .B(G303), .ZN(n926) );
  XNOR2_X1 U1025 ( .A(G1341), .B(n924), .ZN(n925) );
  NOR2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1027 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1028 ( .A1(n930), .A2(n929), .ZN(n931) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(KEYINPUT125), .B(n933), .ZN(n934) );
  NAND2_X1 U1031 ( .A1(n935), .A2(n934), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n937), .A2(n936), .ZN(n1011) );
  XOR2_X1 U1033 ( .A(G2090), .B(G35), .Z(n951) );
  XOR2_X1 U1034 ( .A(KEYINPUT53), .B(KEYINPUT118), .Z(n949) );
  XNOR2_X1 U1035 ( .A(G1996), .B(G32), .ZN(n939) );
  XNOR2_X1 U1036 ( .A(G33), .B(G2072), .ZN(n938) );
  NOR2_X1 U1037 ( .A1(n939), .A2(n938), .ZN(n944) );
  XOR2_X1 U1038 ( .A(G2067), .B(G26), .Z(n940) );
  NAND2_X1 U1039 ( .A1(n940), .A2(G28), .ZN(n942) );
  XNOR2_X1 U1040 ( .A(G25), .B(G1991), .ZN(n941) );
  NOR2_X1 U1041 ( .A1(n942), .A2(n941), .ZN(n943) );
  NAND2_X1 U1042 ( .A1(n944), .A2(n943), .ZN(n947) );
  XOR2_X1 U1043 ( .A(G27), .B(n945), .Z(n946) );
  NOR2_X1 U1044 ( .A1(n947), .A2(n946), .ZN(n948) );
  XNOR2_X1 U1045 ( .A(n949), .B(n948), .ZN(n950) );
  NAND2_X1 U1046 ( .A1(n951), .A2(n950), .ZN(n954) );
  XNOR2_X1 U1047 ( .A(G34), .B(G2084), .ZN(n952) );
  XNOR2_X1 U1048 ( .A(KEYINPUT54), .B(n952), .ZN(n953) );
  NOR2_X1 U1049 ( .A1(n954), .A2(n953), .ZN(n955) );
  XOR2_X1 U1050 ( .A(KEYINPUT119), .B(n955), .Z(n956) );
  NOR2_X1 U1051 ( .A1(G29), .A2(n956), .ZN(n957) );
  XNOR2_X1 U1052 ( .A(KEYINPUT55), .B(n957), .ZN(n958) );
  NAND2_X1 U1053 ( .A1(n958), .A2(G11), .ZN(n1009) );
  XNOR2_X1 U1054 ( .A(n959), .B(G5), .ZN(n969) );
  XNOR2_X1 U1055 ( .A(G1971), .B(G22), .ZN(n961) );
  XNOR2_X1 U1056 ( .A(G23), .B(G1976), .ZN(n960) );
  NOR2_X1 U1057 ( .A1(n961), .A2(n960), .ZN(n962) );
  XOR2_X1 U1058 ( .A(KEYINPUT126), .B(n962), .Z(n964) );
  XNOR2_X1 U1059 ( .A(G1986), .B(G24), .ZN(n963) );
  NOR2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  XOR2_X1 U1061 ( .A(KEYINPUT58), .B(n965), .Z(n967) );
  XNOR2_X1 U1062 ( .A(G1966), .B(G21), .ZN(n966) );
  NOR2_X1 U1063 ( .A1(n967), .A2(n966), .ZN(n968) );
  NAND2_X1 U1064 ( .A1(n969), .A2(n968), .ZN(n979) );
  XOR2_X1 U1065 ( .A(G1348), .B(KEYINPUT59), .Z(n970) );
  XNOR2_X1 U1066 ( .A(G4), .B(n970), .ZN(n972) );
  XNOR2_X1 U1067 ( .A(G20), .B(G1956), .ZN(n971) );
  NOR2_X1 U1068 ( .A1(n972), .A2(n971), .ZN(n976) );
  XNOR2_X1 U1069 ( .A(G1341), .B(G19), .ZN(n974) );
  XNOR2_X1 U1070 ( .A(G6), .B(G1981), .ZN(n973) );
  NOR2_X1 U1071 ( .A1(n974), .A2(n973), .ZN(n975) );
  NAND2_X1 U1072 ( .A1(n976), .A2(n975), .ZN(n977) );
  XNOR2_X1 U1073 ( .A(KEYINPUT60), .B(n977), .ZN(n978) );
  NOR2_X1 U1074 ( .A1(n979), .A2(n978), .ZN(n980) );
  XOR2_X1 U1075 ( .A(KEYINPUT61), .B(n980), .Z(n981) );
  NOR2_X1 U1076 ( .A1(G16), .A2(n981), .ZN(n982) );
  XNOR2_X1 U1077 ( .A(KEYINPUT127), .B(n982), .ZN(n1007) );
  XOR2_X1 U1078 ( .A(G2072), .B(n983), .Z(n985) );
  XOR2_X1 U1079 ( .A(G164), .B(G2078), .Z(n984) );
  NOR2_X1 U1080 ( .A1(n985), .A2(n984), .ZN(n986) );
  XOR2_X1 U1081 ( .A(KEYINPUT50), .B(n986), .Z(n987) );
  NOR2_X1 U1082 ( .A1(n988), .A2(n987), .ZN(n1001) );
  XNOR2_X1 U1083 ( .A(G160), .B(G2084), .ZN(n990) );
  NAND2_X1 U1084 ( .A1(n990), .A2(n989), .ZN(n991) );
  NOR2_X1 U1085 ( .A1(n992), .A2(n991), .ZN(n994) );
  NAND2_X1 U1086 ( .A1(n994), .A2(n993), .ZN(n999) );
  XOR2_X1 U1087 ( .A(G2090), .B(G162), .Z(n995) );
  NOR2_X1 U1088 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1089 ( .A(n997), .B(KEYINPUT51), .ZN(n998) );
  NOR2_X1 U1090 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1091 ( .A1(n1001), .A2(n1000), .ZN(n1002) );
  NOR2_X1 U1092 ( .A1(n1003), .A2(n1002), .ZN(n1004) );
  XOR2_X1 U1093 ( .A(KEYINPUT52), .B(n1004), .Z(n1005) );
  NAND2_X1 U1094 ( .A1(n1005), .A2(G29), .ZN(n1006) );
  NAND2_X1 U1095 ( .A1(n1007), .A2(n1006), .ZN(n1008) );
  NOR2_X1 U1096 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  NAND2_X1 U1097 ( .A1(n1011), .A2(n1010), .ZN(n1012) );
  XOR2_X1 U1098 ( .A(KEYINPUT62), .B(n1012), .Z(G311) );
  INV_X1 U1099 ( .A(G311), .ZN(G150) );
endmodule

