//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 1 1 1 1 0 0 1 1 0 1 1 0 1 1 1 1 0 0 0 1 1 1 0 0 0 0 0 0 0 1 0 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:15:18 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n682, new_n683, new_n684, new_n685,
    new_n687, new_n688, new_n689, new_n691, new_n692, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n754, new_n755, new_n756,
    new_n757, new_n759, new_n760, new_n761, new_n763, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n835, new_n836, new_n838, new_n839, new_n841, new_n842, new_n843,
    new_n844, new_n845, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n904, new_n905, new_n906, new_n907, new_n909, new_n910,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n919,
    new_n920, new_n921, new_n922, new_n924, new_n925, new_n926, new_n927,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n957, new_n958;
  INV_X1    g000(.A(KEYINPUT91), .ZN(new_n202));
  XNOR2_X1  g001(.A(G1gat), .B(G29gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n203), .B(KEYINPUT0), .ZN(new_n204));
  XNOR2_X1  g003(.A(G57gat), .B(G85gat), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n204), .B(new_n205), .Z(new_n206));
  XOR2_X1   g005(.A(KEYINPUT78), .B(KEYINPUT5), .Z(new_n207));
  NAND2_X1  g006(.A1(G155gat), .A2(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n209), .A2(new_n210), .ZN(new_n211));
  OAI21_X1  g010(.A(new_n208), .B1(new_n211), .B2(KEYINPUT2), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT75), .ZN(new_n213));
  INV_X1    g012(.A(G148gat), .ZN(new_n214));
  OAI21_X1  g013(.A(new_n213), .B1(new_n214), .B2(G141gat), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n214), .A2(G141gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(G141gat), .ZN(new_n218));
  NAND2_X1  g017(.A1(new_n218), .A2(G148gat), .ZN(new_n219));
  NOR2_X1   g018(.A1(new_n219), .A2(new_n213), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n212), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT76), .ZN(new_n222));
  XNOR2_X1  g021(.A(new_n221), .B(new_n222), .ZN(new_n223));
  AOI22_X1  g022(.A1(new_n216), .A2(new_n219), .B1(KEYINPUT2), .B2(new_n208), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n211), .A2(new_n208), .ZN(new_n225));
  AOI21_X1  g024(.A(new_n224), .B1(KEYINPUT74), .B2(new_n225), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(KEYINPUT74), .B2(new_n225), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n223), .A2(new_n227), .ZN(new_n228));
  XOR2_X1   g027(.A(G127gat), .B(G134gat), .Z(new_n229));
  XNOR2_X1  g028(.A(G113gat), .B(G120gat), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g030(.A(new_n231), .B(KEYINPUT68), .ZN(new_n232));
  XNOR2_X1  g031(.A(KEYINPUT69), .B(G113gat), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n233), .A2(G120gat), .ZN(new_n234));
  INV_X1    g033(.A(G120gat), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(G113gat), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n234), .A2(KEYINPUT70), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n229), .A2(KEYINPUT1), .ZN(new_n238));
  OAI211_X1 g037(.A(new_n237), .B(new_n238), .C1(KEYINPUT70), .C2(new_n234), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n232), .A2(new_n239), .ZN(new_n240));
  XNOR2_X1  g039(.A(new_n228), .B(new_n240), .ZN(new_n241));
  NAND2_X1  g040(.A1(G225gat), .A2(G233gat), .ZN(new_n242));
  INV_X1    g041(.A(new_n242), .ZN(new_n243));
  AOI21_X1  g042(.A(new_n207), .B1(new_n241), .B2(new_n243), .ZN(new_n244));
  OR3_X1    g043(.A1(new_n228), .A2(new_n240), .A3(KEYINPUT4), .ZN(new_n245));
  OAI21_X1  g044(.A(KEYINPUT4), .B1(new_n228), .B2(new_n240), .ZN(new_n246));
  AND3_X1   g045(.A1(new_n245), .A2(KEYINPUT77), .A3(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n228), .A2(KEYINPUT3), .ZN(new_n248));
  INV_X1    g047(.A(KEYINPUT3), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n223), .A2(new_n249), .A3(new_n227), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n248), .A2(new_n240), .A3(new_n250), .ZN(new_n251));
  OAI211_X1 g050(.A(new_n251), .B(new_n242), .C1(KEYINPUT77), .C2(new_n246), .ZN(new_n252));
  OAI21_X1  g051(.A(new_n244), .B1(new_n247), .B2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n245), .A2(new_n246), .ZN(new_n254));
  NAND4_X1  g053(.A1(new_n254), .A2(new_n242), .A3(new_n251), .A4(new_n207), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n206), .B1(new_n253), .B2(new_n255), .ZN(new_n256));
  INV_X1    g055(.A(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT6), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n253), .A2(new_n255), .A3(new_n206), .ZN(new_n259));
  NAND3_X1  g058(.A1(new_n257), .A2(new_n258), .A3(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n259), .A2(new_n258), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n261), .A2(new_n256), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  XNOR2_X1  g062(.A(G8gat), .B(G36gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(G64gat), .B(G92gat), .ZN(new_n265));
  XOR2_X1   g064(.A(new_n264), .B(new_n265), .Z(new_n266));
  XNOR2_X1  g065(.A(G197gat), .B(G204gat), .ZN(new_n267));
  INV_X1    g066(.A(KEYINPUT22), .ZN(new_n268));
  INV_X1    g067(.A(G211gat), .ZN(new_n269));
  INV_X1    g068(.A(G218gat), .ZN(new_n270));
  OAI21_X1  g069(.A(new_n268), .B1(new_n269), .B2(new_n270), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n267), .A2(new_n271), .ZN(new_n272));
  XOR2_X1   g071(.A(G211gat), .B(G218gat), .Z(new_n273));
  NAND2_X1  g072(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(new_n273), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n275), .A2(new_n267), .A3(new_n271), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT71), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n272), .A2(new_n273), .ZN(new_n279));
  NOR2_X1   g078(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n280));
  OAI21_X1  g079(.A(new_n274), .B1(new_n278), .B2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G226gat), .A2(G233gat), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NOR2_X1   g082(.A1(new_n283), .A2(KEYINPUT29), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  XOR2_X1   g084(.A(KEYINPUT66), .B(G190gat), .Z(new_n286));
  INV_X1    g085(.A(G183gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g087(.A(KEYINPUT24), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n289), .A2(G183gat), .A3(G190gat), .ZN(new_n290));
  INV_X1    g089(.A(G190gat), .ZN(new_n291));
  NOR2_X1   g090(.A1(new_n287), .A2(new_n291), .ZN(new_n292));
  OAI21_X1  g091(.A(new_n290), .B1(new_n292), .B2(new_n289), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  NOR2_X1   g093(.A1(G169gat), .A2(G176gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n295), .A2(KEYINPUT23), .ZN(new_n296));
  NAND2_X1  g095(.A1(G169gat), .A2(G176gat), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n297), .A2(KEYINPUT23), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(G169gat), .B2(G176gat), .ZN(new_n299));
  NAND4_X1  g098(.A1(new_n294), .A2(KEYINPUT25), .A3(new_n296), .A4(new_n299), .ZN(new_n300));
  OAI21_X1  g099(.A(new_n293), .B1(G183gat), .B2(G190gat), .ZN(new_n301));
  NAND3_X1  g100(.A1(new_n295), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT65), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n296), .A2(new_n303), .ZN(new_n304));
  AND4_X1   g103(.A1(new_n301), .A2(new_n302), .A3(new_n299), .A4(new_n304), .ZN(new_n305));
  XNOR2_X1  g104(.A(KEYINPUT64), .B(KEYINPUT25), .ZN(new_n306));
  OAI21_X1  g105(.A(new_n300), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  XNOR2_X1  g106(.A(KEYINPUT27), .B(G183gat), .ZN(new_n308));
  AOI21_X1  g107(.A(KEYINPUT67), .B1(new_n286), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT28), .ZN(new_n310));
  XNOR2_X1  g109(.A(new_n309), .B(new_n310), .ZN(new_n311));
  AND2_X1   g110(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n295), .A2(KEYINPUT26), .ZN(new_n313));
  AOI211_X1 g112(.A(new_n292), .B(new_n312), .C1(new_n297), .C2(new_n313), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n311), .A2(new_n314), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n307), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT73), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n307), .A2(new_n315), .A3(KEYINPUT73), .ZN(new_n319));
  AOI21_X1  g118(.A(new_n285), .B1(new_n318), .B2(new_n319), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n316), .A2(new_n282), .ZN(new_n321));
  OAI21_X1  g120(.A(new_n281), .B1(new_n320), .B2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n318), .A2(new_n283), .A3(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n276), .A2(new_n277), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n279), .A2(KEYINPUT71), .ZN(new_n325));
  AOI22_X1  g124(.A1(new_n324), .A2(new_n325), .B1(new_n273), .B2(new_n272), .ZN(new_n326));
  XNOR2_X1  g125(.A(KEYINPUT72), .B(KEYINPUT29), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n316), .A2(new_n282), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n323), .A2(new_n326), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n266), .B1(new_n322), .B2(new_n329), .ZN(new_n330));
  INV_X1    g129(.A(new_n330), .ZN(new_n331));
  NAND3_X1  g130(.A1(new_n322), .A2(new_n329), .A3(new_n266), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n331), .A2(new_n332), .A3(KEYINPUT30), .ZN(new_n333));
  INV_X1    g132(.A(KEYINPUT30), .ZN(new_n334));
  NAND4_X1  g133(.A1(new_n322), .A2(new_n334), .A3(new_n329), .A4(new_n266), .ZN(new_n335));
  NAND2_X1  g134(.A1(new_n333), .A2(new_n335), .ZN(new_n336));
  NAND2_X1  g135(.A1(new_n263), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n250), .A2(new_n327), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(new_n326), .ZN(new_n339));
  INV_X1    g138(.A(KEYINPUT81), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n340), .B1(new_n278), .B2(new_n280), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n324), .A2(KEYINPUT81), .A3(new_n325), .ZN(new_n342));
  XNOR2_X1  g141(.A(new_n274), .B(KEYINPUT82), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(new_n342), .A3(new_n343), .ZN(new_n344));
  AOI21_X1  g143(.A(KEYINPUT3), .B1(new_n344), .B2(new_n327), .ZN(new_n345));
  INV_X1    g144(.A(new_n228), .ZN(new_n346));
  OAI21_X1  g145(.A(new_n339), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT83), .ZN(new_n348));
  AND2_X1   g147(.A1(G228gat), .A2(G233gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n349), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n347), .A2(new_n348), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n347), .B2(new_n350), .ZN(new_n352));
  INV_X1    g151(.A(KEYINPUT84), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n353), .B1(new_n326), .B2(KEYINPUT29), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n354), .A2(new_n249), .ZN(new_n355));
  NOR3_X1   g154(.A1(new_n326), .A2(new_n353), .A3(KEYINPUT29), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n228), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n350), .B1(new_n338), .B2(new_n326), .ZN(new_n358));
  AND3_X1   g157(.A1(new_n357), .A2(KEYINPUT85), .A3(new_n358), .ZN(new_n359));
  AOI21_X1  g158(.A(KEYINPUT85), .B1(new_n357), .B2(new_n358), .ZN(new_n360));
  OAI22_X1  g159(.A1(new_n351), .A2(new_n352), .B1(new_n359), .B2(new_n360), .ZN(new_n361));
  NOR2_X1   g160(.A1(new_n361), .A2(G22gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(G78gat), .B(G106gat), .ZN(new_n363));
  XNOR2_X1  g162(.A(new_n363), .B(KEYINPUT79), .ZN(new_n364));
  XNOR2_X1  g163(.A(KEYINPUT31), .B(G50gat), .ZN(new_n365));
  XNOR2_X1  g164(.A(new_n364), .B(new_n365), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n362), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n361), .A2(G22gat), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT87), .ZN(new_n369));
  NAND2_X1  g168(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(KEYINPUT87), .A3(G22gat), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(new_n370), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(G22gat), .ZN(new_n373));
  OAI221_X1 g172(.A(new_n373), .B1(new_n359), .B2(new_n360), .C1(new_n351), .C2(new_n352), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n368), .A2(new_n374), .ZN(new_n375));
  XOR2_X1   g174(.A(new_n366), .B(KEYINPUT80), .Z(new_n376));
  INV_X1    g175(.A(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(KEYINPUT86), .B1(new_n375), .B2(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT86), .ZN(new_n379));
  AOI211_X1 g178(.A(new_n379), .B(new_n376), .C1(new_n368), .C2(new_n374), .ZN(new_n380));
  OAI211_X1 g179(.A(new_n337), .B(new_n372), .C1(new_n378), .C2(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT36), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n316), .B(new_n240), .ZN(new_n383));
  AND2_X1   g182(.A1(G227gat), .A2(G233gat), .ZN(new_n384));
  NOR3_X1   g183(.A1(new_n383), .A2(KEYINPUT34), .A3(new_n384), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OAI21_X1  g185(.A(KEYINPUT34), .B1(new_n383), .B2(new_n384), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT33), .B1(new_n383), .B2(new_n384), .ZN(new_n388));
  XOR2_X1   g187(.A(G15gat), .B(G43gat), .Z(new_n389));
  XNOR2_X1  g188(.A(G71gat), .B(G99gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n389), .B(new_n390), .ZN(new_n391));
  INV_X1    g190(.A(new_n391), .ZN(new_n392));
  OAI211_X1 g191(.A(new_n386), .B(new_n387), .C1(new_n388), .C2(new_n392), .ZN(new_n393));
  NOR2_X1   g192(.A1(new_n388), .A2(new_n392), .ZN(new_n394));
  INV_X1    g193(.A(new_n387), .ZN(new_n395));
  OAI21_X1  g194(.A(new_n394), .B1(new_n395), .B2(new_n385), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n383), .A2(new_n384), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n397), .A2(KEYINPUT32), .ZN(new_n398));
  INV_X1    g197(.A(new_n398), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n393), .A2(new_n396), .A3(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(new_n400), .ZN(new_n401));
  AOI21_X1  g200(.A(new_n399), .B1(new_n393), .B2(new_n396), .ZN(new_n402));
  OAI21_X1  g201(.A(new_n382), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n393), .A2(new_n396), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n404), .A2(new_n398), .ZN(new_n405));
  NAND3_X1  g204(.A1(new_n405), .A2(KEYINPUT36), .A3(new_n400), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT88), .ZN(new_n408));
  AND3_X1   g207(.A1(new_n381), .A2(new_n407), .A3(new_n408), .ZN(new_n409));
  AOI21_X1  g208(.A(new_n408), .B1(new_n381), .B2(new_n407), .ZN(new_n410));
  OAI21_X1  g209(.A(new_n326), .B1(new_n320), .B2(new_n321), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n323), .A2(new_n281), .A3(new_n328), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(KEYINPUT37), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT38), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT37), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n266), .A2(new_n415), .ZN(new_n416));
  OAI211_X1 g215(.A(new_n413), .B(new_n414), .C1(new_n330), .C2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n415), .B1(new_n322), .B2(new_n329), .ZN(new_n418));
  INV_X1    g217(.A(new_n416), .ZN(new_n419));
  AOI21_X1  g218(.A(new_n418), .B1(new_n331), .B2(new_n419), .ZN(new_n420));
  OAI211_X1 g219(.A(new_n332), .B(new_n417), .C1(new_n420), .C2(new_n414), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT39), .B1(new_n241), .B2(new_n243), .ZN(new_n422));
  INV_X1    g221(.A(new_n422), .ZN(new_n423));
  AND2_X1   g222(.A1(new_n254), .A2(new_n251), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n423), .B1(new_n424), .B2(new_n242), .ZN(new_n425));
  AOI21_X1  g224(.A(new_n242), .B1(new_n254), .B2(new_n251), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT39), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n425), .A2(KEYINPUT40), .A3(new_n206), .A4(new_n428), .ZN(new_n429));
  XNOR2_X1  g228(.A(new_n429), .B(KEYINPUT89), .ZN(new_n430));
  INV_X1    g229(.A(KEYINPUT40), .ZN(new_n431));
  NAND2_X1  g230(.A1(new_n428), .A2(new_n206), .ZN(new_n432));
  NOR2_X1   g231(.A1(new_n426), .A2(new_n422), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n431), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND4_X1  g233(.A1(new_n333), .A2(new_n335), .A3(new_n434), .A4(new_n257), .ZN(new_n435));
  OAI22_X1  g234(.A1(new_n421), .A2(new_n263), .B1(new_n430), .B2(new_n435), .ZN(new_n436));
  INV_X1    g235(.A(new_n378), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n375), .A2(KEYINPUT86), .A3(new_n377), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g238(.A(new_n436), .B1(new_n439), .B2(new_n372), .ZN(new_n440));
  NOR3_X1   g239(.A1(new_n409), .A2(new_n410), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n405), .A2(new_n400), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n442), .B1(new_n439), .B2(new_n372), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT35), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n337), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n443), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(new_n372), .B1(new_n378), .B2(new_n380), .ZN(new_n447));
  INV_X1    g246(.A(KEYINPUT90), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n448), .B1(new_n401), .B2(new_n402), .ZN(new_n449));
  NAND3_X1  g248(.A1(new_n405), .A2(KEYINPUT90), .A3(new_n400), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n337), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n447), .A2(new_n451), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(new_n444), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n446), .A2(new_n454), .ZN(new_n455));
  OAI21_X1  g254(.A(new_n202), .B1(new_n441), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(new_n410), .ZN(new_n457));
  INV_X1    g256(.A(new_n440), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n381), .A2(new_n408), .A3(new_n407), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n457), .A2(new_n458), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g259(.A1(new_n443), .A2(new_n445), .B1(new_n453), .B2(new_n444), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n460), .A2(KEYINPUT91), .A3(new_n461), .ZN(new_n462));
  XNOR2_X1  g261(.A(G113gat), .B(G141gat), .ZN(new_n463));
  XNOR2_X1  g262(.A(new_n463), .B(G197gat), .ZN(new_n464));
  XOR2_X1   g263(.A(KEYINPUT11), .B(G169gat), .Z(new_n465));
  XNOR2_X1  g264(.A(new_n464), .B(new_n465), .ZN(new_n466));
  XNOR2_X1  g265(.A(new_n466), .B(KEYINPUT12), .ZN(new_n467));
  NAND2_X1  g266(.A1(G229gat), .A2(G233gat), .ZN(new_n468));
  XOR2_X1   g267(.A(new_n468), .B(KEYINPUT13), .Z(new_n469));
  INV_X1    g268(.A(new_n469), .ZN(new_n470));
  XNOR2_X1  g269(.A(G15gat), .B(G22gat), .ZN(new_n471));
  INV_X1    g270(.A(G1gat), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n472), .A2(KEYINPUT16), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n474), .B1(G1gat), .B2(new_n471), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n475), .A2(G8gat), .ZN(new_n476));
  INV_X1    g275(.A(G8gat), .ZN(new_n477));
  OAI211_X1 g276(.A(new_n474), .B(new_n477), .C1(G1gat), .C2(new_n471), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n476), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT94), .ZN(new_n480));
  INV_X1    g279(.A(G50gat), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n480), .B1(new_n481), .B2(G43gat), .ZN(new_n482));
  INV_X1    g281(.A(G43gat), .ZN(new_n483));
  NAND3_X1  g282(.A1(new_n483), .A2(KEYINPUT94), .A3(G50gat), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n481), .A2(G43gat), .ZN(new_n485));
  NAND3_X1  g284(.A1(new_n482), .A2(new_n484), .A3(new_n485), .ZN(new_n486));
  XOR2_X1   g285(.A(KEYINPUT93), .B(KEYINPUT15), .Z(new_n487));
  NAND2_X1  g286(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  OAI21_X1  g287(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT14), .ZN(new_n490));
  INV_X1    g289(.A(G29gat), .ZN(new_n491));
  INV_X1    g290(.A(G36gat), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n490), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(G29gat), .A2(G36gat), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  NAND3_X1  g295(.A1(KEYINPUT92), .A2(G29gat), .A3(G36gat), .ZN(new_n497));
  AOI22_X1  g296(.A1(new_n489), .A2(new_n493), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n483), .A2(G50gat), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n499), .A2(new_n485), .A3(KEYINPUT15), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n488), .A2(KEYINPUT95), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  OR2_X1    g300(.A1(new_n498), .A2(new_n500), .ZN(new_n502));
  NAND2_X1  g301(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n493), .A2(new_n489), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n496), .A2(new_n497), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT95), .B1(new_n506), .B2(new_n488), .ZN(new_n507));
  OAI21_X1  g306(.A(new_n479), .B1(new_n503), .B2(new_n507), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT97), .ZN(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT95), .ZN(new_n511));
  AND2_X1   g310(.A1(new_n486), .A2(new_n487), .ZN(new_n512));
  NAND3_X1  g311(.A1(new_n504), .A2(new_n500), .A3(new_n505), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n514), .A2(new_n502), .A3(new_n501), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n515), .A2(KEYINPUT97), .A3(new_n479), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n510), .A2(new_n516), .ZN(new_n517));
  NOR2_X1   g316(.A1(new_n503), .A2(new_n507), .ZN(new_n518));
  INV_X1    g317(.A(new_n479), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n470), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  AOI21_X1  g320(.A(new_n479), .B1(new_n518), .B2(KEYINPUT17), .ZN(new_n522));
  INV_X1    g321(.A(KEYINPUT96), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT17), .ZN(new_n524));
  OAI211_X1 g323(.A(new_n523), .B(new_n524), .C1(new_n503), .C2(new_n507), .ZN(new_n525));
  INV_X1    g324(.A(new_n525), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n523), .B1(new_n515), .B2(new_n524), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n522), .B1(new_n526), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n528), .A2(new_n468), .A3(new_n517), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT18), .ZN(new_n530));
  AOI21_X1  g329(.A(new_n521), .B1(new_n529), .B2(new_n530), .ZN(new_n531));
  NAND4_X1  g330(.A1(new_n528), .A2(KEYINPUT18), .A3(new_n468), .A4(new_n517), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n467), .B1(new_n531), .B2(new_n532), .ZN(new_n533));
  INV_X1    g332(.A(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n531), .A2(new_n467), .A3(new_n532), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  XOR2_X1   g335(.A(G134gat), .B(G162gat), .Z(new_n537));
  INV_X1    g336(.A(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT7), .ZN(new_n539));
  INV_X1    g338(.A(G85gat), .ZN(new_n540));
  OAI21_X1  g339(.A(G92gat), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G92gat), .ZN(new_n542));
  NAND3_X1  g341(.A1(new_n542), .A2(KEYINPUT7), .A3(G85gat), .ZN(new_n543));
  AOI22_X1  g342(.A1(new_n541), .A2(new_n543), .B1(new_n539), .B2(new_n540), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT8), .ZN(new_n545));
  NAND2_X1  g344(.A1(G99gat), .A2(G106gat), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n545), .B1(new_n546), .B2(KEYINPUT104), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n547), .B1(KEYINPUT104), .B2(new_n546), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n544), .A2(new_n548), .ZN(new_n549));
  XNOR2_X1  g348(.A(G99gat), .B(G106gat), .ZN(new_n550));
  INV_X1    g349(.A(new_n550), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n549), .B(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n552), .B1(new_n515), .B2(new_n524), .ZN(new_n553));
  OAI21_X1  g352(.A(KEYINPUT96), .B1(new_n518), .B2(KEYINPUT17), .ZN(new_n554));
  AOI21_X1  g353(.A(new_n553), .B1(new_n554), .B2(new_n525), .ZN(new_n555));
  XNOR2_X1  g354(.A(new_n549), .B(new_n550), .ZN(new_n556));
  AND2_X1   g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  AOI22_X1  g356(.A1(new_n515), .A2(new_n556), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  OAI21_X1  g358(.A(G190gat), .B1(new_n555), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g359(.A1(new_n526), .A2(new_n527), .ZN(new_n561));
  OAI211_X1 g360(.A(new_n291), .B(new_n558), .C1(new_n561), .C2(new_n553), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n560), .A2(new_n562), .ZN(new_n563));
  AOI21_X1  g362(.A(KEYINPUT103), .B1(new_n563), .B2(new_n270), .ZN(new_n564));
  NOR2_X1   g363(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n565));
  INV_X1    g364(.A(new_n565), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n560), .A2(G218gat), .A3(new_n562), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n566), .B1(new_n564), .B2(new_n567), .ZN(new_n569));
  OAI21_X1  g368(.A(new_n538), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(new_n209), .ZN(new_n572));
  OR2_X1    g371(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n573));
  NAND2_X1  g372(.A1(KEYINPUT100), .A2(G57gat), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n573), .A2(G64gat), .A3(new_n574), .ZN(new_n575));
  INV_X1    g374(.A(G64gat), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n576), .A2(G57gat), .ZN(new_n577));
  INV_X1    g376(.A(G71gat), .ZN(new_n578));
  INV_X1    g377(.A(G78gat), .ZN(new_n579));
  NOR2_X1   g378(.A1(new_n578), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(G71gat), .A2(G78gat), .ZN(new_n582));
  NAND2_X1  g381(.A1(new_n582), .A2(KEYINPUT9), .ZN(new_n583));
  AOI22_X1  g382(.A1(new_n575), .A2(new_n577), .B1(new_n581), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  XNOR2_X1  g384(.A(G57gat), .B(G64gat), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT9), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n581), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND2_X1  g387(.A1(new_n582), .A2(KEYINPUT98), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT98), .ZN(new_n590));
  OAI21_X1  g389(.A(new_n590), .B1(G71gat), .B2(G78gat), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT99), .ZN(new_n593));
  NOR3_X1   g392(.A1(new_n588), .A2(new_n592), .A3(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(G57gat), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(G64gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n577), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n580), .B1(new_n597), .B2(KEYINPUT9), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n589), .A2(new_n591), .ZN(new_n599));
  AOI21_X1  g398(.A(KEYINPUT99), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  OAI21_X1  g399(.A(new_n585), .B1(new_n594), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n593), .B1(new_n588), .B2(new_n592), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n598), .A2(KEYINPUT99), .A3(new_n599), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n606), .A2(KEYINPUT101), .A3(new_n585), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n603), .A2(new_n607), .ZN(new_n608));
  AOI21_X1  g407(.A(new_n479), .B1(new_n608), .B2(KEYINPUT21), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT102), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g411(.A1(new_n609), .A2(new_n610), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n572), .B1(new_n612), .B2(new_n613), .ZN(new_n614));
  INV_X1    g413(.A(new_n613), .ZN(new_n615));
  INV_X1    g414(.A(new_n572), .ZN(new_n616));
  NAND3_X1  g415(.A1(new_n615), .A2(new_n611), .A3(new_n616), .ZN(new_n617));
  NAND2_X1  g416(.A1(new_n614), .A2(new_n617), .ZN(new_n618));
  XNOR2_X1  g417(.A(G183gat), .B(G211gat), .ZN(new_n619));
  INV_X1    g418(.A(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(G127gat), .ZN(new_n621));
  OAI211_X1 g420(.A(G231gat), .B(G233gat), .C1(new_n608), .C2(KEYINPUT21), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(G231gat), .A2(G233gat), .ZN(new_n624));
  NAND4_X1  g423(.A1(new_n603), .A2(new_n623), .A3(new_n607), .A4(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n621), .B1(new_n622), .B2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n622), .A2(new_n621), .A3(new_n625), .ZN(new_n628));
  AOI21_X1  g427(.A(new_n620), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  INV_X1    g428(.A(new_n628), .ZN(new_n630));
  NOR3_X1   g429(.A1(new_n630), .A2(new_n626), .A3(new_n619), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n618), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  OAI21_X1  g431(.A(new_n619), .B1(new_n630), .B2(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n627), .A2(new_n620), .A3(new_n628), .ZN(new_n634));
  NAND4_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n617), .A4(new_n614), .ZN(new_n635));
  AND2_X1   g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(G176gat), .B(G204gat), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n637), .B(new_n638), .Z(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND2_X1  g439(.A1(G230gat), .A2(G233gat), .ZN(new_n641));
  XNOR2_X1  g440(.A(new_n641), .B(KEYINPUT106), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT10), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n556), .B1(new_n603), .B2(new_n607), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n556), .A2(new_n601), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n643), .B1(new_n644), .B2(new_n646), .ZN(new_n647));
  NOR2_X1   g446(.A1(new_n552), .A2(new_n643), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n608), .A2(new_n648), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n642), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  NOR3_X1   g449(.A1(new_n644), .A2(new_n641), .A3(new_n646), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n640), .B1(new_n650), .B2(new_n651), .ZN(new_n652));
  INV_X1    g451(.A(KEYINPUT107), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  OAI211_X1 g453(.A(KEYINPUT107), .B(new_n640), .C1(new_n650), .C2(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT105), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n640), .B1(new_n651), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT101), .B1(new_n606), .B2(new_n585), .ZN(new_n659));
  AOI211_X1 g458(.A(new_n602), .B(new_n584), .C1(new_n604), .C2(new_n605), .ZN(new_n660));
  OAI21_X1  g459(.A(new_n552), .B1(new_n659), .B2(new_n660), .ZN(new_n661));
  AOI21_X1  g460(.A(KEYINPUT10), .B1(new_n661), .B2(new_n645), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n608), .A2(new_n648), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n641), .B1(new_n662), .B2(new_n663), .ZN(new_n664));
  OAI211_X1 g463(.A(new_n658), .B(new_n664), .C1(new_n657), .C2(new_n651), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n656), .A2(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(new_n666), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n563), .A2(new_n270), .ZN(new_n668));
  INV_X1    g467(.A(KEYINPUT103), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n668), .A2(new_n669), .A3(new_n567), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n670), .A2(new_n565), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n564), .A2(new_n566), .A3(new_n567), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n671), .A2(new_n537), .A3(new_n672), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n570), .A2(new_n636), .A3(new_n667), .A4(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g474(.A1(new_n456), .A2(new_n462), .A3(new_n536), .A4(new_n675), .ZN(new_n676));
  OR3_X1    g475(.A1(new_n676), .A2(KEYINPUT109), .A3(new_n263), .ZN(new_n677));
  OAI21_X1  g476(.A(KEYINPUT109), .B1(new_n676), .B2(new_n263), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n677), .A2(new_n678), .ZN(new_n679));
  XNOR2_X1  g478(.A(KEYINPUT108), .B(G1gat), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n679), .B(new_n680), .ZN(G1324gat));
  NOR2_X1   g480(.A1(new_n676), .A2(new_n336), .ZN(new_n682));
  XOR2_X1   g481(.A(KEYINPUT16), .B(G8gat), .Z(new_n683));
  NAND2_X1  g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n684), .B1(new_n477), .B2(new_n682), .ZN(new_n685));
  MUX2_X1   g484(.A(new_n684), .B(new_n685), .S(KEYINPUT42), .Z(G1325gat));
  OAI21_X1  g485(.A(G15gat), .B1(new_n676), .B2(new_n407), .ZN(new_n687));
  INV_X1    g486(.A(new_n451), .ZN(new_n688));
  OR2_X1    g487(.A1(new_n688), .A2(G15gat), .ZN(new_n689));
  OAI21_X1  g488(.A(new_n687), .B1(new_n676), .B2(new_n689), .ZN(G1326gat));
  NOR2_X1   g489(.A1(new_n676), .A2(new_n447), .ZN(new_n691));
  XOR2_X1   g490(.A(KEYINPUT43), .B(G22gat), .Z(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1327gat));
  NAND2_X1  g492(.A1(new_n570), .A2(new_n673), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  NOR2_X1   g495(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n456), .A2(new_n462), .A3(new_n697), .ZN(new_n698));
  NAND2_X1  g497(.A1(new_n381), .A2(new_n407), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n446), .B(new_n454), .C1(new_n699), .C2(new_n440), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n700), .A2(new_n694), .ZN(new_n701));
  NAND2_X1  g500(.A1(new_n701), .A2(new_n696), .ZN(new_n702));
  AND2_X1   g501(.A1(new_n698), .A2(new_n702), .ZN(new_n703));
  INV_X1    g502(.A(new_n536), .ZN(new_n704));
  NOR3_X1   g503(.A1(new_n636), .A2(new_n704), .A3(new_n666), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n703), .A2(new_n705), .ZN(new_n706));
  OAI21_X1  g505(.A(G29gat), .B1(new_n706), .B2(new_n263), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT45), .ZN(new_n708));
  NOR3_X1   g507(.A1(new_n695), .A2(new_n636), .A3(new_n666), .ZN(new_n709));
  NAND4_X1  g508(.A1(new_n456), .A2(new_n462), .A3(new_n536), .A4(new_n709), .ZN(new_n710));
  INV_X1    g509(.A(new_n263), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n491), .ZN(new_n712));
  OAI21_X1  g511(.A(new_n708), .B1(new_n710), .B2(new_n712), .ZN(new_n713));
  OR3_X1    g512(.A1(new_n710), .A2(new_n708), .A3(new_n712), .ZN(new_n714));
  NAND3_X1  g513(.A1(new_n707), .A2(new_n713), .A3(new_n714), .ZN(G1328gat));
  OAI21_X1  g514(.A(G36gat), .B1(new_n706), .B2(new_n336), .ZN(new_n716));
  INV_X1    g515(.A(new_n710), .ZN(new_n717));
  INV_X1    g516(.A(new_n336), .ZN(new_n718));
  NAND2_X1  g517(.A1(KEYINPUT110), .A2(KEYINPUT46), .ZN(new_n719));
  NAND4_X1  g518(.A1(new_n717), .A2(new_n492), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  XNOR2_X1  g519(.A(KEYINPUT110), .B(KEYINPUT46), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n718), .A2(new_n492), .ZN(new_n722));
  OAI21_X1  g521(.A(new_n721), .B1(new_n710), .B2(new_n722), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n716), .A2(new_n720), .A3(new_n723), .ZN(G1329gat));
  NOR2_X1   g523(.A1(new_n688), .A2(G43gat), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT47), .ZN(new_n726));
  AOI22_X1  g525(.A1(new_n717), .A2(new_n725), .B1(KEYINPUT111), .B2(new_n726), .ZN(new_n727));
  INV_X1    g526(.A(new_n407), .ZN(new_n728));
  NAND4_X1  g527(.A1(new_n698), .A2(new_n728), .A3(new_n702), .A4(new_n705), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(G43gat), .ZN(new_n730));
  NAND2_X1  g529(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  OR2_X1    g530(.A1(new_n726), .A2(KEYINPUT111), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n731), .B(new_n732), .ZN(G1330gat));
  INV_X1    g532(.A(new_n447), .ZN(new_n734));
  NAND2_X1  g533(.A1(new_n734), .A2(new_n481), .ZN(new_n735));
  XOR2_X1   g534(.A(new_n735), .B(KEYINPUT112), .Z(new_n736));
  NOR2_X1   g535(.A1(new_n710), .A2(new_n736), .ZN(new_n737));
  NAND4_X1  g536(.A1(new_n698), .A2(new_n734), .A3(new_n702), .A4(new_n705), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n737), .B1(G50gat), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(KEYINPUT113), .ZN(new_n740));
  AOI21_X1  g539(.A(new_n740), .B1(new_n738), .B2(G50gat), .ZN(new_n741));
  INV_X1    g540(.A(KEYINPUT48), .ZN(new_n742));
  NOR3_X1   g541(.A1(new_n739), .A2(new_n741), .A3(new_n742), .ZN(new_n743));
  AOI221_X4 g542(.A(new_n737), .B1(new_n740), .B2(KEYINPUT48), .C1(G50gat), .C2(new_n738), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n743), .A2(new_n744), .ZN(G1331gat));
  AND3_X1   g544(.A1(new_n570), .A2(new_n636), .A3(new_n673), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n704), .A3(new_n666), .ZN(new_n747));
  XOR2_X1   g546(.A(new_n747), .B(KEYINPUT114), .Z(new_n748));
  NAND2_X1  g547(.A1(new_n700), .A2(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(new_n711), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n573), .A2(new_n574), .ZN(new_n752));
  XNOR2_X1  g551(.A(new_n751), .B(new_n752), .ZN(G1332gat));
  NOR2_X1   g552(.A1(new_n749), .A2(new_n336), .ZN(new_n754));
  NOR2_X1   g553(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n755));
  AND2_X1   g554(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n756));
  OAI21_X1  g555(.A(new_n754), .B1(new_n755), .B2(new_n756), .ZN(new_n757));
  OAI21_X1  g556(.A(new_n757), .B1(new_n754), .B2(new_n755), .ZN(G1333gat));
  NOR3_X1   g557(.A1(new_n749), .A2(G71gat), .A3(new_n688), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n750), .A2(new_n728), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n759), .B1(G71gat), .B2(new_n760), .ZN(new_n761));
  XNOR2_X1  g560(.A(new_n761), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g561(.A1(new_n749), .A2(new_n447), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n763), .B(new_n579), .ZN(G1335gat));
  NOR2_X1   g563(.A1(new_n636), .A2(new_n536), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n765), .A2(new_n666), .ZN(new_n766));
  XOR2_X1   g565(.A(new_n766), .B(KEYINPUT115), .Z(new_n767));
  NAND2_X1  g566(.A1(new_n703), .A2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(G85gat), .B1(new_n768), .B2(new_n263), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n700), .A2(new_n694), .A3(new_n765), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT51), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g571(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n694), .A4(new_n765), .ZN(new_n773));
  AOI21_X1  g572(.A(new_n667), .B1(new_n772), .B2(new_n773), .ZN(new_n774));
  NAND3_X1  g573(.A1(new_n774), .A2(new_n540), .A3(new_n711), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n769), .A2(new_n775), .ZN(G1336gat));
  NAND3_X1  g575(.A1(new_n774), .A2(new_n542), .A3(new_n718), .ZN(new_n777));
  NAND4_X1  g576(.A1(new_n698), .A2(new_n718), .A3(new_n702), .A4(new_n767), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G92gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(new_n780));
  XNOR2_X1  g579(.A(new_n780), .B(KEYINPUT52), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n768), .A2(new_n782), .A3(new_n407), .ZN(new_n783));
  AOI21_X1  g582(.A(G99gat), .B1(new_n774), .B2(new_n451), .ZN(new_n784));
  NOR2_X1   g583(.A1(new_n783), .A2(new_n784), .ZN(G1338gat));
  NOR2_X1   g584(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n786));
  AND2_X1   g585(.A1(KEYINPUT116), .A2(KEYINPUT53), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n698), .A2(new_n734), .A3(new_n702), .A4(new_n767), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n788), .A2(G106gat), .ZN(new_n789));
  OR2_X1    g588(.A1(new_n447), .A2(G106gat), .ZN(new_n790));
  INV_X1    g589(.A(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n774), .A2(new_n791), .ZN(new_n792));
  AOI211_X1 g591(.A(new_n786), .B(new_n787), .C1(new_n789), .C2(new_n792), .ZN(new_n793));
  AND4_X1   g592(.A1(KEYINPUT116), .A2(new_n789), .A3(new_n792), .A4(KEYINPUT53), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n793), .A2(new_n794), .ZN(G1339gat));
  AOI21_X1  g594(.A(new_n468), .B1(new_n528), .B2(new_n517), .ZN(new_n796));
  AND2_X1   g595(.A1(new_n796), .A2(KEYINPUT118), .ZN(new_n797));
  NAND3_X1  g596(.A1(new_n517), .A2(new_n520), .A3(new_n470), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n798), .B1(new_n796), .B2(KEYINPUT118), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n466), .B1(new_n797), .B2(new_n799), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n535), .ZN(new_n801));
  NAND3_X1  g600(.A1(new_n647), .A2(new_n649), .A3(new_n642), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n664), .A2(new_n802), .A3(KEYINPUT54), .ZN(new_n803));
  INV_X1    g602(.A(KEYINPUT54), .ZN(new_n804));
  INV_X1    g603(.A(new_n642), .ZN(new_n805));
  OAI211_X1 g604(.A(new_n804), .B(new_n805), .C1(new_n662), .C2(new_n663), .ZN(new_n806));
  NAND4_X1  g605(.A1(new_n803), .A2(KEYINPUT55), .A3(new_n640), .A4(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n807), .A2(new_n665), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n639), .B1(new_n650), .B2(new_n804), .ZN(new_n809));
  AOI21_X1  g608(.A(KEYINPUT55), .B1(new_n809), .B2(new_n803), .ZN(new_n810));
  NOR3_X1   g609(.A1(new_n801), .A2(new_n808), .A3(new_n810), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n694), .A2(new_n811), .ZN(new_n812));
  AND3_X1   g611(.A1(new_n531), .A2(new_n467), .A3(new_n532), .ZN(new_n813));
  OAI211_X1 g612(.A(new_n807), .B(new_n665), .C1(new_n813), .C2(new_n533), .ZN(new_n814));
  NOR2_X1   g613(.A1(new_n814), .A2(new_n810), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n801), .B1(new_n665), .B2(new_n656), .ZN(new_n816));
  NOR2_X1   g615(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n812), .B1(new_n817), .B2(new_n694), .ZN(new_n818));
  INV_X1    g617(.A(new_n636), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT117), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n746), .A2(new_n821), .A3(new_n704), .A4(new_n667), .ZN(new_n822));
  OAI21_X1  g621(.A(KEYINPUT117), .B1(new_n674), .B2(new_n536), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n822), .A2(new_n823), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n820), .A2(new_n824), .ZN(new_n825));
  INV_X1    g624(.A(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n826), .A2(new_n263), .ZN(new_n827));
  AND3_X1   g626(.A1(new_n827), .A2(new_n336), .A3(new_n443), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n828), .A2(new_n233), .A3(new_n536), .ZN(new_n829));
  NOR2_X1   g628(.A1(new_n734), .A2(new_n688), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n825), .A2(new_n830), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n831), .A2(new_n711), .A3(new_n336), .ZN(new_n832));
  OAI21_X1  g631(.A(G113gat), .B1(new_n832), .B2(new_n704), .ZN(new_n833));
  NAND2_X1  g632(.A1(new_n829), .A2(new_n833), .ZN(G1340gat));
  NOR3_X1   g633(.A1(new_n832), .A2(new_n235), .A3(new_n667), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n828), .A2(new_n666), .ZN(new_n836));
  AOI21_X1  g635(.A(new_n835), .B1(new_n836), .B2(new_n235), .ZN(G1341gat));
  NAND3_X1  g636(.A1(new_n828), .A2(new_n621), .A3(new_n636), .ZN(new_n838));
  OAI21_X1  g637(.A(G127gat), .B1(new_n832), .B2(new_n819), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n838), .A2(new_n839), .ZN(G1342gat));
  INV_X1    g639(.A(G134gat), .ZN(new_n841));
  NAND3_X1  g640(.A1(new_n828), .A2(new_n841), .A3(new_n694), .ZN(new_n842));
  OR2_X1    g641(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n843));
  OAI21_X1  g642(.A(G134gat), .B1(new_n832), .B2(new_n695), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n842), .A2(KEYINPUT56), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(G1343gat));
  NAND2_X1  g645(.A1(new_n734), .A2(new_n407), .ZN(new_n847));
  NOR2_X1   g646(.A1(new_n847), .A2(new_n718), .ZN(new_n848));
  NAND2_X1  g647(.A1(new_n827), .A2(new_n848), .ZN(new_n849));
  NOR3_X1   g648(.A1(new_n849), .A2(G141gat), .A3(new_n704), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n263), .B(new_n718), .C1(new_n403), .C2(new_n406), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(KEYINPUT119), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n852), .A2(new_n853), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT57), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n855), .B1(new_n826), .B2(new_n447), .ZN(new_n856));
  INV_X1    g655(.A(new_n824), .ZN(new_n857));
  NAND2_X1  g656(.A1(new_n809), .A2(new_n803), .ZN(new_n858));
  INV_X1    g657(.A(KEYINPUT55), .ZN(new_n859));
  AOI21_X1  g658(.A(KEYINPUT120), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT120), .ZN(new_n861));
  AOI211_X1 g660(.A(new_n861), .B(KEYINPUT55), .C1(new_n809), .C2(new_n803), .ZN(new_n862));
  NOR3_X1   g661(.A1(new_n814), .A2(new_n860), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(KEYINPUT121), .B1(new_n863), .B2(new_n816), .ZN(new_n864));
  INV_X1    g663(.A(new_n801), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n666), .ZN(new_n866));
  INV_X1    g665(.A(KEYINPUT121), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n858), .A2(new_n859), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n868), .A2(new_n861), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n810), .A2(KEYINPUT120), .ZN(new_n870));
  NAND2_X1  g669(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  OAI211_X1 g670(.A(new_n866), .B(new_n867), .C1(new_n871), .C2(new_n814), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n864), .A2(new_n695), .A3(new_n872), .ZN(new_n873));
  AOI21_X1  g672(.A(new_n636), .B1(new_n873), .B2(new_n812), .ZN(new_n874));
  OAI211_X1 g673(.A(KEYINPUT57), .B(new_n734), .C1(new_n857), .C2(new_n874), .ZN(new_n875));
  AOI21_X1  g674(.A(new_n854), .B1(new_n856), .B2(new_n875), .ZN(new_n876));
  NAND2_X1  g675(.A1(new_n876), .A2(new_n536), .ZN(new_n877));
  AOI21_X1  g676(.A(new_n850), .B1(G141gat), .B2(new_n877), .ZN(new_n878));
  XOR2_X1   g677(.A(new_n878), .B(KEYINPUT58), .Z(G1344gat));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n880));
  NOR2_X1   g679(.A1(new_n214), .A2(KEYINPUT59), .ZN(new_n881));
  INV_X1    g680(.A(new_n881), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(new_n876), .B2(new_n666), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n734), .A2(KEYINPUT57), .ZN(new_n884));
  AOI21_X1  g683(.A(new_n884), .B1(new_n820), .B2(new_n824), .ZN(new_n885));
  NOR2_X1   g684(.A1(new_n674), .A2(new_n536), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n734), .B1(new_n874), .B2(new_n886), .ZN(new_n887));
  AOI21_X1  g686(.A(new_n885), .B1(new_n887), .B2(new_n855), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n852), .A2(new_n666), .A3(new_n853), .ZN(new_n889));
  OAI21_X1  g688(.A(G148gat), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT59), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT122), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT122), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT59), .ZN(new_n894));
  AOI21_X1  g693(.A(new_n883), .B1(new_n892), .B2(new_n894), .ZN(new_n895));
  NOR3_X1   g694(.A1(new_n849), .A2(G148gat), .A3(new_n667), .ZN(new_n896));
  OAI21_X1  g695(.A(new_n880), .B1(new_n895), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(new_n896), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n890), .A2(new_n893), .A3(KEYINPUT59), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n893), .B1(new_n890), .B2(KEYINPUT59), .ZN(new_n900));
  NOR2_X1   g699(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  OAI211_X1 g700(.A(KEYINPUT123), .B(new_n898), .C1(new_n901), .C2(new_n883), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n897), .A2(new_n902), .ZN(G1345gat));
  INV_X1    g702(.A(new_n849), .ZN(new_n904));
  AOI21_X1  g703(.A(G155gat), .B1(new_n904), .B2(new_n636), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n636), .A2(G155gat), .ZN(new_n906));
  XNOR2_X1  g705(.A(new_n906), .B(KEYINPUT124), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n905), .B1(new_n876), .B2(new_n907), .ZN(G1346gat));
  NAND3_X1  g707(.A1(new_n904), .A2(new_n210), .A3(new_n694), .ZN(new_n909));
  AND2_X1   g708(.A1(new_n876), .A2(new_n694), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n910), .B2(new_n210), .ZN(G1347gat));
  AOI21_X1  g710(.A(new_n711), .B1(new_n820), .B2(new_n824), .ZN(new_n912));
  AND3_X1   g711(.A1(new_n912), .A2(new_n718), .A3(new_n443), .ZN(new_n913));
  AOI21_X1  g712(.A(G169gat), .B1(new_n913), .B2(new_n536), .ZN(new_n914));
  NOR2_X1   g713(.A1(new_n711), .A2(new_n336), .ZN(new_n915));
  AND2_X1   g714(.A1(new_n831), .A2(new_n915), .ZN(new_n916));
  AND2_X1   g715(.A1(new_n536), .A2(G169gat), .ZN(new_n917));
  AOI21_X1  g716(.A(new_n914), .B1(new_n916), .B2(new_n917), .ZN(G1348gat));
  NOR3_X1   g717(.A1(new_n667), .A2(new_n336), .A3(G176gat), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n912), .A2(new_n443), .A3(new_n919), .ZN(new_n920));
  AND2_X1   g719(.A1(new_n916), .A2(new_n666), .ZN(new_n921));
  INV_X1    g720(.A(G176gat), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n920), .B1(new_n921), .B2(new_n922), .ZN(G1349gat));
  NAND4_X1  g722(.A1(new_n825), .A2(new_n830), .A3(new_n636), .A4(new_n915), .ZN(new_n924));
  OR2_X1    g723(.A1(new_n924), .A2(KEYINPUT125), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n287), .B1(new_n924), .B2(KEYINPUT125), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n913), .A2(new_n308), .A3(new_n636), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n927), .A2(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(KEYINPUT127), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT127), .ZN(new_n931));
  NAND3_X1  g730(.A1(new_n927), .A2(new_n931), .A3(new_n928), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g732(.A(KEYINPUT60), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n934), .A2(KEYINPUT126), .ZN(new_n935));
  XNOR2_X1  g734(.A(new_n933), .B(new_n935), .ZN(G1350gat));
  AOI21_X1  g735(.A(new_n291), .B1(new_n916), .B2(new_n694), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT61), .Z(new_n938));
  NAND3_X1  g737(.A1(new_n913), .A2(new_n286), .A3(new_n694), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n938), .A2(new_n939), .ZN(G1351gat));
  NAND3_X1  g739(.A1(new_n912), .A2(new_n734), .A3(new_n407), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n941), .A2(new_n336), .ZN(new_n942));
  AOI21_X1  g741(.A(G197gat), .B1(new_n942), .B2(new_n536), .ZN(new_n943));
  NOR4_X1   g742(.A1(new_n888), .A2(new_n711), .A3(new_n336), .A4(new_n728), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n536), .A2(G197gat), .ZN(new_n945));
  AOI21_X1  g744(.A(new_n943), .B1(new_n944), .B2(new_n945), .ZN(G1352gat));
  NOR4_X1   g745(.A1(new_n941), .A2(G204gat), .A3(new_n336), .A4(new_n667), .ZN(new_n947));
  XNOR2_X1  g746(.A(new_n947), .B(KEYINPUT62), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n944), .A2(new_n666), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(G204gat), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n948), .A2(new_n950), .ZN(G1353gat));
  NAND3_X1  g750(.A1(new_n942), .A2(new_n269), .A3(new_n636), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n944), .A2(new_n636), .ZN(new_n953));
  AND3_X1   g752(.A1(new_n953), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n954));
  AOI21_X1  g753(.A(KEYINPUT63), .B1(new_n953), .B2(G211gat), .ZN(new_n955));
  OAI21_X1  g754(.A(new_n952), .B1(new_n954), .B2(new_n955), .ZN(G1354gat));
  NAND3_X1  g755(.A1(new_n942), .A2(new_n270), .A3(new_n694), .ZN(new_n957));
  AND2_X1   g756(.A1(new_n944), .A2(new_n694), .ZN(new_n958));
  OAI21_X1  g757(.A(new_n957), .B1(new_n958), .B2(new_n270), .ZN(G1355gat));
endmodule


