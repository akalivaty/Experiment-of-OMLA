//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0 1 0 1 0 0 0 1 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 0 1 0 1 1 0 0 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:24 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n454, new_n458,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n555, new_n556, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n583, new_n584, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n609, new_n611, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n855, new_n856,
    new_n857, new_n858, new_n859, new_n860, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n866, new_n868, new_n869, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1209, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1216, new_n1217, new_n1218,
    new_n1219, new_n1220, new_n1221, new_n1222, new_n1223, new_n1224,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  INV_X1    g026(.A(new_n451), .ZN(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n453));
  INV_X1    g028(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g029(.A1(new_n452), .A2(new_n454), .ZN(G325));
  INV_X1    g030(.A(G325), .ZN(G261));
  AOI22_X1  g031(.A1(new_n452), .A2(G2106), .B1(G567), .B2(new_n454), .ZN(G319));
  INV_X1    g032(.A(G125), .ZN(new_n458));
  OR2_X1    g033(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n459));
  NAND2_X1  g034(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n460));
  AOI21_X1  g035(.A(new_n458), .B1(new_n459), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT65), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT65), .ZN(new_n464));
  NAND3_X1  g039(.A1(new_n464), .A2(G113), .A3(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g041(.A(G2105), .B1(new_n461), .B2(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(G2105), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  INV_X1    g044(.A(G101), .ZN(new_n470));
  NOR2_X1   g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n459), .B2(new_n460), .ZN(new_n472));
  AOI21_X1  g047(.A(new_n471), .B1(new_n472), .B2(G137), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n467), .A2(new_n473), .ZN(new_n474));
  INV_X1    g049(.A(new_n474), .ZN(G160));
  AOI21_X1  g050(.A(new_n468), .B1(new_n459), .B2(new_n460), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n476), .A2(G124), .ZN(new_n477));
  OR2_X1    g052(.A1(G100), .A2(G2105), .ZN(new_n478));
  OAI211_X1 g053(.A(new_n478), .B(G2104), .C1(G112), .C2(new_n468), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n477), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g055(.A(new_n480), .B1(G136), .B2(new_n472), .ZN(G162));
  INV_X1    g056(.A(KEYINPUT66), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n482), .B1(new_n468), .B2(G114), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n484), .A2(KEYINPUT66), .A3(G2105), .ZN(new_n485));
  INV_X1    g060(.A(G102), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(new_n468), .ZN(new_n487));
  NAND4_X1  g062(.A1(new_n483), .A2(new_n485), .A3(G2104), .A4(new_n487), .ZN(new_n488));
  AND2_X1   g063(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n489));
  NOR2_X1   g064(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n490));
  OAI211_X1 g065(.A(G126), .B(G2105), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n488), .A2(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI21_X1  g069(.A(new_n494), .B1(new_n489), .B2(new_n490), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(KEYINPUT4), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  OAI211_X1 g072(.A(new_n494), .B(new_n497), .C1(new_n490), .C2(new_n489), .ZN(new_n498));
  AOI21_X1  g073(.A(new_n492), .B1(new_n496), .B2(new_n498), .ZN(G164));
  XNOR2_X1  g074(.A(KEYINPUT6), .B(G651), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n500), .A2(G543), .ZN(new_n501));
  INV_X1    g076(.A(G50), .ZN(new_n502));
  NOR2_X1   g077(.A1(KEYINPUT5), .A2(G543), .ZN(new_n503));
  AND2_X1   g078(.A1(KEYINPUT5), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(KEYINPUT6), .A2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  OAI22_X1  g081(.A1(new_n503), .A2(new_n504), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g082(.A(G88), .ZN(new_n508));
  OAI22_X1  g083(.A1(new_n501), .A2(new_n502), .B1(new_n507), .B2(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G651), .ZN(new_n510));
  INV_X1    g085(.A(KEYINPUT5), .ZN(new_n511));
  INV_X1    g086(.A(G543), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(KEYINPUT5), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n515), .A2(G62), .ZN(new_n516));
  NAND2_X1  g091(.A1(G75), .A2(G543), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT67), .ZN(new_n518));
  XNOR2_X1  g093(.A(new_n517), .B(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n510), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  OR2_X1    g095(.A1(new_n509), .A2(new_n520), .ZN(G303));
  INV_X1    g096(.A(G303), .ZN(G166));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  XNOR2_X1  g098(.A(new_n523), .B(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(G51), .ZN(new_n525));
  OAI21_X1  g100(.A(new_n524), .B1(new_n501), .B2(new_n525), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n504), .A2(new_n503), .ZN(new_n527));
  NAND2_X1  g102(.A1(new_n500), .A2(G89), .ZN(new_n528));
  NAND2_X1  g103(.A1(G63), .A2(G651), .ZN(new_n529));
  AOI21_X1  g104(.A(new_n527), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n526), .A2(new_n530), .ZN(G168));
  AOI22_X1  g106(.A1(new_n515), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n532), .A2(new_n510), .ZN(new_n533));
  INV_X1    g108(.A(G52), .ZN(new_n534));
  INV_X1    g109(.A(G90), .ZN(new_n535));
  OAI22_X1  g110(.A1(new_n501), .A2(new_n534), .B1(new_n507), .B2(new_n535), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n533), .A2(new_n536), .ZN(G171));
  NAND2_X1  g112(.A1(G68), .A2(G543), .ZN(new_n538));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  OAI21_X1  g114(.A(new_n538), .B1(new_n527), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n540), .A2(G651), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT68), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(new_n507), .ZN(new_n544));
  NOR2_X1   g119(.A1(new_n505), .A2(new_n506), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n545), .A2(new_n512), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n544), .A2(G81), .B1(new_n546), .B2(G43), .ZN(new_n547));
  AND2_X1   g122(.A1(new_n543), .A2(new_n547), .ZN(new_n548));
  NOR2_X1   g123(.A1(new_n541), .A2(new_n542), .ZN(new_n549));
  INV_X1    g124(.A(new_n549), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n552), .A2(G860), .ZN(G153));
  NAND4_X1  g128(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND4_X1  g131(.A1(G319), .A2(G483), .A3(G661), .A4(new_n556), .ZN(G188));
  NAND3_X1  g132(.A1(new_n500), .A2(G53), .A3(G543), .ZN(new_n558));
  INV_X1    g133(.A(KEYINPUT9), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(G78), .A2(G543), .ZN(new_n561));
  INV_X1    g136(.A(G65), .ZN(new_n562));
  OAI21_X1  g137(.A(new_n561), .B1(new_n527), .B2(new_n562), .ZN(new_n563));
  NAND2_X1  g138(.A1(new_n563), .A2(G651), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n544), .A2(G91), .ZN(new_n565));
  NAND2_X1  g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NOR2_X1   g141(.A1(new_n560), .A2(new_n566), .ZN(new_n567));
  INV_X1    g142(.A(new_n567), .ZN(G299));
  INV_X1    g143(.A(G171), .ZN(G301));
  INV_X1    g144(.A(G168), .ZN(G286));
  OAI21_X1  g145(.A(G651), .B1(new_n515), .B2(G74), .ZN(new_n571));
  INV_X1    g146(.A(G87), .ZN(new_n572));
  INV_X1    g147(.A(G49), .ZN(new_n573));
  OAI221_X1 g148(.A(new_n571), .B1(new_n507), .B2(new_n572), .C1(new_n573), .C2(new_n501), .ZN(G288));
  OAI211_X1 g149(.A(G48), .B(G543), .C1(new_n505), .C2(new_n506), .ZN(new_n575));
  INV_X1    g150(.A(G86), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n507), .B2(new_n576), .ZN(new_n577));
  OAI21_X1  g152(.A(G61), .B1(new_n504), .B2(new_n503), .ZN(new_n578));
  NAND2_X1  g153(.A1(G73), .A2(G543), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n510), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  NOR2_X1   g155(.A1(new_n577), .A2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G305));
  AOI22_X1  g157(.A1(new_n544), .A2(G85), .B1(new_n546), .B2(G47), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n515), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n584));
  OAI21_X1  g159(.A(new_n583), .B1(new_n510), .B2(new_n584), .ZN(G290));
  NAND2_X1  g160(.A1(G301), .A2(G868), .ZN(new_n586));
  INV_X1    g161(.A(KEYINPUT69), .ZN(new_n587));
  OR2_X1    g162(.A1(new_n587), .A2(G66), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(G66), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n515), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(G79), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n590), .B1(new_n591), .B2(new_n512), .ZN(new_n592));
  INV_X1    g167(.A(KEYINPUT70), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  OAI211_X1 g169(.A(new_n590), .B(KEYINPUT70), .C1(new_n591), .C2(new_n512), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n594), .A2(G651), .A3(new_n595), .ZN(new_n596));
  NAND3_X1  g171(.A1(new_n544), .A2(KEYINPUT10), .A3(G92), .ZN(new_n597));
  INV_X1    g172(.A(KEYINPUT10), .ZN(new_n598));
  INV_X1    g173(.A(G92), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n598), .B1(new_n507), .B2(new_n599), .ZN(new_n600));
  AOI22_X1  g175(.A1(new_n597), .A2(new_n600), .B1(G54), .B2(new_n546), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n596), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n586), .B1(new_n603), .B2(G868), .ZN(G284));
  OAI21_X1  g179(.A(new_n586), .B1(new_n603), .B2(G868), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  OAI21_X1  g181(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G297));
  OAI21_X1  g182(.A(new_n606), .B1(new_n567), .B2(G868), .ZN(G280));
  INV_X1    g183(.A(G559), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n603), .B1(new_n609), .B2(G860), .ZN(G148));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n551), .A2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n602), .A2(G559), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n612), .B1(new_n613), .B2(new_n611), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT71), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  XNOR2_X1  g191(.A(KEYINPUT3), .B(G2104), .ZN(new_n617));
  INV_X1    g192(.A(new_n469), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n619), .B(KEYINPUT12), .ZN(new_n620));
  XNOR2_X1  g195(.A(new_n620), .B(KEYINPUT13), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2100), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n472), .A2(G135), .ZN(new_n623));
  NAND2_X1  g198(.A1(new_n476), .A2(G123), .ZN(new_n624));
  NOR2_X1   g199(.A1(new_n468), .A2(G111), .ZN(new_n625));
  OAI21_X1  g200(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n626));
  OAI211_X1 g201(.A(new_n623), .B(new_n624), .C1(new_n625), .C2(new_n626), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT72), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2096), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n622), .A2(new_n629), .ZN(G156));
  INV_X1    g205(.A(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2427), .B(G2438), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(G2430), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT15), .B(G2435), .ZN(new_n634));
  AOI21_X1  g209(.A(new_n631), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  OAI21_X1  g210(.A(new_n635), .B1(new_n634), .B2(new_n633), .ZN(new_n636));
  XNOR2_X1  g211(.A(G2451), .B(G2454), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(KEYINPUT16), .ZN(new_n638));
  XOR2_X1   g213(.A(G1341), .B(G1348), .Z(new_n639));
  XNOR2_X1  g214(.A(new_n638), .B(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n636), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2443), .B(G2446), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(new_n643));
  AND2_X1   g218(.A1(new_n641), .A2(new_n643), .ZN(new_n644));
  OAI21_X1  g219(.A(G14), .B1(new_n641), .B2(new_n643), .ZN(new_n645));
  NOR2_X1   g220(.A1(new_n644), .A2(new_n645), .ZN(G401));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  XNOR2_X1  g222(.A(G2072), .B(G2078), .ZN(new_n648));
  XNOR2_X1  g223(.A(G2067), .B(G2678), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n648), .A3(new_n649), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT73), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n651), .B(KEYINPUT18), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(KEYINPUT74), .ZN(new_n653));
  INV_X1    g228(.A(new_n648), .ZN(new_n654));
  NAND2_X1  g229(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g230(.A(new_n647), .ZN(new_n656));
  XOR2_X1   g231(.A(KEYINPUT75), .B(KEYINPUT17), .Z(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(new_n648), .ZN(new_n658));
  OAI211_X1 g233(.A(new_n655), .B(new_n656), .C1(new_n653), .C2(new_n658), .ZN(new_n659));
  NAND3_X1  g234(.A1(new_n658), .A2(new_n647), .A3(new_n653), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n652), .A2(new_n659), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2096), .B(G2100), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g238(.A1(new_n661), .A2(new_n663), .ZN(new_n664));
  NAND4_X1  g239(.A1(new_n652), .A2(new_n659), .A3(new_n660), .A4(new_n662), .ZN(new_n665));
  NAND2_X1  g240(.A1(new_n664), .A2(new_n665), .ZN(G227));
  XNOR2_X1  g241(.A(G1981), .B(G1986), .ZN(new_n667));
  INV_X1    g242(.A(new_n667), .ZN(new_n668));
  XNOR2_X1  g243(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1971), .B(G1976), .ZN(new_n671));
  INV_X1    g246(.A(KEYINPUT19), .ZN(new_n672));
  OR2_X1    g247(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n671), .A2(new_n672), .ZN(new_n674));
  NAND2_X1  g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(G1956), .B(G2474), .ZN(new_n676));
  XNOR2_X1  g251(.A(G1961), .B(G1966), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n676), .A2(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(KEYINPUT76), .B(KEYINPUT20), .Z(new_n679));
  AND3_X1   g254(.A1(new_n675), .A2(new_n678), .A3(new_n679), .ZN(new_n680));
  AOI21_X1  g255(.A(new_n679), .B1(new_n675), .B2(new_n678), .ZN(new_n681));
  NOR2_X1   g256(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  NAND3_X1  g257(.A1(new_n673), .A2(new_n678), .A3(new_n674), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n676), .A2(new_n677), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT77), .ZN(new_n685));
  OAI211_X1 g260(.A(new_n683), .B(new_n684), .C1(new_n675), .C2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n671), .B(KEYINPUT19), .ZN(new_n687));
  INV_X1    g262(.A(new_n684), .ZN(new_n688));
  OAI211_X1 g263(.A(new_n687), .B(KEYINPUT77), .C1(new_n688), .C2(new_n678), .ZN(new_n689));
  NAND2_X1  g264(.A1(new_n686), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(KEYINPUT78), .ZN(new_n691));
  AND3_X1   g266(.A1(new_n682), .A2(new_n690), .A3(new_n691), .ZN(new_n692));
  AOI21_X1  g267(.A(new_n691), .B1(new_n682), .B2(new_n690), .ZN(new_n693));
  OAI21_X1  g268(.A(new_n670), .B1(new_n692), .B2(new_n693), .ZN(new_n694));
  NAND2_X1  g269(.A1(new_n682), .A2(new_n690), .ZN(new_n695));
  NAND2_X1  g270(.A1(new_n695), .A2(KEYINPUT78), .ZN(new_n696));
  NAND3_X1  g271(.A1(new_n682), .A2(new_n690), .A3(new_n691), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n696), .A2(new_n697), .A3(new_n669), .ZN(new_n698));
  XNOR2_X1  g273(.A(G1991), .B(G1996), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT79), .Z(new_n700));
  INV_X1    g275(.A(new_n700), .ZN(new_n701));
  AND3_X1   g276(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n701), .B1(new_n694), .B2(new_n698), .ZN(new_n703));
  OAI21_X1  g278(.A(new_n668), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n694), .A2(new_n698), .ZN(new_n705));
  NAND2_X1  g280(.A1(new_n705), .A2(new_n700), .ZN(new_n706));
  NAND3_X1  g281(.A1(new_n694), .A2(new_n698), .A3(new_n701), .ZN(new_n707));
  NAND3_X1  g282(.A1(new_n706), .A2(new_n667), .A3(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n704), .A2(new_n708), .ZN(G229));
  XOR2_X1   g284(.A(KEYINPUT27), .B(G1996), .Z(new_n710));
  INV_X1    g285(.A(G29), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n711), .A2(G32), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n472), .A2(G141), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT90), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n713), .B(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n476), .A2(G129), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n716), .B(KEYINPUT91), .ZN(new_n717));
  NAND3_X1  g292(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT26), .ZN(new_n719));
  OR2_X1    g294(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n718), .A2(new_n719), .ZN(new_n721));
  AOI22_X1  g296(.A1(new_n720), .A2(new_n721), .B1(G105), .B2(new_n618), .ZN(new_n722));
  NAND3_X1  g297(.A1(new_n715), .A2(new_n717), .A3(new_n722), .ZN(new_n723));
  INV_X1    g298(.A(new_n723), .ZN(new_n724));
  OAI21_X1  g299(.A(new_n712), .B1(new_n724), .B2(new_n711), .ZN(new_n725));
  XOR2_X1   g300(.A(new_n725), .B(KEYINPUT92), .Z(new_n726));
  AND2_X1   g301(.A1(new_n711), .A2(G33), .ZN(new_n727));
  XOR2_X1   g302(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n728));
  NAND3_X1  g303(.A1(new_n468), .A2(G103), .A3(G2104), .ZN(new_n729));
  XNOR2_X1  g304(.A(new_n728), .B(new_n729), .ZN(new_n730));
  NAND2_X1  g305(.A1(new_n472), .A2(G139), .ZN(new_n731));
  AOI22_X1  g306(.A1(new_n617), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n730), .B(new_n731), .C1(new_n468), .C2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(KEYINPUT88), .ZN(new_n734));
  XNOR2_X1  g309(.A(new_n733), .B(new_n734), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(G29), .ZN(new_n736));
  INV_X1    g311(.A(G2072), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n736), .A2(new_n737), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n738), .A2(KEYINPUT89), .ZN(new_n739));
  OR2_X1    g314(.A1(new_n738), .A2(KEYINPUT89), .ZN(new_n740));
  AOI22_X1  g315(.A1(new_n710), .A2(new_n726), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(new_n710), .B2(new_n726), .ZN(new_n742));
  INV_X1    g317(.A(G16), .ZN(new_n743));
  NAND2_X1  g318(.A1(new_n743), .A2(G19), .ZN(new_n744));
  OAI21_X1  g319(.A(new_n744), .B1(new_n552), .B2(new_n743), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n745), .B(G1341), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n711), .A2(G27), .ZN(new_n747));
  OAI21_X1  g322(.A(new_n747), .B1(G164), .B2(new_n711), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n748), .B(KEYINPUT93), .ZN(new_n749));
  INV_X1    g324(.A(G2078), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n749), .B(new_n750), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT31), .B(G11), .Z(new_n752));
  INV_X1    g327(.A(G28), .ZN(new_n753));
  OR2_X1    g328(.A1(new_n753), .A2(KEYINPUT30), .ZN(new_n754));
  AOI21_X1  g329(.A(G29), .B1(new_n753), .B2(KEYINPUT30), .ZN(new_n755));
  AOI21_X1  g330(.A(new_n752), .B1(new_n754), .B2(new_n755), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT24), .ZN(new_n757));
  INV_X1    g332(.A(G34), .ZN(new_n758));
  AOI21_X1  g333(.A(G29), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  OAI21_X1  g334(.A(new_n759), .B1(new_n757), .B2(new_n758), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G160), .B2(new_n711), .ZN(new_n761));
  OAI221_X1 g336(.A(new_n756), .B1(new_n711), .B2(new_n627), .C1(new_n761), .C2(G2084), .ZN(new_n762));
  NAND2_X1  g337(.A1(new_n711), .A2(G26), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT28), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n472), .A2(G140), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n476), .A2(G128), .ZN(new_n766));
  OR2_X1    g341(.A1(G104), .A2(G2105), .ZN(new_n767));
  OAI211_X1 g342(.A(new_n767), .B(G2104), .C1(G116), .C2(new_n468), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n765), .A2(new_n766), .A3(new_n768), .ZN(new_n769));
  INV_X1    g344(.A(new_n769), .ZN(new_n770));
  OAI21_X1  g345(.A(new_n764), .B1(new_n770), .B2(new_n711), .ZN(new_n771));
  XOR2_X1   g346(.A(KEYINPUT86), .B(G2067), .Z(new_n772));
  NOR2_X1   g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G2084), .B2(new_n761), .ZN(new_n774));
  NAND2_X1  g349(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NOR2_X1   g350(.A1(G171), .A2(new_n743), .ZN(new_n776));
  AOI21_X1  g351(.A(new_n776), .B1(G5), .B2(new_n743), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  OAI211_X1 g353(.A(new_n774), .B(new_n775), .C1(new_n778), .C2(G1961), .ZN(new_n779));
  OR4_X1    g354(.A1(new_n746), .A2(new_n751), .A3(new_n762), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n743), .A2(G20), .ZN(new_n781));
  XOR2_X1   g356(.A(new_n781), .B(KEYINPUT23), .Z(new_n782));
  AOI21_X1  g357(.A(new_n782), .B1(G299), .B2(G16), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(G1956), .ZN(new_n784));
  NOR2_X1   g359(.A1(G29), .A2(G35), .ZN(new_n785));
  AOI21_X1  g360(.A(new_n785), .B1(G162), .B2(G29), .ZN(new_n786));
  XNOR2_X1  g361(.A(KEYINPUT94), .B(KEYINPUT29), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  INV_X1    g363(.A(G2090), .ZN(new_n789));
  OAI221_X1 g364(.A(new_n784), .B1(new_n737), .B2(new_n736), .C1(new_n788), .C2(new_n789), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n603), .A2(G16), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n791), .B1(G4), .B2(G16), .ZN(new_n792));
  INV_X1    g367(.A(G1348), .ZN(new_n793));
  AOI22_X1  g368(.A1(new_n792), .A2(new_n793), .B1(new_n789), .B2(new_n788), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n743), .A2(G21), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(G168), .B2(new_n743), .ZN(new_n796));
  NOR2_X1   g371(.A1(new_n796), .A2(G1966), .ZN(new_n797));
  AND2_X1   g372(.A1(new_n796), .A2(G1966), .ZN(new_n798));
  AOI211_X1 g373(.A(new_n797), .B(new_n798), .C1(new_n778), .C2(G1961), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n794), .B(new_n799), .C1(new_n793), .C2(new_n792), .ZN(new_n800));
  NOR4_X1   g375(.A1(new_n742), .A2(new_n780), .A3(new_n790), .A4(new_n800), .ZN(new_n801));
  INV_X1    g376(.A(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n743), .A2(G22), .ZN(new_n803));
  INV_X1    g378(.A(new_n803), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n804), .B1(G303), .B2(G16), .ZN(new_n805));
  INV_X1    g380(.A(G1971), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g382(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g383(.A1(new_n805), .A2(new_n806), .ZN(new_n809));
  OAI21_X1  g384(.A(KEYINPUT83), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n809), .ZN(new_n811));
  INV_X1    g386(.A(KEYINPUT83), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n811), .A2(new_n812), .A3(new_n807), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n743), .A2(G23), .ZN(new_n814));
  INV_X1    g389(.A(G288), .ZN(new_n815));
  OAI21_X1  g390(.A(new_n814), .B1(new_n815), .B2(new_n743), .ZN(new_n816));
  XNOR2_X1  g391(.A(KEYINPUT33), .B(G1976), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(KEYINPUT82), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n816), .B(new_n818), .Z(new_n819));
  NAND3_X1  g394(.A1(new_n810), .A2(new_n813), .A3(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n581), .A2(G16), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n821), .B1(G6), .B2(G16), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n822), .A2(KEYINPUT32), .ZN(new_n823));
  INV_X1    g398(.A(KEYINPUT32), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n824), .C1(G6), .C2(G16), .ZN(new_n825));
  NAND2_X1  g400(.A1(new_n823), .A2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(G1981), .ZN(new_n827));
  XNOR2_X1  g402(.A(new_n826), .B(new_n827), .ZN(new_n828));
  OAI21_X1  g403(.A(KEYINPUT84), .B1(new_n820), .B2(new_n828), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n816), .B(new_n818), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n811), .A2(new_n807), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n830), .B1(new_n831), .B2(KEYINPUT83), .ZN(new_n832));
  XNOR2_X1  g407(.A(new_n826), .B(G1981), .ZN(new_n833));
  INV_X1    g408(.A(KEYINPUT84), .ZN(new_n834));
  NAND4_X1  g409(.A1(new_n832), .A2(new_n833), .A3(new_n834), .A4(new_n813), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n829), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(KEYINPUT34), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(KEYINPUT85), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n743), .A2(G24), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT81), .Z(new_n841));
  AOI21_X1  g416(.A(new_n841), .B1(G290), .B2(G16), .ZN(new_n842));
  XOR2_X1   g417(.A(new_n842), .B(G1986), .Z(new_n843));
  NAND2_X1  g418(.A1(new_n711), .A2(G25), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(KEYINPUT80), .Z(new_n845));
  NAND2_X1  g420(.A1(new_n472), .A2(G131), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n476), .A2(G119), .ZN(new_n847));
  OR2_X1    g422(.A1(G95), .A2(G2105), .ZN(new_n848));
  OAI211_X1 g423(.A(new_n848), .B(G2104), .C1(G107), .C2(new_n468), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n846), .A2(new_n847), .A3(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  OAI21_X1  g426(.A(new_n845), .B1(new_n851), .B2(new_n711), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT35), .B(G1991), .Z(new_n853));
  XOR2_X1   g428(.A(new_n852), .B(new_n853), .Z(new_n854));
  NOR2_X1   g429(.A1(new_n843), .A2(new_n854), .ZN(new_n855));
  NAND3_X1  g430(.A1(new_n838), .A2(new_n839), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g431(.A(KEYINPUT34), .B1(new_n829), .B2(new_n835), .ZN(new_n857));
  INV_X1    g432(.A(new_n855), .ZN(new_n858));
  OAI21_X1  g433(.A(KEYINPUT85), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n856), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n836), .A2(new_n837), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n860), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n863), .A2(KEYINPUT36), .ZN(new_n864));
  INV_X1    g439(.A(KEYINPUT36), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n860), .A2(new_n865), .A3(new_n862), .ZN(new_n866));
  AOI21_X1  g441(.A(new_n802), .B1(new_n864), .B2(new_n866), .ZN(G311));
  AOI21_X1  g442(.A(new_n865), .B1(new_n860), .B2(new_n862), .ZN(new_n868));
  AOI211_X1 g443(.A(KEYINPUT36), .B(new_n861), .C1(new_n856), .C2(new_n859), .ZN(new_n869));
  OAI21_X1  g444(.A(new_n801), .B1(new_n868), .B2(new_n869), .ZN(G150));
  AOI22_X1  g445(.A1(new_n515), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n871));
  NOR2_X1   g446(.A1(new_n871), .A2(new_n510), .ZN(new_n872));
  INV_X1    g447(.A(G55), .ZN(new_n873));
  XOR2_X1   g448(.A(KEYINPUT95), .B(G93), .Z(new_n874));
  OAI22_X1  g449(.A1(new_n501), .A2(new_n873), .B1(new_n507), .B2(new_n874), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n872), .A2(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n877), .A2(G860), .ZN(new_n878));
  XOR2_X1   g453(.A(new_n878), .B(KEYINPUT37), .Z(new_n879));
  NAND2_X1  g454(.A1(new_n603), .A2(G559), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(KEYINPUT38), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n548), .A2(new_n550), .A3(new_n876), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n543), .A2(new_n547), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n877), .B1(new_n883), .B2(new_n549), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(new_n881), .B(new_n886), .ZN(new_n887));
  NOR2_X1   g462(.A1(new_n887), .A2(KEYINPUT39), .ZN(new_n888));
  INV_X1    g463(.A(KEYINPUT96), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n888), .B(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G860), .B1(new_n887), .B2(KEYINPUT39), .ZN(new_n891));
  AND3_X1   g466(.A1(new_n890), .A2(KEYINPUT97), .A3(new_n891), .ZN(new_n892));
  AOI21_X1  g467(.A(KEYINPUT97), .B1(new_n890), .B2(new_n891), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n879), .B1(new_n892), .B2(new_n893), .ZN(G145));
  XOR2_X1   g469(.A(KEYINPUT98), .B(G37), .Z(new_n895));
  NAND2_X1  g470(.A1(new_n472), .A2(G142), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n476), .A2(G130), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n468), .A2(G118), .ZN(new_n898));
  OAI21_X1  g473(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n899));
  OAI211_X1 g474(.A(new_n896), .B(new_n897), .C1(new_n898), .C2(new_n899), .ZN(new_n900));
  XNOR2_X1  g475(.A(new_n620), .B(new_n900), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n901), .B(new_n851), .ZN(new_n902));
  INV_X1    g477(.A(new_n902), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n496), .A2(new_n498), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n488), .A2(new_n491), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR2_X1   g481(.A1(new_n770), .A2(new_n906), .ZN(new_n907));
  NOR2_X1   g482(.A1(G164), .A2(new_n769), .ZN(new_n908));
  NOR2_X1   g483(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n909), .A2(new_n724), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n723), .B1(new_n907), .B2(new_n908), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n910), .A2(new_n733), .A3(new_n911), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  AOI21_X1  g488(.A(new_n735), .B1(new_n910), .B2(new_n911), .ZN(new_n914));
  OAI21_X1  g489(.A(new_n903), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  AND2_X1   g490(.A1(new_n910), .A2(new_n911), .ZN(new_n916));
  OAI211_X1 g491(.A(new_n902), .B(new_n912), .C1(new_n916), .C2(new_n735), .ZN(new_n917));
  XOR2_X1   g492(.A(new_n627), .B(new_n474), .Z(new_n918));
  XNOR2_X1  g493(.A(new_n918), .B(G162), .ZN(new_n919));
  AND3_X1   g494(.A1(new_n915), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n919), .B1(new_n915), .B2(new_n917), .ZN(new_n921));
  OAI21_X1  g496(.A(new_n895), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n922), .A2(KEYINPUT99), .ZN(new_n923));
  INV_X1    g498(.A(KEYINPUT99), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n924), .B(new_n895), .C1(new_n920), .C2(new_n921), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n926), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g502(.A(KEYINPUT102), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n928), .B1(new_n876), .B2(G868), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n885), .A2(new_n613), .ZN(new_n930));
  OAI211_X1 g505(.A(new_n882), .B(new_n884), .C1(G559), .C2(new_n602), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT100), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n602), .A2(G299), .A3(new_n933), .ZN(new_n934));
  AND2_X1   g509(.A1(new_n564), .A2(new_n565), .ZN(new_n935));
  XNOR2_X1  g510(.A(new_n558), .B(KEYINPUT9), .ZN(new_n936));
  NAND3_X1  g511(.A1(new_n935), .A2(KEYINPUT100), .A3(new_n936), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n933), .B1(new_n560), .B2(new_n566), .ZN(new_n938));
  NAND4_X1  g513(.A1(new_n937), .A2(new_n938), .A3(new_n596), .A4(new_n601), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n934), .A2(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT41), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  NAND3_X1  g517(.A1(new_n934), .A2(new_n939), .A3(KEYINPUT41), .ZN(new_n943));
  NAND4_X1  g518(.A1(new_n932), .A2(new_n942), .A3(KEYINPUT101), .A4(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n940), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n945), .A2(new_n930), .A3(new_n931), .ZN(new_n946));
  AND2_X1   g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  INV_X1    g522(.A(KEYINPUT42), .ZN(new_n948));
  INV_X1    g523(.A(new_n943), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT41), .B1(new_n934), .B2(new_n939), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n949), .A2(new_n950), .ZN(new_n951));
  AND2_X1   g526(.A1(new_n951), .A2(new_n932), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n947), .B(new_n948), .C1(new_n952), .C2(KEYINPUT101), .ZN(new_n953));
  AOI21_X1  g528(.A(KEYINPUT101), .B1(new_n951), .B2(new_n932), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n944), .A2(new_n946), .ZN(new_n955));
  OAI21_X1  g530(.A(KEYINPUT42), .B1(new_n954), .B2(new_n955), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  XNOR2_X1  g532(.A(new_n815), .B(G303), .ZN(new_n958));
  XNOR2_X1  g533(.A(G290), .B(new_n581), .ZN(new_n959));
  XOR2_X1   g534(.A(new_n958), .B(new_n959), .Z(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n611), .B1(new_n957), .B2(new_n961), .ZN(new_n962));
  NAND3_X1  g537(.A1(new_n953), .A2(new_n956), .A3(new_n960), .ZN(new_n963));
  AOI21_X1  g538(.A(new_n929), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AND2_X1   g539(.A1(new_n962), .A2(new_n963), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n964), .B1(KEYINPUT102), .B2(new_n965), .ZN(G295));
  AOI21_X1  g541(.A(new_n964), .B1(KEYINPUT102), .B2(new_n965), .ZN(G331));
  NAND2_X1  g542(.A1(G301), .A2(G286), .ZN(new_n968));
  NAND2_X1  g543(.A1(G171), .A2(G168), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n885), .A2(new_n970), .ZN(new_n971));
  NAND4_X1  g546(.A1(new_n882), .A2(new_n884), .A3(new_n968), .A4(new_n969), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n971), .A2(KEYINPUT104), .A3(new_n972), .ZN(new_n973));
  INV_X1    g548(.A(new_n970), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT104), .ZN(new_n975));
  NAND4_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n884), .A4(new_n882), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n943), .A3(new_n942), .A4(new_n976), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT105), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n979));
  NAND4_X1  g554(.A1(new_n951), .A2(new_n979), .A3(new_n976), .A4(new_n973), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n945), .A2(new_n972), .A3(new_n971), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(new_n960), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT43), .ZN(new_n984));
  INV_X1    g559(.A(new_n895), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n971), .A2(new_n972), .ZN(new_n986));
  AND3_X1   g561(.A1(new_n986), .A2(new_n942), .A3(new_n943), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n940), .B1(new_n973), .B2(new_n976), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n987), .A2(new_n988), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n985), .B1(new_n989), .B2(new_n961), .ZN(new_n990));
  NAND3_X1  g565(.A1(new_n983), .A2(new_n984), .A3(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n951), .A2(new_n986), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n973), .A2(new_n976), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n992), .B(new_n961), .C1(new_n993), .C2(new_n940), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n960), .B1(new_n987), .B2(new_n988), .ZN(new_n995));
  INV_X1    g570(.A(G37), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n994), .A2(new_n995), .A3(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n991), .A2(new_n998), .ZN(new_n999));
  XNOR2_X1  g574(.A(KEYINPUT103), .B(KEYINPUT44), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  AOI21_X1  g576(.A(new_n984), .B1(new_n983), .B2(new_n990), .ZN(new_n1002));
  OAI21_X1  g577(.A(KEYINPUT44), .B1(new_n997), .B2(KEYINPUT43), .ZN(new_n1003));
  OAI21_X1  g578(.A(new_n1001), .B1(new_n1002), .B2(new_n1003), .ZN(G397));
  XNOR2_X1  g579(.A(new_n769), .B(G2067), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1005), .B(KEYINPUT107), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1006), .A2(new_n724), .ZN(new_n1007));
  INV_X1    g582(.A(KEYINPUT45), .ZN(new_n1008));
  XOR2_X1   g583(.A(KEYINPUT106), .B(G1384), .Z(new_n1009));
  OAI21_X1  g584(.A(new_n1008), .B1(G164), .B2(new_n1009), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n467), .A2(new_n473), .A3(G40), .ZN(new_n1011));
  NOR2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1007), .A2(new_n1012), .ZN(new_n1013));
  XNOR2_X1  g588(.A(new_n1013), .B(KEYINPUT125), .ZN(new_n1014));
  INV_X1    g589(.A(G1996), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1012), .A2(new_n1015), .ZN(new_n1016));
  XNOR2_X1  g591(.A(new_n1016), .B(KEYINPUT46), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1014), .A2(new_n1017), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT47), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n723), .A2(G1996), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n724), .A2(new_n1015), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1006), .A2(new_n1020), .A3(new_n1021), .ZN(new_n1022));
  XOR2_X1   g597(.A(new_n850), .B(new_n853), .Z(new_n1023));
  OAI21_X1  g598(.A(new_n1012), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  NOR2_X1   g599(.A1(G290), .A2(G1986), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n1012), .A2(new_n1025), .ZN(new_n1026));
  XNOR2_X1  g601(.A(new_n1026), .B(KEYINPUT48), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1024), .A2(new_n1027), .ZN(new_n1028));
  NAND2_X1  g603(.A1(new_n851), .A2(new_n853), .ZN(new_n1029));
  XNOR2_X1  g604(.A(new_n1029), .B(KEYINPUT124), .ZN(new_n1030));
  OAI22_X1  g605(.A1(new_n1022), .A2(new_n1030), .B1(G2067), .B2(new_n769), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n1012), .ZN(new_n1032));
  AND3_X1   g607(.A1(new_n1019), .A2(new_n1028), .A3(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1008), .B1(G164), .B2(G1384), .ZN(new_n1034));
  INV_X1    g609(.A(new_n1009), .ZN(new_n1035));
  NAND3_X1  g610(.A1(new_n906), .A2(KEYINPUT45), .A3(new_n1035), .ZN(new_n1036));
  AND3_X1   g611(.A1(new_n467), .A2(new_n473), .A3(G40), .ZN(new_n1037));
  NAND4_X1  g612(.A1(new_n1034), .A2(new_n1015), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1038));
  AOI21_X1  g613(.A(G1384), .B1(new_n904), .B2(new_n905), .ZN(new_n1039));
  NAND2_X1  g614(.A1(new_n1039), .A2(new_n1037), .ZN(new_n1040));
  XOR2_X1   g615(.A(KEYINPUT58), .B(G1341), .Z(new_n1041));
  NAND2_X1  g616(.A1(new_n1040), .A2(new_n1041), .ZN(new_n1042));
  AOI21_X1  g617(.A(new_n551), .B1(new_n1038), .B2(new_n1042), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT59), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n560), .A2(new_n566), .A3(KEYINPUT57), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT57), .ZN(new_n1046));
  AOI21_X1  g621(.A(new_n1046), .B1(new_n935), .B2(new_n936), .ZN(new_n1047));
  OR2_X1    g622(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1048));
  INV_X1    g623(.A(G1384), .ZN(new_n1049));
  INV_X1    g624(.A(new_n498), .ZN(new_n1050));
  AOI21_X1  g625(.A(new_n497), .B1(new_n617), .B2(new_n494), .ZN(new_n1051));
  NOR2_X1   g626(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1049), .B1(new_n1052), .B2(new_n492), .ZN(new_n1053));
  AOI21_X1  g628(.A(new_n1011), .B1(new_n1053), .B2(KEYINPUT50), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT50), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n906), .A2(new_n1055), .A3(new_n1049), .ZN(new_n1056));
  AOI21_X1  g631(.A(G1956), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n1037), .B1(new_n1039), .B2(KEYINPUT45), .ZN(new_n1058));
  AOI211_X1 g633(.A(new_n1008), .B(new_n1009), .C1(new_n904), .C2(new_n905), .ZN(new_n1059));
  XNOR2_X1  g634(.A(KEYINPUT56), .B(G2072), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n1058), .A2(new_n1059), .A3(new_n1061), .ZN(new_n1062));
  OAI21_X1  g637(.A(new_n1048), .B1(new_n1057), .B2(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n1064), .A2(new_n1037), .A3(new_n1056), .ZN(new_n1065));
  INV_X1    g640(.A(G1956), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1067));
  NOR2_X1   g642(.A1(new_n1045), .A2(new_n1047), .ZN(new_n1068));
  AOI21_X1  g643(.A(new_n1011), .B1(new_n1053), .B2(new_n1008), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1069), .A2(new_n1036), .A3(new_n1060), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1067), .A2(new_n1068), .A3(new_n1070), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT61), .B1(new_n1063), .B2(new_n1071), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1044), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g648(.A(new_n1068), .B1(new_n1067), .B2(new_n1070), .ZN(new_n1074));
  OAI21_X1  g649(.A(new_n1071), .B1(new_n1074), .B2(KEYINPUT117), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT117), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1067), .A2(new_n1070), .A3(new_n1068), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n1075), .A2(KEYINPUT61), .A3(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(G2067), .ZN(new_n1079));
  AND3_X1   g654(.A1(new_n1039), .A2(new_n1037), .A3(new_n1079), .ZN(new_n1080));
  AOI211_X1 g655(.A(KEYINPUT115), .B(new_n1080), .C1(new_n1065), .C2(new_n793), .ZN(new_n1081));
  INV_X1    g656(.A(KEYINPUT115), .ZN(new_n1082));
  OAI21_X1  g657(.A(new_n1037), .B1(new_n1039), .B2(new_n1055), .ZN(new_n1083));
  NOR3_X1   g658(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n793), .B1(new_n1083), .B2(new_n1084), .ZN(new_n1085));
  INV_X1    g660(.A(new_n1080), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1082), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g662(.A(KEYINPUT60), .B1(new_n1081), .B2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(G1348), .B1(new_n1054), .B2(new_n1056), .ZN(new_n1089));
  OAI21_X1  g664(.A(KEYINPUT115), .B1(new_n1089), .B2(new_n1080), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT60), .ZN(new_n1091));
  NAND3_X1  g666(.A1(new_n1085), .A2(new_n1082), .A3(new_n1086), .ZN(new_n1092));
  NAND3_X1  g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1088), .A2(new_n603), .A3(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(KEYINPUT60), .B(new_n602), .C1(new_n1081), .C2(new_n1087), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1073), .A2(new_n1078), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1090), .A2(new_n603), .A3(new_n1092), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(new_n1063), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1098), .A2(new_n1071), .ZN(new_n1099));
  INV_X1    g674(.A(KEYINPUT116), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1098), .A2(KEYINPUT116), .A3(new_n1071), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1096), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(G1966), .ZN(new_n1104));
  NOR3_X1   g679(.A1(G164), .A2(new_n1008), .A3(G1384), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1104), .B1(new_n1058), .B2(new_n1105), .ZN(new_n1106));
  INV_X1    g681(.A(G2084), .ZN(new_n1107));
  NAND4_X1  g682(.A1(new_n1064), .A2(new_n1107), .A3(new_n1056), .A4(new_n1037), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1106), .A2(G168), .A3(new_n1108), .ZN(new_n1109));
  AND2_X1   g684(.A1(KEYINPUT118), .A2(G8), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g686(.A1(new_n1111), .A2(KEYINPUT51), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT51), .ZN(new_n1113));
  NAND3_X1  g688(.A1(new_n1109), .A2(new_n1113), .A3(new_n1110), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1106), .A2(new_n1108), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1115), .A2(G8), .A3(G286), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1112), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT54), .ZN(new_n1118));
  NOR2_X1   g693(.A1(new_n1058), .A2(new_n1105), .ZN(new_n1119));
  AND2_X1   g694(.A1(new_n750), .A2(KEYINPUT53), .ZN(new_n1120));
  XOR2_X1   g695(.A(KEYINPUT119), .B(G1961), .Z(new_n1121));
  AOI22_X1  g696(.A1(new_n1119), .A2(new_n1120), .B1(new_n1065), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1034), .A2(new_n750), .A3(new_n1036), .A4(new_n1037), .ZN(new_n1123));
  XNOR2_X1  g698(.A(KEYINPUT120), .B(KEYINPUT53), .ZN(new_n1124));
  NAND2_X1  g699(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(G301), .B1(new_n1122), .B2(new_n1125), .ZN(new_n1126));
  NAND2_X1  g701(.A1(new_n618), .A2(G101), .ZN(new_n1127));
  OAI211_X1 g702(.A(G137), .B(new_n468), .C1(new_n489), .C2(new_n490), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g704(.A(KEYINPUT121), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND3_X1  g706(.A1(new_n1127), .A2(new_n1128), .A3(KEYINPUT121), .ZN(new_n1132));
  AND2_X1   g707(.A1(new_n1120), .A2(G40), .ZN(new_n1133));
  NAND4_X1  g708(.A1(new_n1131), .A2(new_n467), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1009), .B1(new_n904), .B2(new_n905), .ZN(new_n1135));
  AOI21_X1  g710(.A(new_n1134), .B1(KEYINPUT45), .B2(new_n1135), .ZN(new_n1136));
  AOI22_X1  g711(.A1(new_n1065), .A2(new_n1121), .B1(new_n1136), .B2(new_n1010), .ZN(new_n1137));
  AND3_X1   g712(.A1(new_n1137), .A2(G301), .A3(new_n1125), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1118), .B1(new_n1126), .B2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1137), .A2(KEYINPUT122), .A3(new_n1125), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT122), .B1(new_n1137), .B2(new_n1125), .ZN(new_n1141));
  NOR3_X1   g716(.A1(new_n1140), .A2(new_n1141), .A3(G301), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1122), .A2(G301), .A3(new_n1125), .ZN(new_n1143));
  NAND2_X1  g718(.A1(new_n1143), .A2(KEYINPUT54), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1117), .B(new_n1139), .C1(new_n1142), .C2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g720(.A1(G303), .A2(G8), .ZN(new_n1146));
  XNOR2_X1  g721(.A(new_n1146), .B(KEYINPUT55), .ZN(new_n1147));
  XOR2_X1   g722(.A(KEYINPUT109), .B(G1971), .Z(new_n1148));
  AOI21_X1  g723(.A(new_n1148), .B1(new_n1069), .B2(new_n1036), .ZN(new_n1149));
  AOI21_X1  g724(.A(G2090), .B1(new_n1065), .B2(KEYINPUT112), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT112), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1054), .A2(new_n1151), .A3(new_n1056), .ZN(new_n1152));
  AOI21_X1  g727(.A(new_n1149), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  INV_X1    g728(.A(G8), .ZN(new_n1154));
  OAI21_X1  g729(.A(new_n1147), .B1(new_n1153), .B2(new_n1154), .ZN(new_n1155));
  INV_X1    g730(.A(new_n1147), .ZN(new_n1156));
  NAND3_X1  g731(.A1(new_n1054), .A2(new_n789), .A3(new_n1056), .ZN(new_n1157));
  OAI21_X1  g732(.A(new_n1157), .B1(new_n1149), .B2(KEYINPUT110), .ZN(new_n1158));
  NOR2_X1   g733(.A1(new_n1058), .A2(new_n1059), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT110), .ZN(new_n1160));
  NOR3_X1   g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n1148), .ZN(new_n1161));
  OAI211_X1 g736(.A(G8), .B(new_n1156), .C1(new_n1158), .C2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g737(.A(G1981), .B1(new_n577), .B2(new_n580), .ZN(new_n1163));
  INV_X1    g738(.A(G61), .ZN(new_n1164));
  AOI21_X1  g739(.A(new_n1164), .B1(new_n513), .B2(new_n514), .ZN(new_n1165));
  INV_X1    g740(.A(new_n579), .ZN(new_n1166));
  OAI21_X1  g741(.A(G651), .B1(new_n1165), .B2(new_n1166), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n515), .A2(new_n500), .A3(G86), .ZN(new_n1168));
  NAND4_X1  g743(.A1(new_n1167), .A2(new_n827), .A3(new_n1168), .A4(new_n575), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1163), .A2(KEYINPUT49), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1154), .B1(new_n1039), .B2(new_n1037), .ZN(new_n1171));
  NAND2_X1  g746(.A1(new_n1163), .A2(new_n1169), .ZN(new_n1172));
  INV_X1    g747(.A(KEYINPUT49), .ZN(new_n1173));
  AOI21_X1  g748(.A(KEYINPUT111), .B1(new_n1172), .B2(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT111), .ZN(new_n1175));
  AOI211_X1 g750(.A(new_n1175), .B(KEYINPUT49), .C1(new_n1163), .C2(new_n1169), .ZN(new_n1176));
  OAI211_X1 g751(.A(new_n1170), .B(new_n1171), .C1(new_n1174), .C2(new_n1176), .ZN(new_n1177));
  INV_X1    g752(.A(G1976), .ZN(new_n1178));
  AOI21_X1  g753(.A(KEYINPUT52), .B1(G288), .B2(new_n1178), .ZN(new_n1179));
  OAI211_X1 g754(.A(new_n1171), .B(new_n1179), .C1(new_n1178), .C2(G288), .ZN(new_n1180));
  OAI211_X1 g755(.A(new_n1040), .B(G8), .C1(new_n1178), .C2(G288), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1181), .A2(KEYINPUT52), .ZN(new_n1182));
  AND3_X1   g757(.A1(new_n1177), .A2(new_n1180), .A3(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1155), .A2(new_n1162), .A3(new_n1183), .ZN(new_n1184));
  NOR2_X1   g759(.A1(new_n1145), .A2(new_n1184), .ZN(new_n1185));
  NAND2_X1  g760(.A1(new_n1103), .A2(new_n1185), .ZN(new_n1186));
  AND3_X1   g761(.A1(new_n1155), .A2(new_n1162), .A3(new_n1183), .ZN(new_n1187));
  INV_X1    g762(.A(KEYINPUT62), .ZN(new_n1188));
  NAND4_X1  g763(.A1(new_n1112), .A2(new_n1114), .A3(new_n1188), .A4(new_n1116), .ZN(new_n1189));
  NAND4_X1  g764(.A1(new_n1187), .A2(KEYINPUT123), .A3(new_n1126), .A4(new_n1189), .ZN(new_n1190));
  INV_X1    g765(.A(KEYINPUT123), .ZN(new_n1191));
  INV_X1    g766(.A(new_n1189), .ZN(new_n1192));
  NAND4_X1  g767(.A1(new_n1155), .A2(new_n1162), .A3(new_n1183), .A4(new_n1126), .ZN(new_n1193));
  OAI21_X1  g768(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1117), .A2(KEYINPUT62), .ZN(new_n1195));
  NAND3_X1  g770(.A1(new_n1190), .A2(new_n1194), .A3(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1186), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g772(.A1(new_n1115), .A2(G8), .A3(G168), .ZN(new_n1198));
  INV_X1    g773(.A(new_n1198), .ZN(new_n1199));
  NAND4_X1  g774(.A1(new_n1155), .A2(new_n1162), .A3(new_n1199), .A4(new_n1183), .ZN(new_n1200));
  INV_X1    g775(.A(KEYINPUT63), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1200), .A2(new_n1201), .ZN(new_n1202));
  NAND4_X1  g777(.A1(new_n1177), .A2(KEYINPUT63), .A3(new_n1182), .A4(new_n1180), .ZN(new_n1203));
  NOR2_X1   g778(.A1(new_n1203), .A2(new_n1198), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1204), .A2(new_n1162), .ZN(new_n1205));
  NAND2_X1  g780(.A1(new_n1149), .A2(KEYINPUT110), .ZN(new_n1206));
  OAI21_X1  g781(.A(new_n1160), .B1(new_n1159), .B2(new_n1148), .ZN(new_n1207));
  NAND3_X1  g782(.A1(new_n1206), .A2(new_n1207), .A3(new_n1157), .ZN(new_n1208));
  AOI21_X1  g783(.A(new_n1156), .B1(new_n1208), .B2(G8), .ZN(new_n1209));
  OAI21_X1  g784(.A(KEYINPUT113), .B1(new_n1205), .B2(new_n1209), .ZN(new_n1210));
  NAND2_X1  g785(.A1(new_n1208), .A2(G8), .ZN(new_n1211));
  NAND2_X1  g786(.A1(new_n1211), .A2(new_n1147), .ZN(new_n1212));
  INV_X1    g787(.A(KEYINPUT113), .ZN(new_n1213));
  NAND4_X1  g788(.A1(new_n1212), .A2(new_n1213), .A3(new_n1162), .A4(new_n1204), .ZN(new_n1214));
  NAND3_X1  g789(.A1(new_n1202), .A2(new_n1210), .A3(new_n1214), .ZN(new_n1215));
  INV_X1    g790(.A(KEYINPUT114), .ZN(new_n1216));
  INV_X1    g791(.A(new_n1162), .ZN(new_n1217));
  NAND3_X1  g792(.A1(new_n1177), .A2(new_n1178), .A3(new_n815), .ZN(new_n1218));
  NAND2_X1  g793(.A1(new_n1218), .A2(new_n1169), .ZN(new_n1219));
  AOI22_X1  g794(.A1(new_n1217), .A2(new_n1183), .B1(new_n1171), .B2(new_n1219), .ZN(new_n1220));
  NAND3_X1  g795(.A1(new_n1215), .A2(new_n1216), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g796(.A1(new_n1215), .A2(new_n1220), .ZN(new_n1222));
  NAND2_X1  g797(.A1(new_n1222), .A2(KEYINPUT114), .ZN(new_n1223));
  AOI21_X1  g798(.A(new_n1197), .B1(new_n1221), .B2(new_n1223), .ZN(new_n1224));
  AND2_X1   g799(.A1(G290), .A2(G1986), .ZN(new_n1225));
  OAI21_X1  g800(.A(new_n1012), .B1(new_n1225), .B2(new_n1025), .ZN(new_n1226));
  NAND2_X1  g801(.A1(new_n1024), .A2(new_n1226), .ZN(new_n1227));
  XOR2_X1   g802(.A(new_n1227), .B(KEYINPUT108), .Z(new_n1228));
  OAI21_X1  g803(.A(new_n1033), .B1(new_n1224), .B2(new_n1228), .ZN(G329));
  assign    G231 = 1'b0;
  NAND3_X1  g804(.A1(new_n664), .A2(G319), .A3(new_n665), .ZN(new_n1231));
  NOR2_X1   g805(.A1(G401), .A2(new_n1231), .ZN(new_n1232));
  NAND3_X1  g806(.A1(new_n704), .A2(new_n708), .A3(new_n1232), .ZN(new_n1233));
  INV_X1    g807(.A(KEYINPUT126), .ZN(new_n1234));
  NAND2_X1  g808(.A1(new_n1233), .A2(new_n1234), .ZN(new_n1235));
  NAND4_X1  g809(.A1(new_n704), .A2(new_n708), .A3(KEYINPUT126), .A4(new_n1232), .ZN(new_n1236));
  AOI22_X1  g810(.A1(new_n923), .A2(new_n925), .B1(new_n1235), .B2(new_n1236), .ZN(new_n1237));
  AND3_X1   g811(.A1(new_n1237), .A2(new_n999), .A3(KEYINPUT127), .ZN(new_n1238));
  AOI21_X1  g812(.A(KEYINPUT127), .B1(new_n1237), .B2(new_n999), .ZN(new_n1239));
  NOR2_X1   g813(.A1(new_n1238), .A2(new_n1239), .ZN(G308));
  NAND2_X1  g814(.A1(new_n1237), .A2(new_n999), .ZN(G225));
endmodule


