

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759;

  XNOR2_X1 U368 ( .A(n488), .B(n489), .ZN(n743) );
  XNOR2_X1 U369 ( .A(n474), .B(n473), .ZN(n488) );
  XNOR2_X1 U370 ( .A(n357), .B(n461), .ZN(n742) );
  XOR2_X1 U371 ( .A(G104), .B(G113), .Z(n454) );
  XNOR2_X1 U372 ( .A(n438), .B(KEYINPUT89), .ZN(n440) );
  XNOR2_X1 U373 ( .A(G140), .B(KEYINPUT10), .ZN(n461) );
  XNOR2_X1 U374 ( .A(G146), .B(G125), .ZN(n357) );
  INV_X1 U375 ( .A(G953), .ZN(n745) );
  INV_X2 U376 ( .A(G143), .ZN(n433) );
  BUF_X2 U377 ( .A(n382), .Z(n721) );
  NAND2_X1 U378 ( .A1(n527), .A2(n482), .ZN(n485) );
  NOR2_X1 U379 ( .A1(n623), .A2(n407), .ZN(n382) );
  AND2_X2 U380 ( .A1(n614), .A2(n651), .ZN(n576) );
  NOR2_X2 U381 ( .A1(n668), .A2(n616), .ZN(n615) );
  NOR2_X2 U382 ( .A1(n674), .A2(n577), .ZN(n571) );
  XNOR2_X2 U383 ( .A(n526), .B(KEYINPUT65), .ZN(n674) );
  XNOR2_X2 U384 ( .A(n470), .B(n345), .ZN(n513) );
  AND2_X2 U385 ( .A1(n351), .A2(n352), .ZN(n394) );
  XNOR2_X2 U386 ( .A(G902), .B(KEYINPUT15), .ZN(n616) );
  XNOR2_X2 U387 ( .A(n483), .B(KEYINPUT22), .ZN(n484) );
  NAND2_X1 U388 ( .A1(n409), .A2(n410), .ZN(n408) );
  XNOR2_X2 U389 ( .A(G146), .B(G125), .ZN(n462) );
  XOR2_X1 U390 ( .A(KEYINPUT11), .B(KEYINPUT12), .Z(n456) );
  XNOR2_X1 U391 ( .A(G116), .B(G107), .ZN(n466) );
  NOR2_X1 U392 ( .A1(n581), .A2(n596), .ZN(n582) );
  XNOR2_X2 U393 ( .A(n587), .B(n586), .ZN(n754) );
  OR2_X2 U394 ( .A1(n591), .A2(n673), .ZN(n586) );
  AND2_X2 U395 ( .A1(n414), .A2(n365), .ZN(n409) );
  XNOR2_X2 U396 ( .A(G101), .B(G107), .ZN(n438) );
  XNOR2_X2 U397 ( .A(n423), .B(KEYINPUT0), .ZN(n527) );
  NOR2_X1 U398 ( .A1(n623), .A2(n356), .ZN(n724) );
  XNOR2_X2 U399 ( .A(n730), .B(KEYINPUT71), .ZN(n505) );
  XNOR2_X2 U400 ( .A(n440), .B(n439), .ZN(n730) );
  XNOR2_X2 U401 ( .A(n499), .B(n498), .ZN(n569) );
  OR2_X1 U402 ( .A1(n615), .A2(KEYINPUT82), .ZN(n428) );
  XNOR2_X1 U403 ( .A(n542), .B(n541), .ZN(n635) );
  XNOR2_X1 U404 ( .A(n418), .B(n572), .ZN(n603) );
  NAND2_X1 U405 ( .A1(n361), .A2(n419), .ZN(n418) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n345) );
  XNOR2_X1 U407 ( .A(n406), .B(n549), .ZN(n561) );
  NOR2_X1 U408 ( .A1(n635), .A2(n548), .ZN(n406) );
  XNOR2_X1 U409 ( .A(n402), .B(n558), .ZN(n758) );
  XNOR2_X1 U410 ( .A(n574), .B(KEYINPUT39), .ZN(n614) );
  AND2_X1 U411 ( .A1(n571), .A2(n420), .ZN(n419) );
  XOR2_X1 U412 ( .A(n632), .B(n633), .Z(n368) );
  XNOR2_X1 U413 ( .A(n525), .B(n524), .ZN(n677) );
  XNOR2_X1 U414 ( .A(n629), .B(n628), .ZN(n367) );
  XNOR2_X1 U415 ( .A(KEYINPUT62), .B(n624), .ZN(n369) );
  NOR2_X1 U416 ( .A1(n725), .A2(G902), .ZN(n525) );
  XNOR2_X1 U417 ( .A(n743), .B(G146), .ZN(n506) );
  NAND2_X1 U418 ( .A1(n513), .A2(G221), .ZN(n514) );
  XNOR2_X1 U419 ( .A(KEYINPUT78), .B(KEYINPUT18), .ZN(n379) );
  XNOR2_X1 U420 ( .A(KEYINPUT77), .B(KEYINPUT4), .ZN(n380) );
  NOR2_X1 U421 ( .A1(n677), .A2(n678), .ZN(n526) );
  NAND2_X1 U422 ( .A1(n617), .A2(n429), .ZN(n427) );
  XNOR2_X2 U423 ( .A(n347), .B(KEYINPUT45), .ZN(n617) );
  AND2_X2 U424 ( .A1(n666), .A2(n622), .ZN(n407) );
  NAND2_X1 U425 ( .A1(n346), .A2(n417), .ZN(n416) );
  XNOR2_X1 U426 ( .A(n588), .B(KEYINPUT46), .ZN(n346) );
  NAND2_X1 U427 ( .A1(n565), .A2(n564), .ZN(n347) );
  AND2_X1 U428 ( .A1(n394), .A2(n412), .ZN(n348) );
  NAND2_X1 U429 ( .A1(n410), .A2(n409), .ZN(n349) );
  XNOR2_X2 U430 ( .A(n576), .B(n575), .ZN(n759) );
  NAND2_X1 U431 ( .A1(n543), .A2(n350), .ZN(n542) );
  AND2_X1 U432 ( .A1(n501), .A2(n539), .ZN(n350) );
  NAND2_X1 U433 ( .A1(n511), .A2(n354), .ZN(n351) );
  OR2_X1 U434 ( .A1(n353), .A2(n364), .ZN(n352) );
  INV_X1 U435 ( .A(KEYINPUT100), .ZN(n353) );
  AND2_X1 U436 ( .A1(n425), .A2(KEYINPUT100), .ZN(n354) );
  NAND2_X1 U437 ( .A1(n374), .A2(n373), .ZN(n372) );
  AND2_X1 U438 ( .A1(n374), .A2(n373), .ZN(n355) );
  XNOR2_X2 U439 ( .A(n538), .B(KEYINPUT83), .ZN(n511) );
  XNOR2_X2 U440 ( .A(n485), .B(n484), .ZN(n543) );
  AND2_X2 U441 ( .A1(n666), .A2(n622), .ZN(n356) );
  BUF_X2 U442 ( .A(n617), .Z(n666) );
  NOR2_X1 U443 ( .A1(n617), .A2(KEYINPUT82), .ZN(n359) );
  INV_X1 U444 ( .A(KEYINPUT86), .ZN(n549) );
  NAND2_X1 U445 ( .A1(n397), .A2(n604), .ZN(n396) );
  INV_X1 U446 ( .A(n431), .ZN(n397) );
  XNOR2_X1 U447 ( .A(n379), .B(n381), .ZN(n377) );
  XNOR2_X1 U448 ( .A(n416), .B(n415), .ZN(n621) );
  INV_X1 U449 ( .A(KEYINPUT48), .ZN(n415) );
  AND2_X1 U450 ( .A1(n605), .A2(n606), .ZN(n417) );
  INV_X1 U451 ( .A(n534), .ZN(n554) );
  NAND2_X1 U452 ( .A1(n495), .A2(n358), .ZN(n373) );
  XOR2_X1 U453 ( .A(G110), .B(G104), .Z(n439) );
  XNOR2_X1 U454 ( .A(G128), .B(G110), .ZN(n516) );
  XOR2_X1 U455 ( .A(G119), .B(G137), .Z(n515) );
  INV_X1 U456 ( .A(G134), .ZN(n473) );
  NOR2_X1 U457 ( .A1(n596), .A2(n595), .ZN(n607) );
  INV_X1 U458 ( .A(KEYINPUT87), .ZN(n399) );
  INV_X1 U459 ( .A(KEYINPUT36), .ZN(n598) );
  OR2_X1 U460 ( .A1(n675), .A2(n512), .ZN(n424) );
  NAND2_X1 U461 ( .A1(n401), .A2(n400), .ZN(n405) );
  INV_X1 U462 ( .A(KEYINPUT44), .ZN(n400) );
  NAND2_X1 U463 ( .A1(n758), .A2(KEYINPUT85), .ZN(n401) );
  XNOR2_X1 U464 ( .A(KEYINPUT4), .B(G131), .ZN(n486) );
  XOR2_X1 U465 ( .A(KEYINPUT66), .B(G137), .Z(n487) );
  XNOR2_X1 U466 ( .A(G122), .B(KEYINPUT94), .ZN(n455) );
  NOR2_X1 U467 ( .A1(G953), .A2(G237), .ZN(n490) );
  NOR2_X1 U468 ( .A1(n359), .A2(n426), .ZN(n623) );
  XNOR2_X1 U469 ( .A(n573), .B(KEYINPUT38), .ZN(n689) );
  INV_X1 U470 ( .A(n578), .ZN(n420) );
  XNOR2_X1 U471 ( .A(G119), .B(G116), .ZN(n435) );
  XNOR2_X1 U472 ( .A(G122), .B(KEYINPUT7), .ZN(n467) );
  XNOR2_X1 U473 ( .A(n474), .B(n434), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n551), .B(n366), .ZN(n699) );
  BUF_X1 U475 ( .A(n569), .Z(n395) );
  XNOR2_X1 U476 ( .A(n478), .B(n477), .ZN(n534) );
  XNOR2_X1 U477 ( .A(n355), .B(n731), .ZN(n733) );
  XNOR2_X1 U478 ( .A(n520), .B(n519), .ZN(n725) );
  XNOR2_X1 U479 ( .A(n742), .B(n518), .ZN(n519) );
  XNOR2_X1 U480 ( .A(n599), .B(n398), .ZN(n600) );
  XNOR2_X1 U481 ( .A(n598), .B(n399), .ZN(n398) );
  NAND2_X1 U482 ( .A1(n413), .A2(n371), .ZN(n412) );
  NAND2_X1 U483 ( .A1(n413), .A2(KEYINPUT84), .ZN(n410) );
  XNOR2_X1 U484 ( .A(n723), .B(n722), .ZN(n384) );
  INV_X1 U485 ( .A(KEYINPUT60), .ZN(n388) );
  INV_X1 U486 ( .A(KEYINPUT56), .ZN(n386) );
  XOR2_X1 U487 ( .A(KEYINPUT16), .B(G122), .Z(n358) );
  AND2_X1 U488 ( .A1(n428), .A2(n370), .ZN(n360) );
  XOR2_X1 U489 ( .A(KEYINPUT30), .B(n570), .Z(n361) );
  XOR2_X1 U490 ( .A(KEYINPUT9), .B(KEYINPUT95), .Z(n362) );
  AND2_X1 U491 ( .A1(n443), .A2(G210), .ZN(n363) );
  AND2_X1 U492 ( .A1(n424), .A2(n544), .ZN(n364) );
  AND2_X1 U493 ( .A1(n364), .A2(n353), .ZN(n365) );
  XNOR2_X1 U494 ( .A(KEYINPUT33), .B(KEYINPUT72), .ZN(n366) );
  INV_X1 U495 ( .A(KEYINPUT84), .ZN(n512) );
  OR2_X1 U496 ( .A1(n616), .A2(n667), .ZN(n370) );
  AND2_X1 U497 ( .A1(KEYINPUT84), .A2(KEYINPUT100), .ZN(n371) );
  AND2_X1 U498 ( .A1(n626), .A2(G953), .ZN(n729) );
  INV_X1 U499 ( .A(n729), .ZN(n391) );
  XNOR2_X1 U500 ( .A(n372), .B(n437), .ZN(n441) );
  OR2_X2 U501 ( .A1(n495), .A2(n358), .ZN(n374) );
  XNOR2_X2 U502 ( .A(n375), .B(n435), .ZN(n495) );
  XNOR2_X2 U503 ( .A(n436), .B(KEYINPUT3), .ZN(n375) );
  XNOR2_X1 U504 ( .A(n376), .B(n403), .ZN(n437) );
  XNOR2_X1 U505 ( .A(n378), .B(n377), .ZN(n376) );
  XNOR2_X1 U506 ( .A(n380), .B(n462), .ZN(n378) );
  INV_X1 U507 ( .A(KEYINPUT17), .ZN(n381) );
  NOR2_X1 U508 ( .A1(n561), .A2(n560), .ZN(n422) );
  NAND2_X1 U509 ( .A1(n348), .A2(n349), .ZN(n383) );
  NAND2_X1 U510 ( .A1(n411), .A2(n408), .ZN(n636) );
  NAND2_X1 U511 ( .A1(n427), .A2(n360), .ZN(n426) );
  NOR2_X1 U512 ( .A1(n384), .A2(n729), .ZN(G63) );
  XNOR2_X1 U513 ( .A(n385), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U514 ( .A1(n393), .A2(n391), .ZN(n385) );
  XNOR2_X1 U515 ( .A(n387), .B(n386), .ZN(G51) );
  NAND2_X1 U516 ( .A1(n390), .A2(n391), .ZN(n387) );
  XNOR2_X1 U517 ( .A(n389), .B(n388), .ZN(G60) );
  NAND2_X1 U518 ( .A1(n392), .A2(n391), .ZN(n389) );
  XNOR2_X1 U519 ( .A(n634), .B(n368), .ZN(n390) );
  XNOR2_X1 U520 ( .A(n630), .B(n367), .ZN(n392) );
  XNOR2_X1 U521 ( .A(n625), .B(n369), .ZN(n393) );
  AND2_X2 U522 ( .A1(n394), .A2(n412), .ZN(n411) );
  NAND2_X1 U523 ( .A1(n557), .A2(n556), .ZN(n402) );
  NOR2_X1 U524 ( .A1(n660), .A2(n396), .ZN(n605) );
  XNOR2_X2 U525 ( .A(n433), .B(G128), .ZN(n474) );
  NAND2_X1 U526 ( .A1(n404), .A2(n563), .ZN(n421) );
  NAND2_X1 U527 ( .A1(n561), .A2(n405), .ZN(n404) );
  NOR2_X1 U528 ( .A1(n672), .A2(n356), .ZN(n710) );
  INV_X1 U529 ( .A(n511), .ZN(n413) );
  NAND2_X1 U530 ( .A1(n511), .A2(n425), .ZN(n414) );
  NAND2_X1 U531 ( .A1(n621), .A2(n432), .ZN(n668) );
  NAND2_X1 U532 ( .A1(n603), .A2(n689), .ZN(n574) );
  NOR2_X1 U533 ( .A1(n422), .A2(n421), .ZN(n564) );
  NOR2_X2 U534 ( .A1(n589), .A2(n452), .ZN(n423) );
  XNOR2_X1 U535 ( .A(n597), .B(KEYINPUT19), .ZN(n589) );
  NOR2_X2 U536 ( .A1(n759), .A2(n754), .ZN(n588) );
  AND2_X1 U537 ( .A1(n675), .A2(n512), .ZN(n425) );
  AND2_X1 U538 ( .A1(n615), .A2(KEYINPUT82), .ZN(n429) );
  INV_X1 U539 ( .A(n444), .ZN(n573) );
  XNOR2_X2 U540 ( .A(n430), .B(n363), .ZN(n444) );
  NAND2_X1 U541 ( .A1(n631), .A2(n616), .ZN(n430) );
  XNOR2_X1 U542 ( .A(n441), .B(n505), .ZN(n631) );
  AND2_X1 U543 ( .A1(n603), .A2(n602), .ZN(n431) );
  AND2_X1 U544 ( .A1(n757), .A2(n662), .ZN(n432) );
  XNOR2_X1 U545 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U546 ( .A(n505), .B(n504), .ZN(n507) );
  INV_X1 U547 ( .A(KEYINPUT76), .ZN(n572) );
  INV_X1 U548 ( .A(n668), .ZN(n744) );
  NOR2_X1 U549 ( .A1(n675), .A2(n600), .ZN(n660) );
  NAND2_X1 U550 ( .A1(G224), .A2(n745), .ZN(n434) );
  XNOR2_X2 U551 ( .A(G113), .B(KEYINPUT70), .ZN(n436) );
  INV_X1 U552 ( .A(G902), .ZN(n497) );
  INV_X1 U553 ( .A(G237), .ZN(n442) );
  NAND2_X1 U554 ( .A1(n497), .A2(n442), .ZN(n443) );
  NAND2_X1 U555 ( .A1(n443), .A2(G214), .ZN(n688) );
  NAND2_X1 U556 ( .A1(n444), .A2(n688), .ZN(n446) );
  INV_X1 U557 ( .A(KEYINPUT88), .ZN(n445) );
  XNOR2_X1 U558 ( .A(n446), .B(n445), .ZN(n597) );
  NAND2_X1 U559 ( .A1(G234), .A2(G237), .ZN(n447) );
  XNOR2_X1 U560 ( .A(n447), .B(KEYINPUT14), .ZN(n706) );
  NAND2_X1 U561 ( .A1(G952), .A2(n745), .ZN(n449) );
  NAND2_X1 U562 ( .A1(G953), .A2(G902), .ZN(n448) );
  NAND2_X1 U563 ( .A1(n449), .A2(n448), .ZN(n450) );
  NAND2_X1 U564 ( .A1(n706), .A2(n450), .ZN(n566) );
  AND2_X1 U565 ( .A1(G953), .A2(G898), .ZN(n451) );
  OR2_X1 U566 ( .A1(n566), .A2(n451), .ZN(n452) );
  XNOR2_X1 U567 ( .A(KEYINPUT13), .B(G475), .ZN(n465) );
  XNOR2_X1 U568 ( .A(G143), .B(G131), .ZN(n453) );
  XNOR2_X1 U569 ( .A(n454), .B(n453), .ZN(n458) );
  XNOR2_X1 U570 ( .A(n456), .B(n455), .ZN(n457) );
  XOR2_X1 U571 ( .A(n458), .B(n457), .Z(n460) );
  NAND2_X1 U572 ( .A1(G214), .A2(n490), .ZN(n459) );
  XNOR2_X1 U573 ( .A(n460), .B(n459), .ZN(n463) );
  XNOR2_X1 U574 ( .A(n463), .B(n742), .ZN(n627) );
  NOR2_X1 U575 ( .A1(G902), .A2(n627), .ZN(n464) );
  XOR2_X1 U576 ( .A(n465), .B(n464), .Z(n555) );
  XNOR2_X1 U577 ( .A(n466), .B(KEYINPUT96), .ZN(n469) );
  XNOR2_X1 U578 ( .A(n362), .B(n467), .ZN(n468) );
  XOR2_X1 U579 ( .A(n469), .B(n468), .Z(n472) );
  NAND2_X1 U580 ( .A1(G234), .A2(n745), .ZN(n470) );
  NAND2_X1 U581 ( .A1(G217), .A2(n513), .ZN(n471) );
  XNOR2_X1 U582 ( .A(n472), .B(n471), .ZN(n475) );
  XOR2_X1 U583 ( .A(n475), .B(n488), .Z(n722) );
  NOR2_X1 U584 ( .A1(n722), .A2(G902), .ZN(n478) );
  XNOR2_X1 U585 ( .A(G478), .B(KEYINPUT97), .ZN(n476) );
  XNOR2_X1 U586 ( .A(n476), .B(KEYINPUT98), .ZN(n477) );
  NAND2_X1 U587 ( .A1(n555), .A2(n554), .ZN(n691) );
  NAND2_X1 U588 ( .A1(n616), .A2(G234), .ZN(n479) );
  XNOR2_X1 U589 ( .A(n479), .B(KEYINPUT20), .ZN(n521) );
  NAND2_X1 U590 ( .A1(G221), .A2(n521), .ZN(n480) );
  XNOR2_X1 U591 ( .A(KEYINPUT21), .B(n480), .ZN(n678) );
  NOR2_X1 U592 ( .A1(n691), .A2(n678), .ZN(n481) );
  XOR2_X1 U593 ( .A(n481), .B(KEYINPUT99), .Z(n482) );
  INV_X1 U594 ( .A(KEYINPUT74), .ZN(n483) );
  XNOR2_X1 U595 ( .A(n487), .B(n486), .ZN(n489) );
  NAND2_X1 U596 ( .A1(n490), .A2(G210), .ZN(n491) );
  XNOR2_X1 U597 ( .A(n491), .B(G101), .ZN(n493) );
  XOR2_X1 U598 ( .A(KEYINPUT5), .B(KEYINPUT91), .Z(n492) );
  XNOR2_X1 U599 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U600 ( .A(n495), .B(n494), .ZN(n496) );
  XNOR2_X1 U601 ( .A(n506), .B(n496), .ZN(n624) );
  NAND2_X1 U602 ( .A1(n624), .A2(n497), .ZN(n499) );
  XOR2_X1 U603 ( .A(G472), .B(KEYINPUT73), .Z(n498) );
  INV_X1 U604 ( .A(KEYINPUT6), .ZN(n500) );
  XNOR2_X1 U605 ( .A(n569), .B(n500), .ZN(n594) );
  INV_X1 U606 ( .A(n594), .ZN(n501) );
  NAND2_X1 U607 ( .A1(n543), .A2(n501), .ZN(n538) );
  NAND2_X1 U608 ( .A1(n745), .A2(G227), .ZN(n503) );
  INV_X1 U609 ( .A(G140), .ZN(n502) );
  XNOR2_X1 U610 ( .A(n506), .B(n507), .ZN(n715) );
  NOR2_X1 U611 ( .A1(G902), .A2(n715), .ZN(n510) );
  XNOR2_X1 U612 ( .A(G469), .B(KEYINPUT68), .ZN(n508) );
  XOR2_X1 U613 ( .A(n508), .B(KEYINPUT69), .Z(n509) );
  XNOR2_X2 U614 ( .A(n510), .B(n509), .ZN(n577) );
  XNOR2_X2 U615 ( .A(n577), .B(KEYINPUT1), .ZN(n675) );
  XNOR2_X1 U616 ( .A(n515), .B(n514), .ZN(n520) );
  XOR2_X1 U617 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n517) );
  XNOR2_X1 U618 ( .A(n517), .B(n516), .ZN(n518) );
  NAND2_X1 U619 ( .A1(n521), .A2(G217), .ZN(n523) );
  XOR2_X1 U620 ( .A(KEYINPUT90), .B(KEYINPUT25), .Z(n522) );
  XNOR2_X1 U621 ( .A(n523), .B(n522), .ZN(n524) );
  NOR2_X1 U622 ( .A1(n675), .A2(n674), .ZN(n550) );
  INV_X1 U623 ( .A(n395), .ZN(n581) );
  NAND2_X1 U624 ( .A1(n550), .A2(n395), .ZN(n683) );
  BUF_X1 U625 ( .A(n527), .Z(n528) );
  INV_X1 U626 ( .A(n528), .ZN(n533) );
  OR2_X1 U627 ( .A1(n683), .A2(n533), .ZN(n531) );
  XNOR2_X1 U628 ( .A(KEYINPUT93), .B(KEYINPUT31), .ZN(n529) );
  XNOR2_X1 U629 ( .A(n529), .B(KEYINPUT92), .ZN(n530) );
  XNOR2_X1 U630 ( .A(n531), .B(n530), .ZN(n657) );
  NAND2_X1 U631 ( .A1(n571), .A2(n581), .ZN(n532) );
  OR2_X1 U632 ( .A1(n533), .A2(n532), .ZN(n641) );
  NAND2_X1 U633 ( .A1(n657), .A2(n641), .ZN(n535) );
  NOR2_X1 U634 ( .A1(n555), .A2(n534), .ZN(n651) );
  NAND2_X1 U635 ( .A1(n555), .A2(n534), .ZN(n656) );
  INV_X1 U636 ( .A(n656), .ZN(n646) );
  OR2_X1 U637 ( .A1(n651), .A2(n646), .ZN(n692) );
  NAND2_X1 U638 ( .A1(n535), .A2(n692), .ZN(n536) );
  NAND2_X1 U639 ( .A1(n636), .A2(n536), .ZN(n537) );
  XNOR2_X1 U640 ( .A(n537), .B(KEYINPUT101), .ZN(n565) );
  INV_X1 U641 ( .A(n677), .ZN(n544) );
  NOR2_X1 U642 ( .A1(n675), .A2(n544), .ZN(n539) );
  XNOR2_X1 U643 ( .A(KEYINPUT79), .B(KEYINPUT32), .ZN(n540) );
  XNOR2_X1 U644 ( .A(n540), .B(KEYINPUT64), .ZN(n541) );
  BUF_X1 U645 ( .A(n543), .Z(n547) );
  NOR2_X1 U646 ( .A1(n395), .A2(n544), .ZN(n545) );
  AND2_X1 U647 ( .A1(n675), .A2(n545), .ZN(n546) );
  NAND2_X1 U648 ( .A1(n547), .A2(n546), .ZN(n645) );
  INV_X1 U649 ( .A(n645), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n550), .A2(n594), .ZN(n551) );
  NAND2_X1 U651 ( .A1(n699), .A2(n528), .ZN(n553) );
  INV_X1 U652 ( .A(KEYINPUT34), .ZN(n552) );
  XNOR2_X1 U653 ( .A(n553), .B(n552), .ZN(n557) );
  OR2_X1 U654 ( .A1(n555), .A2(n554), .ZN(n601) );
  INV_X1 U655 ( .A(n601), .ZN(n556) );
  INV_X1 U656 ( .A(KEYINPUT35), .ZN(n558) );
  NOR2_X1 U657 ( .A1(KEYINPUT85), .A2(KEYINPUT44), .ZN(n559) );
  NAND2_X1 U658 ( .A1(n758), .A2(n559), .ZN(n560) );
  INV_X1 U659 ( .A(n758), .ZN(n562) );
  NAND2_X1 U660 ( .A1(n562), .A2(KEYINPUT44), .ZN(n563) );
  INV_X1 U661 ( .A(n566), .ZN(n568) );
  NAND2_X1 U662 ( .A1(G953), .A2(G900), .ZN(n567) );
  NAND2_X1 U663 ( .A1(n568), .A2(n567), .ZN(n578) );
  NAND2_X1 U664 ( .A1(n569), .A2(n688), .ZN(n570) );
  XOR2_X1 U665 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n575) );
  XOR2_X1 U666 ( .A(KEYINPUT106), .B(KEYINPUT42), .Z(n587) );
  XOR2_X1 U667 ( .A(n577), .B(KEYINPUT104), .Z(n584) );
  NOR2_X1 U668 ( .A1(n678), .A2(n578), .ZN(n579) );
  NAND2_X1 U669 ( .A1(n677), .A2(n579), .ZN(n580) );
  XOR2_X1 U670 ( .A(n580), .B(KEYINPUT67), .Z(n596) );
  XNOR2_X1 U671 ( .A(n582), .B(KEYINPUT28), .ZN(n583) );
  NAND2_X1 U672 ( .A1(n584), .A2(n583), .ZN(n591) );
  NAND2_X1 U673 ( .A1(n689), .A2(n688), .ZN(n693) );
  NOR2_X1 U674 ( .A1(n691), .A2(n693), .ZN(n585) );
  XNOR2_X1 U675 ( .A(KEYINPUT41), .B(n585), .ZN(n673) );
  NOR2_X1 U676 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n593) );
  BUF_X1 U677 ( .A(n589), .Z(n590) );
  NOR2_X1 U678 ( .A1(n591), .A2(n590), .ZN(n652) );
  NAND2_X1 U679 ( .A1(n652), .A2(n692), .ZN(n592) );
  XNOR2_X1 U680 ( .A(n593), .B(n592), .ZN(n606) );
  NAND2_X1 U681 ( .A1(KEYINPUT47), .A2(KEYINPUT75), .ZN(n604) );
  NAND2_X1 U682 ( .A1(n594), .A2(n651), .ZN(n595) );
  AND2_X1 U683 ( .A1(n597), .A2(n607), .ZN(n599) );
  NOR2_X1 U684 ( .A1(n573), .A2(n601), .ZN(n602) );
  NAND2_X1 U685 ( .A1(n607), .A2(n688), .ZN(n608) );
  XOR2_X1 U686 ( .A(KEYINPUT102), .B(n608), .Z(n609) );
  NAND2_X1 U687 ( .A1(n609), .A2(n675), .ZN(n610) );
  XOR2_X1 U688 ( .A(KEYINPUT43), .B(n610), .Z(n612) );
  INV_X1 U689 ( .A(n573), .ZN(n611) );
  NOR2_X1 U690 ( .A1(n612), .A2(n611), .ZN(n613) );
  XNOR2_X1 U691 ( .A(n613), .B(KEYINPUT103), .ZN(n757) );
  NAND2_X1 U692 ( .A1(n614), .A2(n646), .ZN(n662) );
  INV_X1 U693 ( .A(KEYINPUT2), .ZN(n667) );
  NAND2_X1 U694 ( .A1(KEYINPUT2), .A2(n662), .ZN(n618) );
  XOR2_X1 U695 ( .A(KEYINPUT80), .B(n618), .Z(n619) );
  AND2_X1 U696 ( .A1(n757), .A2(n619), .ZN(n620) );
  AND2_X1 U697 ( .A1(n621), .A2(n620), .ZN(n622) );
  NAND2_X1 U698 ( .A1(n724), .A2(G472), .ZN(n625) );
  INV_X1 U699 ( .A(G952), .ZN(n626) );
  NAND2_X1 U700 ( .A1(n382), .A2(G475), .ZN(n630) );
  XOR2_X1 U701 ( .A(KEYINPUT121), .B(KEYINPUT59), .Z(n629) );
  XNOR2_X1 U702 ( .A(n627), .B(KEYINPUT120), .ZN(n628) );
  NAND2_X1 U703 ( .A1(n724), .A2(G210), .ZN(n634) );
  BUF_X1 U704 ( .A(n631), .Z(n632) );
  XNOR2_X1 U705 ( .A(KEYINPUT54), .B(KEYINPUT55), .ZN(n633) );
  XOR2_X1 U706 ( .A(n635), .B(G119), .Z(G21) );
  XNOR2_X1 U707 ( .A(n383), .B(G101), .ZN(G3) );
  INV_X1 U708 ( .A(n651), .ZN(n654) );
  NOR2_X1 U709 ( .A1(n641), .A2(n654), .ZN(n638) );
  XNOR2_X1 U710 ( .A(G104), .B(KEYINPUT107), .ZN(n637) );
  XNOR2_X1 U711 ( .A(n638), .B(n637), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n640) );
  XNOR2_X1 U713 ( .A(G107), .B(KEYINPUT108), .ZN(n639) );
  XNOR2_X1 U714 ( .A(n640), .B(n639), .ZN(n643) );
  NOR2_X1 U715 ( .A1(n641), .A2(n656), .ZN(n642) );
  XOR2_X1 U716 ( .A(n643), .B(n642), .Z(G9) );
  XOR2_X1 U717 ( .A(G110), .B(KEYINPUT109), .Z(n644) );
  XNOR2_X1 U718 ( .A(n645), .B(n644), .ZN(G12) );
  XOR2_X1 U719 ( .A(KEYINPUT110), .B(KEYINPUT29), .Z(n648) );
  NAND2_X1 U720 ( .A1(n652), .A2(n646), .ZN(n647) );
  XNOR2_X1 U721 ( .A(n648), .B(n647), .ZN(n649) );
  XNOR2_X1 U722 ( .A(G128), .B(n649), .ZN(G30) );
  XNOR2_X1 U723 ( .A(G143), .B(n431), .ZN(n650) );
  XNOR2_X1 U724 ( .A(n650), .B(KEYINPUT111), .ZN(G45) );
  NAND2_X1 U725 ( .A1(n652), .A2(n651), .ZN(n653) );
  XNOR2_X1 U726 ( .A(G146), .B(n653), .ZN(G48) );
  NOR2_X1 U727 ( .A1(n657), .A2(n654), .ZN(n655) );
  XOR2_X1 U728 ( .A(G113), .B(n655), .Z(G15) );
  NOR2_X1 U729 ( .A1(n657), .A2(n656), .ZN(n658) );
  XOR2_X1 U730 ( .A(KEYINPUT112), .B(n658), .Z(n659) );
  XNOR2_X1 U731 ( .A(G116), .B(n659), .ZN(G18) );
  XNOR2_X1 U732 ( .A(G125), .B(n660), .ZN(n661) );
  XNOR2_X1 U733 ( .A(n661), .B(KEYINPUT37), .ZN(G27) );
  INV_X1 U734 ( .A(n662), .ZN(n663) );
  XOR2_X1 U735 ( .A(G134), .B(n663), .Z(G36) );
  XOR2_X1 U736 ( .A(KEYINPUT118), .B(KEYINPUT53), .Z(n714) );
  INV_X1 U737 ( .A(n699), .ZN(n664) );
  NOR2_X1 U738 ( .A1(n664), .A2(n673), .ZN(n665) );
  NOR2_X1 U739 ( .A1(G953), .A2(n665), .ZN(n712) );
  INV_X1 U740 ( .A(n666), .ZN(n734) );
  NAND2_X1 U741 ( .A1(n734), .A2(n667), .ZN(n671) );
  NOR2_X1 U742 ( .A1(KEYINPUT2), .A2(n744), .ZN(n669) );
  XNOR2_X1 U743 ( .A(n669), .B(KEYINPUT81), .ZN(n670) );
  NAND2_X1 U744 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n705) );
  INV_X1 U746 ( .A(n673), .ZN(n687) );
  NAND2_X1 U747 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U748 ( .A(n676), .B(KEYINPUT50), .ZN(n682) );
  AND2_X1 U749 ( .A1(n678), .A2(n677), .ZN(n679) );
  XOR2_X1 U750 ( .A(KEYINPUT49), .B(n679), .Z(n680) );
  NOR2_X1 U751 ( .A1(n395), .A2(n680), .ZN(n681) );
  NAND2_X1 U752 ( .A1(n682), .A2(n681), .ZN(n684) );
  NAND2_X1 U753 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U754 ( .A(KEYINPUT51), .B(n685), .Z(n686) );
  NAND2_X1 U755 ( .A1(n687), .A2(n686), .ZN(n702) );
  NOR2_X1 U756 ( .A1(n689), .A2(n688), .ZN(n690) );
  NOR2_X1 U757 ( .A1(n691), .A2(n690), .ZN(n697) );
  INV_X1 U758 ( .A(n692), .ZN(n694) );
  NOR2_X1 U759 ( .A1(n694), .A2(n693), .ZN(n695) );
  XNOR2_X1 U760 ( .A(n695), .B(KEYINPUT114), .ZN(n696) );
  NOR2_X1 U761 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U762 ( .A(n698), .B(KEYINPUT115), .ZN(n700) );
  NAND2_X1 U763 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U764 ( .A1(n702), .A2(n701), .ZN(n703) );
  XNOR2_X1 U765 ( .A(n703), .B(KEYINPUT52), .ZN(n704) );
  XNOR2_X1 U766 ( .A(n705), .B(n704), .ZN(n708) );
  NAND2_X1 U767 ( .A1(n706), .A2(G952), .ZN(n707) );
  NOR2_X1 U768 ( .A1(n708), .A2(n707), .ZN(n709) );
  NOR2_X1 U769 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U770 ( .A1(n712), .A2(n711), .ZN(n713) );
  XNOR2_X1 U771 ( .A(n714), .B(n713), .ZN(G75) );
  NAND2_X1 U772 ( .A1(n721), .A2(G469), .ZN(n719) );
  XNOR2_X1 U773 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n717) );
  XNOR2_X1 U774 ( .A(n715), .B(KEYINPUT57), .ZN(n716) );
  XNOR2_X1 U775 ( .A(n717), .B(n716), .ZN(n718) );
  XNOR2_X1 U776 ( .A(n719), .B(n718), .ZN(n720) );
  NOR2_X1 U777 ( .A1(n729), .A2(n720), .ZN(G54) );
  NAND2_X1 U778 ( .A1(n721), .A2(G478), .ZN(n723) );
  NAND2_X1 U779 ( .A1(n721), .A2(G217), .ZN(n727) );
  XNOR2_X1 U780 ( .A(n725), .B(KEYINPUT122), .ZN(n726) );
  XNOR2_X1 U781 ( .A(n727), .B(n726), .ZN(n728) );
  NOR2_X1 U782 ( .A1(n729), .A2(n728), .ZN(G66) );
  XNOR2_X1 U783 ( .A(n730), .B(KEYINPUT124), .ZN(n731) );
  NOR2_X1 U784 ( .A1(G898), .A2(n745), .ZN(n732) );
  NOR2_X1 U785 ( .A1(n733), .A2(n732), .ZN(n741) );
  NOR2_X1 U786 ( .A1(n734), .A2(G953), .ZN(n735) );
  XNOR2_X1 U787 ( .A(n735), .B(KEYINPUT123), .ZN(n739) );
  NAND2_X1 U788 ( .A1(G953), .A2(G224), .ZN(n736) );
  XNOR2_X1 U789 ( .A(KEYINPUT61), .B(n736), .ZN(n737) );
  NAND2_X1 U790 ( .A1(n737), .A2(G898), .ZN(n738) );
  NAND2_X1 U791 ( .A1(n739), .A2(n738), .ZN(n740) );
  XNOR2_X1 U792 ( .A(n741), .B(n740), .ZN(G69) );
  XOR2_X1 U793 ( .A(n743), .B(n742), .Z(n747) );
  XNOR2_X1 U794 ( .A(n744), .B(n747), .ZN(n746) );
  NAND2_X1 U795 ( .A1(n746), .A2(n745), .ZN(n753) );
  XNOR2_X1 U796 ( .A(n747), .B(G227), .ZN(n748) );
  XNOR2_X1 U797 ( .A(n748), .B(KEYINPUT125), .ZN(n749) );
  NAND2_X1 U798 ( .A1(n749), .A2(G900), .ZN(n750) );
  XNOR2_X1 U799 ( .A(KEYINPUT126), .B(n750), .ZN(n751) );
  NAND2_X1 U800 ( .A1(G953), .A2(n751), .ZN(n752) );
  NAND2_X1 U801 ( .A1(n753), .A2(n752), .ZN(G72) );
  XNOR2_X1 U802 ( .A(G137), .B(n754), .ZN(n755) );
  XNOR2_X1 U803 ( .A(n755), .B(KEYINPUT127), .ZN(G39) );
  XOR2_X1 U804 ( .A(G140), .B(KEYINPUT113), .Z(n756) );
  XNOR2_X1 U805 ( .A(n757), .B(n756), .ZN(G42) );
  XNOR2_X1 U806 ( .A(G122), .B(n758), .ZN(G24) );
  XOR2_X1 U807 ( .A(n759), .B(G131), .Z(G33) );
endmodule

