//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 1 1 0 0 0 1 1 1 1 1 1 0 0 0 0 0 1 1 1 1 0 1 1 0 1 0 1 0 0 1 1 1 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 1 0 0 0 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:48 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n714, new_n715, new_n716, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n741, new_n742,
    new_n743, new_n744, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n851, new_n852, new_n854, new_n855, new_n856, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n935, new_n936, new_n937, new_n939, new_n940, new_n941, new_n943,
    new_n944, new_n945, new_n946, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  XOR2_X1   g001(.A(G197gat), .B(G204gat), .Z(new_n203));
  NAND2_X1  g002(.A1(KEYINPUT69), .A2(KEYINPUT22), .ZN(new_n204));
  INV_X1    g003(.A(KEYINPUT69), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT22), .ZN(new_n206));
  AOI22_X1  g005(.A1(new_n205), .A2(new_n206), .B1(G211gat), .B2(G218gat), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n203), .B1(new_n204), .B2(new_n207), .ZN(new_n208));
  XOR2_X1   g007(.A(G211gat), .B(G218gat), .Z(new_n209));
  NAND2_X1  g008(.A1(new_n209), .A2(KEYINPUT70), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n208), .B(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(G148gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n212), .A2(G141gat), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT74), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n212), .A2(KEYINPUT74), .A3(G141gat), .ZN(new_n216));
  INV_X1    g015(.A(G141gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(G148gat), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n215), .A2(new_n216), .A3(new_n218), .ZN(new_n219));
  NAND2_X1  g018(.A1(G155gat), .A2(G162gat), .ZN(new_n220));
  INV_X1    g019(.A(G155gat), .ZN(new_n221));
  INV_X1    g020(.A(G162gat), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  OAI21_X1  g022(.A(new_n220), .B1(new_n223), .B2(KEYINPUT2), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  XOR2_X1   g024(.A(KEYINPUT73), .B(KEYINPUT2), .Z(new_n226));
  NAND2_X1  g025(.A1(new_n213), .A2(new_n218), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT72), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND3_X1  g028(.A1(new_n213), .A2(new_n218), .A3(KEYINPUT72), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n226), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n223), .A2(new_n220), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n225), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT3), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g035(.A(KEYINPUT29), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n211), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n208), .A2(new_n209), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n208), .A2(new_n209), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n239), .A2(new_n237), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g040(.A(new_n234), .B1(new_n241), .B2(new_n235), .ZN(new_n242));
  INV_X1    g041(.A(G228gat), .ZN(new_n243));
  INV_X1    g042(.A(G233gat), .ZN(new_n244));
  OAI22_X1  g043(.A1(new_n238), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n245), .B(KEYINPUT79), .ZN(new_n246));
  INV_X1    g045(.A(G22gat), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n211), .A2(new_n237), .ZN(new_n248));
  AOI21_X1  g047(.A(new_n234), .B1(new_n248), .B2(new_n235), .ZN(new_n249));
  OR4_X1    g048(.A1(new_n243), .A2(new_n249), .A3(new_n238), .A4(new_n244), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n246), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(new_n247), .B1(new_n246), .B2(new_n250), .ZN(new_n253));
  OAI21_X1  g052(.A(G78gat), .B1(new_n252), .B2(new_n253), .ZN(new_n254));
  INV_X1    g053(.A(new_n253), .ZN(new_n255));
  INV_X1    g054(.A(G78gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n255), .A2(new_n256), .A3(new_n251), .ZN(new_n257));
  XNOR2_X1  g056(.A(KEYINPUT31), .B(G50gat), .ZN(new_n258));
  XOR2_X1   g057(.A(new_n258), .B(G106gat), .Z(new_n259));
  NAND3_X1  g058(.A1(new_n254), .A2(new_n257), .A3(new_n259), .ZN(new_n260));
  INV_X1    g059(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g060(.A(new_n259), .B1(new_n254), .B2(new_n257), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n202), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n254), .A2(new_n257), .ZN(new_n264));
  INV_X1    g063(.A(new_n259), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n266), .A2(KEYINPUT80), .A3(new_n260), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n263), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n233), .A2(KEYINPUT3), .ZN(new_n269));
  OR2_X1    g068(.A1(new_n269), .A2(KEYINPUT75), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n269), .A2(KEYINPUT75), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  XNOR2_X1  g071(.A(G127gat), .B(G134gat), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT64), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n273), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(G113gat), .ZN(new_n276));
  INV_X1    g075(.A(G120gat), .ZN(new_n277));
  AOI21_X1  g076(.A(KEYINPUT1), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n278), .B1(new_n276), .B2(new_n277), .ZN(new_n279));
  NAND2_X1  g078(.A1(new_n275), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g079(.A(KEYINPUT65), .B(G113gat), .Z(new_n281));
  OAI211_X1 g080(.A(new_n278), .B(new_n273), .C1(new_n281), .C2(new_n277), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n280), .A2(new_n282), .ZN(new_n283));
  NAND3_X1  g082(.A1(new_n272), .A2(new_n283), .A3(new_n236), .ZN(new_n284));
  NOR2_X1   g083(.A1(new_n283), .A2(new_n233), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT4), .ZN(new_n286));
  XNOR2_X1  g085(.A(new_n285), .B(new_n286), .ZN(new_n287));
  NAND2_X1  g086(.A1(G225gat), .A2(G233gat), .ZN(new_n288));
  XOR2_X1   g087(.A(KEYINPUT76), .B(KEYINPUT5), .Z(new_n289));
  INV_X1    g088(.A(new_n289), .ZN(new_n290));
  NAND4_X1  g089(.A1(new_n284), .A2(new_n287), .A3(new_n288), .A4(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(G1gat), .B(G29gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n292), .B(KEYINPUT0), .ZN(new_n293));
  XNOR2_X1  g092(.A(G57gat), .B(G85gat), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  INV_X1    g094(.A(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n236), .A2(new_n283), .ZN(new_n297));
  AOI21_X1  g096(.A(new_n297), .B1(new_n271), .B2(new_n270), .ZN(new_n298));
  XNOR2_X1  g097(.A(new_n285), .B(KEYINPUT4), .ZN(new_n299));
  INV_X1    g098(.A(new_n288), .ZN(new_n300));
  NOR3_X1   g099(.A1(new_n298), .A2(new_n299), .A3(new_n300), .ZN(new_n301));
  XNOR2_X1  g100(.A(new_n283), .B(new_n233), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n289), .B1(new_n302), .B2(new_n300), .ZN(new_n303));
  OAI211_X1 g102(.A(new_n291), .B(new_n296), .C1(new_n301), .C2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT6), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  AND2_X1   g105(.A1(new_n304), .A2(new_n305), .ZN(new_n307));
  OAI21_X1  g106(.A(new_n291), .B1(new_n301), .B2(new_n303), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT77), .ZN(new_n309));
  AND3_X1   g108(.A1(new_n308), .A2(new_n309), .A3(new_n295), .ZN(new_n310));
  AOI21_X1  g109(.A(new_n309), .B1(new_n308), .B2(new_n295), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n307), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT78), .ZN(new_n313));
  AOI21_X1  g112(.A(new_n306), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  OAI211_X1 g113(.A(new_n307), .B(KEYINPUT78), .C1(new_n310), .C2(new_n311), .ZN(new_n315));
  NAND2_X1  g114(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(G226gat), .A2(G233gat), .ZN(new_n318));
  INV_X1    g117(.A(G169gat), .ZN(new_n319));
  INV_X1    g118(.A(G176gat), .ZN(new_n320));
  NOR2_X1   g119(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NOR2_X1   g120(.A1(G169gat), .A2(G176gat), .ZN(new_n322));
  OR3_X1    g121(.A1(new_n321), .A2(KEYINPUT26), .A3(new_n322), .ZN(new_n323));
  AOI22_X1  g122(.A1(new_n322), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n324));
  XNOR2_X1  g123(.A(KEYINPUT27), .B(G183gat), .ZN(new_n325));
  INV_X1    g124(.A(G190gat), .ZN(new_n326));
  AND3_X1   g125(.A1(new_n325), .A2(KEYINPUT28), .A3(new_n326), .ZN(new_n327));
  AOI21_X1  g126(.A(KEYINPUT28), .B1(new_n325), .B2(new_n326), .ZN(new_n328));
  OAI211_X1 g127(.A(new_n323), .B(new_n324), .C1(new_n327), .C2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT23), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n322), .B(new_n330), .ZN(new_n331));
  NAND2_X1  g130(.A1(G183gat), .A2(G190gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n332), .A2(KEYINPUT24), .ZN(new_n333));
  NOR2_X1   g132(.A1(new_n333), .A2(new_n321), .ZN(new_n334));
  OR2_X1    g133(.A1(G183gat), .A2(G190gat), .ZN(new_n335));
  NAND3_X1  g134(.A1(new_n335), .A2(KEYINPUT24), .A3(new_n332), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n331), .A2(new_n334), .A3(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT25), .ZN(new_n338));
  AND2_X1   g137(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  NOR2_X1   g138(.A1(new_n337), .A2(new_n338), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n329), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(new_n341), .ZN(new_n342));
  OAI21_X1  g141(.A(new_n318), .B1(new_n342), .B2(KEYINPUT29), .ZN(new_n343));
  NAND3_X1  g142(.A1(new_n341), .A2(G226gat), .A3(G233gat), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  INV_X1    g144(.A(new_n211), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n345), .A2(new_n346), .ZN(new_n347));
  XOR2_X1   g146(.A(G8gat), .B(G36gat), .Z(new_n348));
  XNOR2_X1  g147(.A(new_n348), .B(KEYINPUT71), .ZN(new_n349));
  XNOR2_X1  g148(.A(G64gat), .B(G92gat), .ZN(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  NAND3_X1  g150(.A1(new_n343), .A2(new_n211), .A3(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n347), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g152(.A(new_n353), .ZN(new_n354));
  OR2_X1    g153(.A1(new_n354), .A2(KEYINPUT30), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n354), .A2(KEYINPUT30), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n347), .A2(new_n352), .ZN(new_n357));
  INV_X1    g156(.A(new_n351), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NAND3_X1  g158(.A1(new_n355), .A2(new_n356), .A3(new_n359), .ZN(new_n360));
  OAI21_X1  g159(.A(new_n268), .B1(new_n317), .B2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n283), .ZN(new_n362));
  NAND2_X1  g161(.A1(new_n341), .A2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G227gat), .ZN(new_n364));
  NOR2_X1   g163(.A1(new_n364), .A2(new_n244), .ZN(new_n365));
  OAI211_X1 g164(.A(new_n283), .B(new_n329), .C1(new_n339), .C2(new_n340), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n363), .A2(new_n365), .A3(new_n366), .ZN(new_n367));
  XOR2_X1   g166(.A(G71gat), .B(G99gat), .Z(new_n368));
  XNOR2_X1  g167(.A(G15gat), .B(G43gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(new_n368), .B(new_n369), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n370), .A2(KEYINPUT33), .ZN(new_n371));
  NAND3_X1  g170(.A1(new_n367), .A2(KEYINPUT32), .A3(new_n371), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT66), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  NAND4_X1  g173(.A1(new_n367), .A2(KEYINPUT66), .A3(KEYINPUT32), .A4(new_n371), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT34), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n363), .A2(new_n366), .ZN(new_n378));
  INV_X1    g177(.A(new_n365), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI211_X1 g179(.A(KEYINPUT34), .B(new_n365), .C1(new_n363), .C2(new_n366), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n367), .A2(KEYINPUT32), .ZN(new_n383));
  INV_X1    g182(.A(new_n367), .ZN(new_n384));
  OAI211_X1 g183(.A(new_n383), .B(new_n370), .C1(new_n384), .C2(KEYINPUT33), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n376), .A2(new_n382), .A3(new_n385), .ZN(new_n386));
  NAND2_X1  g185(.A1(new_n386), .A2(KEYINPUT67), .ZN(new_n387));
  AOI21_X1  g186(.A(new_n382), .B1(new_n376), .B2(new_n385), .ZN(new_n388));
  NOR2_X1   g187(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  AOI211_X1 g188(.A(KEYINPUT67), .B(new_n382), .C1(new_n376), .C2(new_n385), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT36), .B1(new_n389), .B2(new_n390), .ZN(new_n391));
  NOR2_X1   g190(.A1(new_n388), .A2(KEYINPUT68), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(new_n386), .ZN(new_n393));
  INV_X1    g192(.A(KEYINPUT36), .ZN(new_n394));
  NAND4_X1  g193(.A1(new_n376), .A2(KEYINPUT68), .A3(new_n382), .A4(new_n385), .ZN(new_n395));
  NAND3_X1  g194(.A1(new_n393), .A2(new_n394), .A3(new_n395), .ZN(new_n396));
  AND2_X1   g195(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n266), .A2(new_n260), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n300), .B1(new_n298), .B2(new_n299), .ZN(new_n399));
  OAI211_X1 g198(.A(new_n399), .B(KEYINPUT39), .C1(new_n300), .C2(new_n302), .ZN(new_n400));
  OAI211_X1 g199(.A(new_n400), .B(new_n295), .C1(KEYINPUT39), .C2(new_n399), .ZN(new_n401));
  NOR2_X1   g200(.A1(KEYINPUT81), .A2(KEYINPUT40), .ZN(new_n402));
  OR2_X1    g201(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n402), .ZN(new_n404));
  AND4_X1   g203(.A1(new_n304), .A2(new_n403), .A3(new_n360), .A4(new_n404), .ZN(new_n405));
  NOR2_X1   g204(.A1(new_n398), .A2(new_n405), .ZN(new_n406));
  INV_X1    g205(.A(new_n306), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n312), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT38), .ZN(new_n409));
  NOR2_X1   g208(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n357), .A2(KEYINPUT37), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n411), .A2(new_n358), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT82), .ZN(new_n413));
  AOI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  NAND3_X1  g213(.A1(new_n411), .A2(KEYINPUT82), .A3(new_n358), .ZN(new_n415));
  AOI21_X1  g214(.A(new_n409), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  NOR3_X1   g215(.A1(new_n412), .A2(KEYINPUT38), .A3(new_n410), .ZN(new_n417));
  OR4_X1    g216(.A1(new_n354), .A2(new_n408), .A3(new_n416), .A4(new_n417), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n397), .B1(new_n406), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n361), .A2(new_n419), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n261), .A2(new_n262), .ZN(new_n421));
  OR2_X1    g220(.A1(new_n389), .A2(new_n390), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  INV_X1    g222(.A(new_n360), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n316), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g224(.A(KEYINPUT35), .B1(new_n423), .B2(new_n425), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n393), .A2(new_n395), .ZN(new_n427));
  NOR2_X1   g226(.A1(new_n360), .A2(KEYINPUT35), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n421), .A2(new_n408), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n426), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n420), .A2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n432));
  INV_X1    g231(.A(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT98), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  INV_X1    g234(.A(G71gat), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n436), .B(new_n256), .C1(new_n434), .C2(KEYINPUT9), .ZN(new_n437));
  NAND2_X1  g236(.A1(G71gat), .A2(G78gat), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  XOR2_X1   g238(.A(G57gat), .B(G64gat), .Z(new_n440));
  NAND3_X1  g239(.A1(new_n435), .A2(new_n439), .A3(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n440), .A2(new_n433), .ZN(new_n442));
  INV_X1    g241(.A(KEYINPUT96), .ZN(new_n443));
  NOR3_X1   g242(.A1(new_n443), .A2(G71gat), .A3(G78gat), .ZN(new_n444));
  AOI21_X1  g243(.A(KEYINPUT96), .B1(new_n436), .B2(new_n256), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n438), .B1(new_n444), .B2(new_n445), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT97), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n442), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  NAND3_X1  g247(.A1(new_n436), .A2(new_n256), .A3(KEYINPUT96), .ZN(new_n449));
  OAI21_X1  g248(.A(new_n443), .B1(G71gat), .B2(G78gat), .ZN(new_n450));
  AOI22_X1  g249(.A1(new_n449), .A2(new_n450), .B1(G71gat), .B2(G78gat), .ZN(new_n451));
  NOR2_X1   g250(.A1(new_n451), .A2(KEYINPUT97), .ZN(new_n452));
  OAI21_X1  g251(.A(new_n441), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT21), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  NAND2_X1  g254(.A1(G231gat), .A2(G233gat), .ZN(new_n456));
  XNOR2_X1  g255(.A(new_n455), .B(new_n456), .ZN(new_n457));
  XNOR2_X1  g256(.A(new_n457), .B(G127gat), .ZN(new_n458));
  XOR2_X1   g257(.A(KEYINPUT90), .B(G8gat), .Z(new_n459));
  XNOR2_X1  g258(.A(G15gat), .B(G22gat), .ZN(new_n460));
  INV_X1    g259(.A(G1gat), .ZN(new_n461));
  AND2_X1   g260(.A1(new_n461), .A2(KEYINPUT16), .ZN(new_n462));
  AND2_X1   g261(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  NOR2_X1   g262(.A1(new_n460), .A2(new_n461), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n459), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT91), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n460), .A2(new_n462), .ZN(new_n468));
  OAI211_X1 g267(.A(new_n468), .B(G8gat), .C1(new_n461), .C2(new_n460), .ZN(new_n469));
  OAI211_X1 g268(.A(KEYINPUT91), .B(new_n459), .C1(new_n463), .C2(new_n464), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n467), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(KEYINPUT92), .ZN(new_n472));
  INV_X1    g271(.A(KEYINPUT92), .ZN(new_n473));
  NAND4_X1  g272(.A1(new_n467), .A2(new_n473), .A3(new_n469), .A4(new_n470), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n472), .A2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n454), .B2(new_n453), .ZN(new_n476));
  XNOR2_X1  g275(.A(new_n458), .B(new_n476), .ZN(new_n477));
  XNOR2_X1  g276(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n478), .B(new_n221), .ZN(new_n479));
  XOR2_X1   g278(.A(G183gat), .B(G211gat), .Z(new_n480));
  XNOR2_X1  g279(.A(new_n479), .B(new_n480), .ZN(new_n481));
  INV_X1    g280(.A(new_n481), .ZN(new_n482));
  XNOR2_X1  g281(.A(new_n477), .B(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(G232gat), .A2(G233gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n484), .B(KEYINPUT99), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT41), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  XOR2_X1   g286(.A(G134gat), .B(G162gat), .Z(new_n488));
  XNOR2_X1  g287(.A(new_n487), .B(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g289(.A1(G85gat), .A2(G92gat), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT100), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT100), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(G85gat), .A3(G92gat), .ZN(new_n494));
  NAND3_X1  g293(.A1(new_n492), .A2(new_n494), .A3(KEYINPUT7), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT7), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n491), .A2(KEYINPUT100), .A3(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(G99gat), .A2(G106gat), .ZN(new_n498));
  INV_X1    g297(.A(G85gat), .ZN(new_n499));
  INV_X1    g298(.A(G92gat), .ZN(new_n500));
  AOI22_X1  g299(.A1(KEYINPUT8), .A2(new_n498), .B1(new_n499), .B2(new_n500), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n495), .A2(new_n497), .A3(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G99gat), .B(G106gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND4_X1  g304(.A1(new_n495), .A2(new_n503), .A3(new_n497), .A4(new_n501), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(KEYINPUT101), .A3(new_n506), .ZN(new_n507));
  AND2_X1   g306(.A1(new_n501), .A2(new_n497), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT101), .ZN(new_n509));
  NAND4_X1  g308(.A1(new_n508), .A2(new_n509), .A3(new_n503), .A4(new_n495), .ZN(new_n510));
  NAND2_X1  g309(.A1(new_n507), .A2(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  INV_X1    g311(.A(KEYINPUT87), .ZN(new_n513));
  INV_X1    g312(.A(G43gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n513), .B1(new_n514), .B2(G50gat), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n514), .A2(G50gat), .ZN(new_n516));
  INV_X1    g315(.A(G50gat), .ZN(new_n517));
  NAND3_X1  g316(.A1(new_n517), .A2(KEYINPUT87), .A3(G43gat), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n515), .A2(new_n516), .A3(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT15), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT88), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n520), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT83), .ZN(new_n526));
  NOR2_X1   g325(.A1(new_n514), .A2(G50gat), .ZN(new_n527));
  NOR2_X1   g326(.A1(new_n517), .A2(G43gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n526), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n517), .A2(G43gat), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n530), .A2(new_n516), .A3(KEYINPUT83), .ZN(new_n531));
  NAND3_X1  g330(.A1(new_n529), .A2(KEYINPUT15), .A3(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G36gat), .ZN(new_n533));
  OR2_X1    g332(.A1(KEYINPUT86), .A2(G29gat), .ZN(new_n534));
  NAND2_X1  g333(.A1(KEYINPUT86), .A2(G29gat), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n533), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT84), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g339(.A(KEYINPUT84), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  INV_X1    g341(.A(KEYINPUT14), .ZN(new_n543));
  INV_X1    g342(.A(G29gat), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n543), .A2(new_n544), .A3(new_n533), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n542), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n532), .A2(new_n537), .A3(new_n546), .ZN(new_n547));
  NOR2_X1   g346(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n548), .A2(KEYINPUT85), .A3(new_n533), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  AOI21_X1  g349(.A(KEYINPUT85), .B1(new_n548), .B2(new_n533), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  AOI21_X1  g351(.A(new_n536), .B1(new_n552), .B2(new_n542), .ZN(new_n553));
  OAI22_X1  g352(.A1(new_n525), .A2(new_n547), .B1(new_n553), .B2(new_n532), .ZN(new_n554));
  INV_X1    g353(.A(KEYINPUT17), .ZN(new_n555));
  OAI21_X1  g354(.A(new_n512), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  INV_X1    g355(.A(KEYINPUT89), .ZN(new_n557));
  XNOR2_X1  g356(.A(G43gat), .B(G50gat), .ZN(new_n558));
  AOI21_X1  g357(.A(new_n520), .B1(new_n558), .B2(KEYINPUT83), .ZN(new_n559));
  AOI21_X1  g358(.A(new_n536), .B1(new_n559), .B2(new_n529), .ZN(new_n560));
  NAND4_X1  g359(.A1(new_n560), .A2(new_n523), .A3(new_n546), .A4(new_n524), .ZN(new_n561));
  INV_X1    g360(.A(new_n542), .ZN(new_n562));
  INV_X1    g361(.A(KEYINPUT85), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n545), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n564), .A2(new_n549), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n537), .B1(new_n562), .B2(new_n565), .ZN(new_n566));
  INV_X1    g365(.A(new_n532), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  AOI211_X1 g367(.A(new_n557), .B(KEYINPUT17), .C1(new_n561), .C2(new_n568), .ZN(new_n569));
  INV_X1    g368(.A(new_n569), .ZN(new_n570));
  AOI21_X1  g369(.A(KEYINPUT89), .B1(new_n554), .B2(new_n555), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  AOI21_X1  g371(.A(new_n556), .B1(new_n570), .B2(new_n572), .ZN(new_n573));
  XNOR2_X1  g372(.A(G190gat), .B(G218gat), .ZN(new_n574));
  XOR2_X1   g373(.A(new_n574), .B(KEYINPUT102), .Z(new_n575));
  AND3_X1   g374(.A1(new_n532), .A2(new_n537), .A3(new_n546), .ZN(new_n576));
  AND3_X1   g375(.A1(new_n519), .A2(KEYINPUT88), .A3(new_n520), .ZN(new_n577));
  AOI21_X1  g376(.A(KEYINPUT88), .B1(new_n519), .B2(new_n520), .ZN(new_n578));
  NOR2_X1   g377(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  AOI22_X1  g378(.A1(new_n576), .A2(new_n579), .B1(new_n566), .B2(new_n567), .ZN(new_n580));
  OAI22_X1  g379(.A1(new_n512), .A2(new_n580), .B1(new_n486), .B2(new_n485), .ZN(new_n581));
  NOR3_X1   g380(.A1(new_n573), .A2(new_n575), .A3(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n575), .ZN(new_n583));
  INV_X1    g382(.A(new_n556), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n584), .B1(new_n569), .B2(new_n571), .ZN(new_n585));
  INV_X1    g384(.A(new_n581), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n583), .B1(new_n585), .B2(new_n586), .ZN(new_n587));
  OAI21_X1  g386(.A(new_n490), .B1(new_n582), .B2(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n575), .B1(new_n573), .B2(new_n581), .ZN(new_n589));
  NAND3_X1  g388(.A1(new_n585), .A2(new_n583), .A3(new_n586), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n589), .A2(new_n590), .A3(new_n489), .ZN(new_n591));
  AND2_X1   g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n483), .A2(new_n592), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n471), .B1(new_n580), .B2(KEYINPUT17), .ZN(new_n594));
  OAI21_X1  g393(.A(new_n594), .B1(new_n569), .B2(new_n571), .ZN(new_n595));
  NAND2_X1  g394(.A1(G229gat), .A2(G233gat), .ZN(new_n596));
  NAND3_X1  g395(.A1(new_n472), .A2(new_n474), .A3(new_n554), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n595), .A2(new_n596), .A3(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT93), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(KEYINPUT18), .ZN(new_n601));
  NAND4_X1  g400(.A1(new_n595), .A2(KEYINPUT93), .A3(new_n596), .A4(new_n597), .ZN(new_n602));
  NAND3_X1  g401(.A1(new_n600), .A2(new_n601), .A3(new_n602), .ZN(new_n603));
  NAND4_X1  g402(.A1(new_n595), .A2(KEYINPUT18), .A3(new_n596), .A4(new_n597), .ZN(new_n604));
  XNOR2_X1  g403(.A(KEYINPUT94), .B(KEYINPUT13), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n605), .B(new_n596), .ZN(new_n606));
  INV_X1    g405(.A(new_n597), .ZN(new_n607));
  AOI21_X1  g406(.A(new_n554), .B1(new_n472), .B2(new_n474), .ZN(new_n608));
  OAI21_X1  g407(.A(new_n606), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  INV_X1    g409(.A(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n603), .A2(new_n611), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT95), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n603), .A2(new_n613), .ZN(new_n614));
  XNOR2_X1  g413(.A(G113gat), .B(G141gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n615), .B(G197gat), .ZN(new_n616));
  XOR2_X1   g415(.A(KEYINPUT11), .B(G169gat), .Z(new_n617));
  XNOR2_X1  g416(.A(new_n616), .B(new_n617), .ZN(new_n618));
  XOR2_X1   g417(.A(new_n618), .B(KEYINPUT12), .Z(new_n619));
  NAND3_X1  g418(.A1(new_n612), .A2(new_n614), .A3(new_n619), .ZN(new_n620));
  AOI21_X1  g419(.A(KEYINPUT18), .B1(new_n598), .B2(new_n599), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n610), .B1(new_n621), .B2(new_n602), .ZN(new_n622));
  AOI21_X1  g421(.A(KEYINPUT95), .B1(new_n621), .B2(new_n602), .ZN(new_n623));
  INV_X1    g422(.A(new_n619), .ZN(new_n624));
  OAI21_X1  g423(.A(new_n622), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n620), .A2(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n511), .A2(new_n453), .ZN(new_n628));
  INV_X1    g427(.A(KEYINPUT103), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n506), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n630), .A2(new_n505), .ZN(new_n631));
  NAND3_X1  g430(.A1(new_n502), .A2(new_n629), .A3(new_n504), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  INV_X1    g432(.A(new_n441), .ZN(new_n634));
  AOI22_X1  g433(.A1(new_n451), .A2(KEYINPUT97), .B1(new_n433), .B2(new_n440), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n446), .A2(new_n447), .ZN(new_n636));
  AOI21_X1  g435(.A(new_n634), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n633), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g437(.A1(G230gat), .A2(G233gat), .ZN(new_n639));
  INV_X1    g438(.A(new_n639), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n628), .A2(new_n638), .A3(new_n640), .ZN(new_n641));
  AND3_X1   g440(.A1(new_n511), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n628), .A2(new_n638), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT10), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  XOR2_X1   g444(.A(new_n639), .B(KEYINPUT105), .Z(new_n646));
  OAI21_X1  g445(.A(new_n641), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g446(.A(G120gat), .B(G148gat), .Z(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT104), .ZN(new_n649));
  XNOR2_X1  g448(.A(G176gat), .B(G204gat), .ZN(new_n650));
  XOR2_X1   g449(.A(new_n649), .B(new_n650), .Z(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n647), .A2(new_n652), .ZN(new_n653));
  AOI21_X1  g452(.A(new_n453), .B1(new_n631), .B2(new_n632), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n635), .A2(new_n636), .ZN(new_n655));
  AOI22_X1  g454(.A1(new_n507), .A2(new_n510), .B1(new_n655), .B2(new_n441), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n644), .B1(new_n654), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g456(.A1(new_n511), .A2(KEYINPUT10), .A3(new_n637), .ZN(new_n658));
  NAND2_X1  g457(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n659), .A2(new_n639), .ZN(new_n660));
  AND2_X1   g459(.A1(new_n641), .A2(new_n651), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n653), .A2(new_n662), .ZN(new_n663));
  NOR3_X1   g462(.A1(new_n593), .A2(new_n627), .A3(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n431), .A2(new_n664), .ZN(new_n665));
  NOR2_X1   g464(.A1(new_n665), .A2(new_n316), .ZN(new_n666));
  XNOR2_X1  g465(.A(new_n666), .B(new_n461), .ZN(G1324gat));
  NOR2_X1   g466(.A1(new_n665), .A2(new_n424), .ZN(new_n668));
  OR2_X1    g467(.A1(new_n668), .A2(KEYINPUT106), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n668), .A2(KEYINPUT106), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(G8gat), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g470(.A(KEYINPUT16), .B(G8gat), .ZN(new_n672));
  INV_X1    g471(.A(KEYINPUT42), .ZN(new_n673));
  NOR2_X1   g472(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  AOI21_X1  g474(.A(new_n672), .B1(new_n669), .B2(new_n670), .ZN(new_n676));
  OAI211_X1 g475(.A(new_n671), .B(new_n675), .C1(new_n676), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g476(.A(new_n665), .ZN(new_n678));
  AOI21_X1  g477(.A(G15gat), .B1(new_n678), .B2(new_n427), .ZN(new_n679));
  OR2_X1    g478(.A1(new_n679), .A2(KEYINPUT107), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n679), .A2(KEYINPUT107), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT108), .ZN(new_n682));
  AND3_X1   g481(.A1(new_n391), .A2(new_n396), .A3(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n682), .B1(new_n391), .B2(new_n396), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(G15gat), .ZN(new_n686));
  XNOR2_X1  g485(.A(new_n686), .B(KEYINPUT109), .ZN(new_n687));
  AOI22_X1  g486(.A1(new_n680), .A2(new_n681), .B1(new_n678), .B2(new_n687), .ZN(G1326gat));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n678), .A2(new_n268), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(KEYINPUT110), .ZN(new_n692));
  INV_X1    g491(.A(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n691), .A2(KEYINPUT110), .ZN(new_n694));
  OAI21_X1  g493(.A(new_n690), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NAND3_X1  g495(.A1(new_n696), .A2(new_n692), .A3(new_n689), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n695), .A2(new_n697), .ZN(G1327gat));
  AOI22_X1  g497(.A1(new_n419), .A2(new_n361), .B1(new_n426), .B2(new_n429), .ZN(new_n699));
  NOR2_X1   g498(.A1(new_n699), .A2(new_n592), .ZN(new_n700));
  NOR3_X1   g499(.A1(new_n627), .A2(new_n483), .A3(new_n663), .ZN(new_n701));
  AND2_X1   g500(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n534), .A2(new_n535), .ZN(new_n703));
  INV_X1    g502(.A(new_n703), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n702), .A2(new_n317), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT45), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n700), .A2(KEYINPUT44), .ZN(new_n707));
  INV_X1    g506(.A(KEYINPUT44), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n708), .B1(new_n699), .B2(new_n592), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n710), .A2(new_n317), .A3(new_n701), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n711), .A2(new_n703), .ZN(new_n712));
  NAND2_X1  g511(.A1(new_n706), .A2(new_n712), .ZN(G1328gat));
  NAND4_X1  g512(.A1(new_n700), .A2(new_n533), .A3(new_n360), .A4(new_n701), .ZN(new_n714));
  XOR2_X1   g513(.A(new_n714), .B(KEYINPUT46), .Z(new_n715));
  AND3_X1   g514(.A1(new_n710), .A2(new_n360), .A3(new_n701), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n715), .B1(new_n716), .B2(new_n533), .ZN(G1329gat));
  NAND4_X1  g516(.A1(new_n707), .A2(new_n709), .A3(new_n397), .A4(new_n701), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(G43gat), .ZN(new_n719));
  AOI21_X1  g518(.A(G43gat), .B1(new_n393), .B2(new_n395), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n702), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g520(.A1(new_n719), .A2(KEYINPUT47), .A3(new_n721), .ZN(new_n722));
  NAND4_X1  g521(.A1(new_n707), .A2(new_n709), .A3(new_n685), .A4(new_n701), .ZN(new_n723));
  AOI22_X1  g522(.A1(new_n723), .A2(G43gat), .B1(new_n702), .B2(new_n720), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n722), .B1(new_n724), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND4_X1  g524(.A1(new_n707), .A2(new_n709), .A3(new_n398), .A4(new_n701), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n726), .A2(G50gat), .ZN(new_n727));
  INV_X1    g526(.A(new_n268), .ZN(new_n728));
  NOR2_X1   g527(.A1(new_n728), .A2(G50gat), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n702), .A2(new_n729), .ZN(new_n730));
  NAND3_X1  g529(.A1(new_n727), .A2(KEYINPUT48), .A3(new_n730), .ZN(new_n731));
  NAND4_X1  g530(.A1(new_n707), .A2(new_n709), .A3(new_n268), .A4(new_n701), .ZN(new_n732));
  AOI22_X1  g531(.A1(new_n732), .A2(G50gat), .B1(new_n702), .B2(new_n729), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n731), .B1(KEYINPUT48), .B2(new_n733), .ZN(G1331gat));
  INV_X1    g533(.A(new_n663), .ZN(new_n735));
  NOR3_X1   g534(.A1(new_n593), .A2(new_n626), .A3(new_n735), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n431), .A2(new_n736), .ZN(new_n737));
  NOR2_X1   g536(.A1(new_n737), .A2(new_n316), .ZN(new_n738));
  XOR2_X1   g537(.A(KEYINPUT111), .B(G57gat), .Z(new_n739));
  XNOR2_X1  g538(.A(new_n738), .B(new_n739), .ZN(G1332gat));
  NOR2_X1   g539(.A1(new_n737), .A2(new_n424), .ZN(new_n741));
  NOR2_X1   g540(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n742));
  AND2_X1   g541(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n741), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(new_n744), .B1(new_n741), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g544(.A(new_n685), .ZN(new_n746));
  OAI21_X1  g545(.A(G71gat), .B1(new_n737), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n427), .A2(new_n436), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n747), .B1(new_n737), .B2(new_n748), .ZN(new_n749));
  XOR2_X1   g548(.A(new_n749), .B(KEYINPUT50), .Z(G1334gat));
  NOR2_X1   g549(.A1(new_n737), .A2(new_n728), .ZN(new_n751));
  XNOR2_X1  g550(.A(new_n751), .B(new_n256), .ZN(G1335gat));
  NOR2_X1   g551(.A1(new_n483), .A2(new_n626), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n700), .A2(KEYINPUT51), .A3(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n592), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n431), .A2(new_n755), .A3(new_n753), .ZN(new_n756));
  INV_X1    g555(.A(KEYINPUT51), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  INV_X1    g557(.A(KEYINPUT113), .ZN(new_n759));
  NAND3_X1  g558(.A1(new_n754), .A2(new_n758), .A3(new_n759), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n756), .A2(KEYINPUT113), .A3(new_n757), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n317), .A2(new_n499), .A3(new_n663), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT114), .ZN(new_n763));
  NAND3_X1  g562(.A1(new_n760), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n753), .A2(new_n663), .ZN(new_n765));
  XNOR2_X1  g564(.A(new_n765), .B(KEYINPUT112), .ZN(new_n766));
  AND3_X1   g565(.A1(new_n710), .A2(new_n317), .A3(new_n766), .ZN(new_n767));
  OAI21_X1  g566(.A(new_n764), .B1(new_n767), .B2(new_n499), .ZN(G1336gat));
  NAND4_X1  g567(.A1(new_n707), .A2(new_n709), .A3(new_n360), .A4(new_n766), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n769), .A2(G92gat), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT52), .ZN(new_n771));
  NAND2_X1  g570(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NOR3_X1   g571(.A1(new_n424), .A2(G92gat), .A3(new_n735), .ZN(new_n773));
  AND3_X1   g572(.A1(new_n760), .A2(new_n761), .A3(new_n773), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n754), .A2(new_n758), .ZN(new_n775));
  AOI22_X1  g574(.A1(G92gat), .A2(new_n769), .B1(new_n775), .B2(new_n773), .ZN(new_n776));
  OAI22_X1  g575(.A1(new_n772), .A2(new_n774), .B1(new_n776), .B2(new_n771), .ZN(G1337gat));
  NAND3_X1  g576(.A1(new_n710), .A2(new_n685), .A3(new_n766), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n778), .A2(G99gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n427), .A2(new_n663), .ZN(new_n780));
  NOR2_X1   g579(.A1(new_n780), .A2(G99gat), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n760), .A2(new_n761), .A3(new_n781), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n779), .A2(new_n782), .ZN(G1338gat));
  NAND4_X1  g582(.A1(new_n707), .A2(new_n709), .A3(new_n398), .A4(new_n766), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n784), .A2(G106gat), .ZN(new_n785));
  INV_X1    g584(.A(KEYINPUT53), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR3_X1   g586(.A1(new_n421), .A2(G106gat), .A3(new_n735), .ZN(new_n788));
  AND3_X1   g587(.A1(new_n760), .A2(new_n761), .A3(new_n788), .ZN(new_n789));
  NAND4_X1  g588(.A1(new_n707), .A2(new_n709), .A3(new_n268), .A4(new_n766), .ZN(new_n790));
  AOI22_X1  g589(.A1(G106gat), .A2(new_n790), .B1(new_n775), .B2(new_n788), .ZN(new_n791));
  OAI22_X1  g590(.A1(new_n787), .A2(new_n789), .B1(new_n791), .B2(new_n786), .ZN(G1339gat));
  NAND3_X1  g591(.A1(new_n657), .A2(new_n646), .A3(new_n658), .ZN(new_n793));
  OAI211_X1 g592(.A(new_n793), .B(KEYINPUT54), .C1(new_n645), .C2(new_n640), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n794), .A2(KEYINPUT55), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT54), .ZN(new_n796));
  INV_X1    g595(.A(new_n646), .ZN(new_n797));
  AOI21_X1  g596(.A(KEYINPUT10), .B1(new_n628), .B2(new_n638), .ZN(new_n798));
  OAI211_X1 g597(.A(new_n796), .B(new_n797), .C1(new_n798), .C2(new_n642), .ZN(new_n799));
  INV_X1    g598(.A(KEYINPUT115), .ZN(new_n800));
  NAND3_X1  g599(.A1(new_n799), .A2(new_n800), .A3(new_n652), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n799), .A2(new_n652), .ZN(new_n802));
  NAND2_X1  g601(.A1(new_n802), .A2(KEYINPUT115), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n801), .B2(new_n803), .ZN(new_n804));
  INV_X1    g603(.A(new_n662), .ZN(new_n805));
  OAI21_X1  g604(.A(KEYINPUT116), .B1(new_n804), .B2(new_n805), .ZN(new_n806));
  INV_X1    g605(.A(KEYINPUT55), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n796), .B1(new_n659), .B2(new_n639), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n807), .B1(new_n808), .B2(new_n793), .ZN(new_n809));
  AND3_X1   g608(.A1(new_n799), .A2(new_n800), .A3(new_n652), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n800), .B1(new_n799), .B2(new_n652), .ZN(new_n811));
  OAI21_X1  g610(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  INV_X1    g611(.A(KEYINPUT116), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n812), .A2(new_n813), .A3(new_n662), .ZN(new_n814));
  NAND2_X1  g613(.A1(new_n806), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n603), .A2(new_n611), .A3(new_n624), .ZN(new_n816));
  AOI21_X1  g615(.A(new_n596), .B1(new_n595), .B2(new_n597), .ZN(new_n817));
  NOR3_X1   g616(.A1(new_n607), .A2(new_n608), .A3(new_n606), .ZN(new_n818));
  OAI21_X1  g617(.A(new_n618), .B1(new_n817), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g618(.A1(new_n816), .A2(new_n819), .ZN(new_n820));
  OAI21_X1  g619(.A(new_n794), .B1(new_n810), .B2(new_n811), .ZN(new_n821));
  AOI22_X1  g620(.A1(new_n821), .A2(new_n807), .B1(new_n588), .B2(new_n591), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n815), .A2(new_n820), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n816), .A2(new_n663), .A3(new_n819), .ZN(new_n824));
  INV_X1    g623(.A(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n803), .A2(new_n801), .ZN(new_n826));
  AOI21_X1  g625(.A(KEYINPUT55), .B1(new_n826), .B2(new_n794), .ZN(new_n827));
  AOI21_X1  g626(.A(new_n827), .B1(new_n620), .B2(new_n625), .ZN(new_n828));
  AOI21_X1  g627(.A(new_n825), .B1(new_n828), .B2(new_n815), .ZN(new_n829));
  OAI21_X1  g628(.A(new_n823), .B1(new_n829), .B2(new_n755), .ZN(new_n830));
  INV_X1    g629(.A(new_n483), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NOR3_X1   g631(.A1(new_n593), .A2(new_n626), .A3(new_n663), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n832), .A2(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(new_n728), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n317), .A2(new_n424), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(new_n427), .ZN(new_n839));
  OAI21_X1  g638(.A(G113gat), .B1(new_n839), .B2(new_n627), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n833), .B1(new_n830), .B2(new_n831), .ZN(new_n841));
  NOR2_X1   g640(.A1(new_n841), .A2(new_n316), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n423), .A2(new_n360), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n845), .A2(new_n281), .A3(new_n626), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n840), .A2(new_n846), .ZN(G1340gat));
  AOI21_X1  g646(.A(G120gat), .B1(new_n845), .B2(new_n663), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n780), .A2(new_n277), .ZN(new_n849));
  AOI21_X1  g648(.A(new_n848), .B1(new_n838), .B2(new_n849), .ZN(G1341gat));
  OAI21_X1  g649(.A(G127gat), .B1(new_n839), .B2(new_n831), .ZN(new_n851));
  OR2_X1    g650(.A1(new_n831), .A2(G127gat), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n851), .B1(new_n844), .B2(new_n852), .ZN(G1342gat));
  NOR3_X1   g652(.A1(new_n844), .A2(G134gat), .A3(new_n592), .ZN(new_n854));
  XNOR2_X1  g653(.A(new_n854), .B(KEYINPUT56), .ZN(new_n855));
  OAI21_X1  g654(.A(G134gat), .B1(new_n839), .B2(new_n592), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n855), .A2(new_n856), .ZN(G1343gat));
  NAND2_X1  g656(.A1(new_n812), .A2(new_n662), .ZN(new_n858));
  AOI211_X1 g657(.A(new_n858), .B(new_n827), .C1(new_n620), .C2(new_n625), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT117), .ZN(new_n860));
  NAND2_X1  g659(.A1(new_n824), .A2(new_n860), .ZN(new_n861));
  NAND4_X1  g660(.A1(new_n816), .A2(KEYINPUT117), .A3(new_n663), .A4(new_n819), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n861), .A2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n592), .B1(new_n859), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(new_n823), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n831), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n728), .B1(new_n866), .B2(new_n834), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT57), .ZN(new_n868));
  OR2_X1    g667(.A1(new_n867), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n841), .A2(KEYINPUT57), .A3(new_n421), .ZN(new_n870));
  INV_X1    g669(.A(new_n870), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n837), .A2(new_n397), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n869), .A2(new_n871), .A3(new_n872), .ZN(new_n873));
  OAI21_X1  g672(.A(G141gat), .B1(new_n873), .B2(new_n627), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT58), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n626), .A2(new_n217), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n685), .A2(new_n421), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n842), .A2(new_n877), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT119), .ZN(new_n879));
  AOI21_X1  g678(.A(new_n360), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n842), .A2(KEYINPUT119), .A3(new_n877), .ZN(new_n881));
  NAND2_X1  g680(.A1(new_n880), .A2(new_n881), .ZN(new_n882));
  OAI211_X1 g681(.A(new_n874), .B(new_n875), .C1(new_n876), .C2(new_n882), .ZN(new_n883));
  NOR3_X1   g682(.A1(new_n878), .A2(new_n360), .A3(new_n876), .ZN(new_n884));
  NAND4_X1  g683(.A1(new_n869), .A2(KEYINPUT118), .A3(new_n871), .A4(new_n872), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT118), .ZN(new_n886));
  OAI21_X1  g685(.A(new_n872), .B1(new_n867), .B2(new_n868), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n886), .B1(new_n887), .B2(new_n870), .ZN(new_n888));
  NAND3_X1  g687(.A1(new_n885), .A2(new_n626), .A3(new_n888), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n889), .B2(G141gat), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n883), .B1(new_n890), .B2(new_n875), .ZN(G1344gat));
  NAND4_X1  g690(.A1(new_n880), .A2(new_n212), .A3(new_n663), .A4(new_n881), .ZN(new_n892));
  XOR2_X1   g691(.A(new_n892), .B(KEYINPUT120), .Z(new_n893));
  INV_X1    g692(.A(KEYINPUT59), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n894), .A2(G148gat), .ZN(new_n895));
  AND2_X1   g694(.A1(new_n885), .A2(new_n888), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n895), .B1(new_n896), .B2(new_n663), .ZN(new_n897));
  OAI21_X1  g696(.A(KEYINPUT57), .B1(new_n841), .B2(new_n421), .ZN(new_n898));
  AOI21_X1  g697(.A(KEYINPUT57), .B1(new_n263), .B2(new_n267), .ZN(new_n899));
  AND3_X1   g698(.A1(new_n812), .A2(new_n813), .A3(new_n662), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n813), .B1(new_n812), .B2(new_n662), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n822), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n902), .A2(KEYINPUT121), .ZN(new_n903));
  INV_X1    g702(.A(KEYINPUT121), .ZN(new_n904));
  NAND3_X1  g703(.A1(new_n815), .A2(new_n904), .A3(new_n822), .ZN(new_n905));
  NAND3_X1  g704(.A1(new_n903), .A2(new_n905), .A3(new_n820), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n483), .B1(new_n906), .B2(new_n864), .ZN(new_n907));
  OAI21_X1  g706(.A(new_n899), .B1(new_n907), .B2(new_n833), .ZN(new_n908));
  AND2_X1   g707(.A1(new_n898), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g708(.A1(new_n909), .A2(new_n663), .A3(new_n872), .ZN(new_n910));
  AOI21_X1  g709(.A(new_n894), .B1(new_n910), .B2(G148gat), .ZN(new_n911));
  OAI21_X1  g710(.A(new_n893), .B1(new_n897), .B2(new_n911), .ZN(G1345gat));
  NOR3_X1   g711(.A1(new_n882), .A2(KEYINPUT122), .A3(new_n831), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n913), .A2(G155gat), .ZN(new_n914));
  OAI21_X1  g713(.A(KEYINPUT122), .B1(new_n882), .B2(new_n831), .ZN(new_n915));
  NOR2_X1   g714(.A1(new_n831), .A2(new_n221), .ZN(new_n916));
  AOI22_X1  g715(.A1(new_n914), .A2(new_n915), .B1(new_n896), .B2(new_n916), .ZN(G1346gat));
  NOR2_X1   g716(.A1(new_n592), .A2(new_n222), .ZN(new_n918));
  NAND3_X1  g717(.A1(new_n880), .A2(new_n755), .A3(new_n881), .ZN(new_n919));
  AOI22_X1  g718(.A1(new_n896), .A2(new_n918), .B1(new_n222), .B2(new_n919), .ZN(G1347gat));
  AOI21_X1  g719(.A(new_n424), .B1(new_n314), .B2(new_n315), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n835), .A2(new_n728), .A3(new_n427), .A4(new_n921), .ZN(new_n922));
  NOR3_X1   g721(.A1(new_n922), .A2(new_n319), .A3(new_n627), .ZN(new_n923));
  NOR2_X1   g722(.A1(new_n841), .A2(new_n317), .ZN(new_n924));
  INV_X1    g723(.A(KEYINPUT123), .ZN(new_n925));
  XNOR2_X1  g724(.A(new_n924), .B(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(new_n423), .A2(new_n424), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  INV_X1    g727(.A(new_n928), .ZN(new_n929));
  NAND2_X1  g728(.A1(new_n929), .A2(new_n626), .ZN(new_n930));
  AOI21_X1  g729(.A(new_n923), .B1(new_n930), .B2(new_n319), .ZN(G1348gat));
  NOR3_X1   g730(.A1(new_n922), .A2(new_n320), .A3(new_n735), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n663), .ZN(new_n933));
  AOI21_X1  g732(.A(new_n932), .B1(new_n933), .B2(new_n320), .ZN(G1349gat));
  OAI21_X1  g733(.A(G183gat), .B1(new_n922), .B2(new_n831), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n483), .A2(new_n325), .ZN(new_n936));
  OAI21_X1  g735(.A(new_n935), .B1(new_n928), .B2(new_n936), .ZN(new_n937));
  XNOR2_X1  g736(.A(new_n937), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g737(.A(G190gat), .B1(new_n922), .B2(new_n592), .ZN(new_n939));
  XNOR2_X1  g738(.A(new_n939), .B(KEYINPUT61), .ZN(new_n940));
  NAND2_X1  g739(.A1(new_n755), .A2(new_n326), .ZN(new_n941));
  OAI21_X1  g740(.A(new_n940), .B1(new_n928), .B2(new_n941), .ZN(G1351gat));
  OAI21_X1  g741(.A(new_n921), .B1(new_n683), .B2(new_n684), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT124), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  OAI211_X1 g744(.A(new_n921), .B(KEYINPUT124), .C1(new_n683), .C2(new_n684), .ZN(new_n946));
  NAND2_X1  g745(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n909), .A2(new_n947), .ZN(new_n948));
  INV_X1    g747(.A(G197gat), .ZN(new_n949));
  NOR3_X1   g748(.A1(new_n948), .A2(new_n949), .A3(new_n627), .ZN(new_n950));
  NOR3_X1   g749(.A1(new_n685), .A2(new_n424), .A3(new_n421), .ZN(new_n951));
  NAND3_X1  g750(.A1(new_n926), .A2(new_n626), .A3(new_n951), .ZN(new_n952));
  AOI21_X1  g751(.A(new_n950), .B1(new_n949), .B2(new_n952), .ZN(G1352gat));
  NOR2_X1   g752(.A1(new_n735), .A2(G204gat), .ZN(new_n954));
  NAND3_X1  g753(.A1(new_n926), .A2(new_n951), .A3(new_n954), .ZN(new_n955));
  OR2_X1    g754(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n956));
  OAI21_X1  g755(.A(G204gat), .B1(new_n948), .B2(new_n735), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n955), .A2(KEYINPUT62), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n956), .A2(new_n957), .A3(new_n958), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(KEYINPUT125), .ZN(new_n960));
  INV_X1    g759(.A(KEYINPUT125), .ZN(new_n961));
  NAND4_X1  g760(.A1(new_n956), .A2(new_n961), .A3(new_n957), .A4(new_n958), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n960), .A2(new_n962), .ZN(G1353gat));
  INV_X1    g762(.A(KEYINPUT63), .ZN(new_n964));
  NAND4_X1  g763(.A1(new_n898), .A2(new_n483), .A3(new_n908), .A4(new_n947), .ZN(new_n965));
  AND2_X1   g764(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n966));
  OAI21_X1  g765(.A(G211gat), .B1(new_n965), .B2(KEYINPUT126), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n964), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  INV_X1    g767(.A(KEYINPUT126), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n909), .A2(new_n969), .A3(new_n483), .A4(new_n947), .ZN(new_n970));
  NAND2_X1  g769(.A1(new_n965), .A2(KEYINPUT126), .ZN(new_n971));
  NAND4_X1  g770(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n971), .ZN(new_n972));
  NAND2_X1  g771(.A1(new_n968), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n926), .A2(new_n951), .ZN(new_n974));
  OR3_X1    g773(.A1(new_n974), .A2(G211gat), .A3(new_n831), .ZN(new_n975));
  NAND2_X1  g774(.A1(new_n973), .A2(new_n975), .ZN(new_n976));
  NAND2_X1  g775(.A1(new_n976), .A2(KEYINPUT127), .ZN(new_n977));
  INV_X1    g776(.A(KEYINPUT127), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n973), .A2(new_n975), .A3(new_n978), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n977), .A2(new_n979), .ZN(G1354gat));
  OAI21_X1  g779(.A(G218gat), .B1(new_n948), .B2(new_n592), .ZN(new_n981));
  OR2_X1    g780(.A1(new_n592), .A2(G218gat), .ZN(new_n982));
  OAI21_X1  g781(.A(new_n981), .B1(new_n974), .B2(new_n982), .ZN(G1355gat));
endmodule


