

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762,
         n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773,
         n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
         n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795,
         n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
         n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817,
         n818, n819, n820, n821, n822, n823, n824, n825, n826, n827, n828,
         n829, n830, n831, n832, n833, n834, n835, n836, n837, n838, n839,
         n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
         n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861,
         n862, n863, n864, n865, n866, n867, n868, n869, n870, n871, n872,
         n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883,
         n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, n894,
         n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905,
         n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
         n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
         n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938,
         n939, n940, n941, n942, n943, n944, n945, n946, n947, n948, n949,
         n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
         n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
         n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982,
         n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993,
         n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  OR2_X1 U552 ( .A1(n962), .A2(n707), .ZN(n706) );
  XNOR2_X1 U553 ( .A(n761), .B(KEYINPUT103), .ZN(n762) );
  NOR2_X1 U554 ( .A1(G651), .A2(n646), .ZN(n651) );
  NOR2_X1 U555 ( .A1(G2104), .A2(G2105), .ZN(n517) );
  XOR2_X2 U556 ( .A(KEYINPUT17), .B(n517), .Z(n881) );
  NAND2_X1 U557 ( .A1(n881), .A2(G137), .ZN(n518) );
  XNOR2_X1 U558 ( .A(n518), .B(KEYINPUT68), .ZN(n521) );
  AND2_X1 U559 ( .A1(G2104), .A2(G2105), .ZN(n887) );
  NAND2_X1 U560 ( .A1(n887), .A2(G113), .ZN(n519) );
  XOR2_X1 U561 ( .A(KEYINPUT67), .B(n519), .Z(n520) );
  NAND2_X1 U562 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U563 ( .A(n522), .B(KEYINPUT69), .ZN(n524) );
  INV_X1 U564 ( .A(G2105), .ZN(n525) );
  NOR2_X1 U565 ( .A1(G2104), .A2(n525), .ZN(n886) );
  NAND2_X1 U566 ( .A1(G125), .A2(n886), .ZN(n523) );
  NAND2_X1 U567 ( .A1(n524), .A2(n523), .ZN(n529) );
  AND2_X1 U568 ( .A1(n525), .A2(G2104), .ZN(n882) );
  NAND2_X1 U569 ( .A1(G101), .A2(n882), .ZN(n526) );
  XNOR2_X1 U570 ( .A(n526), .B(KEYINPUT66), .ZN(n527) );
  XNOR2_X1 U571 ( .A(n527), .B(KEYINPUT23), .ZN(n528) );
  NOR2_X4 U572 ( .A1(n529), .A2(n528), .ZN(G160) );
  XOR2_X1 U573 ( .A(G543), .B(KEYINPUT0), .Z(n646) );
  NAND2_X1 U574 ( .A1(G52), .A2(n651), .ZN(n532) );
  INV_X1 U575 ( .A(G651), .ZN(n536) );
  NOR2_X1 U576 ( .A1(G543), .A2(n536), .ZN(n530) );
  XOR2_X1 U577 ( .A(KEYINPUT1), .B(n530), .Z(n650) );
  NAND2_X1 U578 ( .A1(G64), .A2(n650), .ZN(n531) );
  NAND2_X1 U579 ( .A1(n532), .A2(n531), .ZN(n533) );
  XOR2_X1 U580 ( .A(KEYINPUT71), .B(n533), .Z(n541) );
  NOR2_X1 U581 ( .A1(G543), .A2(G651), .ZN(n534) );
  XOR2_X1 U582 ( .A(KEYINPUT65), .B(n534), .Z(n637) );
  NAND2_X1 U583 ( .A1(n637), .A2(G90), .ZN(n535) );
  XNOR2_X1 U584 ( .A(n535), .B(KEYINPUT72), .ZN(n538) );
  NOR2_X1 U585 ( .A1(n646), .A2(n536), .ZN(n638) );
  NAND2_X1 U586 ( .A1(G77), .A2(n638), .ZN(n537) );
  NAND2_X1 U587 ( .A1(n538), .A2(n537), .ZN(n539) );
  XOR2_X1 U588 ( .A(KEYINPUT9), .B(n539), .Z(n540) );
  NOR2_X1 U589 ( .A1(n541), .A2(n540), .ZN(G171) );
  INV_X1 U590 ( .A(G171), .ZN(G301) );
  XOR2_X1 U591 ( .A(G2443), .B(G2446), .Z(n543) );
  XNOR2_X1 U592 ( .A(G2427), .B(G2451), .ZN(n542) );
  XNOR2_X1 U593 ( .A(n543), .B(n542), .ZN(n549) );
  XOR2_X1 U594 ( .A(G2430), .B(G2454), .Z(n545) );
  XNOR2_X1 U595 ( .A(G1341), .B(G1348), .ZN(n544) );
  XNOR2_X1 U596 ( .A(n545), .B(n544), .ZN(n547) );
  XOR2_X1 U597 ( .A(G2435), .B(G2438), .Z(n546) );
  XNOR2_X1 U598 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U599 ( .A(n549), .B(n548), .Z(n550) );
  AND2_X1 U600 ( .A1(G14), .A2(n550), .ZN(G401) );
  AND2_X1 U601 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U602 ( .A(G132), .ZN(G219) );
  INV_X1 U603 ( .A(G82), .ZN(G220) );
  INV_X1 U604 ( .A(G108), .ZN(G238) );
  NAND2_X1 U605 ( .A1(G50), .A2(n651), .ZN(n552) );
  NAND2_X1 U606 ( .A1(G62), .A2(n650), .ZN(n551) );
  NAND2_X1 U607 ( .A1(n552), .A2(n551), .ZN(n553) );
  XNOR2_X1 U608 ( .A(KEYINPUT87), .B(n553), .ZN(n557) );
  NAND2_X1 U609 ( .A1(G88), .A2(n637), .ZN(n555) );
  NAND2_X1 U610 ( .A1(G75), .A2(n638), .ZN(n554) );
  AND2_X1 U611 ( .A1(n555), .A2(n554), .ZN(n556) );
  NAND2_X1 U612 ( .A1(n557), .A2(n556), .ZN(G303) );
  NAND2_X1 U613 ( .A1(n637), .A2(G89), .ZN(n558) );
  XNOR2_X1 U614 ( .A(n558), .B(KEYINPUT4), .ZN(n560) );
  NAND2_X1 U615 ( .A1(G76), .A2(n638), .ZN(n559) );
  NAND2_X1 U616 ( .A1(n560), .A2(n559), .ZN(n561) );
  XNOR2_X1 U617 ( .A(n561), .B(KEYINPUT5), .ZN(n567) );
  XNOR2_X1 U618 ( .A(KEYINPUT6), .B(KEYINPUT79), .ZN(n565) );
  NAND2_X1 U619 ( .A1(G51), .A2(n651), .ZN(n563) );
  NAND2_X1 U620 ( .A1(G63), .A2(n650), .ZN(n562) );
  NAND2_X1 U621 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U622 ( .A(n565), .B(n564), .ZN(n566) );
  NAND2_X1 U623 ( .A1(n567), .A2(n566), .ZN(n568) );
  XNOR2_X1 U624 ( .A(KEYINPUT7), .B(n568), .ZN(G168) );
  XOR2_X1 U625 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  XOR2_X1 U626 ( .A(KEYINPUT11), .B(KEYINPUT76), .Z(n572) );
  XOR2_X1 U627 ( .A(KEYINPUT75), .B(KEYINPUT10), .Z(n570) );
  NAND2_X1 U628 ( .A1(G7), .A2(G661), .ZN(n569) );
  XOR2_X1 U629 ( .A(n570), .B(n569), .Z(n829) );
  NAND2_X1 U630 ( .A1(G567), .A2(n829), .ZN(n571) );
  XNOR2_X1 U631 ( .A(n572), .B(n571), .ZN(G234) );
  NAND2_X1 U632 ( .A1(n637), .A2(G81), .ZN(n573) );
  XNOR2_X1 U633 ( .A(n573), .B(KEYINPUT12), .ZN(n575) );
  NAND2_X1 U634 ( .A1(G68), .A2(n638), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(n576) );
  XNOR2_X1 U636 ( .A(n576), .B(KEYINPUT13), .ZN(n578) );
  NAND2_X1 U637 ( .A1(G43), .A2(n651), .ZN(n577) );
  NAND2_X1 U638 ( .A1(n578), .A2(n577), .ZN(n581) );
  NAND2_X1 U639 ( .A1(n650), .A2(G56), .ZN(n579) );
  XOR2_X1 U640 ( .A(KEYINPUT14), .B(n579), .Z(n580) );
  NOR2_X1 U641 ( .A1(n581), .A2(n580), .ZN(n980) );
  NAND2_X1 U642 ( .A1(n980), .A2(G860), .ZN(G153) );
  NAND2_X1 U643 ( .A1(G868), .A2(G301), .ZN(n592) );
  NAND2_X1 U644 ( .A1(G92), .A2(n637), .ZN(n583) );
  NAND2_X1 U645 ( .A1(G66), .A2(n650), .ZN(n582) );
  NAND2_X1 U646 ( .A1(n583), .A2(n582), .ZN(n584) );
  XNOR2_X1 U647 ( .A(n584), .B(KEYINPUT77), .ZN(n586) );
  NAND2_X1 U648 ( .A1(G79), .A2(n638), .ZN(n585) );
  NAND2_X1 U649 ( .A1(n586), .A2(n585), .ZN(n589) );
  NAND2_X1 U650 ( .A1(n651), .A2(G54), .ZN(n587) );
  XOR2_X1 U651 ( .A(KEYINPUT78), .B(n587), .Z(n588) );
  NOR2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  XOR2_X1 U653 ( .A(KEYINPUT15), .B(n590), .Z(n899) );
  INV_X1 U654 ( .A(n899), .ZN(n962) );
  INV_X1 U655 ( .A(G868), .ZN(n665) );
  NAND2_X1 U656 ( .A1(n962), .A2(n665), .ZN(n591) );
  NAND2_X1 U657 ( .A1(n592), .A2(n591), .ZN(G284) );
  NAND2_X1 U658 ( .A1(n651), .A2(G53), .ZN(n595) );
  NAND2_X1 U659 ( .A1(G78), .A2(n638), .ZN(n593) );
  XOR2_X1 U660 ( .A(KEYINPUT73), .B(n593), .Z(n594) );
  NAND2_X1 U661 ( .A1(n595), .A2(n594), .ZN(n599) );
  NAND2_X1 U662 ( .A1(G91), .A2(n637), .ZN(n597) );
  NAND2_X1 U663 ( .A1(G65), .A2(n650), .ZN(n596) );
  NAND2_X1 U664 ( .A1(n597), .A2(n596), .ZN(n598) );
  NOR2_X1 U665 ( .A1(n599), .A2(n598), .ZN(n964) );
  XOR2_X1 U666 ( .A(n964), .B(KEYINPUT74), .Z(G299) );
  NOR2_X1 U667 ( .A1(G868), .A2(G299), .ZN(n601) );
  NOR2_X1 U668 ( .A1(G286), .A2(n665), .ZN(n600) );
  NOR2_X1 U669 ( .A1(n601), .A2(n600), .ZN(G297) );
  INV_X1 U670 ( .A(G860), .ZN(n602) );
  NAND2_X1 U671 ( .A1(n602), .A2(G559), .ZN(n603) );
  NAND2_X1 U672 ( .A1(n603), .A2(n899), .ZN(n604) );
  XNOR2_X1 U673 ( .A(n604), .B(KEYINPUT16), .ZN(G148) );
  NAND2_X1 U674 ( .A1(n980), .A2(n665), .ZN(n605) );
  XOR2_X1 U675 ( .A(KEYINPUT80), .B(n605), .Z(n608) );
  NAND2_X1 U676 ( .A1(G868), .A2(n899), .ZN(n606) );
  NOR2_X1 U677 ( .A1(G559), .A2(n606), .ZN(n607) );
  NOR2_X1 U678 ( .A1(n608), .A2(n607), .ZN(G282) );
  NAND2_X1 U679 ( .A1(G123), .A2(n886), .ZN(n609) );
  XOR2_X1 U680 ( .A(KEYINPUT18), .B(n609), .Z(n610) );
  XNOR2_X1 U681 ( .A(n610), .B(KEYINPUT81), .ZN(n612) );
  NAND2_X1 U682 ( .A1(G111), .A2(n887), .ZN(n611) );
  NAND2_X1 U683 ( .A1(n612), .A2(n611), .ZN(n616) );
  NAND2_X1 U684 ( .A1(G135), .A2(n881), .ZN(n614) );
  NAND2_X1 U685 ( .A1(G99), .A2(n882), .ZN(n613) );
  NAND2_X1 U686 ( .A1(n614), .A2(n613), .ZN(n615) );
  NOR2_X1 U687 ( .A1(n616), .A2(n615), .ZN(n918) );
  XOR2_X1 U688 ( .A(G2096), .B(n918), .Z(n617) );
  NOR2_X1 U689 ( .A1(G2100), .A2(n617), .ZN(n618) );
  XOR2_X1 U690 ( .A(KEYINPUT82), .B(n618), .Z(G156) );
  NAND2_X1 U691 ( .A1(G55), .A2(n651), .ZN(n620) );
  NAND2_X1 U692 ( .A1(G67), .A2(n650), .ZN(n619) );
  NAND2_X1 U693 ( .A1(n620), .A2(n619), .ZN(n624) );
  NAND2_X1 U694 ( .A1(G93), .A2(n637), .ZN(n622) );
  NAND2_X1 U695 ( .A1(G80), .A2(n638), .ZN(n621) );
  NAND2_X1 U696 ( .A1(n622), .A2(n621), .ZN(n623) );
  NOR2_X1 U697 ( .A1(n624), .A2(n623), .ZN(n666) );
  NAND2_X1 U698 ( .A1(n899), .A2(G559), .ZN(n663) );
  XOR2_X1 U699 ( .A(n980), .B(n663), .Z(n625) );
  NOR2_X1 U700 ( .A1(G860), .A2(n625), .ZN(n626) );
  XNOR2_X1 U701 ( .A(n666), .B(n626), .ZN(G145) );
  NAND2_X1 U702 ( .A1(G61), .A2(n650), .ZN(n627) );
  XNOR2_X1 U703 ( .A(n627), .B(KEYINPUT84), .ZN(n636) );
  NAND2_X1 U704 ( .A1(G73), .A2(n638), .ZN(n628) );
  XNOR2_X1 U705 ( .A(n628), .B(KEYINPUT86), .ZN(n629) );
  XNOR2_X1 U706 ( .A(n629), .B(KEYINPUT2), .ZN(n631) );
  NAND2_X1 U707 ( .A1(G48), .A2(n651), .ZN(n630) );
  NAND2_X1 U708 ( .A1(n631), .A2(n630), .ZN(n634) );
  NAND2_X1 U709 ( .A1(G86), .A2(n637), .ZN(n632) );
  XNOR2_X1 U710 ( .A(KEYINPUT85), .B(n632), .ZN(n633) );
  NOR2_X1 U711 ( .A1(n634), .A2(n633), .ZN(n635) );
  NAND2_X1 U712 ( .A1(n636), .A2(n635), .ZN(G305) );
  NAND2_X1 U713 ( .A1(G85), .A2(n637), .ZN(n640) );
  NAND2_X1 U714 ( .A1(G72), .A2(n638), .ZN(n639) );
  NAND2_X1 U715 ( .A1(n640), .A2(n639), .ZN(n643) );
  NAND2_X1 U716 ( .A1(G47), .A2(n651), .ZN(n641) );
  XOR2_X1 U717 ( .A(KEYINPUT70), .B(n641), .Z(n642) );
  NOR2_X1 U718 ( .A1(n643), .A2(n642), .ZN(n645) );
  NAND2_X1 U719 ( .A1(n650), .A2(G60), .ZN(n644) );
  NAND2_X1 U720 ( .A1(n645), .A2(n644), .ZN(G290) );
  NAND2_X1 U721 ( .A1(G87), .A2(n646), .ZN(n648) );
  NAND2_X1 U722 ( .A1(G74), .A2(G651), .ZN(n647) );
  NAND2_X1 U723 ( .A1(n648), .A2(n647), .ZN(n649) );
  NOR2_X1 U724 ( .A1(n650), .A2(n649), .ZN(n654) );
  NAND2_X1 U725 ( .A1(G49), .A2(n651), .ZN(n652) );
  XOR2_X1 U726 ( .A(KEYINPUT83), .B(n652), .Z(n653) );
  NAND2_X1 U727 ( .A1(n654), .A2(n653), .ZN(G288) );
  XNOR2_X1 U728 ( .A(KEYINPUT19), .B(KEYINPUT88), .ZN(n656) );
  XNOR2_X1 U729 ( .A(G305), .B(KEYINPUT89), .ZN(n655) );
  XNOR2_X1 U730 ( .A(n656), .B(n655), .ZN(n657) );
  XOR2_X1 U731 ( .A(n657), .B(n666), .Z(n659) );
  XOR2_X1 U732 ( .A(G303), .B(G299), .Z(n658) );
  XNOR2_X1 U733 ( .A(n659), .B(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(G290), .ZN(n661) );
  XNOR2_X1 U735 ( .A(n661), .B(G288), .ZN(n662) );
  XNOR2_X1 U736 ( .A(n980), .B(n662), .ZN(n900) );
  XOR2_X1 U737 ( .A(n900), .B(n663), .Z(n664) );
  NOR2_X1 U738 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U739 ( .A1(G868), .A2(n666), .ZN(n667) );
  NOR2_X1 U740 ( .A1(n668), .A2(n667), .ZN(n669) );
  XOR2_X1 U741 ( .A(KEYINPUT90), .B(n669), .Z(G295) );
  NAND2_X1 U742 ( .A1(G2078), .A2(G2084), .ZN(n670) );
  XOR2_X1 U743 ( .A(KEYINPUT20), .B(n670), .Z(n671) );
  NAND2_X1 U744 ( .A1(G2090), .A2(n671), .ZN(n672) );
  XNOR2_X1 U745 ( .A(KEYINPUT21), .B(n672), .ZN(n673) );
  NAND2_X1 U746 ( .A1(n673), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U747 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NAND2_X1 U748 ( .A1(G69), .A2(G120), .ZN(n674) );
  XOR2_X1 U749 ( .A(KEYINPUT92), .B(n674), .Z(n675) );
  NAND2_X1 U750 ( .A1(G57), .A2(n675), .ZN(n676) );
  NOR2_X1 U751 ( .A1(G238), .A2(n676), .ZN(n677) );
  XNOR2_X1 U752 ( .A(KEYINPUT93), .B(n677), .ZN(n834) );
  NAND2_X1 U753 ( .A1(G567), .A2(n834), .ZN(n678) );
  XNOR2_X1 U754 ( .A(n678), .B(KEYINPUT94), .ZN(n684) );
  NOR2_X1 U755 ( .A1(G220), .A2(G219), .ZN(n679) );
  XOR2_X1 U756 ( .A(KEYINPUT22), .B(n679), .Z(n680) );
  NOR2_X1 U757 ( .A1(G218), .A2(n680), .ZN(n681) );
  NAND2_X1 U758 ( .A1(G96), .A2(n681), .ZN(n835) );
  NAND2_X1 U759 ( .A1(G2106), .A2(n835), .ZN(n682) );
  XOR2_X1 U760 ( .A(KEYINPUT91), .B(n682), .Z(n683) );
  NAND2_X1 U761 ( .A1(n684), .A2(n683), .ZN(n685) );
  XOR2_X1 U762 ( .A(n685), .B(KEYINPUT95), .Z(n833) );
  NAND2_X1 U763 ( .A1(G661), .A2(G483), .ZN(n686) );
  NOR2_X1 U764 ( .A1(n833), .A2(n686), .ZN(n832) );
  NAND2_X1 U765 ( .A1(n832), .A2(G36), .ZN(G176) );
  NAND2_X1 U766 ( .A1(G138), .A2(n881), .ZN(n688) );
  NAND2_X1 U767 ( .A1(G102), .A2(n882), .ZN(n687) );
  NAND2_X1 U768 ( .A1(n688), .A2(n687), .ZN(n692) );
  NAND2_X1 U769 ( .A1(G126), .A2(n886), .ZN(n690) );
  NAND2_X1 U770 ( .A1(G114), .A2(n887), .ZN(n689) );
  NAND2_X1 U771 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U772 ( .A1(n692), .A2(n691), .ZN(G164) );
  NOR2_X1 U773 ( .A1(G164), .A2(G1384), .ZN(n767) );
  AND2_X1 U774 ( .A1(n767), .A2(G40), .ZN(n695) );
  AND2_X1 U775 ( .A1(G1996), .A2(n695), .ZN(n693) );
  NAND2_X1 U776 ( .A1(G160), .A2(n693), .ZN(n694) );
  XNOR2_X1 U777 ( .A(n694), .B(KEYINPUT26), .ZN(n697) );
  NAND2_X1 U778 ( .A1(G160), .A2(n695), .ZN(n733) );
  NAND2_X1 U779 ( .A1(G1341), .A2(n733), .ZN(n696) );
  NAND2_X1 U780 ( .A1(n697), .A2(n696), .ZN(n698) );
  XNOR2_X1 U781 ( .A(n698), .B(KEYINPUT99), .ZN(n699) );
  NAND2_X1 U782 ( .A1(n699), .A2(n980), .ZN(n700) );
  XNOR2_X1 U783 ( .A(KEYINPUT64), .B(n700), .ZN(n707) );
  INV_X1 U784 ( .A(n733), .ZN(n721) );
  NAND2_X1 U785 ( .A1(G2067), .A2(n721), .ZN(n701) );
  XNOR2_X1 U786 ( .A(n701), .B(KEYINPUT100), .ZN(n703) );
  NAND2_X1 U787 ( .A1(G1348), .A2(n733), .ZN(n702) );
  NAND2_X1 U788 ( .A1(n703), .A2(n702), .ZN(n704) );
  XOR2_X1 U789 ( .A(KEYINPUT101), .B(n704), .Z(n705) );
  NAND2_X1 U790 ( .A1(n706), .A2(n705), .ZN(n709) );
  NAND2_X1 U791 ( .A1(n707), .A2(n962), .ZN(n708) );
  NAND2_X1 U792 ( .A1(n709), .A2(n708), .ZN(n714) );
  NAND2_X1 U793 ( .A1(n721), .A2(G2072), .ZN(n710) );
  XNOR2_X1 U794 ( .A(n710), .B(KEYINPUT27), .ZN(n712) );
  INV_X1 U795 ( .A(G1956), .ZN(n963) );
  NOR2_X1 U796 ( .A1(n963), .A2(n721), .ZN(n711) );
  NOR2_X1 U797 ( .A1(n712), .A2(n711), .ZN(n715) );
  NAND2_X1 U798 ( .A1(n964), .A2(n715), .ZN(n713) );
  NAND2_X1 U799 ( .A1(n714), .A2(n713), .ZN(n718) );
  NOR2_X1 U800 ( .A1(n964), .A2(n715), .ZN(n716) );
  XOR2_X1 U801 ( .A(n716), .B(KEYINPUT28), .Z(n717) );
  NAND2_X1 U802 ( .A1(n718), .A2(n717), .ZN(n719) );
  XOR2_X1 U803 ( .A(n719), .B(KEYINPUT29), .Z(n725) );
  NOR2_X1 U804 ( .A1(n721), .A2(G1961), .ZN(n720) );
  XOR2_X1 U805 ( .A(KEYINPUT98), .B(n720), .Z(n723) );
  XNOR2_X1 U806 ( .A(G2078), .B(KEYINPUT25), .ZN(n936) );
  NAND2_X1 U807 ( .A1(n721), .A2(n936), .ZN(n722) );
  NAND2_X1 U808 ( .A1(n723), .A2(n722), .ZN(n729) );
  NAND2_X1 U809 ( .A1(G171), .A2(n729), .ZN(n724) );
  NAND2_X1 U810 ( .A1(n725), .A2(n724), .ZN(n745) );
  NAND2_X1 U811 ( .A1(G8), .A2(n733), .ZN(n786) );
  NOR2_X1 U812 ( .A1(G1966), .A2(n786), .ZN(n747) );
  NOR2_X1 U813 ( .A1(G2084), .A2(n733), .ZN(n746) );
  NOR2_X1 U814 ( .A1(n747), .A2(n746), .ZN(n726) );
  NAND2_X1 U815 ( .A1(G8), .A2(n726), .ZN(n727) );
  XNOR2_X1 U816 ( .A(KEYINPUT30), .B(n727), .ZN(n728) );
  NOR2_X1 U817 ( .A1(G168), .A2(n728), .ZN(n731) );
  NOR2_X1 U818 ( .A1(G171), .A2(n729), .ZN(n730) );
  NOR2_X1 U819 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U820 ( .A(KEYINPUT31), .B(n732), .Z(n744) );
  NOR2_X1 U821 ( .A1(G1971), .A2(n786), .ZN(n735) );
  NOR2_X1 U822 ( .A1(G2090), .A2(n733), .ZN(n734) );
  NOR2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n736) );
  NAND2_X1 U824 ( .A1(n736), .A2(G303), .ZN(n738) );
  AND2_X1 U825 ( .A1(n744), .A2(n738), .ZN(n737) );
  NAND2_X1 U826 ( .A1(n745), .A2(n737), .ZN(n742) );
  INV_X1 U827 ( .A(n738), .ZN(n739) );
  OR2_X1 U828 ( .A1(n739), .A2(G286), .ZN(n740) );
  AND2_X1 U829 ( .A1(G8), .A2(n740), .ZN(n741) );
  NAND2_X1 U830 ( .A1(n742), .A2(n741), .ZN(n743) );
  XNOR2_X1 U831 ( .A(n743), .B(KEYINPUT32), .ZN(n752) );
  AND2_X1 U832 ( .A1(n745), .A2(n744), .ZN(n750) );
  AND2_X1 U833 ( .A1(G8), .A2(n746), .ZN(n748) );
  OR2_X1 U834 ( .A1(n748), .A2(n747), .ZN(n749) );
  OR2_X1 U835 ( .A1(n750), .A2(n749), .ZN(n751) );
  NAND2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n782) );
  NOR2_X1 U837 ( .A1(G1976), .A2(G288), .ZN(n969) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n975) );
  NOR2_X1 U839 ( .A1(n969), .A2(n975), .ZN(n754) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n753) );
  AND2_X1 U841 ( .A1(n754), .A2(n753), .ZN(n755) );
  NAND2_X1 U842 ( .A1(n782), .A2(n755), .ZN(n760) );
  NAND2_X1 U843 ( .A1(G288), .A2(G1976), .ZN(n756) );
  XNOR2_X1 U844 ( .A(n756), .B(KEYINPUT102), .ZN(n971) );
  INV_X1 U845 ( .A(n971), .ZN(n757) );
  NOR2_X1 U846 ( .A1(n757), .A2(n786), .ZN(n758) );
  OR2_X1 U847 ( .A1(KEYINPUT33), .A2(n758), .ZN(n759) );
  NAND2_X1 U848 ( .A1(n760), .A2(n759), .ZN(n761) );
  INV_X1 U849 ( .A(n762), .ZN(n765) );
  NAND2_X1 U850 ( .A1(n969), .A2(KEYINPUT33), .ZN(n763) );
  NOR2_X1 U851 ( .A1(n786), .A2(n763), .ZN(n764) );
  NOR2_X1 U852 ( .A1(n765), .A2(n764), .ZN(n779) );
  XOR2_X1 U853 ( .A(G1981), .B(G305), .Z(n959) );
  NAND2_X1 U854 ( .A1(G160), .A2(G40), .ZN(n766) );
  NOR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n823) );
  XNOR2_X1 U856 ( .A(KEYINPUT37), .B(G2067), .ZN(n821) );
  NAND2_X1 U857 ( .A1(G140), .A2(n881), .ZN(n769) );
  NAND2_X1 U858 ( .A1(G104), .A2(n882), .ZN(n768) );
  NAND2_X1 U859 ( .A1(n769), .A2(n768), .ZN(n770) );
  XNOR2_X1 U860 ( .A(KEYINPUT34), .B(n770), .ZN(n776) );
  NAND2_X1 U861 ( .A1(G128), .A2(n886), .ZN(n772) );
  NAND2_X1 U862 ( .A1(G116), .A2(n887), .ZN(n771) );
  NAND2_X1 U863 ( .A1(n772), .A2(n771), .ZN(n773) );
  XOR2_X1 U864 ( .A(KEYINPUT35), .B(n773), .Z(n774) );
  XNOR2_X1 U865 ( .A(KEYINPUT96), .B(n774), .ZN(n775) );
  NOR2_X1 U866 ( .A1(n776), .A2(n775), .ZN(n777) );
  XNOR2_X1 U867 ( .A(KEYINPUT36), .B(n777), .ZN(n877) );
  NOR2_X1 U868 ( .A1(n821), .A2(n877), .ZN(n931) );
  NAND2_X1 U869 ( .A1(n823), .A2(n931), .ZN(n820) );
  AND2_X1 U870 ( .A1(n959), .A2(n820), .ZN(n778) );
  NAND2_X1 U871 ( .A1(n779), .A2(n778), .ZN(n791) );
  NOR2_X1 U872 ( .A1(G2090), .A2(G303), .ZN(n780) );
  NAND2_X1 U873 ( .A1(G8), .A2(n780), .ZN(n781) );
  NAND2_X1 U874 ( .A1(n782), .A2(n781), .ZN(n783) );
  NAND2_X1 U875 ( .A1(n783), .A2(n786), .ZN(n788) );
  NOR2_X1 U876 ( .A1(G1981), .A2(G305), .ZN(n784) );
  XOR2_X1 U877 ( .A(n784), .B(KEYINPUT24), .Z(n785) );
  OR2_X1 U878 ( .A1(n786), .A2(n785), .ZN(n787) );
  NAND2_X1 U879 ( .A1(n788), .A2(n787), .ZN(n789) );
  NAND2_X1 U880 ( .A1(n820), .A2(n789), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(n810) );
  NAND2_X1 U882 ( .A1(G141), .A2(n881), .ZN(n793) );
  NAND2_X1 U883 ( .A1(G129), .A2(n886), .ZN(n792) );
  NAND2_X1 U884 ( .A1(n793), .A2(n792), .ZN(n796) );
  NAND2_X1 U885 ( .A1(n882), .A2(G105), .ZN(n794) );
  XOR2_X1 U886 ( .A(KEYINPUT38), .B(n794), .Z(n795) );
  NOR2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n798) );
  NAND2_X1 U888 ( .A1(n887), .A2(G117), .ZN(n797) );
  NAND2_X1 U889 ( .A1(n798), .A2(n797), .ZN(n894) );
  NAND2_X1 U890 ( .A1(G1996), .A2(n894), .ZN(n807) );
  NAND2_X1 U891 ( .A1(G131), .A2(n881), .ZN(n800) );
  NAND2_X1 U892 ( .A1(G119), .A2(n886), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n803) );
  NAND2_X1 U894 ( .A1(G95), .A2(n882), .ZN(n801) );
  XNOR2_X1 U895 ( .A(KEYINPUT97), .B(n801), .ZN(n802) );
  NOR2_X1 U896 ( .A1(n803), .A2(n802), .ZN(n805) );
  NAND2_X1 U897 ( .A1(n887), .A2(G107), .ZN(n804) );
  NAND2_X1 U898 ( .A1(n805), .A2(n804), .ZN(n873) );
  NAND2_X1 U899 ( .A1(G1991), .A2(n873), .ZN(n806) );
  NAND2_X1 U900 ( .A1(n807), .A2(n806), .ZN(n923) );
  NAND2_X1 U901 ( .A1(n823), .A2(n923), .ZN(n814) );
  XNOR2_X1 U902 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U903 ( .A1(n823), .A2(n966), .ZN(n808) );
  AND2_X1 U904 ( .A1(n814), .A2(n808), .ZN(n809) );
  NAND2_X1 U905 ( .A1(n810), .A2(n809), .ZN(n811) );
  XNOR2_X1 U906 ( .A(n811), .B(KEYINPUT104), .ZN(n826) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n873), .ZN(n919) );
  NOR2_X1 U908 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U909 ( .A1(n919), .A2(n812), .ZN(n813) );
  XNOR2_X1 U910 ( .A(n813), .B(KEYINPUT105), .ZN(n815) );
  NAND2_X1 U911 ( .A1(n815), .A2(n814), .ZN(n816) );
  OR2_X1 U912 ( .A1(n894), .A2(G1996), .ZN(n916) );
  NAND2_X1 U913 ( .A1(n816), .A2(n916), .ZN(n818) );
  XOR2_X1 U914 ( .A(KEYINPUT106), .B(KEYINPUT39), .Z(n817) );
  XNOR2_X1 U915 ( .A(n818), .B(n817), .ZN(n819) );
  NAND2_X1 U916 ( .A1(n820), .A2(n819), .ZN(n822) );
  NAND2_X1 U917 ( .A1(n821), .A2(n877), .ZN(n928) );
  NAND2_X1 U918 ( .A1(n822), .A2(n928), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n824), .A2(n823), .ZN(n825) );
  NAND2_X1 U920 ( .A1(n826), .A2(n825), .ZN(n827) );
  XNOR2_X1 U921 ( .A(n827), .B(KEYINPUT40), .ZN(G329) );
  INV_X1 U922 ( .A(G303), .ZN(G166) );
  NAND2_X1 U923 ( .A1(n829), .A2(G2106), .ZN(n828) );
  XOR2_X1 U924 ( .A(KEYINPUT107), .B(n828), .Z(G217) );
  INV_X1 U925 ( .A(n829), .ZN(G223) );
  AND2_X1 U926 ( .A1(G15), .A2(G2), .ZN(n830) );
  NAND2_X1 U927 ( .A1(G661), .A2(n830), .ZN(G259) );
  NAND2_X1 U928 ( .A1(G3), .A2(G1), .ZN(n831) );
  NAND2_X1 U929 ( .A1(n832), .A2(n831), .ZN(G188) );
  INV_X1 U930 ( .A(n833), .ZN(G319) );
  XOR2_X1 U931 ( .A(G120), .B(KEYINPUT108), .Z(G236) );
  INV_X1 U933 ( .A(G96), .ZN(G221) );
  INV_X1 U934 ( .A(G69), .ZN(G235) );
  INV_X1 U935 ( .A(G57), .ZN(G237) );
  NOR2_X1 U936 ( .A1(n835), .A2(n834), .ZN(G325) );
  INV_X1 U937 ( .A(G325), .ZN(G261) );
  XOR2_X1 U938 ( .A(G2100), .B(G2096), .Z(n837) );
  XNOR2_X1 U939 ( .A(KEYINPUT42), .B(G2678), .ZN(n836) );
  XNOR2_X1 U940 ( .A(n837), .B(n836), .ZN(n841) );
  XOR2_X1 U941 ( .A(KEYINPUT43), .B(G2090), .Z(n839) );
  XNOR2_X1 U942 ( .A(G2067), .B(G2072), .ZN(n838) );
  XNOR2_X1 U943 ( .A(n839), .B(n838), .ZN(n840) );
  XOR2_X1 U944 ( .A(n841), .B(n840), .Z(n843) );
  XNOR2_X1 U945 ( .A(G2078), .B(G2084), .ZN(n842) );
  XNOR2_X1 U946 ( .A(n843), .B(n842), .ZN(G227) );
  XOR2_X1 U947 ( .A(KEYINPUT110), .B(G1976), .Z(n845) );
  XNOR2_X1 U948 ( .A(G1986), .B(G1971), .ZN(n844) );
  XNOR2_X1 U949 ( .A(n845), .B(n844), .ZN(n846) );
  XOR2_X1 U950 ( .A(n846), .B(KEYINPUT41), .Z(n848) );
  XNOR2_X1 U951 ( .A(G1996), .B(G1991), .ZN(n847) );
  XNOR2_X1 U952 ( .A(n848), .B(n847), .ZN(n852) );
  XNOR2_X1 U953 ( .A(G1981), .B(n963), .ZN(n850) );
  XNOR2_X1 U954 ( .A(G1966), .B(G1961), .ZN(n849) );
  XNOR2_X1 U955 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U956 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U957 ( .A(KEYINPUT109), .B(G2474), .ZN(n853) );
  XNOR2_X1 U958 ( .A(n854), .B(n853), .ZN(G229) );
  NAND2_X1 U959 ( .A1(G124), .A2(n886), .ZN(n855) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n855), .Z(n856) );
  XNOR2_X1 U961 ( .A(n856), .B(KEYINPUT44), .ZN(n858) );
  NAND2_X1 U962 ( .A1(G112), .A2(n887), .ZN(n857) );
  NAND2_X1 U963 ( .A1(n858), .A2(n857), .ZN(n862) );
  NAND2_X1 U964 ( .A1(G136), .A2(n881), .ZN(n860) );
  NAND2_X1 U965 ( .A1(G100), .A2(n882), .ZN(n859) );
  NAND2_X1 U966 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U967 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U968 ( .A(KEYINPUT114), .B(KEYINPUT46), .Z(n864) );
  XNOR2_X1 U969 ( .A(KEYINPUT115), .B(KEYINPUT48), .ZN(n863) );
  XNOR2_X1 U970 ( .A(n864), .B(n863), .ZN(n865) );
  XOR2_X1 U971 ( .A(G164), .B(n865), .Z(n876) );
  NAND2_X1 U972 ( .A1(G130), .A2(n886), .ZN(n867) );
  NAND2_X1 U973 ( .A1(G118), .A2(n887), .ZN(n866) );
  NAND2_X1 U974 ( .A1(n867), .A2(n866), .ZN(n872) );
  NAND2_X1 U975 ( .A1(G142), .A2(n881), .ZN(n869) );
  NAND2_X1 U976 ( .A1(G106), .A2(n882), .ZN(n868) );
  NAND2_X1 U977 ( .A1(n869), .A2(n868), .ZN(n870) );
  XOR2_X1 U978 ( .A(n870), .B(KEYINPUT45), .Z(n871) );
  NOR2_X1 U979 ( .A1(n872), .A2(n871), .ZN(n874) );
  XNOR2_X1 U980 ( .A(n874), .B(n873), .ZN(n875) );
  XNOR2_X1 U981 ( .A(n876), .B(n875), .ZN(n879) );
  XNOR2_X1 U982 ( .A(n877), .B(n918), .ZN(n878) );
  XNOR2_X1 U983 ( .A(n879), .B(n878), .ZN(n880) );
  XOR2_X1 U984 ( .A(n880), .B(G162), .Z(n896) );
  NAND2_X1 U985 ( .A1(G139), .A2(n881), .ZN(n884) );
  NAND2_X1 U986 ( .A1(G103), .A2(n882), .ZN(n883) );
  NAND2_X1 U987 ( .A1(n884), .A2(n883), .ZN(n885) );
  XNOR2_X1 U988 ( .A(KEYINPUT112), .B(n885), .ZN(n893) );
  NAND2_X1 U989 ( .A1(G127), .A2(n886), .ZN(n889) );
  NAND2_X1 U990 ( .A1(G115), .A2(n887), .ZN(n888) );
  NAND2_X1 U991 ( .A1(n889), .A2(n888), .ZN(n890) );
  XNOR2_X1 U992 ( .A(KEYINPUT113), .B(n890), .ZN(n891) );
  XNOR2_X1 U993 ( .A(KEYINPUT47), .B(n891), .ZN(n892) );
  NOR2_X1 U994 ( .A1(n893), .A2(n892), .ZN(n909) );
  XOR2_X1 U995 ( .A(n894), .B(n909), .Z(n895) );
  XNOR2_X1 U996 ( .A(n896), .B(n895), .ZN(n897) );
  XOR2_X1 U997 ( .A(G160), .B(n897), .Z(n898) );
  NOR2_X1 U998 ( .A1(G37), .A2(n898), .ZN(G395) );
  XOR2_X1 U999 ( .A(G286), .B(n899), .Z(n901) );
  XNOR2_X1 U1000 ( .A(n901), .B(n900), .ZN(n902) );
  XOR2_X1 U1001 ( .A(n902), .B(G301), .Z(n903) );
  NOR2_X1 U1002 ( .A1(G37), .A2(n903), .ZN(G397) );
  NOR2_X1 U1003 ( .A1(G227), .A2(G229), .ZN(n904) );
  XNOR2_X1 U1004 ( .A(KEYINPUT49), .B(n904), .ZN(n905) );
  NOR2_X1 U1005 ( .A1(G401), .A2(n905), .ZN(n906) );
  AND2_X1 U1006 ( .A1(G319), .A2(n906), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G395), .A2(G397), .ZN(n907) );
  NAND2_X1 U1008 ( .A1(n908), .A2(n907), .ZN(G225) );
  INV_X1 U1009 ( .A(G225), .ZN(G308) );
  INV_X1 U1010 ( .A(KEYINPUT55), .ZN(n957) );
  XNOR2_X1 U1011 ( .A(KEYINPUT118), .B(KEYINPUT52), .ZN(n933) );
  XOR2_X1 U1012 ( .A(G2072), .B(n909), .Z(n911) );
  XOR2_X1 U1013 ( .A(G164), .B(G2078), .Z(n910) );
  NOR2_X1 U1014 ( .A1(n911), .A2(n910), .ZN(n912) );
  XNOR2_X1 U1015 ( .A(n912), .B(KEYINPUT50), .ZN(n913) );
  XNOR2_X1 U1016 ( .A(n913), .B(KEYINPUT117), .ZN(n927) );
  XNOR2_X1 U1017 ( .A(G160), .B(G2084), .ZN(n925) );
  XNOR2_X1 U1018 ( .A(G2090), .B(G162), .ZN(n914) );
  XNOR2_X1 U1019 ( .A(n914), .B(KEYINPUT116), .ZN(n915) );
  NAND2_X1 U1020 ( .A1(n916), .A2(n915), .ZN(n917) );
  XNOR2_X1 U1021 ( .A(n917), .B(KEYINPUT51), .ZN(n921) );
  NOR2_X1 U1022 ( .A1(n919), .A2(n918), .ZN(n920) );
  NAND2_X1 U1023 ( .A1(n921), .A2(n920), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n926) );
  NOR2_X1 U1026 ( .A1(n927), .A2(n926), .ZN(n929) );
  NAND2_X1 U1027 ( .A1(n929), .A2(n928), .ZN(n930) );
  NOR2_X1 U1028 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1029 ( .A(n933), .B(n932), .ZN(n934) );
  NAND2_X1 U1030 ( .A1(n957), .A2(n934), .ZN(n935) );
  NAND2_X1 U1031 ( .A1(n935), .A2(G29), .ZN(n1020) );
  XOR2_X1 U1032 ( .A(G2090), .B(G35), .Z(n952) );
  XNOR2_X1 U1033 ( .A(G27), .B(n936), .ZN(n940) );
  XNOR2_X1 U1034 ( .A(G2067), .B(G26), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(G33), .B(G2072), .ZN(n937) );
  NOR2_X1 U1036 ( .A1(n938), .A2(n937), .ZN(n939) );
  NAND2_X1 U1037 ( .A1(n940), .A2(n939), .ZN(n943) );
  XNOR2_X1 U1038 ( .A(KEYINPUT120), .B(G1996), .ZN(n941) );
  XNOR2_X1 U1039 ( .A(G32), .B(n941), .ZN(n942) );
  NOR2_X1 U1040 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1041 ( .A(KEYINPUT121), .B(n944), .ZN(n948) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n945) );
  NAND2_X1 U1043 ( .A1(G28), .A2(n945), .ZN(n946) );
  XOR2_X1 U1044 ( .A(n946), .B(KEYINPUT119), .Z(n947) );
  NOR2_X1 U1045 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1046 ( .A(KEYINPUT122), .B(n949), .Z(n950) );
  XNOR2_X1 U1047 ( .A(n950), .B(KEYINPUT53), .ZN(n951) );
  NAND2_X1 U1048 ( .A1(n952), .A2(n951), .ZN(n955) );
  XNOR2_X1 U1049 ( .A(G34), .B(G2084), .ZN(n953) );
  XNOR2_X1 U1050 ( .A(KEYINPUT54), .B(n953), .ZN(n954) );
  NOR2_X1 U1051 ( .A1(n955), .A2(n954), .ZN(n956) );
  XNOR2_X1 U1052 ( .A(n957), .B(n956), .ZN(n958) );
  NOR2_X1 U1053 ( .A1(G29), .A2(n958), .ZN(n1016) );
  INV_X1 U1054 ( .A(G16), .ZN(n1012) );
  XOR2_X1 U1055 ( .A(n1012), .B(KEYINPUT56), .Z(n989) );
  XNOR2_X1 U1056 ( .A(G1966), .B(G168), .ZN(n960) );
  NAND2_X1 U1057 ( .A1(n960), .A2(n959), .ZN(n961) );
  XNOR2_X1 U1058 ( .A(KEYINPUT57), .B(n961), .ZN(n987) );
  XOR2_X1 U1059 ( .A(n962), .B(G1348), .Z(n968) );
  XNOR2_X1 U1060 ( .A(n964), .B(n963), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n979) );
  INV_X1 U1063 ( .A(n969), .ZN(n970) );
  NAND2_X1 U1064 ( .A1(n971), .A2(n970), .ZN(n972) );
  XNOR2_X1 U1065 ( .A(n972), .B(KEYINPUT123), .ZN(n974) );
  NAND2_X1 U1066 ( .A1(G1971), .A2(G303), .ZN(n973) );
  NAND2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n976) );
  NOR2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  XOR2_X1 U1069 ( .A(KEYINPUT124), .B(n977), .Z(n978) );
  NOR2_X1 U1070 ( .A1(n979), .A2(n978), .ZN(n984) );
  XOR2_X1 U1071 ( .A(n980), .B(G1341), .Z(n982) );
  XNOR2_X1 U1072 ( .A(G301), .B(G1961), .ZN(n981) );
  NOR2_X1 U1073 ( .A1(n982), .A2(n981), .ZN(n983) );
  NAND2_X1 U1074 ( .A1(n984), .A2(n983), .ZN(n985) );
  XNOR2_X1 U1075 ( .A(KEYINPUT125), .B(n985), .ZN(n986) );
  NAND2_X1 U1076 ( .A1(n987), .A2(n986), .ZN(n988) );
  NAND2_X1 U1077 ( .A1(n989), .A2(n988), .ZN(n1014) );
  XOR2_X1 U1078 ( .A(G20), .B(G1956), .Z(n993) );
  XNOR2_X1 U1079 ( .A(G1341), .B(G19), .ZN(n991) );
  XNOR2_X1 U1080 ( .A(G6), .B(G1981), .ZN(n990) );
  NOR2_X1 U1081 ( .A1(n991), .A2(n990), .ZN(n992) );
  NAND2_X1 U1082 ( .A1(n993), .A2(n992), .ZN(n996) );
  XOR2_X1 U1083 ( .A(KEYINPUT59), .B(G1348), .Z(n994) );
  XNOR2_X1 U1084 ( .A(G4), .B(n994), .ZN(n995) );
  NOR2_X1 U1085 ( .A1(n996), .A2(n995), .ZN(n997) );
  XNOR2_X1 U1086 ( .A(KEYINPUT60), .B(n997), .ZN(n1001) );
  XNOR2_X1 U1087 ( .A(G1966), .B(G21), .ZN(n999) );
  XNOR2_X1 U1088 ( .A(G1961), .B(G5), .ZN(n998) );
  NOR2_X1 U1089 ( .A1(n999), .A2(n998), .ZN(n1000) );
  NAND2_X1 U1090 ( .A1(n1001), .A2(n1000), .ZN(n1009) );
  XNOR2_X1 U1091 ( .A(G1971), .B(G22), .ZN(n1003) );
  XNOR2_X1 U1092 ( .A(G23), .B(G1976), .ZN(n1002) );
  NOR2_X1 U1093 ( .A1(n1003), .A2(n1002), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(G1986), .B(KEYINPUT126), .Z(n1004) );
  XNOR2_X1 U1095 ( .A(G24), .B(n1004), .ZN(n1005) );
  NAND2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  XNOR2_X1 U1097 ( .A(KEYINPUT58), .B(n1007), .ZN(n1008) );
  NOR2_X1 U1098 ( .A1(n1009), .A2(n1008), .ZN(n1010) );
  XNOR2_X1 U1099 ( .A(KEYINPUT61), .B(n1010), .ZN(n1011) );
  NAND2_X1 U1100 ( .A1(n1012), .A2(n1011), .ZN(n1013) );
  NAND2_X1 U1101 ( .A1(n1014), .A2(n1013), .ZN(n1015) );
  NOR2_X1 U1102 ( .A1(n1016), .A2(n1015), .ZN(n1017) );
  NAND2_X1 U1103 ( .A1(G11), .A2(n1017), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(KEYINPUT127), .B(n1018), .ZN(n1019) );
  NAND2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT62), .B(n1021), .ZN(G150) );
  INV_X1 U1107 ( .A(G150), .ZN(G311) );
endmodule

