

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, n346,
         n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357,
         n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368,
         n369, n370, n371, n372, n373, n374, n375, n376, n377, n378, n379,
         n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, n390,
         n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401,
         n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412,
         n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
         n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434,
         n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
         n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456,
         n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467,
         n468, n469, n470, n471, n472, n473, n474, n475, n476, n477, n478,
         n479, n480, n481, n482, n483, n484, n485, n486, n487, n488, n489,
         n490, n491, n492, n493, n494, n495, n496, n497, n498, n499, n500,
         n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, n511,
         n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
         n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533,
         n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544,
         n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555,
         n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566,
         n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
         n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588,
         n589, n590, n591, n592, n593, n594, n595, n596, n597;

  XNOR2_X1 U324 ( .A(KEYINPUT47), .B(KEYINPUT111), .ZN(n470) );
  XNOR2_X1 U325 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U326 ( .A(n431), .B(n294), .ZN(n390) );
  INV_X1 U327 ( .A(KEYINPUT68), .ZN(n326) );
  XNOR2_X1 U328 ( .A(n474), .B(KEYINPUT48), .ZN(n555) );
  XNOR2_X1 U329 ( .A(n471), .B(n470), .ZN(n472) );
  XNOR2_X1 U330 ( .A(n481), .B(KEYINPUT119), .ZN(n575) );
  XNOR2_X1 U331 ( .A(n369), .B(n368), .ZN(n567) );
  XNOR2_X1 U332 ( .A(n398), .B(n397), .ZN(n400) );
  XNOR2_X1 U333 ( .A(n396), .B(n293), .ZN(n397) );
  XOR2_X1 U334 ( .A(n396), .B(n322), .Z(n292) );
  XOR2_X1 U335 ( .A(G204GAT), .B(G92GAT), .Z(n293) );
  AND2_X1 U336 ( .A1(G226GAT), .A2(G233GAT), .ZN(n294) );
  NOR2_X1 U337 ( .A1(n478), .A2(n533), .ZN(n295) );
  XOR2_X1 U338 ( .A(KEYINPUT45), .B(n464), .Z(n296) );
  INV_X1 U339 ( .A(KEYINPUT23), .ZN(n427) );
  INV_X1 U340 ( .A(KEYINPUT73), .ZN(n350) );
  XNOR2_X1 U341 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U342 ( .A(n351), .B(n350), .ZN(n352) );
  XNOR2_X1 U343 ( .A(n430), .B(n429), .ZN(n432) );
  XNOR2_X1 U344 ( .A(n353), .B(n352), .ZN(n356) );
  INV_X1 U345 ( .A(n437), .ZN(n438) );
  XNOR2_X1 U346 ( .A(KEYINPUT100), .B(KEYINPUT36), .ZN(n370) );
  XNOR2_X1 U347 ( .A(n327), .B(n326), .ZN(n328) );
  XNOR2_X1 U348 ( .A(n439), .B(n438), .ZN(n440) );
  XNOR2_X1 U349 ( .A(n550), .B(n370), .ZN(n463) );
  XNOR2_X1 U350 ( .A(n329), .B(n328), .ZN(n330) );
  XNOR2_X1 U351 ( .A(n441), .B(n440), .ZN(n442) );
  NOR2_X1 U352 ( .A1(n480), .A2(n525), .ZN(n481) );
  XNOR2_X1 U353 ( .A(n367), .B(n366), .ZN(n368) );
  NAND2_X1 U354 ( .A1(n445), .A2(n444), .ZN(n541) );
  INV_X1 U355 ( .A(G190GAT), .ZN(n482) );
  INV_X1 U356 ( .A(KEYINPUT120), .ZN(n492) );
  XOR2_X1 U357 ( .A(KEYINPUT108), .B(n458), .Z(n537) );
  XNOR2_X1 U358 ( .A(n483), .B(n482), .ZN(n484) );
  XNOR2_X1 U359 ( .A(G106GAT), .B(KEYINPUT44), .ZN(n460) );
  XNOR2_X1 U360 ( .A(n489), .B(n298), .ZN(n490) );
  XNOR2_X1 U361 ( .A(n485), .B(n484), .ZN(G1351GAT) );
  XNOR2_X1 U362 ( .A(n491), .B(n490), .ZN(G1328GAT) );
  INV_X1 U363 ( .A(G43GAT), .ZN(n297) );
  NAND2_X1 U364 ( .A1(G29GAT), .A2(n297), .ZN(n300) );
  INV_X1 U365 ( .A(G29GAT), .ZN(n298) );
  NAND2_X1 U366 ( .A1(n298), .A2(G43GAT), .ZN(n299) );
  NAND2_X1 U367 ( .A1(n300), .A2(n299), .ZN(n302) );
  XNOR2_X1 U368 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n301) );
  XNOR2_X1 U369 ( .A(n302), .B(n301), .ZN(n353) );
  XOR2_X1 U370 ( .A(G1GAT), .B(KEYINPUT66), .Z(n337) );
  XOR2_X1 U371 ( .A(n353), .B(n337), .Z(n304) );
  NAND2_X1 U372 ( .A1(G229GAT), .A2(G233GAT), .ZN(n303) );
  XNOR2_X1 U373 ( .A(n304), .B(n303), .ZN(n308) );
  XOR2_X1 U374 ( .A(KEYINPUT30), .B(KEYINPUT65), .Z(n306) );
  XNOR2_X1 U375 ( .A(G8GAT), .B(KEYINPUT29), .ZN(n305) );
  XNOR2_X1 U376 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U377 ( .A(n308), .B(n307), .Z(n316) );
  XOR2_X1 U378 ( .A(G15GAT), .B(G36GAT), .Z(n310) );
  XNOR2_X1 U379 ( .A(G169GAT), .B(G50GAT), .ZN(n309) );
  XNOR2_X1 U380 ( .A(n310), .B(n309), .ZN(n314) );
  XOR2_X1 U381 ( .A(G141GAT), .B(G197GAT), .Z(n312) );
  XNOR2_X1 U382 ( .A(G113GAT), .B(G22GAT), .ZN(n311) );
  XNOR2_X1 U383 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U384 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U385 ( .A(n316), .B(n315), .Z(n557) );
  XOR2_X1 U386 ( .A(G78GAT), .B(G148GAT), .Z(n318) );
  XNOR2_X1 U387 ( .A(KEYINPUT67), .B(G204GAT), .ZN(n317) );
  XNOR2_X1 U388 ( .A(n318), .B(n317), .ZN(n430) );
  XNOR2_X1 U389 ( .A(G71GAT), .B(G57GAT), .ZN(n319) );
  XNOR2_X1 U390 ( .A(n319), .B(KEYINPUT13), .ZN(n343) );
  XNOR2_X1 U391 ( .A(n430), .B(n343), .ZN(n331) );
  XOR2_X1 U392 ( .A(G176GAT), .B(G64GAT), .Z(n396) );
  XOR2_X1 U393 ( .A(KEYINPUT31), .B(KEYINPUT32), .Z(n321) );
  XNOR2_X1 U394 ( .A(G120GAT), .B(KEYINPUT33), .ZN(n320) );
  XNOR2_X1 U395 ( .A(n321), .B(n320), .ZN(n322) );
  NAND2_X1 U396 ( .A1(G230GAT), .A2(G233GAT), .ZN(n323) );
  XNOR2_X1 U397 ( .A(n292), .B(n323), .ZN(n329) );
  XOR2_X1 U398 ( .A(G92GAT), .B(G85GAT), .Z(n325) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G106GAT), .ZN(n324) );
  XNOR2_X1 U400 ( .A(n325), .B(n324), .ZN(n363) );
  XNOR2_X1 U401 ( .A(n363), .B(KEYINPUT69), .ZN(n327) );
  XNOR2_X1 U402 ( .A(n331), .B(n330), .ZN(n462) );
  XOR2_X1 U403 ( .A(KEYINPUT41), .B(n462), .Z(n559) );
  INV_X1 U404 ( .A(n559), .ZN(n570) );
  NOR2_X1 U405 ( .A1(n557), .A2(n570), .ZN(n519) );
  XOR2_X1 U406 ( .A(KEYINPUT12), .B(KEYINPUT77), .Z(n333) );
  XNOR2_X1 U407 ( .A(KEYINPUT79), .B(KEYINPUT76), .ZN(n332) );
  XNOR2_X1 U408 ( .A(n333), .B(n332), .ZN(n349) );
  XOR2_X1 U409 ( .A(G22GAT), .B(G155GAT), .Z(n435) );
  XOR2_X1 U410 ( .A(G64GAT), .B(n435), .Z(n335) );
  XOR2_X1 U411 ( .A(G15GAT), .B(G127GAT), .Z(n379) );
  XNOR2_X1 U412 ( .A(n379), .B(G78GAT), .ZN(n334) );
  XNOR2_X1 U413 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U414 ( .A(n337), .B(n336), .ZN(n347) );
  XOR2_X1 U415 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n339) );
  NAND2_X1 U416 ( .A1(G231GAT), .A2(G233GAT), .ZN(n338) );
  XNOR2_X1 U417 ( .A(n339), .B(n338), .ZN(n340) );
  XOR2_X1 U418 ( .A(n340), .B(KEYINPUT78), .Z(n345) );
  XOR2_X1 U419 ( .A(KEYINPUT75), .B(G211GAT), .Z(n342) );
  XNOR2_X1 U420 ( .A(G8GAT), .B(G183GAT), .ZN(n341) );
  XNOR2_X1 U421 ( .A(n342), .B(n341), .ZN(n391) );
  XNOR2_X1 U422 ( .A(n391), .B(n343), .ZN(n344) );
  XNOR2_X1 U423 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U424 ( .A(n347), .B(n346), .ZN(n348) );
  XOR2_X1 U425 ( .A(n349), .B(n348), .Z(n495) );
  NAND2_X1 U426 ( .A1(G232GAT), .A2(G233GAT), .ZN(n351) );
  INV_X1 U427 ( .A(n356), .ZN(n355) );
  INV_X1 U428 ( .A(KEYINPUT64), .ZN(n354) );
  NAND2_X1 U429 ( .A1(n355), .A2(n354), .ZN(n358) );
  NAND2_X1 U430 ( .A1(n356), .A2(KEYINPUT64), .ZN(n357) );
  NAND2_X1 U431 ( .A1(n358), .A2(n357), .ZN(n360) );
  XOR2_X1 U432 ( .A(G50GAT), .B(G162GAT), .Z(n436) );
  XOR2_X1 U433 ( .A(n436), .B(KEYINPUT10), .Z(n359) );
  XNOR2_X1 U434 ( .A(n360), .B(n359), .ZN(n369) );
  XOR2_X1 U435 ( .A(KEYINPUT72), .B(G218GAT), .Z(n362) );
  XNOR2_X1 U436 ( .A(G36GAT), .B(G190GAT), .ZN(n361) );
  XNOR2_X1 U437 ( .A(n362), .B(n361), .ZN(n393) );
  XNOR2_X1 U438 ( .A(n393), .B(n363), .ZN(n367) );
  XOR2_X1 U439 ( .A(KEYINPUT9), .B(KEYINPUT71), .Z(n365) );
  XNOR2_X1 U440 ( .A(G134GAT), .B(KEYINPUT11), .ZN(n364) );
  XOR2_X1 U441 ( .A(n365), .B(n364), .Z(n366) );
  XOR2_X1 U442 ( .A(n567), .B(KEYINPUT74), .Z(n550) );
  XOR2_X1 U443 ( .A(KEYINPUT82), .B(KEYINPUT17), .Z(n372) );
  XNOR2_X1 U444 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n371) );
  XNOR2_X1 U445 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U446 ( .A(G169GAT), .B(n373), .ZN(n399) );
  XOR2_X1 U447 ( .A(KEYINPUT20), .B(KEYINPUT81), .Z(n375) );
  XNOR2_X1 U448 ( .A(G183GAT), .B(G176GAT), .ZN(n374) );
  XNOR2_X1 U449 ( .A(n375), .B(n374), .ZN(n388) );
  XOR2_X1 U450 ( .A(KEYINPUT80), .B(G190GAT), .Z(n377) );
  XNOR2_X1 U451 ( .A(G43GAT), .B(G99GAT), .ZN(n376) );
  XNOR2_X1 U452 ( .A(n377), .B(n376), .ZN(n378) );
  XOR2_X1 U453 ( .A(n379), .B(n378), .Z(n381) );
  NAND2_X1 U454 ( .A1(G227GAT), .A2(G233GAT), .ZN(n380) );
  XNOR2_X1 U455 ( .A(n381), .B(n380), .ZN(n382) );
  XOR2_X1 U456 ( .A(n382), .B(G71GAT), .Z(n386) );
  XOR2_X1 U457 ( .A(G120GAT), .B(KEYINPUT0), .Z(n384) );
  XNOR2_X1 U458 ( .A(G113GAT), .B(G134GAT), .ZN(n383) );
  XNOR2_X1 U459 ( .A(n384), .B(n383), .ZN(n418) );
  XNOR2_X1 U460 ( .A(n418), .B(KEYINPUT83), .ZN(n385) );
  XNOR2_X1 U461 ( .A(n386), .B(n385), .ZN(n387) );
  XOR2_X1 U462 ( .A(n388), .B(n387), .Z(n389) );
  XOR2_X1 U463 ( .A(n399), .B(n389), .Z(n539) );
  XOR2_X1 U464 ( .A(G197GAT), .B(KEYINPUT21), .Z(n431) );
  XOR2_X1 U465 ( .A(n392), .B(KEYINPUT92), .Z(n395) );
  XNOR2_X1 U466 ( .A(n393), .B(KEYINPUT91), .ZN(n394) );
  XNOR2_X1 U467 ( .A(n395), .B(n394), .ZN(n398) );
  XOR2_X1 U468 ( .A(n400), .B(n399), .Z(n401) );
  XNOR2_X1 U469 ( .A(n401), .B(KEYINPUT93), .ZN(n402) );
  XOR2_X1 U470 ( .A(KEYINPUT27), .B(n402), .Z(n448) );
  INV_X1 U471 ( .A(n448), .ZN(n445) );
  XOR2_X1 U472 ( .A(KEYINPUT6), .B(KEYINPUT86), .Z(n404) );
  XNOR2_X1 U473 ( .A(G148GAT), .B(G155GAT), .ZN(n403) );
  XNOR2_X1 U474 ( .A(n404), .B(n403), .ZN(n408) );
  XOR2_X1 U475 ( .A(KEYINPUT90), .B(G57GAT), .Z(n406) );
  XNOR2_X1 U476 ( .A(G1GAT), .B(KEYINPUT1), .ZN(n405) );
  XNOR2_X1 U477 ( .A(n406), .B(n405), .ZN(n407) );
  XOR2_X1 U478 ( .A(n408), .B(n407), .Z(n415) );
  XOR2_X1 U479 ( .A(KEYINPUT84), .B(KEYINPUT3), .Z(n410) );
  XNOR2_X1 U480 ( .A(G141GAT), .B(KEYINPUT2), .ZN(n409) );
  XNOR2_X1 U481 ( .A(n410), .B(n409), .ZN(n437) );
  XOR2_X1 U482 ( .A(G85GAT), .B(n437), .Z(n412) );
  XNOR2_X1 U483 ( .A(G29GAT), .B(G162GAT), .ZN(n411) );
  XNOR2_X1 U484 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U485 ( .A(G127GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U486 ( .A(n415), .B(n414), .ZN(n424) );
  XOR2_X1 U487 ( .A(KEYINPUT88), .B(KEYINPUT87), .Z(n417) );
  XNOR2_X1 U488 ( .A(KEYINPUT5), .B(KEYINPUT89), .ZN(n416) );
  XNOR2_X1 U489 ( .A(n417), .B(n416), .ZN(n422) );
  XOR2_X1 U490 ( .A(n418), .B(KEYINPUT4), .Z(n420) );
  NAND2_X1 U491 ( .A1(G225GAT), .A2(G233GAT), .ZN(n419) );
  XNOR2_X1 U492 ( .A(n420), .B(n419), .ZN(n421) );
  XOR2_X1 U493 ( .A(n422), .B(n421), .Z(n423) );
  XOR2_X1 U494 ( .A(n424), .B(n423), .Z(n533) );
  XOR2_X1 U495 ( .A(KEYINPUT24), .B(KEYINPUT22), .Z(n426) );
  XNOR2_X1 U496 ( .A(G211GAT), .B(KEYINPUT85), .ZN(n425) );
  XNOR2_X1 U497 ( .A(n426), .B(n425), .ZN(n443) );
  NAND2_X1 U498 ( .A1(G228GAT), .A2(G233GAT), .ZN(n428) );
  XOR2_X1 U499 ( .A(n432), .B(n431), .Z(n434) );
  XNOR2_X1 U500 ( .A(G218GAT), .B(G106GAT), .ZN(n433) );
  XNOR2_X1 U501 ( .A(n434), .B(n433), .ZN(n441) );
  XNOR2_X1 U502 ( .A(n436), .B(n435), .ZN(n439) );
  XOR2_X1 U503 ( .A(n443), .B(n442), .Z(n478) );
  XOR2_X1 U504 ( .A(n478), .B(KEYINPUT28), .Z(n529) );
  AND2_X1 U505 ( .A1(n533), .A2(n529), .ZN(n444) );
  XNOR2_X1 U506 ( .A(n541), .B(KEYINPUT94), .ZN(n446) );
  NOR2_X1 U507 ( .A1(n539), .A2(n446), .ZN(n455) );
  INV_X1 U508 ( .A(n539), .ZN(n525) );
  NAND2_X1 U509 ( .A1(n478), .A2(n525), .ZN(n447) );
  XNOR2_X1 U510 ( .A(n447), .B(KEYINPUT26), .ZN(n581) );
  NOR2_X1 U511 ( .A1(n581), .A2(n448), .ZN(n554) );
  NOR2_X1 U512 ( .A1(n525), .A2(n401), .ZN(n449) );
  NOR2_X1 U513 ( .A1(n478), .A2(n449), .ZN(n450) );
  XNOR2_X1 U514 ( .A(n450), .B(KEYINPUT95), .ZN(n451) );
  XNOR2_X1 U515 ( .A(n451), .B(KEYINPUT25), .ZN(n452) );
  NOR2_X1 U516 ( .A1(n554), .A2(n452), .ZN(n453) );
  NOR2_X1 U517 ( .A1(n533), .A2(n453), .ZN(n454) );
  NOR2_X1 U518 ( .A1(n455), .A2(n454), .ZN(n497) );
  NOR2_X1 U519 ( .A1(n463), .A2(n497), .ZN(n456) );
  NAND2_X1 U520 ( .A1(n495), .A2(n456), .ZN(n457) );
  XNOR2_X1 U521 ( .A(KEYINPUT37), .B(n457), .ZN(n487) );
  NAND2_X1 U522 ( .A1(n519), .A2(n487), .ZN(n458) );
  INV_X1 U523 ( .A(n529), .ZN(n459) );
  NAND2_X1 U524 ( .A1(n537), .A2(n459), .ZN(n461) );
  XNOR2_X1 U525 ( .A(n461), .B(n460), .ZN(G1339GAT) );
  NOR2_X1 U526 ( .A1(n495), .A2(n463), .ZN(n464) );
  NOR2_X1 U527 ( .A1(n462), .A2(n296), .ZN(n465) );
  INV_X1 U528 ( .A(n557), .ZN(n582) );
  NAND2_X1 U529 ( .A1(n465), .A2(n582), .ZN(n473) );
  XNOR2_X1 U530 ( .A(KEYINPUT46), .B(KEYINPUT110), .ZN(n467) );
  NOR2_X1 U531 ( .A1(n582), .A2(n570), .ZN(n466) );
  XNOR2_X1 U532 ( .A(n467), .B(n466), .ZN(n468) );
  NOR2_X1 U533 ( .A1(n567), .A2(n468), .ZN(n469) );
  XOR2_X1 U534 ( .A(KEYINPUT109), .B(n495), .Z(n576) );
  NAND2_X1 U535 ( .A1(n469), .A2(n576), .ZN(n471) );
  NAND2_X1 U536 ( .A1(n473), .A2(n472), .ZN(n474) );
  INV_X1 U537 ( .A(n401), .ZN(n535) );
  NAND2_X1 U538 ( .A1(n555), .A2(n535), .ZN(n477) );
  XNOR2_X1 U539 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n475) );
  XNOR2_X1 U540 ( .A(n475), .B(KEYINPUT54), .ZN(n476) );
  XNOR2_X1 U541 ( .A(n477), .B(n476), .ZN(n579) );
  AND2_X1 U542 ( .A1(n579), .A2(n295), .ZN(n479) );
  XNOR2_X1 U543 ( .A(n479), .B(KEYINPUT55), .ZN(n480) );
  NOR2_X1 U544 ( .A1(n550), .A2(n575), .ZN(n485) );
  XNOR2_X1 U545 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n483) );
  NOR2_X1 U546 ( .A1(n462), .A2(n582), .ZN(n486) );
  XNOR2_X1 U547 ( .A(n486), .B(KEYINPUT70), .ZN(n500) );
  NAND2_X1 U548 ( .A1(n487), .A2(n500), .ZN(n488) );
  XNOR2_X1 U549 ( .A(KEYINPUT38), .B(n488), .ZN(n516) );
  INV_X1 U550 ( .A(n533), .ZN(n578) );
  NOR2_X1 U551 ( .A1(n516), .A2(n578), .ZN(n491) );
  XNOR2_X1 U552 ( .A(KEYINPUT99), .B(KEYINPUT39), .ZN(n489) );
  NOR2_X1 U553 ( .A1(n582), .A2(n575), .ZN(n494) );
  XNOR2_X1 U554 ( .A(n492), .B(G169GAT), .ZN(n493) );
  XNOR2_X1 U555 ( .A(n494), .B(n493), .ZN(G1348GAT) );
  INV_X1 U556 ( .A(n495), .ZN(n590) );
  NAND2_X1 U557 ( .A1(n550), .A2(n590), .ZN(n496) );
  XNOR2_X1 U558 ( .A(KEYINPUT16), .B(n496), .ZN(n498) );
  NOR2_X1 U559 ( .A1(n498), .A2(n497), .ZN(n499) );
  XNOR2_X1 U560 ( .A(n499), .B(KEYINPUT96), .ZN(n518) );
  NAND2_X1 U561 ( .A1(n500), .A2(n518), .ZN(n508) );
  NOR2_X1 U562 ( .A1(n578), .A2(n508), .ZN(n501) );
  XOR2_X1 U563 ( .A(G1GAT), .B(n501), .Z(n502) );
  XNOR2_X1 U564 ( .A(KEYINPUT34), .B(n502), .ZN(G1324GAT) );
  NOR2_X1 U565 ( .A1(n401), .A2(n508), .ZN(n504) );
  XNOR2_X1 U566 ( .A(G8GAT), .B(KEYINPUT97), .ZN(n503) );
  XNOR2_X1 U567 ( .A(n504), .B(n503), .ZN(G1325GAT) );
  NOR2_X1 U568 ( .A1(n525), .A2(n508), .ZN(n506) );
  XNOR2_X1 U569 ( .A(KEYINPUT98), .B(KEYINPUT35), .ZN(n505) );
  XNOR2_X1 U570 ( .A(n506), .B(n505), .ZN(n507) );
  XNOR2_X1 U571 ( .A(G15GAT), .B(n507), .ZN(G1326GAT) );
  NOR2_X1 U572 ( .A1(n529), .A2(n508), .ZN(n509) );
  XOR2_X1 U573 ( .A(G22GAT), .B(n509), .Z(G1327GAT) );
  NOR2_X1 U574 ( .A1(n516), .A2(n401), .ZN(n511) );
  XNOR2_X1 U575 ( .A(G36GAT), .B(KEYINPUT101), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1329GAT) );
  XOR2_X1 U577 ( .A(KEYINPUT103), .B(KEYINPUT40), .Z(n513) );
  XNOR2_X1 U578 ( .A(G43GAT), .B(KEYINPUT102), .ZN(n512) );
  XNOR2_X1 U579 ( .A(n513), .B(n512), .ZN(n515) );
  NOR2_X1 U580 ( .A1(n525), .A2(n516), .ZN(n514) );
  XOR2_X1 U581 ( .A(n515), .B(n514), .Z(G1330GAT) );
  NOR2_X1 U582 ( .A1(n516), .A2(n529), .ZN(n517) );
  XOR2_X1 U583 ( .A(G50GAT), .B(n517), .Z(G1331GAT) );
  NAND2_X1 U584 ( .A1(n519), .A2(n518), .ZN(n528) );
  NOR2_X1 U585 ( .A1(n578), .A2(n528), .ZN(n521) );
  XNOR2_X1 U586 ( .A(KEYINPUT104), .B(KEYINPUT42), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n522) );
  XOR2_X1 U588 ( .A(G57GAT), .B(n522), .Z(G1332GAT) );
  NOR2_X1 U589 ( .A1(n401), .A2(n528), .ZN(n524) );
  XNOR2_X1 U590 ( .A(G64GAT), .B(KEYINPUT105), .ZN(n523) );
  XNOR2_X1 U591 ( .A(n524), .B(n523), .ZN(G1333GAT) );
  NOR2_X1 U592 ( .A1(n525), .A2(n528), .ZN(n526) );
  XOR2_X1 U593 ( .A(KEYINPUT106), .B(n526), .Z(n527) );
  XNOR2_X1 U594 ( .A(G71GAT), .B(n527), .ZN(G1334GAT) );
  NOR2_X1 U595 ( .A1(n529), .A2(n528), .ZN(n531) );
  XNOR2_X1 U596 ( .A(KEYINPUT43), .B(KEYINPUT107), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n532) );
  XOR2_X1 U598 ( .A(G78GAT), .B(n532), .Z(G1335GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n533), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(G85GAT), .ZN(G1336GAT) );
  NAND2_X1 U601 ( .A1(n537), .A2(n535), .ZN(n536) );
  XNOR2_X1 U602 ( .A(n536), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U603 ( .A1(n537), .A2(n539), .ZN(n538) );
  XNOR2_X1 U604 ( .A(n538), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U605 ( .A1(n555), .A2(n539), .ZN(n540) );
  NOR2_X1 U606 ( .A1(n541), .A2(n540), .ZN(n545) );
  NAND2_X1 U607 ( .A1(n557), .A2(n545), .ZN(n542) );
  XNOR2_X1 U608 ( .A(n542), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U609 ( .A(G120GAT), .B(KEYINPUT49), .Z(n544) );
  NAND2_X1 U610 ( .A1(n545), .A2(n559), .ZN(n543) );
  XNOR2_X1 U611 ( .A(n544), .B(n543), .ZN(G1341GAT) );
  INV_X1 U612 ( .A(n545), .ZN(n549) );
  NOR2_X1 U613 ( .A1(n576), .A2(n549), .ZN(n547) );
  XNOR2_X1 U614 ( .A(KEYINPUT50), .B(KEYINPUT112), .ZN(n546) );
  XNOR2_X1 U615 ( .A(n547), .B(n546), .ZN(n548) );
  XOR2_X1 U616 ( .A(G127GAT), .B(n548), .Z(G1342GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n552) );
  XNOR2_X1 U618 ( .A(KEYINPUT113), .B(KEYINPUT51), .ZN(n551) );
  XNOR2_X1 U619 ( .A(n552), .B(n551), .ZN(n553) );
  XOR2_X1 U620 ( .A(G134GAT), .B(n553), .Z(G1343GAT) );
  NAND2_X1 U621 ( .A1(n555), .A2(n554), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n578), .A2(n556), .ZN(n568) );
  NAND2_X1 U623 ( .A1(n557), .A2(n568), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n558), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U625 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n563) );
  XOR2_X1 U626 ( .A(KEYINPUT52), .B(KEYINPUT114), .Z(n561) );
  NAND2_X1 U627 ( .A1(n568), .A2(n559), .ZN(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(G1345GAT) );
  XOR2_X1 U630 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n565) );
  NAND2_X1 U631 ( .A1(n568), .A2(n590), .ZN(n564) );
  XNOR2_X1 U632 ( .A(n565), .B(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(G155GAT), .B(n566), .ZN(G1346GAT) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n569), .B(G162GAT), .ZN(G1347GAT) );
  NOR2_X1 U636 ( .A1(n575), .A2(n570), .ZN(n574) );
  XOR2_X1 U637 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n572) );
  XNOR2_X1 U638 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n571) );
  XNOR2_X1 U639 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1349GAT) );
  NOR2_X1 U641 ( .A1(n576), .A2(n575), .ZN(n577) );
  XOR2_X1 U642 ( .A(G183GAT), .B(n577), .Z(G1350GAT) );
  NAND2_X1 U643 ( .A1(n579), .A2(n578), .ZN(n580) );
  NOR2_X1 U644 ( .A1(n581), .A2(n580), .ZN(n591) );
  INV_X1 U645 ( .A(n591), .ZN(n594) );
  NOR2_X1 U646 ( .A1(n594), .A2(n582), .ZN(n586) );
  XOR2_X1 U647 ( .A(KEYINPUT60), .B(KEYINPUT59), .Z(n584) );
  XNOR2_X1 U648 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n583) );
  XNOR2_X1 U649 ( .A(n584), .B(n583), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1352GAT) );
  XOR2_X1 U651 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n588) );
  NAND2_X1 U652 ( .A1(n591), .A2(n462), .ZN(n587) );
  XNOR2_X1 U653 ( .A(n588), .B(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(G204GAT), .B(n589), .ZN(G1353GAT) );
  XOR2_X1 U655 ( .A(G211GAT), .B(KEYINPUT125), .Z(n593) );
  NAND2_X1 U656 ( .A1(n591), .A2(n590), .ZN(n592) );
  XNOR2_X1 U657 ( .A(n593), .B(n592), .ZN(G1354GAT) );
  NOR2_X1 U658 ( .A1(n463), .A2(n594), .ZN(n596) );
  XNOR2_X1 U659 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n595) );
  XNOR2_X1 U660 ( .A(n596), .B(n595), .ZN(n597) );
  XOR2_X1 U661 ( .A(G218GAT), .B(n597), .Z(G1355GAT) );
endmodule

