//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 1 1 1 1 0 1 1 1 1 1 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 1 1 0 1 0 0 0 1 1 0 0 1 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:56 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n724, new_n725, new_n726, new_n728, new_n729,
    new_n730, new_n731, new_n732, new_n734, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n808, new_n809, new_n811, new_n812, new_n814, new_n815,
    new_n816, new_n817, new_n818, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n936, new_n937;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(G15gat), .B(G22gat), .ZN(new_n203));
  INV_X1    g002(.A(G1gat), .ZN(new_n204));
  NAND2_X1  g003(.A1(new_n204), .A2(KEYINPUT16), .ZN(new_n205));
  AND2_X1   g004(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g005(.A1(new_n203), .A2(G1gat), .ZN(new_n207));
  NOR3_X1   g006(.A1(new_n206), .A2(new_n207), .A3(G8gat), .ZN(new_n208));
  INV_X1    g007(.A(G8gat), .ZN(new_n209));
  OR2_X1    g008(.A1(new_n203), .A2(G1gat), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n203), .A2(new_n205), .ZN(new_n211));
  AOI21_X1  g010(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  OR2_X1    g011(.A1(G43gat), .A2(G50gat), .ZN(new_n213));
  NAND2_X1  g012(.A1(G43gat), .A2(G50gat), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND2_X1  g014(.A1(new_n215), .A2(KEYINPUT15), .ZN(new_n216));
  NAND2_X1  g015(.A1(G29gat), .A2(G36gat), .ZN(new_n217));
  XNOR2_X1  g016(.A(new_n217), .B(KEYINPUT95), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT15), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n213), .A2(new_n219), .A3(new_n214), .ZN(new_n220));
  INV_X1    g019(.A(KEYINPUT14), .ZN(new_n221));
  INV_X1    g020(.A(G29gat), .ZN(new_n222));
  INV_X1    g021(.A(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  OAI21_X1  g023(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  AND4_X1   g025(.A1(new_n216), .A2(new_n218), .A3(new_n220), .A4(new_n226), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(KEYINPUT94), .ZN(new_n228));
  INV_X1    g027(.A(KEYINPUT94), .ZN(new_n229));
  OAI211_X1 g028(.A(new_n229), .B(KEYINPUT14), .C1(G29gat), .C2(G36gat), .ZN(new_n230));
  NAND3_X1  g029(.A1(new_n228), .A2(new_n230), .A3(new_n224), .ZN(new_n231));
  AOI21_X1  g030(.A(new_n216), .B1(new_n231), .B2(new_n217), .ZN(new_n232));
  OAI22_X1  g031(.A1(new_n208), .A2(new_n212), .B1(new_n227), .B2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n231), .A2(new_n217), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n234), .A2(KEYINPUT15), .A3(new_n215), .ZN(new_n235));
  NAND4_X1  g034(.A1(new_n216), .A2(new_n218), .A3(new_n220), .A4(new_n226), .ZN(new_n236));
  NAND3_X1  g035(.A1(new_n235), .A2(KEYINPUT17), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n208), .A2(new_n212), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  AOI21_X1  g038(.A(KEYINPUT17), .B1(new_n235), .B2(new_n236), .ZN(new_n240));
  OAI211_X1 g039(.A(new_n202), .B(new_n233), .C1(new_n239), .C2(new_n240), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT18), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n241), .A2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT99), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  XNOR2_X1  g044(.A(G113gat), .B(G141gat), .ZN(new_n246));
  XNOR2_X1  g045(.A(G169gat), .B(G197gat), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT93), .B(KEYINPUT11), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n248), .B(new_n249), .ZN(new_n250));
  XOR2_X1   g049(.A(new_n250), .B(KEYINPUT12), .Z(new_n251));
  NAND2_X1  g050(.A1(new_n245), .A2(new_n251), .ZN(new_n252));
  OAI21_X1  g051(.A(KEYINPUT96), .B1(new_n241), .B2(new_n242), .ZN(new_n253));
  OAI21_X1  g052(.A(G8gat), .B1(new_n206), .B2(new_n207), .ZN(new_n254));
  NAND3_X1  g053(.A1(new_n210), .A2(new_n209), .A3(new_n211), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n254), .A2(new_n255), .ZN(new_n256));
  NOR2_X1   g055(.A1(new_n227), .A2(new_n232), .ZN(new_n257));
  AOI21_X1  g056(.A(new_n256), .B1(new_n257), .B2(KEYINPUT17), .ZN(new_n258));
  INV_X1    g057(.A(new_n240), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n235), .A2(new_n236), .ZN(new_n260));
  AOI22_X1  g059(.A1(new_n258), .A2(new_n259), .B1(new_n260), .B2(new_n256), .ZN(new_n261));
  INV_X1    g060(.A(KEYINPUT96), .ZN(new_n262));
  NAND4_X1  g061(.A1(new_n261), .A2(new_n262), .A3(KEYINPUT18), .A4(new_n202), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n253), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g063(.A1(new_n235), .A2(new_n236), .A3(new_n254), .A4(new_n255), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n233), .A2(new_n265), .A3(KEYINPUT97), .ZN(new_n266));
  XOR2_X1   g065(.A(new_n202), .B(KEYINPUT13), .Z(new_n267));
  INV_X1    g066(.A(KEYINPUT97), .ZN(new_n268));
  NAND3_X1  g067(.A1(new_n260), .A2(new_n268), .A3(new_n256), .ZN(new_n269));
  NAND3_X1  g068(.A1(new_n266), .A2(new_n267), .A3(new_n269), .ZN(new_n270));
  NAND2_X1  g069(.A1(new_n270), .A2(KEYINPUT98), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT98), .ZN(new_n272));
  NAND4_X1  g071(.A1(new_n266), .A2(new_n272), .A3(new_n267), .A4(new_n269), .ZN(new_n273));
  AOI22_X1  g072(.A1(new_n271), .A2(new_n273), .B1(new_n242), .B2(new_n241), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n252), .A2(new_n264), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n252), .B1(new_n264), .B2(new_n274), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  NAND2_X1  g076(.A1(G99gat), .A2(G106gat), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n278), .A2(KEYINPUT8), .ZN(new_n279));
  NAND2_X1  g078(.A1(G85gat), .A2(G92gat), .ZN(new_n280));
  INV_X1    g079(.A(KEYINPUT7), .ZN(new_n281));
  NAND2_X1  g080(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(G85gat), .ZN(new_n283));
  INV_X1    g082(.A(G92gat), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND3_X1  g084(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n286));
  NAND4_X1  g085(.A1(new_n279), .A2(new_n282), .A3(new_n285), .A4(new_n286), .ZN(new_n287));
  XNOR2_X1  g086(.A(G99gat), .B(G106gat), .ZN(new_n288));
  INV_X1    g087(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  AOI22_X1  g089(.A1(KEYINPUT8), .A2(new_n278), .B1(new_n283), .B2(new_n284), .ZN(new_n291));
  NAND4_X1  g090(.A1(new_n291), .A2(new_n288), .A3(new_n282), .A4(new_n286), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n290), .A2(new_n292), .ZN(new_n293));
  NAND3_X1  g092(.A1(new_n259), .A2(new_n237), .A3(new_n293), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n290), .A2(new_n292), .ZN(new_n295));
  AND2_X1   g094(.A1(G232gat), .A2(G233gat), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n260), .A2(new_n295), .B1(KEYINPUT41), .B2(new_n296), .ZN(new_n297));
  AND2_X1   g096(.A1(new_n297), .A2(KEYINPUT103), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n297), .A2(KEYINPUT103), .ZN(new_n299));
  OAI21_X1  g098(.A(new_n294), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(G190gat), .B(G218gat), .Z(new_n301));
  OR2_X1    g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n296), .A2(KEYINPUT41), .ZN(new_n303));
  XNOR2_X1  g102(.A(G134gat), .B(G162gat), .ZN(new_n304));
  XNOR2_X1  g103(.A(new_n303), .B(new_n304), .ZN(new_n305));
  NAND2_X1  g104(.A1(new_n300), .A2(new_n301), .ZN(new_n306));
  AND3_X1   g105(.A1(new_n302), .A2(new_n305), .A3(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n305), .B1(new_n302), .B2(new_n306), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n309), .ZN(new_n310));
  INV_X1    g109(.A(G64gat), .ZN(new_n311));
  NAND3_X1  g110(.A1(new_n311), .A2(KEYINPUT100), .A3(G57gat), .ZN(new_n312));
  INV_X1    g111(.A(KEYINPUT9), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n313), .A2(G71gat), .A3(G78gat), .ZN(new_n314));
  NAND2_X1  g113(.A1(G71gat), .A2(G78gat), .ZN(new_n315));
  INV_X1    g114(.A(new_n315), .ZN(new_n316));
  OAI21_X1  g115(.A(new_n312), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n311), .A2(G57gat), .ZN(new_n318));
  INV_X1    g117(.A(G57gat), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n319), .A2(G64gat), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT100), .ZN(new_n321));
  AND3_X1   g120(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  AOI21_X1  g121(.A(new_n313), .B1(new_n318), .B2(new_n320), .ZN(new_n323));
  OR2_X1    g122(.A1(G71gat), .A2(G78gat), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n324), .A2(new_n315), .ZN(new_n325));
  OAI22_X1  g124(.A1(new_n317), .A2(new_n322), .B1(new_n323), .B2(new_n325), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT21), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  NAND2_X1  g127(.A1(G231gat), .A2(G233gat), .ZN(new_n329));
  XNOR2_X1  g128(.A(new_n328), .B(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(new_n330), .B(G127gat), .ZN(new_n331));
  OAI21_X1  g130(.A(new_n238), .B1(new_n327), .B2(new_n326), .ZN(new_n332));
  OR2_X1    g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n331), .A2(new_n332), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n335), .B(KEYINPUT101), .ZN(new_n336));
  XNOR2_X1  g135(.A(new_n336), .B(G155gat), .ZN(new_n337));
  XNOR2_X1  g136(.A(G183gat), .B(G211gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n338), .B(KEYINPUT102), .ZN(new_n339));
  XNOR2_X1  g138(.A(new_n337), .B(new_n339), .ZN(new_n340));
  AND3_X1   g139(.A1(new_n333), .A2(new_n334), .A3(new_n340), .ZN(new_n341));
  AOI21_X1  g140(.A(new_n340), .B1(new_n333), .B2(new_n334), .ZN(new_n342));
  NOR2_X1   g141(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n293), .A2(new_n326), .ZN(new_n344));
  INV_X1    g143(.A(KEYINPUT10), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n318), .A2(new_n320), .A3(new_n321), .ZN(new_n346));
  OAI211_X1 g145(.A(new_n346), .B(new_n312), .C1(new_n316), .C2(new_n314), .ZN(new_n347));
  XNOR2_X1  g146(.A(G57gat), .B(G64gat), .ZN(new_n348));
  OAI211_X1 g147(.A(new_n315), .B(new_n324), .C1(new_n348), .C2(new_n313), .ZN(new_n349));
  NAND4_X1  g148(.A1(new_n347), .A2(new_n290), .A3(new_n349), .A4(new_n292), .ZN(new_n350));
  NAND3_X1  g149(.A1(new_n344), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  NAND4_X1  g150(.A1(new_n295), .A2(KEYINPUT10), .A3(new_n347), .A4(new_n349), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G230gat), .A2(G233gat), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n344), .A2(new_n350), .ZN(new_n356));
  INV_X1    g155(.A(new_n354), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n355), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G120gat), .B(G148gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(G176gat), .B(G204gat), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  INV_X1    g161(.A(new_n362), .ZN(new_n363));
  NOR2_X1   g162(.A1(new_n359), .A2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n364), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n359), .A2(new_n363), .ZN(new_n366));
  AND2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n310), .A2(new_n343), .A3(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G8gat), .B(G36gat), .ZN(new_n369));
  XNOR2_X1  g168(.A(G64gat), .B(G92gat), .ZN(new_n370));
  XOR2_X1   g169(.A(new_n369), .B(new_n370), .Z(new_n371));
  INV_X1    g170(.A(new_n371), .ZN(new_n372));
  NAND2_X1  g171(.A1(G169gat), .A2(G176gat), .ZN(new_n373));
  XNOR2_X1  g172(.A(new_n373), .B(KEYINPUT66), .ZN(new_n374));
  NOR2_X1   g173(.A1(G169gat), .A2(G176gat), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT23), .ZN(new_n376));
  AND3_X1   g175(.A1(new_n374), .A2(KEYINPUT67), .A3(new_n376), .ZN(new_n377));
  NAND3_X1  g176(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n378));
  OAI21_X1  g177(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n379));
  INV_X1    g178(.A(new_n379), .ZN(new_n380));
  AND2_X1   g179(.A1(G183gat), .A2(G190gat), .ZN(new_n381));
  OAI21_X1  g180(.A(new_n378), .B1(new_n380), .B2(new_n381), .ZN(new_n382));
  AND2_X1   g181(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n383));
  NOR2_X1   g182(.A1(KEYINPUT65), .A2(KEYINPUT23), .ZN(new_n384));
  OAI22_X1  g183(.A1(new_n383), .A2(new_n384), .B1(G169gat), .B2(G176gat), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n382), .A2(new_n385), .A3(KEYINPUT25), .ZN(new_n386));
  AOI21_X1  g185(.A(KEYINPUT67), .B1(new_n374), .B2(new_n376), .ZN(new_n387));
  OR3_X1    g186(.A1(new_n377), .A2(new_n386), .A3(new_n387), .ZN(new_n388));
  INV_X1    g187(.A(KEYINPUT25), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT64), .ZN(new_n390));
  OAI211_X1 g189(.A(new_n382), .B(new_n374), .C1(new_n390), .C2(new_n376), .ZN(new_n391));
  AOI22_X1  g190(.A1(new_n385), .A2(KEYINPUT64), .B1(KEYINPUT23), .B2(new_n375), .ZN(new_n392));
  OAI21_X1  g191(.A(new_n389), .B1(new_n391), .B2(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n388), .A2(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(KEYINPUT27), .B(G183gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(KEYINPUT69), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  INV_X1    g196(.A(G190gat), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n398), .A2(KEYINPUT28), .ZN(new_n399));
  AND2_X1   g198(.A1(new_n395), .A2(new_n398), .ZN(new_n400));
  OAI22_X1  g199(.A1(new_n397), .A2(new_n399), .B1(KEYINPUT28), .B2(new_n400), .ZN(new_n401));
  XNOR2_X1  g200(.A(new_n375), .B(KEYINPUT26), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n381), .B1(new_n402), .B2(new_n374), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n401), .A2(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n394), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT77), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND3_X1  g206(.A1(new_n394), .A2(new_n404), .A3(KEYINPUT77), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n407), .A2(new_n408), .ZN(new_n409));
  AND2_X1   g208(.A1(G226gat), .A2(G233gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n409), .A2(new_n410), .ZN(new_n411));
  XNOR2_X1  g210(.A(KEYINPUT75), .B(G197gat), .ZN(new_n412));
  XNOR2_X1  g211(.A(new_n412), .B(G204gat), .ZN(new_n413));
  INV_X1    g212(.A(G211gat), .ZN(new_n414));
  INV_X1    g213(.A(G218gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  OAI21_X1  g215(.A(new_n413), .B1(KEYINPUT22), .B2(new_n416), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n417), .A2(KEYINPUT76), .ZN(new_n418));
  XOR2_X1   g217(.A(G211gat), .B(G218gat), .Z(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n418), .B(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT68), .ZN(new_n423));
  AND3_X1   g222(.A1(new_n388), .A2(new_n423), .A3(new_n393), .ZN(new_n424));
  AOI21_X1  g223(.A(new_n423), .B1(new_n388), .B2(new_n393), .ZN(new_n425));
  OAI21_X1  g224(.A(new_n404), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  NOR2_X1   g225(.A1(new_n410), .A2(KEYINPUT29), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n426), .A2(new_n427), .ZN(new_n428));
  AND3_X1   g227(.A1(new_n411), .A2(new_n422), .A3(new_n428), .ZN(new_n429));
  NAND3_X1  g228(.A1(new_n407), .A2(new_n408), .A3(new_n427), .ZN(new_n430));
  OAI211_X1 g229(.A(new_n404), .B(new_n410), .C1(new_n424), .C2(new_n425), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n422), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n372), .B1(new_n429), .B2(new_n432), .ZN(new_n433));
  INV_X1    g232(.A(new_n432), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n411), .A2(new_n422), .A3(new_n428), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n371), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n433), .A2(KEYINPUT30), .A3(new_n436), .ZN(new_n437));
  INV_X1    g236(.A(KEYINPUT30), .ZN(new_n438));
  NAND4_X1  g237(.A1(new_n434), .A2(new_n435), .A3(new_n438), .A4(new_n371), .ZN(new_n439));
  AND2_X1   g238(.A1(new_n437), .A2(new_n439), .ZN(new_n440));
  XNOR2_X1  g239(.A(G155gat), .B(G162gat), .ZN(new_n441));
  NAND2_X1  g240(.A1(KEYINPUT82), .A2(G162gat), .ZN(new_n442));
  NAND2_X1  g241(.A1(new_n442), .A2(KEYINPUT2), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(G148gat), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n445), .A2(G141gat), .ZN(new_n446));
  XNOR2_X1  g245(.A(new_n446), .B(KEYINPUT80), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  XNOR2_X1  g247(.A(KEYINPUT78), .B(G141gat), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n449), .A2(G148gat), .ZN(new_n450));
  OR2_X1    g249(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n450), .A2(KEYINPUT79), .ZN(new_n452));
  AOI21_X1  g251(.A(new_n448), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n444), .B1(new_n453), .B2(KEYINPUT81), .ZN(new_n454));
  XNOR2_X1  g253(.A(new_n450), .B(KEYINPUT79), .ZN(new_n455));
  NAND2_X1  g254(.A1(new_n455), .A2(new_n447), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT81), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n454), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n441), .ZN(new_n460));
  XNOR2_X1  g259(.A(G141gat), .B(G148gat), .ZN(new_n461));
  OAI21_X1  g260(.A(new_n460), .B1(new_n461), .B2(KEYINPUT2), .ZN(new_n462));
  XOR2_X1   g261(.A(KEYINPUT83), .B(KEYINPUT3), .Z(new_n463));
  NAND3_X1  g262(.A1(new_n459), .A2(new_n462), .A3(new_n463), .ZN(new_n464));
  XNOR2_X1  g263(.A(KEYINPUT72), .B(KEYINPUT1), .ZN(new_n465));
  XOR2_X1   g264(.A(G127gat), .B(G134gat), .Z(new_n466));
  XNOR2_X1  g265(.A(KEYINPUT71), .B(G113gat), .ZN(new_n467));
  AOI211_X1 g266(.A(new_n465), .B(new_n466), .C1(G120gat), .C2(new_n467), .ZN(new_n468));
  OAI21_X1  g267(.A(new_n468), .B1(G120gat), .B2(new_n467), .ZN(new_n469));
  NOR2_X1   g268(.A1(G127gat), .A2(G134gat), .ZN(new_n470));
  XOR2_X1   g269(.A(KEYINPUT70), .B(G127gat), .Z(new_n471));
  AOI21_X1  g270(.A(new_n470), .B1(new_n471), .B2(G134gat), .ZN(new_n472));
  INV_X1    g271(.A(G113gat), .ZN(new_n473));
  INV_X1    g272(.A(G120gat), .ZN(new_n474));
  AOI21_X1  g273(.A(KEYINPUT1), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OAI21_X1  g274(.A(new_n475), .B1(new_n473), .B2(new_n474), .ZN(new_n476));
  NAND2_X1  g275(.A1(new_n472), .A2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n469), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT3), .ZN(new_n479));
  INV_X1    g278(.A(new_n462), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n480), .B1(new_n454), .B2(new_n458), .ZN(new_n481));
  OAI211_X1 g280(.A(new_n464), .B(new_n478), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  NAND2_X1  g281(.A1(G225gat), .A2(G233gat), .ZN(new_n483));
  INV_X1    g282(.A(new_n478), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n459), .A2(new_n484), .A3(new_n462), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n481), .A2(KEYINPUT4), .A3(new_n484), .ZN(new_n488));
  NAND4_X1  g287(.A1(new_n482), .A2(new_n483), .A3(new_n487), .A4(new_n488), .ZN(new_n489));
  XOR2_X1   g288(.A(KEYINPUT86), .B(KEYINPUT5), .Z(new_n490));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n491));
  NOR2_X1   g290(.A1(new_n490), .A2(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AND2_X1   g292(.A1(new_n487), .A2(new_n488), .ZN(new_n494));
  INV_X1    g293(.A(new_n492), .ZN(new_n495));
  NAND4_X1  g294(.A1(new_n494), .A2(new_n483), .A3(new_n482), .A4(new_n495), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n459), .A2(new_n462), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n498), .A2(new_n478), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n483), .B1(new_n499), .B2(new_n485), .ZN(new_n500));
  INV_X1    g299(.A(KEYINPUT85), .ZN(new_n501));
  AOI21_X1  g300(.A(new_n490), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(new_n481), .B(new_n478), .ZN(new_n503));
  OAI21_X1  g302(.A(KEYINPUT85), .B1(new_n503), .B2(new_n483), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g304(.A1(new_n497), .A2(new_n505), .ZN(new_n506));
  XOR2_X1   g305(.A(G1gat), .B(G29gat), .Z(new_n507));
  XNOR2_X1  g306(.A(G57gat), .B(G85gat), .ZN(new_n508));
  XNOR2_X1  g307(.A(new_n507), .B(new_n508), .ZN(new_n509));
  XNOR2_X1  g308(.A(KEYINPUT87), .B(KEYINPUT0), .ZN(new_n510));
  XNOR2_X1  g309(.A(new_n509), .B(new_n510), .ZN(new_n511));
  INV_X1    g310(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n506), .A2(new_n512), .ZN(new_n513));
  INV_X1    g312(.A(KEYINPUT6), .ZN(new_n514));
  AOI22_X1  g313(.A1(new_n493), .A2(new_n496), .B1(new_n502), .B2(new_n504), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n511), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n514), .B1(new_n515), .B2(new_n511), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n497), .A2(new_n511), .A3(new_n505), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g319(.A(new_n440), .B1(new_n517), .B2(new_n520), .ZN(new_n521));
  INV_X1    g320(.A(KEYINPUT29), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n421), .B1(new_n464), .B2(new_n522), .ZN(new_n523));
  INV_X1    g322(.A(KEYINPUT89), .ZN(new_n524));
  OR2_X1    g323(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n523), .A2(new_n524), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT88), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n419), .B1(new_n417), .B2(new_n527), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n528), .B1(new_n527), .B2(new_n417), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n417), .A2(new_n527), .A3(new_n420), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n530), .A2(new_n522), .ZN(new_n531));
  OAI21_X1  g330(.A(new_n463), .B1(new_n529), .B2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n532), .A2(new_n498), .B1(G228gat), .B2(G233gat), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n525), .A2(new_n526), .A3(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n421), .A2(new_n522), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n481), .B1(new_n535), .B2(new_n479), .ZN(new_n536));
  OAI211_X1 g335(.A(G228gat), .B(G233gat), .C1(new_n536), .C2(new_n523), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n534), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(KEYINPUT31), .B(G50gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n538), .A2(new_n539), .ZN(new_n540));
  XNOR2_X1  g339(.A(G78gat), .B(G106gat), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G22gat), .ZN(new_n542));
  INV_X1    g341(.A(new_n539), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n533), .ZN(new_n544));
  NOR2_X1   g343(.A1(new_n523), .A2(new_n524), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n537), .B(new_n543), .C1(new_n544), .C2(new_n545), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n540), .A2(new_n542), .A3(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(new_n542), .ZN(new_n548));
  INV_X1    g347(.A(new_n546), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n543), .B1(new_n534), .B2(new_n537), .ZN(new_n550));
  OAI21_X1  g349(.A(new_n548), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(KEYINPUT35), .ZN(new_n552));
  AND3_X1   g351(.A1(new_n547), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n521), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n426), .A2(new_n484), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n478), .B(new_n404), .C1(new_n424), .C2(new_n425), .ZN(new_n556));
  NAND4_X1  g355(.A1(new_n555), .A2(G227gat), .A3(G233gat), .A4(new_n556), .ZN(new_n557));
  XOR2_X1   g356(.A(G71gat), .B(G99gat), .Z(new_n558));
  XNOR2_X1  g357(.A(G15gat), .B(G43gat), .ZN(new_n559));
  XNOR2_X1  g358(.A(new_n558), .B(new_n559), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(KEYINPUT33), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n557), .A2(KEYINPUT32), .A3(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n562), .A2(KEYINPUT73), .ZN(new_n563));
  INV_X1    g362(.A(KEYINPUT73), .ZN(new_n564));
  NAND4_X1  g363(.A1(new_n557), .A2(new_n564), .A3(KEYINPUT32), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g364(.A1(new_n563), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n557), .A2(KEYINPUT32), .ZN(new_n567));
  INV_X1    g366(.A(new_n557), .ZN(new_n568));
  OAI211_X1 g367(.A(new_n567), .B(new_n560), .C1(new_n568), .C2(KEYINPUT33), .ZN(new_n569));
  NAND2_X1  g368(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n556), .ZN(new_n571));
  NAND2_X1  g370(.A1(G227gat), .A2(G233gat), .ZN(new_n572));
  NAND2_X1  g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  AND2_X1   g372(.A1(new_n573), .A2(KEYINPUT34), .ZN(new_n574));
  NOR2_X1   g373(.A1(new_n573), .A2(KEYINPUT34), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(new_n576), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n570), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n566), .A3(new_n569), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n578), .A2(KEYINPUT74), .A3(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(KEYINPUT74), .ZN(new_n581));
  NAND4_X1  g380(.A1(new_n576), .A2(new_n566), .A3(new_n581), .A4(new_n569), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n580), .A2(KEYINPUT92), .A3(new_n582), .ZN(new_n583));
  INV_X1    g382(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g383(.A(KEYINPUT92), .B1(new_n580), .B2(new_n582), .ZN(new_n585));
  OAI21_X1  g384(.A(new_n554), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n578), .A2(new_n579), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n547), .A2(new_n551), .ZN(new_n588));
  NOR2_X1   g387(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI21_X1  g388(.A(new_n552), .B1(new_n589), .B2(new_n521), .ZN(new_n590));
  INV_X1    g389(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n586), .A2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(KEYINPUT36), .ZN(new_n593));
  AOI21_X1  g392(.A(new_n593), .B1(new_n578), .B2(new_n579), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n580), .A2(new_n582), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n594), .B1(new_n595), .B2(new_n593), .ZN(new_n596));
  INV_X1    g395(.A(new_n588), .ZN(new_n597));
  NOR2_X1   g396(.A1(KEYINPUT90), .A2(KEYINPUT40), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT39), .ZN(new_n599));
  AOI21_X1  g398(.A(new_n599), .B1(new_n503), .B2(new_n483), .ZN(new_n600));
  INV_X1    g399(.A(new_n600), .ZN(new_n601));
  NAND2_X1  g400(.A1(new_n494), .A2(new_n482), .ZN(new_n602));
  INV_X1    g401(.A(new_n483), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n602), .A2(new_n599), .A3(new_n603), .ZN(new_n605));
  NAND2_X1  g404(.A1(new_n605), .A2(new_n512), .ZN(new_n606));
  OAI21_X1  g405(.A(new_n598), .B1(new_n604), .B2(new_n606), .ZN(new_n607));
  NAND2_X1  g406(.A1(new_n602), .A2(new_n603), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n608), .A2(new_n600), .ZN(new_n609));
  INV_X1    g408(.A(new_n598), .ZN(new_n610));
  NAND4_X1  g409(.A1(new_n609), .A2(new_n512), .A3(new_n610), .A4(new_n605), .ZN(new_n611));
  AND2_X1   g410(.A1(new_n607), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n437), .A2(new_n439), .ZN(new_n613));
  NOR2_X1   g412(.A1(new_n613), .A2(new_n519), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT91), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT37), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n617), .B1(new_n434), .B2(new_n435), .ZN(new_n618));
  OAI21_X1  g417(.A(new_n616), .B1(new_n618), .B2(new_n371), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n434), .A2(new_n617), .A3(new_n435), .ZN(new_n620));
  NAND2_X1  g419(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g420(.A1(new_n618), .A2(new_n616), .A3(new_n371), .ZN(new_n622));
  OAI21_X1  g421(.A(KEYINPUT38), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n411), .A2(new_n421), .A3(new_n428), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n430), .A2(new_n431), .ZN(new_n625));
  OAI211_X1 g424(.A(new_n624), .B(KEYINPUT37), .C1(new_n421), .C2(new_n625), .ZN(new_n626));
  NOR2_X1   g425(.A1(new_n371), .A2(KEYINPUT38), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n626), .A2(new_n620), .A3(new_n627), .ZN(new_n628));
  AND2_X1   g427(.A1(new_n628), .A2(new_n436), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n623), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n517), .A2(new_n520), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n597), .B(new_n615), .C1(new_n630), .C2(new_n631), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n613), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n633), .A2(new_n588), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n596), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  AOI211_X1 g434(.A(new_n277), .B(new_n368), .C1(new_n592), .C2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n631), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  XNOR2_X1  g437(.A(new_n638), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g438(.A1(new_n636), .A2(new_n440), .ZN(new_n640));
  NOR2_X1   g439(.A1(new_n640), .A2(KEYINPUT42), .ZN(new_n641));
  INV_X1    g440(.A(KEYINPUT42), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n642), .A2(KEYINPUT104), .ZN(new_n643));
  XNOR2_X1  g442(.A(new_n643), .B(KEYINPUT16), .ZN(new_n644));
  NAND3_X1  g443(.A1(new_n636), .A2(new_n440), .A3(new_n644), .ZN(new_n645));
  AOI21_X1  g444(.A(new_n641), .B1(G8gat), .B2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n646), .B1(G8gat), .B2(new_n645), .ZN(G1325gat));
  INV_X1    g446(.A(new_n596), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n636), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(new_n585), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n583), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g451(.A1(new_n652), .A2(G15gat), .ZN(new_n653));
  AOI22_X1  g452(.A1(new_n649), .A2(G15gat), .B1(new_n636), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g453(.A(new_n654), .B(KEYINPUT105), .Z(G1326gat));
  NAND2_X1  g454(.A1(new_n636), .A2(new_n588), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT106), .ZN(new_n657));
  XNOR2_X1  g456(.A(new_n656), .B(new_n657), .ZN(new_n658));
  XNOR2_X1  g457(.A(KEYINPUT43), .B(G22gat), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n656), .B(KEYINPUT106), .ZN(new_n661));
  INV_X1    g460(.A(new_n659), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n660), .A2(new_n663), .ZN(G1327gat));
  NAND2_X1  g463(.A1(new_n521), .A2(new_n553), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n665), .B1(new_n650), .B2(new_n583), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n635), .B1(new_n666), .B2(new_n590), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n667), .A2(new_n309), .ZN(new_n668));
  INV_X1    g467(.A(new_n367), .ZN(new_n669));
  NOR3_X1   g468(.A1(new_n277), .A2(new_n343), .A3(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n670), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  NAND3_X1  g471(.A1(new_n672), .A2(new_n222), .A3(new_n637), .ZN(new_n673));
  XNOR2_X1  g472(.A(new_n673), .B(KEYINPUT45), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n668), .A2(KEYINPUT44), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n633), .A2(KEYINPUT107), .A3(new_n588), .ZN(new_n676));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n677));
  OAI21_X1  g476(.A(new_n677), .B1(new_n521), .B2(new_n597), .ZN(new_n678));
  NAND4_X1  g477(.A1(new_n596), .A2(new_n632), .A3(new_n676), .A4(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n310), .B1(new_n592), .B2(new_n679), .ZN(new_n680));
  XOR2_X1   g479(.A(KEYINPUT108), .B(KEYINPUT44), .Z(new_n681));
  NAND2_X1  g480(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n671), .B1(new_n675), .B2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n683), .A2(new_n637), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n674), .B1(new_n222), .B2(new_n684), .ZN(G1328gat));
  NAND2_X1  g484(.A1(new_n675), .A2(new_n682), .ZN(new_n686));
  NAND3_X1  g485(.A1(new_n686), .A2(new_n440), .A3(new_n670), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT109), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n683), .A2(KEYINPUT109), .A3(new_n440), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(G36gat), .A3(new_n690), .ZN(new_n691));
  NOR4_X1   g490(.A1(new_n668), .A2(G36gat), .A3(new_n613), .A4(new_n671), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n692), .B(KEYINPUT46), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n691), .A2(new_n693), .ZN(G1329gat));
  NOR4_X1   g493(.A1(new_n668), .A2(G43gat), .A3(new_n652), .A4(new_n671), .ZN(new_n695));
  INV_X1    g494(.A(new_n681), .ZN(new_n696));
  AOI211_X1 g495(.A(new_n310), .B(new_n696), .C1(new_n592), .C2(new_n679), .ZN(new_n697));
  INV_X1    g496(.A(KEYINPUT44), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n698), .B1(new_n667), .B2(new_n309), .ZN(new_n699));
  OAI211_X1 g498(.A(new_n648), .B(new_n670), .C1(new_n697), .C2(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n695), .B1(new_n700), .B2(G43gat), .ZN(new_n701));
  XNOR2_X1  g500(.A(new_n701), .B(KEYINPUT47), .ZN(G1330gat));
  OAI211_X1 g501(.A(new_n588), .B(new_n670), .C1(new_n697), .C2(new_n699), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n703), .A2(G50gat), .ZN(new_n704));
  NOR2_X1   g503(.A1(new_n597), .A2(G50gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n705), .B(KEYINPUT110), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n672), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n704), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(KEYINPUT48), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND3_X1  g509(.A1(new_n704), .A2(KEYINPUT48), .A3(new_n707), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(G1331gat));
  INV_X1    g511(.A(new_n277), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n310), .A2(new_n343), .A3(new_n669), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n713), .B(new_n714), .C1(new_n592), .C2(new_n679), .ZN(new_n715));
  INV_X1    g514(.A(KEYINPUT111), .ZN(new_n716));
  NOR2_X1   g515(.A1(new_n518), .A2(new_n519), .ZN(new_n717));
  NOR3_X1   g516(.A1(new_n506), .A2(new_n514), .A3(new_n512), .ZN(new_n718));
  OAI21_X1  g517(.A(new_n716), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND3_X1  g518(.A1(new_n517), .A2(new_n520), .A3(KEYINPUT111), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND2_X1  g520(.A1(new_n715), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n722), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g522(.A1(new_n715), .A2(new_n440), .ZN(new_n724));
  OAI21_X1  g523(.A(new_n724), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n725));
  XOR2_X1   g524(.A(KEYINPUT49), .B(G64gat), .Z(new_n726));
  OAI21_X1  g525(.A(new_n725), .B1(new_n724), .B2(new_n726), .ZN(G1333gat));
  NAND3_X1  g526(.A1(new_n715), .A2(G71gat), .A3(new_n648), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT112), .ZN(new_n729));
  XNOR2_X1  g528(.A(new_n651), .B(new_n729), .ZN(new_n730));
  AND2_X1   g529(.A1(new_n715), .A2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n728), .B1(new_n731), .B2(G71gat), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g532(.A1(new_n715), .A2(new_n588), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G78gat), .ZN(G1335gat));
  NOR3_X1   g534(.A1(new_n631), .A2(G85gat), .A3(new_n367), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n713), .A2(new_n343), .ZN(new_n737));
  AND3_X1   g536(.A1(new_n680), .A2(KEYINPUT51), .A3(new_n737), .ZN(new_n738));
  AOI21_X1  g537(.A(KEYINPUT51), .B1(new_n680), .B2(new_n737), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n736), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n737), .A2(new_n669), .ZN(new_n741));
  AOI21_X1  g540(.A(new_n741), .B1(new_n675), .B2(new_n682), .ZN(new_n742));
  AND2_X1   g541(.A1(new_n742), .A2(new_n637), .ZN(new_n743));
  OAI21_X1  g542(.A(new_n740), .B1(new_n743), .B2(new_n283), .ZN(G1336gat));
  INV_X1    g543(.A(new_n741), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n440), .B(new_n745), .C1(new_n697), .C2(new_n699), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n746), .A2(G92gat), .ZN(new_n747));
  NOR3_X1   g546(.A1(new_n613), .A2(G92gat), .A3(new_n367), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n748), .B1(new_n738), .B2(new_n739), .ZN(new_n749));
  XNOR2_X1  g548(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n750));
  AND3_X1   g549(.A1(new_n747), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n750), .B1(new_n747), .B2(new_n749), .ZN(new_n752));
  NOR2_X1   g551(.A1(new_n751), .A2(new_n752), .ZN(G1337gat));
  NAND3_X1  g552(.A1(new_n686), .A2(new_n648), .A3(new_n745), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT114), .ZN(new_n755));
  INV_X1    g554(.A(KEYINPUT114), .ZN(new_n756));
  NAND3_X1  g555(.A1(new_n742), .A2(new_n756), .A3(new_n648), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n755), .A2(G99gat), .A3(new_n757), .ZN(new_n758));
  NOR3_X1   g557(.A1(new_n652), .A2(G99gat), .A3(new_n367), .ZN(new_n759));
  OAI21_X1  g558(.A(new_n759), .B1(new_n738), .B2(new_n739), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n758), .A2(new_n760), .ZN(G1338gat));
  OAI211_X1 g560(.A(new_n588), .B(new_n745), .C1(new_n697), .C2(new_n699), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n762), .A2(G106gat), .ZN(new_n763));
  NOR2_X1   g562(.A1(new_n367), .A2(G106gat), .ZN(new_n764));
  OAI211_X1 g563(.A(new_n588), .B(new_n764), .C1(new_n738), .C2(new_n739), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n766), .A2(KEYINPUT53), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT53), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n763), .A2(new_n765), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n767), .A2(new_n769), .ZN(G1339gat));
  NOR2_X1   g569(.A1(new_n261), .A2(new_n202), .ZN(new_n771));
  AOI21_X1  g570(.A(new_n267), .B1(new_n266), .B2(new_n269), .ZN(new_n772));
  OAI21_X1  g571(.A(new_n250), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n274), .A2(new_n264), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n773), .B1(new_n774), .B2(new_n251), .ZN(new_n775));
  INV_X1    g574(.A(KEYINPUT116), .ZN(new_n776));
  OR2_X1    g575(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  OAI21_X1  g576(.A(new_n363), .B1(new_n355), .B2(KEYINPUT54), .ZN(new_n778));
  NAND3_X1  g577(.A1(new_n351), .A2(new_n352), .A3(new_n357), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n355), .A2(KEYINPUT54), .A3(new_n779), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  NAND2_X1  g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NAND4_X1  g581(.A1(new_n355), .A2(KEYINPUT115), .A3(KEYINPUT54), .A4(new_n779), .ZN(new_n783));
  AOI21_X1  g582(.A(new_n778), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OR2_X1    g583(.A1(new_n784), .A2(KEYINPUT55), .ZN(new_n785));
  AOI21_X1  g584(.A(new_n364), .B1(new_n784), .B2(KEYINPUT55), .ZN(new_n786));
  AND2_X1   g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NAND2_X1  g586(.A1(new_n775), .A2(new_n776), .ZN(new_n788));
  NAND4_X1  g587(.A1(new_n777), .A2(new_n787), .A3(new_n309), .A4(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n775), .A2(new_n367), .ZN(new_n790));
  AOI21_X1  g589(.A(new_n790), .B1(new_n713), .B2(new_n787), .ZN(new_n791));
  OAI21_X1  g590(.A(new_n789), .B1(new_n791), .B2(new_n309), .ZN(new_n792));
  INV_X1    g591(.A(new_n343), .ZN(new_n793));
  NAND2_X1  g592(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n368), .A2(new_n713), .ZN(new_n795));
  INV_X1    g594(.A(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n588), .B1(new_n794), .B2(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n651), .A2(new_n637), .A3(new_n613), .A4(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(G113gat), .B1(new_n798), .B2(new_n277), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n794), .A2(new_n796), .ZN(new_n800));
  NAND2_X1  g599(.A1(new_n800), .A2(new_n721), .ZN(new_n801));
  INV_X1    g600(.A(new_n589), .ZN(new_n802));
  NOR3_X1   g601(.A1(new_n801), .A2(new_n440), .A3(new_n802), .ZN(new_n803));
  INV_X1    g602(.A(new_n803), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n713), .A2(new_n473), .ZN(new_n805));
  XNOR2_X1  g604(.A(new_n805), .B(KEYINPUT117), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n804), .B2(new_n806), .ZN(G1340gat));
  NOR3_X1   g606(.A1(new_n798), .A2(new_n474), .A3(new_n367), .ZN(new_n808));
  AOI21_X1  g607(.A(G120gat), .B1(new_n803), .B2(new_n669), .ZN(new_n809));
  NOR2_X1   g608(.A1(new_n808), .A2(new_n809), .ZN(G1341gat));
  OAI21_X1  g609(.A(new_n471), .B1(new_n798), .B2(new_n793), .ZN(new_n811));
  OR2_X1    g610(.A1(new_n793), .A2(new_n471), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n804), .B2(new_n812), .ZN(G1342gat));
  INV_X1    g612(.A(G134gat), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n803), .A2(new_n814), .A3(new_n309), .ZN(new_n815));
  NAND2_X1  g614(.A1(new_n815), .A2(KEYINPUT56), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(KEYINPUT118), .ZN(new_n817));
  OAI21_X1  g616(.A(G134gat), .B1(new_n798), .B2(new_n310), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n817), .B(new_n818), .C1(KEYINPUT56), .C2(new_n815), .ZN(G1343gat));
  INV_X1    g618(.A(new_n449), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT121), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n800), .A2(new_n588), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT57), .ZN(new_n823));
  AOI21_X1  g622(.A(new_n821), .B1(new_n822), .B2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  INV_X1    g624(.A(KEYINPUT119), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n825), .B1(new_n784), .B2(new_n826), .ZN(new_n827));
  AOI211_X1 g626(.A(KEYINPUT119), .B(new_n778), .C1(new_n782), .C2(new_n783), .ZN(new_n828));
  OAI21_X1  g627(.A(new_n786), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(KEYINPUT120), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  OAI211_X1 g630(.A(KEYINPUT120), .B(new_n786), .C1(new_n827), .C2(new_n828), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n831), .A2(new_n713), .A3(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n790), .ZN(new_n834));
  AOI21_X1  g633(.A(new_n309), .B1(new_n833), .B2(new_n834), .ZN(new_n835));
  INV_X1    g634(.A(new_n789), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n793), .B1(new_n835), .B2(new_n836), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n597), .B1(new_n837), .B2(new_n796), .ZN(new_n838));
  NAND2_X1  g637(.A1(new_n838), .A2(KEYINPUT57), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n824), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n838), .A2(new_n821), .A3(KEYINPUT57), .ZN(new_n841));
  NOR3_X1   g640(.A1(new_n648), .A2(new_n631), .A3(new_n440), .ZN(new_n842));
  NAND3_X1  g641(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n820), .B1(new_n843), .B2(new_n277), .ZN(new_n844));
  NAND2_X1  g643(.A1(new_n596), .A2(new_n588), .ZN(new_n845));
  NOR3_X1   g644(.A1(new_n845), .A2(new_n801), .A3(new_n440), .ZN(new_n846));
  INV_X1    g645(.A(G141gat), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n846), .A2(new_n847), .A3(new_n713), .ZN(new_n848));
  AND2_X1   g647(.A1(new_n844), .A2(new_n848), .ZN(new_n849));
  AOI21_X1  g648(.A(KEYINPUT58), .B1(new_n844), .B2(KEYINPUT122), .ZN(new_n850));
  XNOR2_X1  g649(.A(new_n849), .B(new_n850), .ZN(G1344gat));
  NAND3_X1  g650(.A1(new_n846), .A2(new_n445), .A3(new_n669), .ZN(new_n852));
  NOR2_X1   g651(.A1(new_n843), .A2(new_n367), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n853), .A2(KEYINPUT59), .A3(new_n445), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT59), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n277), .B1(new_n829), .B2(new_n830), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n790), .B1(new_n856), .B2(new_n832), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n789), .B1(new_n857), .B2(new_n309), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n795), .B1(new_n858), .B2(new_n793), .ZN(new_n859));
  OAI21_X1  g658(.A(new_n823), .B1(new_n859), .B2(new_n597), .ZN(new_n860));
  NAND3_X1  g659(.A1(new_n800), .A2(KEYINPUT57), .A3(new_n588), .ZN(new_n861));
  AOI21_X1  g660(.A(new_n367), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n862), .A2(new_n842), .ZN(new_n863));
  AOI21_X1  g662(.A(new_n855), .B1(new_n863), .B2(G148gat), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n852), .B1(new_n854), .B2(new_n864), .ZN(G1345gat));
  OAI21_X1  g664(.A(G155gat), .B1(new_n843), .B2(new_n793), .ZN(new_n866));
  INV_X1    g665(.A(G155gat), .ZN(new_n867));
  NAND3_X1  g666(.A1(new_n846), .A2(new_n867), .A3(new_n343), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n866), .A2(new_n868), .ZN(G1346gat));
  XNOR2_X1  g668(.A(KEYINPUT82), .B(G162gat), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n310), .A2(new_n870), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n846), .A2(new_n871), .ZN(new_n872));
  XOR2_X1   g671(.A(new_n872), .B(KEYINPUT123), .Z(new_n873));
  NAND4_X1  g672(.A1(new_n840), .A2(new_n309), .A3(new_n841), .A4(new_n842), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(KEYINPUT124), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n870), .B1(new_n874), .B2(KEYINPUT124), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n873), .B1(new_n875), .B2(new_n876), .ZN(new_n877));
  INV_X1    g676(.A(KEYINPUT125), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n877), .A2(new_n878), .ZN(new_n879));
  OAI211_X1 g678(.A(new_n873), .B(KEYINPUT125), .C1(new_n875), .C2(new_n876), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n879), .A2(new_n880), .ZN(G1347gat));
  AOI211_X1 g680(.A(new_n613), .B(new_n637), .C1(new_n794), .C2(new_n796), .ZN(new_n882));
  AND2_X1   g681(.A1(new_n882), .A2(new_n589), .ZN(new_n883));
  AOI21_X1  g682(.A(G169gat), .B1(new_n883), .B2(new_n713), .ZN(new_n884));
  AND3_X1   g683(.A1(new_n719), .A2(new_n720), .A3(new_n440), .ZN(new_n885));
  AND2_X1   g684(.A1(new_n797), .A2(new_n885), .ZN(new_n886));
  NAND2_X1  g685(.A1(new_n730), .A2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(new_n887), .ZN(new_n888));
  AND2_X1   g687(.A1(new_n713), .A2(G169gat), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n884), .B1(new_n888), .B2(new_n889), .ZN(G1348gat));
  OAI21_X1  g689(.A(G176gat), .B1(new_n887), .B2(new_n367), .ZN(new_n891));
  INV_X1    g690(.A(G176gat), .ZN(new_n892));
  NAND3_X1  g691(.A1(new_n883), .A2(new_n892), .A3(new_n669), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n891), .A2(new_n893), .ZN(G1349gat));
  NAND2_X1  g693(.A1(new_n888), .A2(new_n343), .ZN(new_n895));
  NOR2_X1   g694(.A1(new_n793), .A2(new_n397), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n895), .A2(G183gat), .B1(new_n883), .B2(new_n896), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT60), .ZN(new_n898));
  XNOR2_X1  g697(.A(new_n897), .B(new_n898), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n883), .A2(new_n398), .A3(new_n309), .ZN(new_n900));
  OAI21_X1  g699(.A(G190gat), .B1(new_n887), .B2(new_n310), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  INV_X1    g703(.A(new_n845), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n882), .ZN(new_n906));
  INV_X1    g705(.A(new_n906), .ZN(new_n907));
  AOI21_X1  g706(.A(G197gat), .B1(new_n907), .B2(new_n713), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n885), .A2(new_n596), .ZN(new_n909));
  AOI21_X1  g708(.A(new_n909), .B1(new_n860), .B2(new_n861), .ZN(new_n910));
  AND2_X1   g709(.A1(new_n713), .A2(G197gat), .ZN(new_n911));
  AOI21_X1  g710(.A(new_n908), .B1(new_n910), .B2(new_n911), .ZN(G1352gat));
  NOR3_X1   g711(.A1(new_n906), .A2(G204gat), .A3(new_n367), .ZN(new_n913));
  XNOR2_X1  g712(.A(new_n913), .B(KEYINPUT62), .ZN(new_n914));
  INV_X1    g713(.A(new_n909), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n862), .A2(new_n915), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n916), .A2(G204gat), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n914), .A2(new_n917), .ZN(G1353gat));
  INV_X1    g717(.A(KEYINPUT63), .ZN(new_n919));
  OAI21_X1  g718(.A(new_n861), .B1(new_n838), .B2(KEYINPUT57), .ZN(new_n920));
  INV_X1    g719(.A(KEYINPUT126), .ZN(new_n921));
  NAND4_X1  g720(.A1(new_n920), .A2(new_n921), .A3(new_n343), .A4(new_n915), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n922), .A2(G211gat), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n921), .B1(new_n910), .B2(new_n343), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n919), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  NAND3_X1  g724(.A1(new_n920), .A2(new_n343), .A3(new_n915), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n926), .A2(KEYINPUT126), .ZN(new_n927));
  NAND4_X1  g726(.A1(new_n927), .A2(KEYINPUT63), .A3(G211gat), .A4(new_n922), .ZN(new_n928));
  NAND2_X1  g727(.A1(new_n925), .A2(new_n928), .ZN(new_n929));
  NAND3_X1  g728(.A1(new_n907), .A2(new_n414), .A3(new_n343), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(KEYINPUT127), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND3_X1  g732(.A1(new_n929), .A2(KEYINPUT127), .A3(new_n930), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(G1354gat));
  NAND3_X1  g734(.A1(new_n907), .A2(new_n415), .A3(new_n309), .ZN(new_n936));
  AND2_X1   g735(.A1(new_n910), .A2(new_n309), .ZN(new_n937));
  OAI21_X1  g736(.A(new_n936), .B1(new_n937), .B2(new_n415), .ZN(G1355gat));
endmodule


