//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 1 1 0 1 0 1 1 0 0 0 1 1 1 0 0 1 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 0 0 0 0 0 0 0 1 0 1 1 0 0 1 0 1 1 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:34:30 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n443, new_n447, new_n449, new_n451, new_n454, new_n455,
    new_n456, new_n457, new_n458, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n517, new_n518, new_n519,
    new_n520, new_n521, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n531, new_n532, new_n533, new_n534, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n544,
    new_n546, new_n547, new_n548, new_n550, new_n551, new_n552, new_n553,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n569, new_n570,
    new_n571, new_n572, new_n573, new_n574, new_n576, new_n577, new_n578,
    new_n579, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n591, new_n594, new_n595, new_n597, new_n598,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n621, new_n622,
    new_n623, new_n624, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n823, new_n824, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1120, new_n1121;
  XOR2_X1   g000(.A(KEYINPUT64), .B(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  XNOR2_X1  g003(.A(KEYINPUT65), .B(G1083), .ZN(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XNOR2_X1  g007(.A(KEYINPUT66), .B(G2066), .ZN(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(new_n443));
  XOR2_X1   g018(.A(new_n443), .B(KEYINPUT67), .Z(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XOR2_X1   g020(.A(KEYINPUT68), .B(G452), .Z(G391));
  NAND2_X1  g021(.A1(G94), .A2(G452), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n447), .B(KEYINPUT69), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT70), .ZN(G234));
  NAND3_X1  g027(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g028(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n454));
  XOR2_X1   g029(.A(new_n454), .B(KEYINPUT2), .Z(new_n455));
  INV_X1    g030(.A(new_n455), .ZN(new_n456));
  NOR4_X1   g031(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n457));
  INV_X1    g032(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g033(.A1(new_n456), .A2(new_n458), .ZN(G325));
  INV_X1    g034(.A(G325), .ZN(G261));
  AOI22_X1  g035(.A1(new_n456), .A2(G2106), .B1(G567), .B2(new_n458), .ZN(G319));
  INV_X1    g036(.A(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(KEYINPUT3), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT3), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G2104), .ZN(new_n465));
  INV_X1    g040(.A(G2105), .ZN(new_n466));
  NAND3_X1  g041(.A1(new_n463), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  INV_X1    g042(.A(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n462), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G137), .B1(G101), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(G113), .A2(G2104), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n463), .A2(new_n465), .ZN(new_n472));
  INV_X1    g047(.A(G125), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n470), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(G160));
  NAND2_X1  g052(.A1(new_n468), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n466), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n472), .A2(new_n466), .ZN(new_n482));
  AOI21_X1  g057(.A(new_n481), .B1(G124), .B2(new_n482), .ZN(G162));
  AND2_X1   g058(.A1(KEYINPUT71), .A2(G114), .ZN(new_n484));
  NOR2_X1   g059(.A1(KEYINPUT71), .A2(G114), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  OAI211_X1 g061(.A(new_n486), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n487));
  INV_X1    g062(.A(KEYINPUT4), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(KEYINPUT72), .ZN(new_n489));
  INV_X1    g064(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g065(.A(G138), .B1(new_n488), .B2(KEYINPUT72), .ZN(new_n491));
  OAI21_X1  g066(.A(new_n490), .B1(new_n467), .B2(new_n491), .ZN(new_n492));
  XNOR2_X1  g067(.A(KEYINPUT3), .B(G2104), .ZN(new_n493));
  NAND3_X1  g068(.A1(new_n493), .A2(G126), .A3(G2105), .ZN(new_n494));
  INV_X1    g069(.A(G138), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT72), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n495), .B1(new_n496), .B2(KEYINPUT4), .ZN(new_n497));
  NAND4_X1  g072(.A1(new_n493), .A2(new_n497), .A3(new_n466), .A4(new_n489), .ZN(new_n498));
  NAND4_X1  g073(.A1(new_n487), .A2(new_n492), .A3(new_n494), .A4(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(G164));
  INV_X1    g075(.A(G543), .ZN(new_n501));
  NAND2_X1  g076(.A1(new_n501), .A2(KEYINPUT5), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT5), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n503), .A2(G543), .ZN(new_n504));
  AND2_X1   g079(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  AOI22_X1  g080(.A1(new_n505), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n506));
  INV_X1    g081(.A(G651), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  XNOR2_X1  g083(.A(KEYINPUT6), .B(G651), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n505), .A2(new_n509), .ZN(new_n510));
  INV_X1    g085(.A(G88), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n509), .A2(G543), .ZN(new_n512));
  INV_X1    g087(.A(G50), .ZN(new_n513));
  OAI22_X1  g088(.A1(new_n510), .A2(new_n511), .B1(new_n512), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g089(.A1(new_n508), .A2(new_n514), .ZN(G303));
  INV_X1    g090(.A(G303), .ZN(G166));
  NAND3_X1  g091(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n517));
  XNOR2_X1  g092(.A(new_n517), .B(KEYINPUT7), .ZN(new_n518));
  INV_X1    g093(.A(G89), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n518), .B1(new_n510), .B2(new_n519), .ZN(new_n520));
  INV_X1    g095(.A(KEYINPUT74), .ZN(new_n521));
  XNOR2_X1  g096(.A(new_n520), .B(new_n521), .ZN(new_n522));
  NAND3_X1  g097(.A1(new_n505), .A2(G63), .A3(G651), .ZN(new_n523));
  INV_X1    g098(.A(G51), .ZN(new_n524));
  OR2_X1    g099(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n525));
  NAND2_X1  g100(.A1(new_n512), .A2(KEYINPUT73), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(new_n527), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n522), .B(new_n523), .C1(new_n524), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AND2_X1   g105(.A1(new_n527), .A2(G52), .ZN(new_n531));
  AOI22_X1  g106(.A1(new_n505), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n532));
  INV_X1    g107(.A(G90), .ZN(new_n533));
  OAI22_X1  g108(.A1(new_n532), .A2(new_n507), .B1(new_n510), .B2(new_n533), .ZN(new_n534));
  NOR2_X1   g109(.A1(new_n531), .A2(new_n534), .ZN(G171));
  AOI22_X1  g110(.A1(new_n505), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n536));
  NOR2_X1   g111(.A1(new_n536), .A2(new_n507), .ZN(new_n537));
  XNOR2_X1  g112(.A(new_n537), .B(KEYINPUT75), .ZN(new_n538));
  INV_X1    g113(.A(new_n510), .ZN(new_n539));
  AOI22_X1  g114(.A1(new_n527), .A2(G43), .B1(G81), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g115(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g116(.A(new_n541), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(G860), .ZN(G153));
  AND3_X1   g118(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G36), .ZN(G176));
  NAND2_X1  g120(.A1(G1), .A2(G3), .ZN(new_n546));
  XNOR2_X1  g121(.A(new_n546), .B(KEYINPUT76), .ZN(new_n547));
  XNOR2_X1  g122(.A(new_n547), .B(KEYINPUT8), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n544), .A2(new_n548), .ZN(G188));
  AND3_X1   g124(.A1(new_n509), .A2(G53), .A3(G543), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT9), .ZN(new_n551));
  NAND2_X1  g126(.A1(G78), .A2(G543), .ZN(new_n552));
  NAND2_X1  g127(.A1(new_n502), .A2(new_n504), .ZN(new_n553));
  XNOR2_X1  g128(.A(KEYINPUT77), .B(G65), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n552), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G651), .ZN(new_n556));
  INV_X1    g131(.A(G91), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n556), .B1(new_n557), .B2(new_n510), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n551), .A2(new_n558), .ZN(new_n559));
  INV_X1    g134(.A(new_n559), .ZN(G299));
  INV_X1    g135(.A(G171), .ZN(G301));
  INV_X1    g136(.A(new_n512), .ZN(new_n562));
  AOI22_X1  g137(.A1(new_n539), .A2(G87), .B1(G49), .B2(new_n562), .ZN(new_n563));
  OAI21_X1  g138(.A(G651), .B1(new_n505), .B2(G74), .ZN(new_n564));
  INV_X1    g139(.A(KEYINPUT78), .ZN(new_n565));
  OR2_X1    g140(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND3_X1  g142(.A1(new_n563), .A2(new_n566), .A3(new_n567), .ZN(G288));
  NAND2_X1  g143(.A1(new_n539), .A2(G86), .ZN(new_n569));
  NAND2_X1  g144(.A1(G73), .A2(G543), .ZN(new_n570));
  INV_X1    g145(.A(G61), .ZN(new_n571));
  OAI21_X1  g146(.A(new_n570), .B1(new_n553), .B2(new_n571), .ZN(new_n572));
  NAND2_X1  g147(.A1(new_n572), .A2(G651), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n562), .A2(G48), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(G305));
  NAND2_X1  g150(.A1(new_n527), .A2(G47), .ZN(new_n576));
  AOI22_X1  g151(.A1(new_n505), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n577));
  NOR2_X1   g152(.A1(new_n577), .A2(new_n507), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n578), .B1(G85), .B2(new_n539), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n576), .A2(new_n579), .ZN(G290));
  NAND2_X1  g155(.A1(new_n527), .A2(G54), .ZN(new_n581));
  AND3_X1   g156(.A1(new_n505), .A2(G92), .A3(new_n509), .ZN(new_n582));
  XNOR2_X1  g157(.A(new_n582), .B(KEYINPUT10), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n505), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n584));
  OR2_X1    g159(.A1(new_n584), .A2(new_n507), .ZN(new_n585));
  NAND3_X1  g160(.A1(new_n581), .A2(new_n583), .A3(new_n585), .ZN(new_n586));
  INV_X1    g161(.A(G868), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n588), .B1(new_n587), .B2(G171), .ZN(G284));
  OAI21_X1  g164(.A(new_n588), .B1(new_n587), .B2(G171), .ZN(G321));
  NAND2_X1  g165(.A1(G299), .A2(new_n587), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n591), .B1(G168), .B2(new_n587), .ZN(G297));
  OAI21_X1  g167(.A(new_n591), .B1(G168), .B2(new_n587), .ZN(G280));
  INV_X1    g168(.A(new_n586), .ZN(new_n594));
  INV_X1    g169(.A(G559), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n595), .B2(G860), .ZN(G148));
  NAND2_X1  g171(.A1(new_n541), .A2(new_n587), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n586), .A2(G559), .ZN(new_n598));
  OAI21_X1  g173(.A(new_n597), .B1(new_n598), .B2(new_n587), .ZN(G323));
  XNOR2_X1  g174(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g175(.A1(new_n482), .A2(G123), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n468), .A2(KEYINPUT79), .A3(G135), .ZN(new_n602));
  OAI21_X1  g177(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n603));
  INV_X1    g178(.A(KEYINPUT80), .ZN(new_n604));
  OR2_X1    g179(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n603), .A2(new_n604), .ZN(new_n606));
  OAI211_X1 g181(.A(new_n605), .B(new_n606), .C1(G111), .C2(new_n466), .ZN(new_n607));
  INV_X1    g182(.A(KEYINPUT79), .ZN(new_n608));
  INV_X1    g183(.A(G135), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n467), .B2(new_n609), .ZN(new_n610));
  AND4_X1   g185(.A1(new_n601), .A2(new_n602), .A3(new_n607), .A4(new_n610), .ZN(new_n611));
  XNOR2_X1  g186(.A(new_n611), .B(KEYINPUT81), .ZN(new_n612));
  OR2_X1    g187(.A1(new_n612), .A2(G2096), .ZN(new_n613));
  NAND2_X1  g188(.A1(new_n493), .A2(new_n469), .ZN(new_n614));
  XNOR2_X1  g189(.A(new_n614), .B(KEYINPUT12), .ZN(new_n615));
  XNOR2_X1  g190(.A(KEYINPUT13), .B(G2100), .ZN(new_n616));
  XNOR2_X1  g191(.A(new_n615), .B(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n612), .A2(G2096), .ZN(new_n618));
  NAND3_X1  g193(.A1(new_n613), .A2(new_n617), .A3(new_n618), .ZN(new_n619));
  XOR2_X1   g194(.A(new_n619), .B(KEYINPUT82), .Z(G156));
  XNOR2_X1  g195(.A(G2427), .B(G2438), .ZN(new_n621));
  XNOR2_X1  g196(.A(new_n621), .B(G2430), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT15), .ZN(new_n623));
  XOR2_X1   g198(.A(new_n623), .B(G2435), .Z(new_n624));
  NAND2_X1  g199(.A1(new_n624), .A2(KEYINPUT14), .ZN(new_n625));
  XNOR2_X1  g200(.A(G2451), .B(G2454), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT84), .ZN(new_n627));
  XNOR2_X1  g202(.A(KEYINPUT83), .B(KEYINPUT16), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XNOR2_X1  g204(.A(G1341), .B(G1348), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT85), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2443), .B(G2446), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n631), .B(new_n632), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n629), .B(new_n633), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n625), .B(new_n634), .Z(new_n635));
  AND2_X1   g210(.A1(new_n635), .A2(G14), .ZN(G401));
  XOR2_X1   g211(.A(G2072), .B(G2078), .Z(new_n637));
  XOR2_X1   g212(.A(G2067), .B(G2678), .Z(new_n638));
  INV_X1    g213(.A(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G2084), .B(G2090), .Z(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  AOI21_X1  g216(.A(new_n637), .B1(new_n641), .B2(KEYINPUT18), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n642), .B(G2096), .ZN(new_n643));
  XNOR2_X1  g218(.A(new_n643), .B(G2100), .ZN(new_n644));
  AND2_X1   g219(.A1(new_n641), .A2(KEYINPUT17), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n639), .A2(new_n640), .ZN(new_n646));
  AOI21_X1  g221(.A(KEYINPUT18), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n644), .B(new_n647), .Z(G227));
  XNOR2_X1  g223(.A(G1971), .B(G1976), .ZN(new_n649));
  XNOR2_X1  g224(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n649), .B(new_n650), .Z(new_n651));
  XOR2_X1   g226(.A(G1956), .B(G2474), .Z(new_n652));
  XOR2_X1   g227(.A(G1961), .B(G1966), .Z(new_n653));
  AND2_X1   g228(.A1(new_n652), .A2(new_n653), .ZN(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n651), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n656), .B(new_n657), .ZN(new_n658));
  NOR2_X1   g233(.A1(new_n652), .A2(new_n653), .ZN(new_n659));
  INV_X1    g234(.A(new_n659), .ZN(new_n660));
  NAND3_X1  g235(.A1(new_n651), .A2(new_n655), .A3(new_n660), .ZN(new_n661));
  OAI211_X1 g236(.A(new_n658), .B(new_n661), .C1(new_n651), .C2(new_n660), .ZN(new_n662));
  XOR2_X1   g237(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n663));
  XOR2_X1   g238(.A(new_n662), .B(new_n663), .Z(new_n664));
  XNOR2_X1  g239(.A(G1991), .B(G1996), .ZN(new_n665));
  INV_X1    g240(.A(G1981), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(G1986), .ZN(new_n668));
  XOR2_X1   g243(.A(new_n664), .B(new_n668), .Z(G229));
  NOR2_X1   g244(.A1(G16), .A2(G23), .ZN(new_n670));
  INV_X1    g245(.A(G288), .ZN(new_n671));
  AOI21_X1  g246(.A(new_n670), .B1(new_n671), .B2(G16), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT33), .B(G1976), .Z(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(new_n675));
  XNOR2_X1  g250(.A(new_n672), .B(new_n675), .ZN(new_n676));
  NOR2_X1   g251(.A1(G16), .A2(G22), .ZN(new_n677));
  AOI21_X1  g252(.A(new_n677), .B1(G166), .B2(G16), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  MUX2_X1   g255(.A(G6), .B(G305), .S(G16), .Z(new_n681));
  XOR2_X1   g256(.A(KEYINPUT32), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(new_n683));
  NAND3_X1  g258(.A1(new_n676), .A2(new_n680), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT91), .B(KEYINPUT34), .ZN(new_n685));
  OR2_X1    g260(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  NOR2_X1   g261(.A1(G16), .A2(G24), .ZN(new_n687));
  INV_X1    g262(.A(G290), .ZN(new_n688));
  AOI21_X1  g263(.A(new_n687), .B1(new_n688), .B2(G16), .ZN(new_n689));
  INV_X1    g264(.A(G1986), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n689), .B(new_n690), .ZN(new_n691));
  NOR2_X1   g266(.A1(G25), .A2(G29), .ZN(new_n692));
  INV_X1    g267(.A(G107), .ZN(new_n693));
  AOI21_X1  g268(.A(new_n462), .B1(new_n693), .B2(G2105), .ZN(new_n694));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n695), .B1(G95), .B2(G2105), .ZN(new_n696));
  INV_X1    g271(.A(G95), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(new_n466), .A3(KEYINPUT88), .ZN(new_n698));
  NAND3_X1  g273(.A1(new_n694), .A2(new_n696), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT89), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n482), .A2(G119), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n468), .A2(G131), .ZN(new_n702));
  NAND3_X1  g277(.A1(new_n700), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  INV_X1    g278(.A(new_n703), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n692), .B1(new_n704), .B2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT90), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n706), .B(new_n707), .ZN(new_n708));
  NAND3_X1  g283(.A1(new_n686), .A2(new_n691), .A3(new_n708), .ZN(new_n709));
  INV_X1    g284(.A(KEYINPUT94), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND4_X1  g286(.A1(new_n686), .A2(KEYINPUT94), .A3(new_n691), .A4(new_n708), .ZN(new_n712));
  NAND2_X1  g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  INV_X1    g288(.A(KEYINPUT96), .ZN(new_n714));
  AOI22_X1  g289(.A1(new_n684), .A2(new_n685), .B1(new_n714), .B2(KEYINPUT36), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g291(.A1(new_n716), .A2(KEYINPUT97), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n714), .B1(KEYINPUT95), .B2(KEYINPUT36), .ZN(new_n718));
  INV_X1    g293(.A(KEYINPUT97), .ZN(new_n719));
  NAND3_X1  g294(.A1(new_n713), .A2(new_n719), .A3(new_n715), .ZN(new_n720));
  NAND3_X1  g295(.A1(new_n717), .A2(new_n718), .A3(new_n720), .ZN(new_n721));
  INV_X1    g296(.A(new_n718), .ZN(new_n722));
  AOI21_X1  g297(.A(new_n719), .B1(new_n713), .B2(new_n715), .ZN(new_n723));
  INV_X1    g298(.A(new_n715), .ZN(new_n724));
  AOI211_X1 g299(.A(KEYINPUT97), .B(new_n724), .C1(new_n711), .C2(new_n712), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n722), .B1(new_n723), .B2(new_n725), .ZN(new_n726));
  AOI22_X1  g301(.A1(G129), .A2(new_n482), .B1(new_n468), .B2(G141), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n469), .A2(G105), .ZN(new_n728));
  XNOR2_X1  g303(.A(KEYINPUT101), .B(KEYINPUT26), .ZN(new_n729));
  NAND3_X1  g304(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n729), .B(new_n730), .Z(new_n731));
  AND3_X1   g306(.A1(new_n727), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G29), .ZN(new_n733));
  INV_X1    g308(.A(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(G29), .ZN(new_n735));
  INV_X1    g310(.A(G32), .ZN(new_n736));
  AOI21_X1  g311(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  XNOR2_X1  g312(.A(KEYINPUT27), .B(G1996), .ZN(new_n738));
  XNOR2_X1  g313(.A(new_n738), .B(KEYINPUT102), .ZN(new_n739));
  NOR2_X1   g314(.A1(new_n737), .A2(new_n739), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n740), .B(KEYINPUT103), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n611), .A2(G29), .ZN(new_n742));
  INV_X1    g317(.A(KEYINPUT31), .ZN(new_n743));
  OAI21_X1  g318(.A(new_n742), .B1(new_n743), .B2(G11), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G35), .ZN(new_n745));
  AOI21_X1  g320(.A(new_n745), .B1(G162), .B2(G29), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n746), .B(KEYINPUT29), .ZN(new_n747));
  XNOR2_X1  g322(.A(new_n747), .B(G2090), .ZN(new_n748));
  AOI211_X1 g323(.A(new_n744), .B(new_n748), .C1(new_n743), .C2(G11), .ZN(new_n749));
  INV_X1    g324(.A(KEYINPUT99), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(G29), .B2(G33), .ZN(new_n751));
  OR3_X1    g326(.A1(new_n750), .A2(G29), .A3(G33), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n469), .A2(G103), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT25), .Z(new_n754));
  NAND2_X1  g329(.A1(new_n468), .A2(G139), .ZN(new_n755));
  AOI22_X1  g330(.A1(new_n493), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n756));
  OAI211_X1 g331(.A(new_n754), .B(new_n755), .C1(new_n466), .C2(new_n756), .ZN(new_n757));
  OAI211_X1 g332(.A(new_n751), .B(new_n752), .C1(new_n757), .C2(new_n735), .ZN(new_n758));
  INV_X1    g333(.A(G2072), .ZN(new_n759));
  OR2_X1    g334(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NOR2_X1   g335(.A1(G164), .A2(new_n735), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n761), .B1(G27), .B2(new_n735), .ZN(new_n762));
  INV_X1    g337(.A(G2078), .ZN(new_n763));
  OR2_X1    g338(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G16), .ZN(new_n765));
  NAND3_X1  g340(.A1(new_n765), .A2(KEYINPUT23), .A3(G20), .ZN(new_n766));
  INV_X1    g341(.A(KEYINPUT23), .ZN(new_n767));
  INV_X1    g342(.A(G20), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n767), .B1(new_n768), .B2(G16), .ZN(new_n769));
  OAI211_X1 g344(.A(new_n766), .B(new_n769), .C1(new_n559), .C2(new_n765), .ZN(new_n770));
  XOR2_X1   g345(.A(new_n770), .B(G1956), .Z(new_n771));
  NAND4_X1  g346(.A1(new_n749), .A2(new_n760), .A3(new_n764), .A4(new_n771), .ZN(new_n772));
  NOR2_X1   g347(.A1(G16), .A2(G21), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(G168), .B2(G16), .ZN(new_n774));
  INV_X1    g349(.A(new_n774), .ZN(new_n775));
  INV_X1    g350(.A(G1966), .ZN(new_n776));
  AOI22_X1  g351(.A1(new_n775), .A2(new_n776), .B1(new_n763), .B2(new_n762), .ZN(new_n777));
  NAND2_X1  g352(.A1(new_n758), .A2(new_n759), .ZN(new_n778));
  XNOR2_X1  g353(.A(KEYINPUT30), .B(G28), .ZN(new_n779));
  AOI22_X1  g354(.A1(new_n774), .A2(G1966), .B1(new_n735), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n765), .A2(G5), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G171), .B2(new_n765), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT104), .B(G1961), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n782), .B(new_n783), .ZN(new_n784));
  NAND4_X1  g359(.A1(new_n777), .A2(new_n778), .A3(new_n780), .A4(new_n784), .ZN(new_n785));
  INV_X1    g360(.A(KEYINPUT28), .ZN(new_n786));
  INV_X1    g361(.A(G26), .ZN(new_n787));
  OAI21_X1  g362(.A(new_n786), .B1(new_n787), .B2(G29), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n787), .A2(G29), .ZN(new_n789));
  NAND2_X1  g364(.A1(new_n482), .A2(G128), .ZN(new_n790));
  NAND2_X1  g365(.A1(new_n468), .A2(G140), .ZN(new_n791));
  OAI21_X1  g366(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n792));
  NOR2_X1   g367(.A1(new_n466), .A2(G116), .ZN(new_n793));
  OAI211_X1 g368(.A(new_n790), .B(new_n791), .C1(new_n792), .C2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G29), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n788), .B1(new_n795), .B2(new_n786), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n796), .A2(G2067), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n542), .A2(G16), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G16), .B2(G19), .ZN(new_n799));
  INV_X1    g374(.A(G1341), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n801), .B1(new_n800), .B2(new_n799), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n765), .A2(G4), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(new_n594), .B2(new_n765), .ZN(new_n804));
  XOR2_X1   g379(.A(new_n804), .B(G1348), .Z(new_n805));
  OAI211_X1 g380(.A(new_n802), .B(new_n805), .C1(G2067), .C2(new_n796), .ZN(new_n806));
  OR2_X1    g381(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n807));
  NAND2_X1  g382(.A1(new_n806), .A2(KEYINPUT98), .ZN(new_n808));
  AOI211_X1 g383(.A(new_n772), .B(new_n785), .C1(new_n807), .C2(new_n808), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n721), .A2(new_n726), .A3(new_n741), .A4(new_n809), .ZN(new_n810));
  INV_X1    g385(.A(new_n737), .ZN(new_n811));
  INV_X1    g386(.A(new_n739), .ZN(new_n812));
  NOR2_X1   g387(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(G34), .ZN(new_n814));
  AND2_X1   g389(.A1(new_n814), .A2(KEYINPUT24), .ZN(new_n815));
  NOR2_X1   g390(.A1(new_n814), .A2(KEYINPUT24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n735), .B1(new_n815), .B2(new_n816), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(G160), .B2(new_n735), .ZN(new_n818));
  XOR2_X1   g393(.A(KEYINPUT100), .B(G2084), .Z(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  INV_X1    g395(.A(new_n820), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n810), .A2(new_n813), .A3(new_n821), .ZN(G311));
  AND3_X1   g397(.A1(new_n721), .A2(new_n726), .A3(new_n809), .ZN(new_n823));
  INV_X1    g398(.A(new_n813), .ZN(new_n824));
  NAND4_X1  g399(.A1(new_n823), .A2(new_n824), .A3(new_n820), .A4(new_n741), .ZN(G150));
  AND2_X1   g400(.A1(new_n527), .A2(G55), .ZN(new_n826));
  AOI22_X1  g401(.A1(new_n505), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n827));
  XNOR2_X1  g402(.A(KEYINPUT105), .B(G93), .ZN(new_n828));
  OAI22_X1  g403(.A1(new_n827), .A2(new_n507), .B1(new_n510), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g404(.A1(new_n826), .A2(new_n829), .ZN(new_n830));
  INV_X1    g405(.A(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n831), .A2(G860), .ZN(new_n832));
  XOR2_X1   g407(.A(new_n832), .B(KEYINPUT37), .Z(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n542), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n830), .A2(new_n541), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n836), .B(KEYINPUT39), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n594), .A2(G559), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT38), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n837), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n833), .B1(new_n840), .B2(G860), .ZN(G145));
  NAND2_X1  g416(.A1(new_n487), .A2(new_n494), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n492), .A2(new_n498), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n843), .A2(KEYINPUT106), .ZN(new_n844));
  INV_X1    g419(.A(KEYINPUT106), .ZN(new_n845));
  NAND3_X1  g420(.A1(new_n492), .A2(new_n845), .A3(new_n498), .ZN(new_n846));
  AOI21_X1  g421(.A(new_n842), .B1(new_n844), .B2(new_n846), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n847), .B(new_n794), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n732), .B(new_n757), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n703), .B(new_n615), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n468), .A2(G142), .ZN(new_n852));
  OAI21_X1  g427(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n466), .A2(G118), .ZN(new_n854));
  OAI21_X1  g429(.A(new_n852), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AOI21_X1  g430(.A(new_n855), .B1(G130), .B2(new_n482), .ZN(new_n856));
  XOR2_X1   g431(.A(new_n851), .B(new_n856), .Z(new_n857));
  NOR2_X1   g432(.A1(new_n850), .A2(new_n857), .ZN(new_n858));
  OR2_X1    g433(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n859));
  NAND2_X1  g434(.A1(new_n858), .A2(KEYINPUT107), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g436(.A1(new_n861), .A2(KEYINPUT108), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n850), .A2(new_n857), .ZN(new_n863));
  INV_X1    g438(.A(KEYINPUT108), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n859), .A2(new_n864), .A3(new_n860), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n863), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(G162), .B(new_n476), .ZN(new_n867));
  XNOR2_X1  g442(.A(new_n867), .B(new_n611), .ZN(new_n868));
  AOI21_X1  g443(.A(G37), .B1(new_n866), .B2(new_n868), .ZN(new_n869));
  INV_X1    g444(.A(new_n868), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n861), .A2(new_n870), .A3(new_n863), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n869), .A2(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g448(.A1(new_n831), .A2(new_n587), .ZN(new_n874));
  XNOR2_X1  g449(.A(new_n836), .B(new_n598), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n594), .A2(new_n559), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n586), .A2(G299), .ZN(new_n877));
  NOR2_X1   g452(.A1(new_n876), .A2(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n875), .A2(new_n878), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(KEYINPUT41), .ZN(new_n880));
  INV_X1    g455(.A(KEYINPUT41), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n881), .B1(new_n876), .B2(new_n877), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n880), .A2(new_n882), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n879), .B1(new_n883), .B2(new_n875), .ZN(new_n884));
  XNOR2_X1  g459(.A(G290), .B(G288), .ZN(new_n885));
  XNOR2_X1  g460(.A(G303), .B(G305), .ZN(new_n886));
  OR2_X1    g461(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n886), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g464(.A1(new_n889), .A2(KEYINPUT42), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT109), .ZN(new_n891));
  INV_X1    g466(.A(new_n888), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n885), .A2(new_n886), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n891), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND3_X1  g469(.A1(new_n887), .A2(KEYINPUT109), .A3(new_n888), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  AOI21_X1  g471(.A(new_n890), .B1(new_n896), .B2(KEYINPUT42), .ZN(new_n897));
  XOR2_X1   g472(.A(new_n884), .B(new_n897), .Z(new_n898));
  OAI21_X1  g473(.A(new_n874), .B1(new_n898), .B2(new_n587), .ZN(G295));
  OAI21_X1  g474(.A(new_n874), .B1(new_n898), .B2(new_n587), .ZN(G331));
  INV_X1    g475(.A(KEYINPUT111), .ZN(new_n901));
  AND2_X1   g476(.A1(new_n894), .A2(new_n895), .ZN(new_n902));
  NAND2_X1  g477(.A1(G168), .A2(G301), .ZN(new_n903));
  NAND2_X1  g478(.A1(G286), .A2(G171), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n903), .A2(new_n834), .A3(new_n835), .A4(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n903), .A2(new_n904), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(new_n836), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n883), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  NAND3_X1  g483(.A1(new_n907), .A2(new_n878), .A3(new_n905), .ZN(new_n909));
  INV_X1    g484(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n902), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(G37), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n905), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(new_n882), .A3(new_n880), .ZN(new_n914));
  NAND3_X1  g489(.A1(new_n914), .A2(new_n896), .A3(new_n909), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n911), .A2(new_n912), .A3(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n901), .B1(new_n916), .B2(KEYINPUT43), .ZN(new_n917));
  NOR2_X1   g492(.A1(new_n916), .A2(KEYINPUT43), .ZN(new_n918));
  INV_X1    g493(.A(KEYINPUT110), .ZN(new_n919));
  AOI21_X1  g494(.A(new_n896), .B1(new_n914), .B2(new_n909), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n919), .B1(new_n920), .B2(G37), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n911), .A2(KEYINPUT110), .A3(new_n912), .ZN(new_n922));
  NAND3_X1  g497(.A1(new_n921), .A2(new_n922), .A3(new_n915), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n918), .B1(new_n923), .B2(KEYINPUT43), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n917), .B1(new_n924), .B2(new_n901), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  NAND2_X1  g501(.A1(new_n925), .A2(new_n926), .ZN(new_n927));
  INV_X1    g502(.A(KEYINPUT43), .ZN(new_n928));
  NOR2_X1   g503(.A1(new_n916), .A2(new_n928), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n929), .B1(new_n923), .B2(new_n928), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n927), .B1(new_n926), .B2(new_n930), .ZN(G397));
  INV_X1    g506(.A(new_n842), .ZN(new_n932));
  AND3_X1   g507(.A1(new_n492), .A2(new_n845), .A3(new_n498), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n845), .B1(new_n492), .B2(new_n498), .ZN(new_n934));
  OAI21_X1  g509(.A(new_n932), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  INV_X1    g510(.A(G1384), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT45), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n470), .A2(new_n475), .A3(G40), .ZN(new_n938));
  INV_X1    g513(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n937), .A2(new_n939), .ZN(new_n940));
  XNOR2_X1  g515(.A(new_n794), .B(G2067), .ZN(new_n941));
  XNOR2_X1  g516(.A(new_n941), .B(KEYINPUT112), .ZN(new_n942));
  XNOR2_X1  g517(.A(new_n732), .B(G1996), .ZN(new_n943));
  AND2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(new_n707), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n944), .A2(new_n945), .A3(new_n704), .ZN(new_n946));
  OR2_X1    g521(.A1(new_n794), .A2(G2067), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n940), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  AOI21_X1  g523(.A(new_n940), .B1(new_n942), .B2(new_n732), .ZN(new_n949));
  AOI21_X1  g524(.A(new_n949), .B1(KEYINPUT125), .B2(KEYINPUT46), .ZN(new_n950));
  NOR2_X1   g525(.A1(new_n940), .A2(G1996), .ZN(new_n951));
  NOR2_X1   g526(.A1(KEYINPUT125), .A2(KEYINPUT46), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AND2_X1   g528(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n950), .B1(new_n953), .B2(new_n954), .ZN(new_n955));
  XOR2_X1   g530(.A(new_n955), .B(KEYINPUT47), .Z(new_n956));
  OAI21_X1  g531(.A(new_n944), .B1(new_n707), .B2(new_n703), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n704), .A2(new_n945), .ZN(new_n958));
  OAI211_X1 g533(.A(new_n939), .B(new_n937), .C1(new_n957), .C2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n688), .A2(new_n690), .ZN(new_n960));
  NOR2_X1   g535(.A1(new_n960), .A2(new_n940), .ZN(new_n961));
  XOR2_X1   g536(.A(new_n961), .B(KEYINPUT48), .Z(new_n962));
  AOI211_X1 g537(.A(new_n948), .B(new_n956), .C1(new_n959), .C2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT114), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n935), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n499), .A2(new_n936), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  AOI21_X1  g542(.A(new_n938), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n965), .A2(new_n968), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(new_n679), .ZN(new_n970));
  INV_X1    g545(.A(new_n970), .ZN(new_n971));
  INV_X1    g546(.A(KEYINPUT50), .ZN(new_n972));
  NAND3_X1  g547(.A1(new_n935), .A2(new_n972), .A3(new_n936), .ZN(new_n973));
  AOI21_X1  g548(.A(new_n938), .B1(new_n966), .B2(KEYINPUT50), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  XNOR2_X1  g550(.A(KEYINPUT113), .B(G2090), .ZN(new_n976));
  NOR2_X1   g551(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n964), .B1(new_n971), .B2(new_n977), .ZN(new_n978));
  OAI211_X1 g553(.A(new_n970), .B(KEYINPUT114), .C1(new_n975), .C2(new_n976), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n978), .A2(G8), .A3(new_n979), .ZN(new_n980));
  NAND2_X1  g555(.A1(G303), .A2(G8), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n981), .B(KEYINPUT55), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n980), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n983), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n671), .A2(G1976), .ZN(new_n985));
  NAND3_X1  g560(.A1(new_n935), .A2(new_n939), .A3(new_n936), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n985), .A2(G8), .A3(new_n986), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT52), .ZN(new_n988));
  AND2_X1   g563(.A1(new_n986), .A2(G8), .ZN(new_n989));
  XNOR2_X1  g564(.A(KEYINPUT115), .B(G1976), .ZN(new_n990));
  AOI21_X1  g565(.A(KEYINPUT52), .B1(G288), .B2(new_n990), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n989), .A2(new_n985), .A3(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(G305), .A2(G1981), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n569), .A2(new_n666), .A3(new_n573), .A4(new_n574), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NOR2_X1   g570(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n996));
  INV_X1    g571(.A(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n995), .A2(new_n997), .ZN(new_n998));
  NAND3_X1  g573(.A1(new_n993), .A2(new_n994), .A3(new_n996), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(KEYINPUT116), .A2(KEYINPUT49), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n989), .A2(new_n1002), .ZN(new_n1003));
  OAI211_X1 g578(.A(new_n988), .B(new_n992), .C1(new_n1001), .C2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n1005));
  XNOR2_X1  g580(.A(new_n1004), .B(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT63), .ZN(new_n1007));
  AOI21_X1  g582(.A(new_n1007), .B1(new_n980), .B2(new_n982), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n984), .A2(new_n1006), .A3(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n975), .A2(G2084), .ZN(new_n1010));
  NOR2_X1   g585(.A1(new_n937), .A2(new_n938), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n499), .A2(KEYINPUT45), .A3(new_n936), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1011), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(new_n1010), .B1(new_n1013), .B2(new_n776), .ZN(new_n1014));
  INV_X1    g589(.A(G8), .ZN(new_n1015));
  NOR3_X1   g590(.A1(new_n1014), .A2(new_n1015), .A3(G286), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1016), .ZN(new_n1017));
  OAI21_X1  g592(.A(KEYINPUT63), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1006), .A2(new_n983), .ZN(new_n1019));
  INV_X1    g594(.A(G1976), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(new_n1001), .B2(new_n1003), .ZN(new_n1021));
  OAI21_X1  g596(.A(new_n994), .B1(new_n1021), .B2(G288), .ZN(new_n1022));
  NAND2_X1  g597(.A1(new_n1022), .A2(new_n989), .ZN(new_n1023));
  NAND3_X1  g598(.A1(new_n1018), .A2(new_n1019), .A3(new_n1023), .ZN(new_n1024));
  AOI21_X1  g599(.A(G1961), .B1(new_n973), .B2(new_n974), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n935), .A2(new_n936), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n967), .ZN(new_n1028));
  NAND4_X1  g603(.A1(new_n1028), .A2(new_n763), .A3(new_n939), .A4(new_n1012), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n1026), .B1(new_n1029), .B2(KEYINPUT123), .ZN(new_n1030));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1011), .A2(new_n1031), .A3(new_n763), .A4(new_n1012), .ZN(new_n1032));
  AOI21_X1  g607(.A(new_n1025), .B1(new_n1030), .B2(new_n1032), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1026), .B1(new_n969), .B2(G2078), .ZN(new_n1034));
  AOI21_X1  g609(.A(G301), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AND2_X1   g610(.A1(new_n1035), .A2(KEYINPUT62), .ZN(new_n1036));
  NAND2_X1  g611(.A1(G286), .A2(G8), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT122), .ZN(new_n1038));
  AOI21_X1  g613(.A(KEYINPUT51), .B1(new_n1037), .B2(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(new_n1014), .ZN(new_n1041));
  OAI211_X1 g616(.A(new_n1040), .B(G8), .C1(new_n1041), .C2(G286), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1037), .B(new_n1039), .C1(new_n1014), .C2(new_n1015), .ZN(new_n1043));
  OR3_X1    g618(.A1(new_n1014), .A2(KEYINPUT121), .A3(new_n1037), .ZN(new_n1044));
  OAI21_X1  g619(.A(KEYINPUT121), .B1(new_n1014), .B2(new_n1037), .ZN(new_n1045));
  AOI22_X1  g620(.A1(new_n1042), .A2(new_n1043), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  AOI22_X1  g621(.A1(new_n1009), .A2(new_n1016), .B1(new_n1036), .B2(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(KEYINPUT62), .B(G301), .C1(new_n1033), .C2(new_n1034), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n559), .A2(KEYINPUT57), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT57), .ZN(new_n1050));
  OAI21_X1  g625(.A(new_n1050), .B1(new_n551), .B2(new_n558), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1049), .A2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1052), .ZN(new_n1053));
  XNOR2_X1  g628(.A(KEYINPUT118), .B(G1956), .ZN(new_n1054));
  INV_X1    g629(.A(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(KEYINPUT50), .B1(new_n847), .B2(G1384), .ZN(new_n1056));
  NAND3_X1  g631(.A1(new_n499), .A2(new_n972), .A3(new_n936), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1057), .A2(new_n939), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1058), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n1055), .B1(new_n1056), .B2(new_n1059), .ZN(new_n1060));
  XNOR2_X1  g635(.A(KEYINPUT119), .B(KEYINPUT56), .ZN(new_n1061));
  XNOR2_X1  g636(.A(new_n1061), .B(G2072), .ZN(new_n1062));
  AND3_X1   g637(.A1(new_n965), .A2(new_n968), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1053), .B1(new_n1060), .B2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n972), .B1(new_n935), .B2(new_n936), .ZN(new_n1065));
  OAI21_X1  g640(.A(new_n1054), .B1(new_n1065), .B2(new_n1058), .ZN(new_n1066));
  NAND3_X1  g641(.A1(new_n965), .A2(new_n968), .A3(new_n1062), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1066), .A2(new_n1052), .A3(new_n1067), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n986), .A2(G2067), .ZN(new_n1069));
  AOI21_X1  g644(.A(G1348), .B1(new_n973), .B2(new_n974), .ZN(new_n1070));
  OAI211_X1 g645(.A(new_n1068), .B(new_n594), .C1(new_n1069), .C2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g646(.A1(new_n1070), .A2(new_n1069), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1072), .A2(KEYINPUT60), .A3(new_n586), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(KEYINPUT60), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1075), .B1(new_n1070), .B2(new_n1069), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1074), .A2(new_n594), .A3(new_n1076), .ZN(new_n1077));
  AND3_X1   g652(.A1(new_n1066), .A2(new_n1052), .A3(new_n1067), .ZN(new_n1078));
  AOI21_X1  g653(.A(new_n1052), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1079));
  NOR3_X1   g654(.A1(new_n1078), .A2(new_n1079), .A3(KEYINPUT61), .ZN(new_n1080));
  INV_X1    g655(.A(KEYINPUT61), .ZN(new_n1081));
  AOI21_X1  g656(.A(new_n1081), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1082));
  OAI211_X1 g657(.A(new_n1073), .B(new_n1077), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  INV_X1    g659(.A(G1996), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n965), .A2(new_n1085), .A3(new_n968), .ZN(new_n1086));
  XOR2_X1   g661(.A(KEYINPUT58), .B(G1341), .Z(new_n1087));
  NAND2_X1  g662(.A1(new_n986), .A2(new_n1087), .ZN(new_n1088));
  AOI21_X1  g663(.A(new_n541), .B1(new_n1086), .B2(new_n1088), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT120), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1084), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1091), .B1(new_n1090), .B2(new_n1089), .ZN(new_n1092));
  OR3_X1    g667(.A1(new_n1089), .A2(new_n1090), .A3(KEYINPUT59), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1092), .A2(new_n1093), .ZN(new_n1094));
  OAI211_X1 g669(.A(new_n1064), .B(new_n1071), .C1(new_n1083), .C2(new_n1094), .ZN(new_n1095));
  AND2_X1   g670(.A1(new_n1034), .A2(G301), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT124), .ZN(new_n1097));
  OR2_X1    g672(.A1(new_n1025), .A2(new_n1097), .ZN(new_n1098));
  NAND4_X1  g673(.A1(new_n1011), .A2(KEYINPUT53), .A3(new_n763), .A4(new_n965), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1025), .A2(new_n1097), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1098), .A2(new_n1099), .A3(new_n1034), .A4(new_n1100), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1033), .A2(new_n1096), .B1(new_n1101), .B2(G171), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT54), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1103), .B1(new_n1101), .B2(G171), .ZN(new_n1104));
  OAI22_X1  g679(.A1(new_n1102), .A2(new_n1103), .B1(new_n1035), .B2(new_n1104), .ZN(new_n1105));
  AOI21_X1  g680(.A(new_n1048), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1106));
  OAI21_X1  g681(.A(new_n1047), .B1(new_n1106), .B2(new_n1046), .ZN(new_n1107));
  NOR3_X1   g682(.A1(new_n1065), .A2(new_n1058), .A3(new_n976), .ZN(new_n1108));
  OAI21_X1  g683(.A(G8), .B1(new_n971), .B2(new_n1108), .ZN(new_n1109));
  AOI211_X1 g684(.A(new_n1004), .B(new_n983), .C1(new_n982), .C2(new_n1109), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1024), .B1(new_n1107), .B2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g686(.A(new_n958), .B(new_n957), .C1(G1986), .C2(G290), .ZN(new_n1112));
  AOI21_X1  g687(.A(new_n940), .B1(new_n1112), .B2(new_n960), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n963), .B1(new_n1111), .B2(new_n1113), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT126), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT126), .ZN(new_n1116));
  OAI211_X1 g691(.A(new_n963), .B(new_n1116), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1115), .A2(new_n1117), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g693(.A(G401), .B(G227), .C1(new_n869), .C2(new_n871), .ZN(new_n1120));
  INV_X1    g694(.A(G229), .ZN(new_n1121));
  AND4_X1   g695(.A1(G319), .A2(new_n925), .A3(new_n1120), .A4(new_n1121), .ZN(G308));
  NAND4_X1  g696(.A1(new_n925), .A2(new_n1120), .A3(G319), .A4(new_n1121), .ZN(G225));
endmodule


