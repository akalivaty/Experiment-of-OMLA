

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790;

  NAND2_X1 U382 ( .A1(n430), .A2(n427), .ZN(n380) );
  XOR2_X1 U383 ( .A(KEYINPUT98), .B(KEYINPUT99), .Z(n361) );
  XNOR2_X2 U384 ( .A(n384), .B(n383), .ZN(n581) );
  XNOR2_X2 U385 ( .A(n514), .B(n513), .ZN(n705) );
  AND2_X1 U386 ( .A1(n710), .A2(n619), .ZN(n448) );
  AND2_X1 U387 ( .A1(n455), .A2(n451), .ZN(n450) );
  AND2_X1 U388 ( .A1(n406), .A2(n636), .ZN(n455) );
  XNOR2_X1 U389 ( .A(n405), .B(KEYINPUT32), .ZN(n391) );
  NOR2_X1 U390 ( .A1(n720), .A2(n626), .ZN(n612) );
  XNOR2_X1 U391 ( .A(n449), .B(n372), .ZN(n720) );
  NAND2_X1 U392 ( .A1(n429), .A2(n428), .ZN(n427) );
  NAND2_X2 U393 ( .A1(n395), .A2(n392), .ZN(n708) );
  XNOR2_X1 U394 ( .A(KEYINPUT107), .B(n492), .ZN(n698) );
  AND2_X1 U395 ( .A1(n397), .A2(n396), .ZN(n395) );
  XNOR2_X1 U396 ( .A(n500), .B(n499), .ZN(n776) );
  XNOR2_X1 U397 ( .A(n423), .B(G101), .ZN(n521) );
  XNOR2_X1 U398 ( .A(n480), .B(G128), .ZN(n545) );
  XNOR2_X1 U399 ( .A(KEYINPUT4), .B(KEYINPUT17), .ZN(n544) );
  XNOR2_X1 U400 ( .A(G137), .B(KEYINPUT79), .ZN(n522) );
  INV_X1 U401 ( .A(G143), .ZN(n480) );
  INV_X1 U402 ( .A(G146), .ZN(n474) );
  NOR2_X2 U403 ( .A1(n743), .A2(n658), .ZN(n362) );
  XNOR2_X1 U404 ( .A(n419), .B(KEYINPUT35), .ZN(n363) );
  BUF_X1 U405 ( .A(n677), .Z(n364) );
  INV_X1 U406 ( .A(n634), .ZN(n365) );
  NOR2_X2 U407 ( .A1(n743), .A2(n658), .ZN(n756) );
  XNOR2_X1 U408 ( .A(n419), .B(KEYINPUT35), .ZN(n637) );
  AND2_X1 U409 ( .A1(n657), .A2(KEYINPUT2), .ZN(n435) );
  NOR2_X1 U410 ( .A1(n786), .A2(n593), .ZN(n594) );
  NOR2_X1 U411 ( .A1(G237), .A2(G902), .ZN(n537) );
  NAND2_X1 U412 ( .A1(n443), .A2(n589), .ZN(n442) );
  INV_X1 U413 ( .A(KEYINPUT6), .ZN(n398) );
  XNOR2_X1 U414 ( .A(n585), .B(n584), .ZN(n600) );
  INV_X1 U415 ( .A(KEYINPUT73), .ZN(n529) );
  XOR2_X1 U416 ( .A(KEYINPUT105), .B(KEYINPUT7), .Z(n482) );
  XNOR2_X1 U417 ( .A(G122), .B(KEYINPUT9), .ZN(n481) );
  XNOR2_X1 U418 ( .A(n420), .B(n421), .ZN(n434) );
  INV_X1 U419 ( .A(KEYINPUT48), .ZN(n421) );
  XNOR2_X1 U420 ( .A(KEYINPUT18), .B(KEYINPUT93), .ZN(n547) );
  XNOR2_X1 U421 ( .A(n766), .B(n389), .ZN(n550) );
  XNOR2_X1 U422 ( .A(n521), .B(KEYINPUT75), .ZN(n389) );
  NAND2_X1 U423 ( .A1(n448), .A2(n709), .ZN(n449) );
  XNOR2_X1 U424 ( .A(n557), .B(n556), .ZN(n603) );
  XNOR2_X1 U425 ( .A(n555), .B(KEYINPUT94), .ZN(n556) );
  NAND2_X1 U426 ( .A1(n536), .A2(n394), .ZN(n393) );
  INV_X1 U427 ( .A(G902), .ZN(n394) );
  XNOR2_X1 U428 ( .A(n775), .B(G146), .ZN(n533) );
  XNOR2_X1 U429 ( .A(n494), .B(G107), .ZN(n766) );
  XNOR2_X1 U430 ( .A(G104), .B(G110), .ZN(n494) );
  XNOR2_X1 U431 ( .A(KEYINPUT16), .B(G122), .ZN(n551) );
  XNOR2_X1 U432 ( .A(n478), .B(n477), .ZN(n672) );
  NOR2_X1 U433 ( .A1(n621), .A2(n366), .ZN(n441) );
  NOR2_X1 U434 ( .A1(n464), .A2(n698), .ZN(n586) );
  INV_X1 U435 ( .A(n619), .ZN(n464) );
  XNOR2_X1 U436 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n445) );
  XNOR2_X1 U437 ( .A(KEYINPUT102), .B(KEYINPUT101), .ZN(n446) );
  XNOR2_X1 U438 ( .A(n569), .B(KEYINPUT46), .ZN(n570) );
  INV_X1 U439 ( .A(KEYINPUT90), .ZN(n453) );
  XNOR2_X1 U440 ( .A(G119), .B(G116), .ZN(n528) );
  XNOR2_X1 U441 ( .A(n493), .B(n468), .ZN(n775) );
  XOR2_X1 U442 ( .A(G131), .B(KEYINPUT4), .Z(n468) );
  XNOR2_X1 U443 ( .A(G128), .B(G110), .ZN(n501) );
  NOR2_X1 U444 ( .A1(G953), .A2(G237), .ZN(n523) );
  XNOR2_X1 U445 ( .A(n447), .B(n444), .ZN(n472) );
  XNOR2_X1 U446 ( .A(n471), .B(KEYINPUT103), .ZN(n447) );
  XNOR2_X1 U447 ( .A(n446), .B(n445), .ZN(n444) );
  XNOR2_X1 U448 ( .A(G131), .B(G140), .ZN(n471) );
  XNOR2_X1 U449 ( .A(G143), .B(G113), .ZN(n469) );
  XOR2_X1 U450 ( .A(G122), .B(G104), .Z(n470) );
  INV_X1 U451 ( .A(KEYINPUT10), .ZN(n475) );
  NOR2_X1 U452 ( .A1(n605), .A2(KEYINPUT80), .ZN(n409) );
  XNOR2_X1 U453 ( .A(G902), .B(KEYINPUT15), .ZN(n647) );
  XOR2_X1 U454 ( .A(G137), .B(G140), .Z(n499) );
  XNOR2_X1 U455 ( .A(n495), .B(n403), .ZN(n402) );
  INV_X1 U456 ( .A(KEYINPUT95), .ZN(n403) );
  NAND2_X1 U457 ( .A1(G234), .A2(G237), .ZN(n516) );
  XNOR2_X1 U458 ( .A(n498), .B(KEYINPUT21), .ZN(n704) );
  INV_X1 U459 ( .A(G469), .ZN(n496) );
  INV_X1 U460 ( .A(KEYINPUT70), .ZN(n423) );
  XNOR2_X1 U461 ( .A(n545), .B(n457), .ZN(n493) );
  INV_X1 U462 ( .A(G134), .ZN(n457) );
  XNOR2_X1 U463 ( .A(G116), .B(G107), .ZN(n484) );
  XOR2_X1 U464 ( .A(KEYINPUT8), .B(KEYINPUT72), .Z(n489) );
  XNOR2_X1 U465 ( .A(n533), .B(n400), .ZN(n750) );
  XNOR2_X1 U466 ( .A(n550), .B(n401), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n456), .B(n402), .ZN(n401) );
  INV_X1 U468 ( .A(n499), .ZN(n456) );
  XNOR2_X1 U469 ( .A(n387), .B(n767), .ZN(n667) );
  INV_X1 U470 ( .A(n739), .ZN(n411) );
  BUF_X1 U471 ( .A(n603), .Z(n425) );
  INV_X1 U472 ( .A(KEYINPUT82), .ZN(n383) );
  NOR2_X2 U473 ( .A1(n603), .A2(n572), .ZN(n458) );
  NAND2_X1 U474 ( .A1(n399), .A2(G902), .ZN(n396) );
  XNOR2_X1 U475 ( .A(n437), .B(n436), .ZN(n580) );
  XNOR2_X1 U476 ( .A(n479), .B(G475), .ZN(n436) );
  OR2_X1 U477 ( .A1(n672), .A2(G902), .ZN(n437) );
  INV_X1 U478 ( .A(n708), .ZN(n629) );
  NOR2_X1 U479 ( .A1(n747), .A2(G953), .ZN(n462) );
  XNOR2_X1 U480 ( .A(n590), .B(KEYINPUT111), .ZN(n786) );
  NAND2_X1 U481 ( .A1(n439), .A2(n438), .ZN(n590) );
  AND2_X1 U482 ( .A1(n440), .A2(n441), .ZN(n439) );
  NAND2_X1 U483 ( .A1(n465), .A2(n463), .ZN(n405) );
  AND2_X1 U484 ( .A1(n620), .A2(n464), .ZN(n463) );
  XNOR2_X1 U485 ( .A(n460), .B(n459), .ZN(G75) );
  INV_X1 U486 ( .A(KEYINPUT53), .ZN(n459) );
  OR2_X1 U487 ( .A1(n748), .A2(n461), .ZN(n460) );
  NAND2_X1 U488 ( .A1(n749), .A2(n462), .ZN(n461) );
  AND2_X1 U489 ( .A1(n442), .A2(n371), .ZN(n366) );
  XNOR2_X1 U490 ( .A(n370), .B(n496), .ZN(n585) );
  AND2_X1 U491 ( .A1(n605), .A2(KEYINPUT80), .ZN(n367) );
  OR2_X1 U492 ( .A1(n442), .A2(n371), .ZN(n368) );
  INV_X1 U493 ( .A(n600), .ZN(n709) );
  OR2_X1 U494 ( .A1(G902), .A2(n757), .ZN(n369) );
  BUF_X1 U495 ( .A(n600), .Z(n621) );
  INV_X1 U496 ( .A(n536), .ZN(n399) );
  XNOR2_X1 U497 ( .A(n535), .B(n534), .ZN(n536) );
  NOR2_X1 U498 ( .A1(n750), .A2(G902), .ZN(n370) );
  INV_X1 U499 ( .A(n698), .ZN(n412) );
  XNOR2_X1 U500 ( .A(KEYINPUT36), .B(KEYINPUT92), .ZN(n371) );
  XOR2_X1 U501 ( .A(KEYINPUT76), .B(KEYINPUT33), .Z(n372) );
  OR2_X1 U502 ( .A1(KEYINPUT44), .A2(KEYINPUT91), .ZN(n373) );
  XOR2_X1 U503 ( .A(n660), .B(n659), .Z(n374) );
  XNOR2_X1 U504 ( .A(n364), .B(KEYINPUT123), .ZN(n375) );
  XNOR2_X1 U505 ( .A(n672), .B(KEYINPUT59), .ZN(n376) );
  XOR2_X1 U506 ( .A(n667), .B(n666), .Z(n377) );
  INV_X1 U507 ( .A(n701), .ZN(n413) );
  NAND2_X1 U508 ( .A1(KEYINPUT44), .A2(KEYINPUT91), .ZN(n378) );
  XNOR2_X1 U509 ( .A(n708), .B(n398), .ZN(n618) );
  XNOR2_X1 U510 ( .A(n424), .B(n533), .ZN(n660) );
  OR2_X1 U511 ( .A1(n660), .A2(n393), .ZN(n392) );
  BUF_X1 U512 ( .A(n743), .Z(n379) );
  NAND2_X1 U513 ( .A1(n390), .A2(n391), .ZN(n639) );
  NAND2_X1 U514 ( .A1(n430), .A2(n427), .ZN(n631) );
  XNOR2_X2 U515 ( .A(n381), .B(KEYINPUT81), .ZN(n743) );
  NAND2_X1 U516 ( .A1(n435), .A2(n433), .ZN(n381) );
  NAND2_X1 U517 ( .A1(n465), .A2(n464), .ZN(n633) );
  INV_X1 U518 ( .A(n623), .ZN(n465) );
  XNOR2_X2 U519 ( .A(n385), .B(KEYINPUT22), .ZN(n623) );
  NAND2_X1 U520 ( .A1(n382), .A2(n635), .ZN(n406) );
  XNOR2_X1 U521 ( .A(n633), .B(KEYINPUT89), .ZN(n382) );
  NAND2_X1 U522 ( .A1(n408), .A2(n407), .ZN(n645) );
  AND2_X2 U523 ( .A1(n541), .A2(n542), .ZN(n384) );
  NOR2_X1 U524 ( .A1(n434), .A2(KEYINPUT80), .ZN(n410) );
  NAND2_X1 U525 ( .A1(n631), .A2(n617), .ZN(n385) );
  XNOR2_X1 U526 ( .A(n386), .B(n549), .ZN(n388) );
  XNOR2_X1 U527 ( .A(n546), .B(n545), .ZN(n386) );
  XNOR2_X1 U528 ( .A(n388), .B(n550), .ZN(n387) );
  NAND2_X1 U529 ( .A1(n404), .A2(n634), .ZN(n390) );
  XNOR2_X1 U530 ( .A(n390), .B(G110), .ZN(G12) );
  XNOR2_X1 U531 ( .A(n391), .B(G119), .ZN(G21) );
  NAND2_X1 U532 ( .A1(n660), .A2(n399), .ZN(n397) );
  NAND2_X1 U533 ( .A1(n639), .A2(n373), .ZN(n451) );
  XNOR2_X1 U534 ( .A(n422), .B(KEYINPUT66), .ZN(n404) );
  XNOR2_X1 U535 ( .A(n406), .B(n683), .ZN(G3) );
  AND2_X2 U536 ( .A1(n434), .A2(n605), .ZN(n433) );
  NAND2_X1 U537 ( .A1(n434), .A2(n367), .ZN(n407) );
  NOR2_X1 U538 ( .A1(n410), .A2(n409), .ZN(n408) );
  NOR2_X1 U539 ( .A1(n433), .A2(n411), .ZN(n740) );
  XNOR2_X1 U540 ( .A(n433), .B(n779), .ZN(n778) );
  NAND2_X1 U541 ( .A1(n414), .A2(n412), .ZN(n559) );
  AND2_X1 U542 ( .A1(n414), .A2(n413), .ZN(n703) );
  XNOR2_X1 U543 ( .A(n558), .B(n415), .ZN(n414) );
  INV_X1 U544 ( .A(KEYINPUT39), .ZN(n415) );
  NAND2_X1 U545 ( .A1(n417), .A2(n416), .ZN(n624) );
  NAND2_X1 U546 ( .A1(n363), .A2(n378), .ZN(n416) );
  NAND2_X1 U547 ( .A1(n418), .A2(KEYINPUT91), .ZN(n417) );
  INV_X1 U548 ( .A(n637), .ZN(n418) );
  NAND2_X1 U549 ( .A1(n615), .A2(n614), .ZN(n419) );
  NAND2_X1 U550 ( .A1(n599), .A2(n598), .ZN(n420) );
  XNOR2_X1 U551 ( .A(n526), .B(n527), .ZN(n532) );
  XNOR2_X2 U552 ( .A(n458), .B(KEYINPUT19), .ZN(n610) );
  XNOR2_X2 U553 ( .A(n426), .B(n644), .ZN(n657) );
  NOR2_X2 U554 ( .A1(n623), .A2(n622), .ZN(n422) );
  XNOR2_X1 U555 ( .A(n532), .B(n552), .ZN(n424) );
  XNOR2_X2 U556 ( .A(n515), .B(KEYINPUT71), .ZN(n710) );
  XNOR2_X2 U557 ( .A(n559), .B(KEYINPUT40), .ZN(n790) );
  NAND2_X1 U558 ( .A1(n452), .A2(n450), .ZN(n454) );
  XNOR2_X1 U559 ( .A(n454), .B(n453), .ZN(n643) );
  XNOR2_X2 U560 ( .A(n474), .B(G125), .ZN(n548) );
  NAND2_X1 U561 ( .A1(n643), .A2(n642), .ZN(n426) );
  NOR2_X1 U562 ( .A1(n609), .A2(n611), .ZN(n428) );
  INV_X1 U563 ( .A(n610), .ZN(n429) );
  AND2_X2 U564 ( .A1(n432), .A2(n431), .ZN(n430) );
  NAND2_X1 U565 ( .A1(n609), .A2(n611), .ZN(n431) );
  NAND2_X1 U566 ( .A1(n610), .A2(n611), .ZN(n432) );
  OR2_X1 U567 ( .A1(n587), .A2(n368), .ZN(n438) );
  NAND2_X1 U568 ( .A1(n587), .A2(n371), .ZN(n440) );
  NOR2_X1 U569 ( .A1(n587), .A2(n588), .ZN(n601) );
  INV_X1 U570 ( .A(n588), .ZN(n443) );
  NAND2_X1 U571 ( .A1(n709), .A2(n710), .ZN(n625) );
  NAND2_X1 U572 ( .A1(n624), .A2(n373), .ZN(n452) );
  XOR2_X1 U573 ( .A(KEYINPUT77), .B(KEYINPUT34), .Z(n466) );
  XOR2_X1 U574 ( .A(KEYINPUT68), .B(KEYINPUT60), .Z(n467) );
  XNOR2_X1 U575 ( .A(n525), .B(n524), .ZN(n526) );
  INV_X1 U576 ( .A(KEYINPUT100), .ZN(n534) );
  XNOR2_X1 U577 ( .A(n506), .B(n505), .ZN(n507) );
  BUF_X1 U578 ( .A(n720), .Z(n745) );
  XNOR2_X1 U579 ( .A(n612), .B(n466), .ZN(n615) );
  XNOR2_X1 U580 ( .A(n508), .B(n507), .ZN(n677) );
  INV_X1 U581 ( .A(n760), .ZN(n674) );
  INV_X1 U582 ( .A(KEYINPUT124), .ZN(n680) );
  XNOR2_X1 U583 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n479) );
  XNOR2_X1 U584 ( .A(n470), .B(n469), .ZN(n473) );
  XOR2_X1 U585 ( .A(n473), .B(n472), .Z(n478) );
  NAND2_X1 U586 ( .A1(G214), .A2(n523), .ZN(n476) );
  XNOR2_X2 U587 ( .A(n548), .B(n475), .ZN(n500) );
  XOR2_X1 U588 ( .A(n476), .B(n500), .Z(n477) );
  INV_X1 U589 ( .A(n493), .ZN(n487) );
  XNOR2_X1 U590 ( .A(n482), .B(n481), .ZN(n483) );
  XOR2_X1 U591 ( .A(n483), .B(KEYINPUT106), .Z(n485) );
  XNOR2_X1 U592 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U593 ( .A(n487), .B(n486), .ZN(n491) );
  INV_X2 U594 ( .A(G953), .ZN(n769) );
  NAND2_X1 U595 ( .A1(G234), .A2(n769), .ZN(n488) );
  XNOR2_X1 U596 ( .A(n489), .B(n488), .ZN(n504) );
  NAND2_X1 U597 ( .A1(G217), .A2(n504), .ZN(n490) );
  XNOR2_X1 U598 ( .A(n491), .B(n490), .ZN(n757) );
  XNOR2_X1 U599 ( .A(G478), .B(n369), .ZN(n574) );
  NOR2_X1 U600 ( .A1(n580), .A2(n574), .ZN(n492) );
  NAND2_X1 U601 ( .A1(G227), .A2(n769), .ZN(n495) );
  NAND2_X1 U602 ( .A1(n647), .A2(G234), .ZN(n497) );
  XNOR2_X1 U603 ( .A(n497), .B(KEYINPUT20), .ZN(n509) );
  AND2_X1 U604 ( .A1(n509), .A2(G221), .ZN(n498) );
  XOR2_X1 U605 ( .A(KEYINPUT24), .B(KEYINPUT74), .Z(n502) );
  XNOR2_X1 U606 ( .A(n502), .B(n501), .ZN(n503) );
  XNOR2_X1 U607 ( .A(n776), .B(n503), .ZN(n508) );
  NAND2_X1 U608 ( .A1(n504), .A2(G221), .ZN(n506) );
  XNOR2_X1 U609 ( .A(G119), .B(KEYINPUT23), .ZN(n505) );
  NOR2_X1 U610 ( .A1(n677), .A2(G902), .ZN(n514) );
  XOR2_X1 U611 ( .A(KEYINPUT25), .B(KEYINPUT97), .Z(n511) );
  NAND2_X1 U612 ( .A1(n509), .A2(G217), .ZN(n510) );
  XNOR2_X1 U613 ( .A(n511), .B(n510), .ZN(n512) );
  XNOR2_X1 U614 ( .A(n512), .B(KEYINPUT96), .ZN(n513) );
  NAND2_X1 U615 ( .A1(n704), .A2(n705), .ZN(n515) );
  NAND2_X1 U616 ( .A1(n585), .A2(n710), .ZN(n628) );
  INV_X1 U617 ( .A(n628), .ZN(n542) );
  XNOR2_X1 U618 ( .A(KEYINPUT14), .B(n516), .ZN(n517) );
  NAND2_X1 U619 ( .A1(G952), .A2(n517), .ZN(n735) );
  NOR2_X1 U620 ( .A1(n735), .A2(G953), .ZN(n607) );
  AND2_X1 U621 ( .A1(G953), .A2(n517), .ZN(n518) );
  NAND2_X1 U622 ( .A1(G902), .A2(n518), .ZN(n606) );
  NOR2_X1 U623 ( .A1(G900), .A2(n606), .ZN(n519) );
  XNOR2_X1 U624 ( .A(n519), .B(KEYINPUT108), .ZN(n520) );
  NOR2_X1 U625 ( .A1(n607), .A2(n520), .ZN(n563) );
  XOR2_X1 U626 ( .A(n521), .B(KEYINPUT5), .Z(n527) );
  XNOR2_X1 U627 ( .A(n361), .B(n522), .ZN(n525) );
  NAND2_X1 U628 ( .A1(G210), .A2(n523), .ZN(n524) );
  XNOR2_X1 U629 ( .A(n528), .B(KEYINPUT3), .ZN(n531) );
  XNOR2_X1 U630 ( .A(n529), .B(G113), .ZN(n530) );
  XNOR2_X1 U631 ( .A(n531), .B(n530), .ZN(n552) );
  INV_X1 U632 ( .A(G472), .ZN(n535) );
  XNOR2_X1 U633 ( .A(n537), .B(KEYINPUT78), .ZN(n554) );
  INV_X1 U634 ( .A(G214), .ZN(n538) );
  OR2_X1 U635 ( .A1(n554), .A2(n538), .ZN(n721) );
  NAND2_X1 U636 ( .A1(n629), .A2(n721), .ZN(n539) );
  XNOR2_X1 U637 ( .A(n539), .B(KEYINPUT30), .ZN(n540) );
  NOR2_X1 U638 ( .A1(n563), .A2(n540), .ZN(n541) );
  NAND2_X1 U639 ( .A1(n769), .A2(G224), .ZN(n543) );
  XNOR2_X1 U640 ( .A(n543), .B(n544), .ZN(n546) );
  XNOR2_X1 U641 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U642 ( .A(n552), .B(n551), .ZN(n767) );
  NAND2_X1 U643 ( .A1(n667), .A2(n647), .ZN(n557) );
  INV_X1 U644 ( .A(G210), .ZN(n553) );
  OR2_X1 U645 ( .A1(n554), .A2(n553), .ZN(n555) );
  XOR2_X1 U646 ( .A(KEYINPUT38), .B(n425), .Z(n560) );
  NOR2_X1 U647 ( .A1(n581), .A2(n560), .ZN(n558) );
  INV_X1 U648 ( .A(n560), .ZN(n722) );
  NAND2_X1 U649 ( .A1(n722), .A2(n721), .ZN(n726) );
  INV_X1 U650 ( .A(n574), .ZN(n579) );
  AND2_X1 U651 ( .A1(n580), .A2(n579), .ZN(n616) );
  INV_X1 U652 ( .A(n616), .ZN(n724) );
  NOR2_X1 U653 ( .A1(n726), .A2(n724), .ZN(n562) );
  XNOR2_X1 U654 ( .A(KEYINPUT41), .B(KEYINPUT110), .ZN(n561) );
  XNOR2_X1 U655 ( .A(n562), .B(n561), .ZN(n746) );
  INV_X1 U656 ( .A(n585), .ZN(n567) );
  NOR2_X1 U657 ( .A1(n705), .A2(n563), .ZN(n564) );
  NAND2_X1 U658 ( .A1(n564), .A2(n704), .ZN(n588) );
  NOR2_X1 U659 ( .A1(n708), .A2(n588), .ZN(n565) );
  XOR2_X1 U660 ( .A(KEYINPUT28), .B(n565), .Z(n566) );
  OR2_X1 U661 ( .A1(n567), .A2(n566), .ZN(n573) );
  NOR2_X1 U662 ( .A1(n746), .A2(n573), .ZN(n568) );
  XOR2_X1 U663 ( .A(KEYINPUT42), .B(n568), .Z(n789) );
  NAND2_X1 U664 ( .A1(n790), .A2(n789), .ZN(n571) );
  XOR2_X1 U665 ( .A(KEYINPUT88), .B(KEYINPUT64), .Z(n569) );
  XNOR2_X1 U666 ( .A(n571), .B(n570), .ZN(n599) );
  INV_X1 U667 ( .A(n721), .ZN(n572) );
  NOR2_X1 U668 ( .A1(n573), .A2(n610), .ZN(n696) );
  NAND2_X1 U669 ( .A1(n696), .A2(KEYINPUT85), .ZN(n578) );
  NAND2_X1 U670 ( .A1(n580), .A2(n574), .ZN(n701) );
  NAND2_X1 U671 ( .A1(n701), .A2(n698), .ZN(n725) );
  OR2_X1 U672 ( .A1(n696), .A2(KEYINPUT85), .ZN(n575) );
  NAND2_X1 U673 ( .A1(n725), .A2(n575), .ZN(n576) );
  NAND2_X1 U674 ( .A1(KEYINPUT47), .A2(n576), .ZN(n577) );
  NAND2_X1 U675 ( .A1(n578), .A2(n577), .ZN(n597) );
  OR2_X1 U676 ( .A1(n580), .A2(n579), .ZN(n613) );
  NOR2_X1 U677 ( .A1(n581), .A2(n425), .ZN(n582) );
  XNOR2_X1 U678 ( .A(n582), .B(KEYINPUT109), .ZN(n583) );
  NOR2_X1 U679 ( .A1(n613), .A2(n583), .ZN(n695) );
  INV_X1 U680 ( .A(n695), .ZN(n595) );
  INV_X1 U681 ( .A(KEYINPUT1), .ZN(n584) );
  NAND2_X1 U682 ( .A1(n586), .A2(n721), .ZN(n587) );
  INV_X1 U683 ( .A(n425), .ZN(n589) );
  AND2_X1 U684 ( .A1(n696), .A2(n725), .ZN(n591) );
  NOR2_X1 U685 ( .A1(KEYINPUT85), .A2(n591), .ZN(n592) );
  NOR2_X1 U686 ( .A1(KEYINPUT47), .A2(n592), .ZN(n593) );
  NAND2_X1 U687 ( .A1(n595), .A2(n594), .ZN(n596) );
  NOR2_X1 U688 ( .A1(n597), .A2(n596), .ZN(n598) );
  NAND2_X1 U689 ( .A1(n621), .A2(n601), .ZN(n602) );
  XNOR2_X1 U690 ( .A(KEYINPUT43), .B(n602), .ZN(n604) );
  AND2_X1 U691 ( .A1(n604), .A2(n425), .ZN(n682) );
  NOR2_X1 U692 ( .A1(n703), .A2(n682), .ZN(n605) );
  NOR2_X1 U693 ( .A1(n606), .A2(G898), .ZN(n608) );
  NOR2_X1 U694 ( .A1(n608), .A2(n607), .ZN(n609) );
  XNOR2_X1 U695 ( .A(KEYINPUT69), .B(KEYINPUT0), .ZN(n611) );
  INV_X1 U696 ( .A(n380), .ZN(n626) );
  INV_X1 U697 ( .A(n613), .ZN(n614) );
  AND2_X1 U698 ( .A1(n616), .A2(n704), .ZN(n617) );
  INV_X1 U699 ( .A(n618), .ZN(n619) );
  NOR2_X1 U700 ( .A1(n621), .A2(n365), .ZN(n620) );
  NAND2_X1 U701 ( .A1(n621), .A2(n708), .ZN(n622) );
  INV_X1 U702 ( .A(n705), .ZN(n634) );
  OR2_X1 U703 ( .A1(n625), .A2(n708), .ZN(n715) );
  NOR2_X1 U704 ( .A1(n715), .A2(n626), .ZN(n627) );
  XNOR2_X1 U705 ( .A(n627), .B(KEYINPUT31), .ZN(n700) );
  NOR2_X1 U706 ( .A1(n629), .A2(n628), .ZN(n630) );
  NAND2_X1 U707 ( .A1(n380), .A2(n630), .ZN(n685) );
  NAND2_X1 U708 ( .A1(n700), .A2(n685), .ZN(n632) );
  NAND2_X1 U709 ( .A1(n632), .A2(n725), .ZN(n636) );
  NOR2_X1 U710 ( .A1(n709), .A2(n634), .ZN(n635) );
  BUF_X1 U711 ( .A(n363), .Z(n638) );
  NOR2_X1 U712 ( .A1(n638), .A2(KEYINPUT44), .ZN(n641) );
  INV_X1 U713 ( .A(n639), .ZN(n640) );
  NAND2_X1 U714 ( .A1(n641), .A2(n640), .ZN(n642) );
  XOR2_X1 U715 ( .A(KEYINPUT65), .B(KEYINPUT45), .Z(n644) );
  BUF_X2 U716 ( .A(n657), .Z(n761) );
  NAND2_X1 U717 ( .A1(n645), .A2(n761), .ZN(n651) );
  INV_X1 U718 ( .A(KEYINPUT67), .ZN(n646) );
  NAND2_X1 U719 ( .A1(n646), .A2(KEYINPUT2), .ZN(n649) );
  INV_X1 U720 ( .A(n647), .ZN(n653) );
  NAND2_X1 U721 ( .A1(n653), .A2(KEYINPUT2), .ZN(n648) );
  NAND2_X1 U722 ( .A1(n648), .A2(KEYINPUT67), .ZN(n652) );
  AND2_X1 U723 ( .A1(n649), .A2(n652), .ZN(n650) );
  NAND2_X1 U724 ( .A1(n651), .A2(n650), .ZN(n656) );
  INV_X1 U725 ( .A(n652), .ZN(n654) );
  OR2_X1 U726 ( .A1(n654), .A2(n653), .ZN(n655) );
  NAND2_X1 U727 ( .A1(n656), .A2(n655), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n756), .A2(G472), .ZN(n661) );
  XNOR2_X1 U729 ( .A(KEYINPUT112), .B(KEYINPUT62), .ZN(n659) );
  XNOR2_X1 U730 ( .A(n661), .B(n374), .ZN(n663) );
  INV_X1 U731 ( .A(G952), .ZN(n662) );
  AND2_X1 U732 ( .A1(n662), .A2(G953), .ZN(n760) );
  NAND2_X1 U733 ( .A1(n663), .A2(n674), .ZN(n664) );
  XNOR2_X1 U734 ( .A(n664), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U735 ( .A1(n756), .A2(G210), .ZN(n668) );
  XOR2_X1 U736 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n665) );
  XNOR2_X1 U737 ( .A(n665), .B(KEYINPUT83), .ZN(n666) );
  XNOR2_X1 U738 ( .A(n668), .B(n377), .ZN(n669) );
  NAND2_X1 U739 ( .A1(n669), .A2(n674), .ZN(n671) );
  INV_X1 U740 ( .A(KEYINPUT56), .ZN(n670) );
  XNOR2_X1 U741 ( .A(n671), .B(n670), .ZN(G51) );
  NAND2_X1 U742 ( .A1(n756), .A2(G475), .ZN(n673) );
  XNOR2_X1 U743 ( .A(n673), .B(n376), .ZN(n675) );
  NAND2_X1 U744 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U745 ( .A(n676), .B(n467), .ZN(G60) );
  NAND2_X1 U746 ( .A1(n362), .A2(G217), .ZN(n678) );
  XNOR2_X1 U747 ( .A(n678), .B(n375), .ZN(n679) );
  NAND2_X1 U748 ( .A1(n679), .A2(n674), .ZN(n681) );
  XNOR2_X1 U749 ( .A(n681), .B(n680), .ZN(G66) );
  XOR2_X1 U750 ( .A(n682), .B(G140), .Z(G42) );
  XOR2_X1 U751 ( .A(n638), .B(G122), .Z(G24) );
  XOR2_X1 U752 ( .A(G101), .B(KEYINPUT113), .Z(n683) );
  NOR2_X1 U753 ( .A1(n698), .A2(n685), .ZN(n684) );
  XOR2_X1 U754 ( .A(G104), .B(n684), .Z(G6) );
  NOR2_X1 U755 ( .A1(n701), .A2(n685), .ZN(n690) );
  XOR2_X1 U756 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n687) );
  XNOR2_X1 U757 ( .A(G107), .B(KEYINPUT26), .ZN(n686) );
  XNOR2_X1 U758 ( .A(n687), .B(n686), .ZN(n688) );
  XNOR2_X1 U759 ( .A(KEYINPUT114), .B(n688), .ZN(n689) );
  XNOR2_X1 U760 ( .A(n690), .B(n689), .ZN(G9) );
  AND2_X1 U761 ( .A1(n696), .A2(n413), .ZN(n694) );
  XOR2_X1 U762 ( .A(KEYINPUT116), .B(KEYINPUT29), .Z(n692) );
  XNOR2_X1 U763 ( .A(G128), .B(KEYINPUT117), .ZN(n691) );
  XNOR2_X1 U764 ( .A(n692), .B(n691), .ZN(n693) );
  XNOR2_X1 U765 ( .A(n694), .B(n693), .ZN(G30) );
  XOR2_X1 U766 ( .A(G143), .B(n695), .Z(G45) );
  NAND2_X1 U767 ( .A1(n696), .A2(n412), .ZN(n697) );
  XNOR2_X1 U768 ( .A(n697), .B(G146), .ZN(G48) );
  NOR2_X1 U769 ( .A1(n698), .A2(n700), .ZN(n699) );
  XOR2_X1 U770 ( .A(G113), .B(n699), .Z(G15) );
  NOR2_X1 U771 ( .A1(n701), .A2(n700), .ZN(n702) );
  XOR2_X1 U772 ( .A(G116), .B(n702), .Z(G18) );
  XOR2_X1 U773 ( .A(G134), .B(n703), .Z(G36) );
  NOR2_X1 U774 ( .A1(n365), .A2(n704), .ZN(n706) );
  XNOR2_X1 U775 ( .A(n706), .B(KEYINPUT49), .ZN(n707) );
  NAND2_X1 U776 ( .A1(n708), .A2(n707), .ZN(n713) );
  NOR2_X1 U777 ( .A1(n710), .A2(n709), .ZN(n711) );
  XNOR2_X1 U778 ( .A(n711), .B(KEYINPUT50), .ZN(n712) );
  NOR2_X1 U779 ( .A1(n713), .A2(n712), .ZN(n714) );
  XNOR2_X1 U780 ( .A(KEYINPUT119), .B(n714), .ZN(n716) );
  NAND2_X1 U781 ( .A1(n716), .A2(n715), .ZN(n717) );
  XNOR2_X1 U782 ( .A(n717), .B(KEYINPUT51), .ZN(n718) );
  XNOR2_X1 U783 ( .A(n718), .B(KEYINPUT120), .ZN(n719) );
  NOR2_X1 U784 ( .A1(n746), .A2(n719), .ZN(n732) );
  NOR2_X1 U785 ( .A1(n722), .A2(n721), .ZN(n723) );
  NOR2_X1 U786 ( .A1(n724), .A2(n723), .ZN(n729) );
  INV_X1 U787 ( .A(n725), .ZN(n727) );
  NOR2_X1 U788 ( .A1(n727), .A2(n726), .ZN(n728) );
  NOR2_X1 U789 ( .A1(n729), .A2(n728), .ZN(n730) );
  NOR2_X1 U790 ( .A1(n745), .A2(n730), .ZN(n731) );
  NOR2_X1 U791 ( .A1(n732), .A2(n731), .ZN(n733) );
  XNOR2_X1 U792 ( .A(n733), .B(KEYINPUT52), .ZN(n734) );
  NOR2_X1 U793 ( .A1(n735), .A2(n734), .ZN(n736) );
  XNOR2_X1 U794 ( .A(KEYINPUT121), .B(n736), .ZN(n749) );
  INV_X1 U795 ( .A(n761), .ZN(n737) );
  XOR2_X1 U796 ( .A(KEYINPUT2), .B(KEYINPUT84), .Z(n739) );
  NAND2_X1 U797 ( .A1(n737), .A2(n739), .ZN(n738) );
  XNOR2_X1 U798 ( .A(n738), .B(KEYINPUT86), .ZN(n742) );
  XNOR2_X1 U799 ( .A(n740), .B(KEYINPUT87), .ZN(n741) );
  NAND2_X1 U800 ( .A1(n742), .A2(n741), .ZN(n744) );
  NOR2_X1 U801 ( .A1(n744), .A2(n379), .ZN(n748) );
  NOR2_X1 U802 ( .A1(n746), .A2(n745), .ZN(n747) );
  XNOR2_X1 U803 ( .A(KEYINPUT58), .B(KEYINPUT122), .ZN(n752) );
  XNOR2_X1 U804 ( .A(n750), .B(KEYINPUT57), .ZN(n751) );
  XNOR2_X1 U805 ( .A(n752), .B(n751), .ZN(n754) );
  NAND2_X1 U806 ( .A1(n362), .A2(G469), .ZN(n753) );
  XOR2_X1 U807 ( .A(n754), .B(n753), .Z(n755) );
  NOR2_X1 U808 ( .A1(n760), .A2(n755), .ZN(G54) );
  NAND2_X1 U809 ( .A1(n362), .A2(G478), .ZN(n758) );
  XNOR2_X1 U810 ( .A(n758), .B(n757), .ZN(n759) );
  NOR2_X1 U811 ( .A1(n760), .A2(n759), .ZN(G63) );
  NAND2_X1 U812 ( .A1(n761), .A2(n769), .ZN(n765) );
  NAND2_X1 U813 ( .A1(G953), .A2(G224), .ZN(n762) );
  XNOR2_X1 U814 ( .A(KEYINPUT61), .B(n762), .ZN(n763) );
  NAND2_X1 U815 ( .A1(n763), .A2(G898), .ZN(n764) );
  NAND2_X1 U816 ( .A1(n765), .A2(n764), .ZN(n773) );
  XOR2_X1 U817 ( .A(n766), .B(G101), .Z(n768) );
  XOR2_X1 U818 ( .A(n768), .B(n767), .Z(n771) );
  NOR2_X1 U819 ( .A1(G898), .A2(n769), .ZN(n770) );
  NOR2_X1 U820 ( .A1(n771), .A2(n770), .ZN(n772) );
  XNOR2_X1 U821 ( .A(n773), .B(n772), .ZN(n774) );
  XOR2_X1 U822 ( .A(KEYINPUT125), .B(n774), .Z(G69) );
  XNOR2_X1 U823 ( .A(KEYINPUT95), .B(n775), .ZN(n777) );
  XNOR2_X1 U824 ( .A(n777), .B(n776), .ZN(n779) );
  NOR2_X1 U825 ( .A1(G953), .A2(n778), .ZN(n784) );
  XNOR2_X1 U826 ( .A(G227), .B(n779), .ZN(n780) );
  NAND2_X1 U827 ( .A1(n780), .A2(G900), .ZN(n781) );
  NAND2_X1 U828 ( .A1(n781), .A2(G953), .ZN(n782) );
  XOR2_X1 U829 ( .A(KEYINPUT126), .B(n782), .Z(n783) );
  NOR2_X1 U830 ( .A1(n784), .A2(n783), .ZN(n785) );
  XNOR2_X1 U831 ( .A(KEYINPUT127), .B(n785), .ZN(G72) );
  XNOR2_X1 U832 ( .A(n786), .B(KEYINPUT118), .ZN(n787) );
  XNOR2_X1 U833 ( .A(n787), .B(KEYINPUT37), .ZN(n788) );
  XNOR2_X1 U834 ( .A(G125), .B(n788), .ZN(G27) );
  XNOR2_X1 U835 ( .A(G137), .B(n789), .ZN(G39) );
  XNOR2_X1 U836 ( .A(n790), .B(G131), .ZN(G33) );
endmodule

