//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 1 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 0 1 1 1 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 1 0 1 1 1 1 0 0 1 1 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:57 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n671, new_n672,
    new_n673, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n756, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n782,
    new_n783, new_n784, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n865, new_n866, new_n867, new_n868, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n937, new_n938, new_n940, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n947, new_n948, new_n949,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n962, new_n963, new_n964,
    new_n965, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n982, new_n983, new_n984, new_n985, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996;
  XNOR2_X1  g000(.A(G8gat), .B(G36gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G64gat), .ZN(new_n203));
  INV_X1    g002(.A(G92gat), .ZN(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  INV_X1    g004(.A(G183gat), .ZN(new_n206));
  INV_X1    g005(.A(G190gat), .ZN(new_n207));
  NAND2_X1  g006(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NAND3_X1  g007(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  AOI21_X1  g009(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  INV_X1    g011(.A(G169gat), .ZN(new_n213));
  INV_X1    g012(.A(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(new_n213), .A2(new_n214), .A3(KEYINPUT23), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT23), .ZN(new_n216));
  OAI21_X1  g015(.A(new_n216), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT25), .ZN(new_n218));
  NAND2_X1  g017(.A1(G169gat), .A2(G176gat), .ZN(new_n219));
  NAND4_X1  g018(.A1(new_n215), .A2(new_n217), .A3(new_n218), .A4(new_n219), .ZN(new_n220));
  NOR2_X1   g019(.A1(new_n212), .A2(new_n220), .ZN(new_n221));
  INV_X1    g020(.A(KEYINPUT66), .ZN(new_n222));
  NAND2_X1  g021(.A1(new_n222), .A2(KEYINPUT28), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT28), .ZN(new_n224));
  AOI21_X1  g023(.A(G190gat), .B1(new_n224), .B2(KEYINPUT66), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n206), .A2(KEYINPUT27), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT27), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n227), .A2(G183gat), .ZN(new_n228));
  AND4_X1   g027(.A1(new_n223), .A2(new_n225), .A3(new_n226), .A4(new_n228), .ZN(new_n229));
  XNOR2_X1  g028(.A(KEYINPUT27), .B(G183gat), .ZN(new_n230));
  AOI21_X1  g029(.A(new_n223), .B1(new_n230), .B2(new_n225), .ZN(new_n231));
  NOR2_X1   g030(.A1(new_n229), .A2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(new_n219), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n213), .A2(new_n214), .ZN(new_n234));
  AOI21_X1  g033(.A(new_n233), .B1(KEYINPUT26), .B2(new_n234), .ZN(new_n235));
  OR3_X1    g034(.A1(KEYINPUT26), .A2(G169gat), .A3(G176gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n235), .A2(new_n236), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  AOI21_X1  g036(.A(new_n221), .B1(new_n232), .B2(new_n237), .ZN(new_n238));
  INV_X1    g037(.A(KEYINPUT64), .ZN(new_n239));
  NOR3_X1   g038(.A1(new_n216), .A2(G169gat), .A3(G176gat), .ZN(new_n240));
  OAI21_X1  g039(.A(new_n239), .B1(new_n240), .B2(new_n233), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n215), .A2(KEYINPUT64), .A3(new_n219), .ZN(new_n242));
  NAND3_X1  g041(.A1(new_n241), .A2(new_n242), .A3(new_n217), .ZN(new_n243));
  OAI211_X1 g042(.A(new_n208), .B(new_n209), .C1(new_n211), .C2(KEYINPUT65), .ZN(new_n244));
  AND2_X1   g043(.A1(new_n211), .A2(KEYINPUT65), .ZN(new_n245));
  NOR2_X1   g044(.A1(new_n244), .A2(new_n245), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n238), .A2(new_n247), .ZN(new_n248));
  INV_X1    g047(.A(G226gat), .ZN(new_n249));
  INV_X1    g048(.A(G233gat), .ZN(new_n250));
  NOR2_X1   g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n248), .A2(new_n251), .ZN(new_n252));
  AOI21_X1  g051(.A(KEYINPUT29), .B1(new_n238), .B2(new_n247), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n251), .B2(new_n253), .ZN(new_n254));
  XNOR2_X1  g053(.A(G197gat), .B(G204gat), .ZN(new_n255));
  INV_X1    g054(.A(KEYINPUT22), .ZN(new_n256));
  INV_X1    g055(.A(G211gat), .ZN(new_n257));
  INV_X1    g056(.A(G218gat), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n256), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n255), .A2(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(G211gat), .B(G218gat), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n260), .A2(new_n262), .ZN(new_n263));
  NAND3_X1  g062(.A1(new_n261), .A2(new_n255), .A3(new_n259), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  NAND2_X1  g065(.A1(new_n254), .A2(new_n266), .ZN(new_n267));
  INV_X1    g066(.A(new_n267), .ZN(new_n268));
  INV_X1    g067(.A(KEYINPUT29), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n248), .A2(new_n269), .ZN(new_n270));
  INV_X1    g069(.A(new_n251), .ZN(new_n271));
  AOI21_X1  g070(.A(KEYINPUT74), .B1(new_n270), .B2(new_n271), .ZN(new_n272));
  AOI21_X1  g071(.A(new_n272), .B1(KEYINPUT74), .B2(new_n254), .ZN(new_n273));
  AOI21_X1  g072(.A(new_n268), .B1(new_n273), .B2(new_n265), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT37), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n205), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(new_n273), .A2(new_n266), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n254), .B2(new_n265), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT38), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  AOI22_X1  g078(.A1(new_n276), .A2(new_n279), .B1(new_n274), .B2(new_n205), .ZN(new_n280));
  XNOR2_X1  g079(.A(G1gat), .B(G29gat), .ZN(new_n281));
  XNOR2_X1  g080(.A(new_n281), .B(KEYINPUT0), .ZN(new_n282));
  XNOR2_X1  g081(.A(new_n282), .B(G57gat), .ZN(new_n283));
  INV_X1    g082(.A(G85gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(new_n283), .B(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(G113gat), .ZN(new_n286));
  INV_X1    g085(.A(G120gat), .ZN(new_n287));
  AOI21_X1  g086(.A(KEYINPUT1), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n288), .B1(new_n286), .B2(new_n287), .ZN(new_n289));
  INV_X1    g088(.A(G127gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(new_n290), .A2(KEYINPUT67), .ZN(new_n291));
  INV_X1    g090(.A(KEYINPUT67), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(G127gat), .ZN(new_n293));
  NAND4_X1  g092(.A1(new_n291), .A2(new_n293), .A3(KEYINPUT68), .A4(G134gat), .ZN(new_n294));
  OR2_X1    g093(.A1(new_n290), .A2(G134gat), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n294), .A2(new_n295), .ZN(new_n296));
  XNOR2_X1  g095(.A(KEYINPUT67), .B(G127gat), .ZN(new_n297));
  AOI21_X1  g096(.A(KEYINPUT68), .B1(new_n297), .B2(G134gat), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n289), .B1(new_n296), .B2(new_n298), .ZN(new_n299));
  AND2_X1   g098(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n300));
  NOR2_X1   g099(.A1(KEYINPUT76), .A2(G155gat), .ZN(new_n301));
  OAI21_X1  g100(.A(G162gat), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(KEYINPUT2), .ZN(new_n303));
  INV_X1    g102(.A(G162gat), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n304), .A2(G155gat), .ZN(new_n305));
  INV_X1    g104(.A(G141gat), .ZN(new_n306));
  INV_X1    g105(.A(G148gat), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(G155gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(G162gat), .ZN(new_n310));
  NAND2_X1  g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311));
  AND4_X1   g110(.A1(new_n305), .A2(new_n308), .A3(new_n310), .A4(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n305), .A2(new_n310), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT2), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n314), .A3(new_n311), .ZN(new_n315));
  AOI22_X1  g114(.A1(new_n303), .A2(new_n312), .B1(new_n313), .B2(new_n315), .ZN(new_n316));
  XOR2_X1   g115(.A(G127gat), .B(G134gat), .Z(new_n317));
  NOR2_X1   g116(.A1(new_n289), .A2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n299), .A2(new_n316), .A3(new_n319), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT4), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND3_X1  g121(.A1(new_n291), .A2(new_n293), .A3(G134gat), .ZN(new_n323));
  INV_X1    g122(.A(KEYINPUT68), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n325), .A2(new_n294), .A3(new_n295), .ZN(new_n326));
  AOI21_X1  g125(.A(new_n318), .B1(new_n326), .B2(new_n289), .ZN(new_n327));
  NAND3_X1  g126(.A1(new_n327), .A2(KEYINPUT4), .A3(new_n316), .ZN(new_n328));
  AOI21_X1  g127(.A(KEYINPUT78), .B1(new_n322), .B2(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(new_n329), .ZN(new_n330));
  NAND3_X1  g129(.A1(new_n320), .A2(KEYINPUT78), .A3(KEYINPUT4), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT77), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n316), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n315), .A2(new_n313), .ZN(new_n334));
  XNOR2_X1  g133(.A(KEYINPUT76), .B(G155gat), .ZN(new_n335));
  AOI21_X1  g134(.A(new_n314), .B1(new_n335), .B2(G162gat), .ZN(new_n336));
  NAND4_X1  g135(.A1(new_n308), .A2(new_n305), .A3(new_n310), .A4(new_n311), .ZN(new_n337));
  OAI21_X1  g136(.A(new_n334), .B1(new_n336), .B2(new_n337), .ZN(new_n338));
  NAND2_X1  g137(.A1(new_n338), .A2(KEYINPUT77), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n333), .A2(new_n339), .A3(KEYINPUT3), .ZN(new_n340));
  INV_X1    g139(.A(KEYINPUT3), .ZN(new_n341));
  AOI22_X1  g140(.A1(new_n299), .A2(new_n319), .B1(new_n316), .B2(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n340), .A2(new_n342), .ZN(new_n343));
  NAND2_X1  g142(.A1(G225gat), .A2(G233gat), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(new_n345), .A2(KEYINPUT5), .ZN(new_n346));
  NAND4_X1  g145(.A1(new_n330), .A2(new_n331), .A3(new_n343), .A4(new_n346), .ZN(new_n347));
  INV_X1    g146(.A(KEYINPUT5), .ZN(new_n348));
  NAND2_X1  g147(.A1(new_n299), .A2(new_n319), .ZN(new_n349));
  NAND3_X1  g148(.A1(new_n349), .A2(new_n333), .A3(new_n339), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n350), .A2(new_n320), .ZN(new_n351));
  AOI21_X1  g150(.A(new_n348), .B1(new_n351), .B2(new_n345), .ZN(new_n352));
  NAND2_X1  g151(.A1(new_n320), .A2(new_n345), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n343), .A2(new_n328), .A3(new_n322), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n285), .B1(new_n347), .B2(new_n355), .ZN(new_n356));
  INV_X1    g155(.A(new_n356), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT6), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n343), .A2(new_n331), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n359), .A2(new_n329), .ZN(new_n360));
  AOI22_X1  g159(.A1(new_n360), .A2(new_n346), .B1(new_n352), .B2(new_n354), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n361), .A2(new_n285), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n357), .A2(new_n358), .A3(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(new_n205), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n254), .A2(KEYINPUT74), .ZN(new_n365));
  INV_X1    g164(.A(new_n272), .ZN(new_n366));
  NAND3_X1  g165(.A1(new_n365), .A2(new_n366), .A3(new_n265), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n267), .ZN(new_n368));
  OAI21_X1  g167(.A(new_n364), .B1(new_n368), .B2(KEYINPUT37), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n275), .B1(new_n367), .B2(new_n267), .ZN(new_n370));
  OAI21_X1  g169(.A(KEYINPUT38), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  NOR4_X1   g170(.A1(new_n361), .A2(KEYINPUT80), .A3(new_n358), .A4(new_n285), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT80), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n373), .B1(new_n356), .B2(KEYINPUT6), .ZN(new_n374));
  NOR2_X1   g173(.A1(new_n372), .A2(new_n374), .ZN(new_n375));
  NAND4_X1  g174(.A1(new_n280), .A2(new_n363), .A3(new_n371), .A4(new_n375), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT75), .ZN(new_n377));
  NAND4_X1  g176(.A1(new_n274), .A2(new_n377), .A3(KEYINPUT30), .A4(new_n205), .ZN(new_n378));
  NAND4_X1  g177(.A1(new_n367), .A2(KEYINPUT30), .A3(new_n267), .A4(new_n205), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n379), .A2(KEYINPUT75), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n367), .A2(new_n267), .A3(new_n205), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT30), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n364), .ZN(new_n384));
  NAND4_X1  g183(.A1(new_n378), .A2(new_n380), .A3(new_n383), .A4(new_n384), .ZN(new_n385));
  NAND3_X1  g184(.A1(new_n350), .A2(new_n320), .A3(new_n344), .ZN(new_n386));
  OAI211_X1 g185(.A(KEYINPUT39), .B(new_n386), .C1(new_n360), .C2(new_n344), .ZN(new_n387));
  INV_X1    g186(.A(KEYINPUT39), .ZN(new_n388));
  OAI211_X1 g187(.A(new_n388), .B(new_n345), .C1(new_n359), .C2(new_n329), .ZN(new_n389));
  NAND3_X1  g188(.A1(new_n387), .A2(new_n285), .A3(new_n389), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT40), .ZN(new_n391));
  OR2_X1    g190(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  AOI21_X1  g191(.A(new_n356), .B1(new_n390), .B2(new_n391), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n385), .A2(new_n392), .A3(new_n393), .ZN(new_n394));
  XNOR2_X1  g193(.A(G78gat), .B(G106gat), .ZN(new_n395));
  XNOR2_X1  g194(.A(new_n395), .B(G22gat), .ZN(new_n396));
  INV_X1    g195(.A(new_n396), .ZN(new_n397));
  XNOR2_X1  g196(.A(KEYINPUT31), .B(G50gat), .ZN(new_n398));
  XNOR2_X1  g197(.A(new_n398), .B(KEYINPUT83), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  INV_X1    g199(.A(G228gat), .ZN(new_n401));
  NOR2_X1   g200(.A1(new_n401), .A2(new_n250), .ZN(new_n402));
  INV_X1    g201(.A(new_n402), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n265), .A2(new_n269), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT81), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(KEYINPUT29), .B1(new_n263), .B2(new_n264), .ZN(new_n407));
  AOI21_X1  g206(.A(KEYINPUT3), .B1(new_n407), .B2(KEYINPUT81), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n316), .B1(new_n406), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n316), .A2(new_n341), .ZN(new_n410));
  AOI21_X1  g209(.A(new_n265), .B1(new_n410), .B2(new_n269), .ZN(new_n411));
  OAI21_X1  g210(.A(new_n403), .B1(new_n409), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g211(.A1(new_n412), .A2(KEYINPUT82), .ZN(new_n413));
  INV_X1    g212(.A(new_n264), .ZN(new_n414));
  AOI21_X1  g213(.A(new_n261), .B1(new_n259), .B2(new_n255), .ZN(new_n415));
  OAI211_X1 g214(.A(KEYINPUT81), .B(new_n269), .C1(new_n414), .C2(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n416), .A2(new_n341), .ZN(new_n417));
  NOR2_X1   g216(.A1(new_n407), .A2(KEYINPUT81), .ZN(new_n418));
  OAI21_X1  g217(.A(new_n338), .B1(new_n417), .B2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n411), .ZN(new_n420));
  NAND2_X1  g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT82), .ZN(new_n422));
  NAND3_X1  g221(.A1(new_n421), .A2(new_n422), .A3(new_n403), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n413), .A2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(new_n411), .A2(new_n403), .ZN(new_n425));
  OAI211_X1 g224(.A(new_n333), .B(new_n339), .C1(KEYINPUT3), .C2(new_n407), .ZN(new_n426));
  NAND2_X1  g225(.A1(new_n425), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n400), .B1(new_n424), .B2(new_n427), .ZN(new_n428));
  INV_X1    g227(.A(new_n427), .ZN(new_n429));
  AOI211_X1 g228(.A(new_n399), .B(new_n429), .C1(new_n413), .C2(new_n423), .ZN(new_n430));
  OAI21_X1  g229(.A(new_n397), .B1(new_n428), .B2(new_n430), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n422), .B1(new_n421), .B2(new_n403), .ZN(new_n432));
  AOI211_X1 g231(.A(KEYINPUT82), .B(new_n402), .C1(new_n419), .C2(new_n420), .ZN(new_n433));
  OAI21_X1  g232(.A(new_n427), .B1(new_n432), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n434), .A2(new_n399), .ZN(new_n435));
  NAND3_X1  g234(.A1(new_n424), .A2(new_n400), .A3(new_n427), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n435), .A2(new_n396), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n431), .A2(new_n437), .ZN(new_n438));
  INV_X1    g237(.A(new_n438), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n376), .A2(new_n394), .A3(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(KEYINPUT79), .ZN(new_n441));
  NAND4_X1  g240(.A1(new_n357), .A2(new_n362), .A3(new_n441), .A4(new_n358), .ZN(new_n442));
  OAI21_X1  g241(.A(new_n358), .B1(new_n361), .B2(new_n285), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n347), .A2(new_n355), .ZN(new_n444));
  INV_X1    g243(.A(new_n285), .ZN(new_n445));
  NOR2_X1   g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  OAI21_X1  g245(.A(KEYINPUT79), .B1(new_n443), .B2(new_n446), .ZN(new_n447));
  NAND3_X1  g246(.A1(new_n375), .A2(new_n442), .A3(new_n447), .ZN(new_n448));
  AND4_X1   g247(.A1(new_n378), .A2(new_n380), .A3(new_n383), .A4(new_n384), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n448), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n450), .A2(new_n438), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n440), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT32), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n453), .A2(KEYINPUT33), .ZN(new_n454));
  INV_X1    g253(.A(KEYINPUT70), .ZN(new_n455));
  NAND2_X1  g254(.A1(G227gat), .A2(G233gat), .ZN(new_n456));
  INV_X1    g255(.A(new_n456), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n238), .A2(new_n327), .A3(new_n247), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n327), .B1(new_n238), .B2(new_n247), .ZN(new_n459));
  OAI21_X1  g258(.A(new_n458), .B1(new_n459), .B2(KEYINPUT69), .ZN(new_n460));
  AND3_X1   g259(.A1(new_n241), .A2(new_n242), .A3(new_n217), .ZN(new_n461));
  INV_X1    g260(.A(new_n246), .ZN(new_n462));
  AOI21_X1  g261(.A(new_n218), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n226), .A2(new_n228), .ZN(new_n464));
  OAI211_X1 g263(.A(new_n222), .B(KEYINPUT28), .C1(new_n464), .C2(G190gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(G183gat), .A2(G190gat), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n234), .A2(KEYINPUT26), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n467), .A2(new_n236), .A3(new_n219), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n230), .A2(new_n223), .A3(new_n225), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n465), .A2(new_n466), .A3(new_n468), .A4(new_n469), .ZN(new_n470));
  OR2_X1    g269(.A1(new_n212), .A2(new_n220), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g271(.A(KEYINPUT69), .B(new_n349), .C1(new_n463), .C2(new_n472), .ZN(new_n473));
  INV_X1    g272(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g273(.A(new_n455), .B(new_n457), .C1(new_n460), .C2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n349), .B1(new_n463), .B2(new_n472), .ZN(new_n477));
  INV_X1    g276(.A(KEYINPUT69), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n477), .A2(new_n478), .ZN(new_n479));
  NAND3_X1  g278(.A1(new_n479), .A2(new_n473), .A3(new_n458), .ZN(new_n480));
  AOI21_X1  g279(.A(new_n455), .B1(new_n480), .B2(new_n457), .ZN(new_n481));
  OAI21_X1  g280(.A(new_n454), .B1(new_n476), .B2(new_n481), .ZN(new_n482));
  XOR2_X1   g281(.A(G71gat), .B(G99gat), .Z(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G43gat), .ZN(new_n484));
  XNOR2_X1  g283(.A(new_n483), .B(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(KEYINPUT71), .ZN(new_n487));
  OAI21_X1  g286(.A(new_n457), .B1(new_n460), .B2(new_n474), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(KEYINPUT70), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n475), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n453), .B1(new_n485), .B2(KEYINPUT33), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  AOI211_X1 g292(.A(KEYINPUT71), .B(new_n493), .C1(new_n489), .C2(new_n475), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n486), .B1(new_n492), .B2(new_n494), .ZN(new_n495));
  INV_X1    g294(.A(KEYINPUT72), .ZN(new_n496));
  OAI21_X1  g295(.A(new_n496), .B1(new_n480), .B2(new_n457), .ZN(new_n497));
  XNOR2_X1  g296(.A(new_n497), .B(KEYINPUT34), .ZN(new_n498));
  INV_X1    g297(.A(new_n498), .ZN(new_n499));
  NAND2_X1  g298(.A1(new_n495), .A2(new_n499), .ZN(new_n500));
  OAI211_X1 g299(.A(new_n498), .B(new_n486), .C1(new_n492), .C2(new_n494), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n500), .A2(KEYINPUT73), .A3(new_n501), .ZN(new_n502));
  INV_X1    g301(.A(KEYINPUT36), .ZN(new_n503));
  INV_X1    g302(.A(KEYINPUT73), .ZN(new_n504));
  NAND3_X1  g303(.A1(new_n495), .A2(new_n504), .A3(new_n499), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n502), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n500), .A2(KEYINPUT36), .A3(new_n501), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n452), .A2(new_n508), .ZN(new_n509));
  NAND3_X1  g308(.A1(new_n439), .A2(new_n500), .A3(new_n501), .ZN(new_n510));
  OAI21_X1  g309(.A(KEYINPUT35), .B1(new_n510), .B2(new_n450), .ZN(new_n511));
  INV_X1    g310(.A(KEYINPUT35), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n431), .A2(new_n437), .A3(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n375), .A2(new_n363), .ZN(new_n514));
  NAND3_X1  g313(.A1(new_n513), .A2(new_n449), .A3(new_n514), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n515), .B1(new_n505), .B2(new_n502), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT84), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n511), .B1(new_n516), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n502), .A2(new_n505), .ZN(new_n519));
  NOR2_X1   g318(.A1(new_n443), .A2(new_n446), .ZN(new_n520));
  NOR3_X1   g319(.A1(new_n520), .A2(new_n372), .A3(new_n374), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n431), .A2(new_n437), .A3(new_n512), .ZN(new_n522));
  NOR3_X1   g321(.A1(new_n521), .A2(new_n522), .A3(new_n385), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n517), .A3(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  OAI21_X1  g324(.A(new_n509), .B1(new_n518), .B2(new_n525), .ZN(new_n526));
  INV_X1    g325(.A(G29gat), .ZN(new_n527));
  INV_X1    g326(.A(G36gat), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n528), .A3(KEYINPUT14), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT14), .ZN(new_n530));
  OAI21_X1  g329(.A(new_n530), .B1(G29gat), .B2(G36gat), .ZN(new_n531));
  OAI211_X1 g330(.A(new_n529), .B(new_n531), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  INV_X1    g331(.A(G43gat), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n533), .A2(G50gat), .ZN(new_n534));
  INV_X1    g333(.A(G50gat), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(G43gat), .ZN(new_n536));
  AND3_X1   g335(.A1(new_n534), .A2(new_n536), .A3(KEYINPUT15), .ZN(new_n537));
  NAND2_X1  g336(.A1(new_n532), .A2(new_n537), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n538), .B(KEYINPUT85), .ZN(new_n539));
  XNOR2_X1  g338(.A(KEYINPUT86), .B(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n534), .B(KEYINPUT87), .ZN(new_n541));
  AOI21_X1  g340(.A(new_n540), .B1(new_n541), .B2(new_n536), .ZN(new_n542));
  OR2_X1    g341(.A1(new_n532), .A2(new_n537), .ZN(new_n543));
  OAI21_X1  g342(.A(new_n539), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  INV_X1    g343(.A(KEYINPUT17), .ZN(new_n545));
  OR2_X1    g344(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  XNOR2_X1  g345(.A(G15gat), .B(G22gat), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT16), .ZN(new_n548));
  OAI21_X1  g347(.A(new_n547), .B1(new_n548), .B2(G1gat), .ZN(new_n549));
  OAI21_X1  g348(.A(new_n549), .B1(G1gat), .B2(new_n547), .ZN(new_n550));
  INV_X1    g349(.A(G8gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n550), .B(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n544), .A2(new_n545), .ZN(new_n553));
  NAND3_X1  g352(.A1(new_n546), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  INV_X1    g353(.A(new_n552), .ZN(new_n555));
  AOI22_X1  g354(.A1(new_n554), .A2(KEYINPUT88), .B1(new_n555), .B2(new_n544), .ZN(new_n556));
  AND2_X1   g355(.A1(new_n546), .A2(new_n553), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT88), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n557), .A2(new_n558), .A3(new_n552), .ZN(new_n559));
  NAND2_X1  g358(.A1(G229gat), .A2(G233gat), .ZN(new_n560));
  NAND3_X1  g359(.A1(new_n556), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g360(.A(KEYINPUT18), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  NAND4_X1  g362(.A1(new_n556), .A2(new_n559), .A3(KEYINPUT18), .A4(new_n560), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n544), .B(new_n552), .ZN(new_n565));
  XOR2_X1   g364(.A(new_n560), .B(KEYINPUT13), .Z(new_n566));
  INV_X1    g365(.A(new_n566), .ZN(new_n567));
  NOR2_X1   g366(.A1(new_n565), .A2(new_n567), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n568), .B(KEYINPUT89), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n563), .A2(new_n564), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g369(.A(G113gat), .B(G141gat), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n571), .B(KEYINPUT11), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(new_n213), .ZN(new_n573));
  XNOR2_X1  g372(.A(new_n573), .B(G197gat), .ZN(new_n574));
  XNOR2_X1  g373(.A(new_n574), .B(KEYINPUT12), .ZN(new_n575));
  INV_X1    g374(.A(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n570), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT90), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n563), .A2(new_n575), .A3(new_n564), .A4(new_n569), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  NAND3_X1  g379(.A1(new_n570), .A2(KEYINPUT90), .A3(new_n576), .ZN(new_n581));
  AND2_X1   g380(.A1(new_n580), .A2(new_n581), .ZN(new_n582));
  INV_X1    g381(.A(new_n582), .ZN(new_n583));
  NAND2_X1  g382(.A1(G85gat), .A2(G92gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n584), .B(KEYINPUT7), .ZN(new_n585));
  NAND2_X1  g384(.A1(G99gat), .A2(G106gat), .ZN(new_n586));
  AOI22_X1  g385(.A1(KEYINPUT8), .A2(new_n586), .B1(new_n284), .B2(new_n204), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n585), .A2(new_n587), .ZN(new_n588));
  XOR2_X1   g387(.A(G99gat), .B(G106gat), .Z(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT93), .ZN(new_n591));
  NAND2_X1  g390(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  OR2_X1    g391(.A1(new_n588), .A2(new_n589), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n592), .B(new_n593), .ZN(new_n594));
  INV_X1    g393(.A(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(new_n544), .ZN(new_n596));
  NAND3_X1  g395(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  INV_X1    g397(.A(KEYINPUT94), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n557), .A2(new_n594), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT41), .ZN(new_n602));
  INV_X1    g401(.A(G232gat), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n602), .B1(new_n603), .B2(new_n250), .ZN(new_n604));
  NAND3_X1  g403(.A1(new_n600), .A2(new_n601), .A3(new_n604), .ZN(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n604), .B1(new_n600), .B2(new_n601), .ZN(new_n607));
  XNOR2_X1  g406(.A(G134gat), .B(G162gat), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n608), .B(KEYINPUT92), .ZN(new_n609));
  XNOR2_X1  g408(.A(G190gat), .B(G218gat), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n609), .B(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n606), .A2(new_n607), .A3(new_n612), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n612), .B1(new_n606), .B2(new_n607), .ZN(new_n614));
  NAND2_X1  g413(.A1(new_n613), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(G230gat), .A2(G233gat), .ZN(new_n616));
  XNOR2_X1  g415(.A(G57gat), .B(G64gat), .ZN(new_n617));
  AOI21_X1  g416(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n618));
  OR2_X1    g417(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  XNOR2_X1  g418(.A(G71gat), .B(G78gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n619), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n594), .A2(new_n622), .ZN(new_n623));
  INV_X1    g422(.A(KEYINPUT10), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n621), .A2(new_n593), .A3(new_n590), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT95), .ZN(new_n627));
  NAND3_X1  g426(.A1(new_n595), .A2(KEYINPUT10), .A3(new_n621), .ZN(new_n628));
  AND3_X1   g427(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n629));
  AOI21_X1  g428(.A(new_n627), .B1(new_n626), .B2(new_n628), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n616), .B1(new_n629), .B2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n623), .A2(new_n625), .ZN(new_n632));
  INV_X1    g431(.A(new_n616), .ZN(new_n633));
  NAND2_X1  g432(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G120gat), .B(G148gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(G176gat), .ZN(new_n636));
  INV_X1    g435(.A(G204gat), .ZN(new_n637));
  XNOR2_X1  g436(.A(new_n636), .B(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n631), .A2(new_n634), .A3(new_n638), .ZN(new_n639));
  INV_X1    g438(.A(new_n638), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n626), .A2(new_n628), .ZN(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  NOR2_X1   g441(.A1(new_n642), .A2(new_n633), .ZN(new_n643));
  INV_X1    g442(.A(new_n634), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n640), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n639), .A2(new_n645), .ZN(new_n646));
  NOR2_X1   g445(.A1(new_n621), .A2(KEYINPUT21), .ZN(new_n647));
  NAND2_X1  g446(.A1(G231gat), .A2(G233gat), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XOR2_X1   g448(.A(G127gat), .B(G155gat), .Z(new_n650));
  XOR2_X1   g449(.A(new_n650), .B(KEYINPUT20), .Z(new_n651));
  XNOR2_X1  g450(.A(new_n649), .B(new_n651), .ZN(new_n652));
  AOI21_X1  g451(.A(new_n555), .B1(KEYINPUT21), .B2(new_n621), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n206), .ZN(new_n654));
  XNOR2_X1  g453(.A(new_n652), .B(new_n654), .ZN(new_n655));
  XNOR2_X1  g454(.A(KEYINPUT91), .B(KEYINPUT19), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n656), .B(G211gat), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n655), .B(new_n657), .Z(new_n658));
  INV_X1    g457(.A(new_n658), .ZN(new_n659));
  NOR4_X1   g458(.A1(new_n583), .A2(new_n615), .A3(new_n646), .A4(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n526), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n661), .A2(new_n448), .ZN(new_n662));
  XOR2_X1   g461(.A(KEYINPUT96), .B(G1gat), .Z(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(G1324gat));
  NOR2_X1   g463(.A1(new_n661), .A2(new_n449), .ZN(new_n665));
  XOR2_X1   g464(.A(KEYINPUT16), .B(G8gat), .Z(new_n666));
  AND2_X1   g465(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  OR2_X1    g466(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n667), .A2(KEYINPUT42), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(new_n669), .C1(new_n551), .C2(new_n665), .ZN(G1325gat));
  OAI21_X1  g469(.A(G15gat), .B1(new_n661), .B2(new_n508), .ZN(new_n671));
  INV_X1    g470(.A(new_n519), .ZN(new_n672));
  OR2_X1    g471(.A1(new_n672), .A2(G15gat), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n671), .B1(new_n661), .B2(new_n673), .ZN(G1326gat));
  NOR2_X1   g473(.A1(new_n661), .A2(new_n439), .ZN(new_n675));
  XOR2_X1   g474(.A(KEYINPUT43), .B(G22gat), .Z(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  INV_X1    g476(.A(new_n615), .ZN(new_n678));
  NAND2_X1  g477(.A1(new_n501), .A2(KEYINPUT73), .ZN(new_n679));
  OAI21_X1  g478(.A(new_n491), .B1(new_n476), .B2(new_n481), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n680), .A2(KEYINPUT71), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n490), .A2(new_n487), .A3(new_n491), .ZN(new_n682));
  NAND2_X1  g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n498), .B1(new_n683), .B2(new_n486), .ZN(new_n684));
  NOR2_X1   g483(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  INV_X1    g484(.A(new_n505), .ZN(new_n686));
  OAI21_X1  g485(.A(new_n523), .B1(new_n685), .B2(new_n686), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n687), .A2(KEYINPUT84), .ZN(new_n688));
  NAND3_X1  g487(.A1(new_n688), .A2(new_n524), .A3(new_n511), .ZN(new_n689));
  AOI21_X1  g488(.A(new_n678), .B1(new_n689), .B2(new_n509), .ZN(new_n690));
  NOR3_X1   g489(.A1(new_n583), .A2(new_n658), .A3(new_n646), .ZN(new_n691));
  AND2_X1   g490(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  INV_X1    g491(.A(new_n448), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n692), .A2(new_n527), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n694), .B(KEYINPUT45), .ZN(new_n695));
  INV_X1    g494(.A(KEYINPUT44), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n690), .B(new_n696), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n697), .A2(new_n691), .ZN(new_n698));
  INV_X1    g497(.A(KEYINPUT97), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n697), .A2(KEYINPUT97), .A3(new_n691), .ZN(new_n701));
  AND3_X1   g500(.A1(new_n700), .A2(new_n693), .A3(new_n701), .ZN(new_n702));
  OAI21_X1  g501(.A(new_n695), .B1(new_n702), .B2(new_n527), .ZN(G1328gat));
  NAND3_X1  g502(.A1(new_n700), .A2(new_n385), .A3(new_n701), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n704), .A2(G36gat), .ZN(new_n705));
  AOI21_X1  g504(.A(G36gat), .B1(KEYINPUT98), .B2(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n692), .A2(new_n385), .A3(new_n706), .ZN(new_n707));
  NOR2_X1   g506(.A1(KEYINPUT98), .A2(KEYINPUT46), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n707), .B(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n705), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n710), .A2(KEYINPUT99), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT99), .ZN(new_n712));
  NAND3_X1  g511(.A1(new_n705), .A2(new_n712), .A3(new_n709), .ZN(new_n713));
  NAND2_X1  g512(.A1(new_n711), .A2(new_n713), .ZN(G1329gat));
  OAI21_X1  g513(.A(G43gat), .B1(new_n698), .B2(new_n508), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n672), .A2(G43gat), .ZN(new_n716));
  NAND2_X1  g515(.A1(new_n692), .A2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n715), .A2(KEYINPUT47), .A3(new_n717), .ZN(new_n718));
  NAND4_X1  g517(.A1(new_n700), .A2(new_n506), .A3(new_n507), .A4(new_n701), .ZN(new_n719));
  AOI22_X1  g518(.A1(new_n719), .A2(G43gat), .B1(new_n692), .B2(new_n716), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n718), .B1(new_n720), .B2(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g520(.A(G50gat), .B1(new_n698), .B2(new_n439), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n692), .A2(new_n535), .A3(new_n438), .ZN(new_n723));
  NAND3_X1  g522(.A1(new_n722), .A2(KEYINPUT48), .A3(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n723), .ZN(new_n725));
  NAND3_X1  g524(.A1(new_n700), .A2(new_n438), .A3(new_n701), .ZN(new_n726));
  AOI21_X1  g525(.A(new_n725), .B1(new_n726), .B2(G50gat), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n724), .B1(new_n727), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND3_X1  g527(.A1(new_n583), .A2(new_n678), .A3(new_n658), .ZN(new_n729));
  INV_X1    g528(.A(new_n646), .ZN(new_n730));
  NOR2_X1   g529(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n526), .ZN(new_n732));
  INV_X1    g531(.A(new_n732), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n733), .A2(new_n693), .ZN(new_n734));
  XNOR2_X1  g533(.A(new_n734), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g534(.A1(new_n732), .A2(new_n449), .ZN(new_n736));
  NOR2_X1   g535(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n737));
  AND2_X1   g536(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n738));
  OAI21_X1  g537(.A(new_n736), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  OAI21_X1  g538(.A(new_n739), .B1(new_n736), .B2(new_n737), .ZN(G1333gat));
  OAI21_X1  g539(.A(G71gat), .B1(new_n732), .B2(new_n508), .ZN(new_n741));
  OR2_X1    g540(.A1(new_n672), .A2(G71gat), .ZN(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n732), .B2(new_n742), .ZN(new_n743));
  XOR2_X1   g542(.A(new_n743), .B(KEYINPUT50), .Z(G1334gat));
  NAND2_X1  g543(.A1(new_n733), .A2(new_n438), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(G78gat), .ZN(G1335gat));
  INV_X1    g545(.A(KEYINPUT51), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n583), .A2(new_n659), .ZN(new_n748));
  INV_X1    g547(.A(new_n748), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT100), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n749), .B1(new_n690), .B2(new_n750), .ZN(new_n751));
  AOI211_X1 g550(.A(KEYINPUT100), .B(new_n678), .C1(new_n689), .C2(new_n509), .ZN(new_n752));
  OAI21_X1  g551(.A(new_n747), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n526), .A2(new_n615), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n754), .A2(KEYINPUT100), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n526), .A2(new_n750), .A3(new_n615), .ZN(new_n756));
  NAND4_X1  g555(.A1(new_n755), .A2(KEYINPUT51), .A3(new_n749), .A4(new_n756), .ZN(new_n757));
  AOI21_X1  g556(.A(new_n730), .B1(new_n753), .B2(new_n757), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n758), .A2(new_n284), .A3(new_n693), .ZN(new_n759));
  NOR2_X1   g558(.A1(new_n748), .A2(new_n730), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n697), .A2(new_n760), .ZN(new_n761));
  OAI21_X1  g560(.A(G85gat), .B1(new_n761), .B2(new_n448), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n759), .A2(new_n762), .ZN(G1336gat));
  INV_X1    g562(.A(KEYINPUT52), .ZN(new_n764));
  NOR2_X1   g563(.A1(new_n754), .A2(KEYINPUT44), .ZN(new_n765));
  NOR2_X1   g564(.A1(new_n690), .A2(new_n696), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n385), .B(new_n760), .C1(new_n765), .C2(new_n766), .ZN(new_n767));
  NAND2_X1  g566(.A1(new_n767), .A2(G92gat), .ZN(new_n768));
  NOR2_X1   g567(.A1(new_n449), .A2(G92gat), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n758), .A2(new_n769), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n770), .A2(KEYINPUT103), .ZN(new_n771));
  NOR2_X1   g570(.A1(new_n770), .A2(KEYINPUT103), .ZN(new_n772));
  OAI211_X1 g571(.A(new_n764), .B(new_n768), .C1(new_n771), .C2(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT101), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n768), .A2(new_n774), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n767), .A2(KEYINPUT101), .A3(G92gat), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n770), .A2(new_n775), .A3(new_n776), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT102), .ZN(new_n778));
  AND3_X1   g577(.A1(new_n777), .A2(new_n778), .A3(KEYINPUT52), .ZN(new_n779));
  AOI21_X1  g578(.A(new_n778), .B1(new_n777), .B2(KEYINPUT52), .ZN(new_n780));
  OAI21_X1  g579(.A(new_n773), .B1(new_n779), .B2(new_n780), .ZN(G1337gat));
  INV_X1    g580(.A(G99gat), .ZN(new_n782));
  NOR3_X1   g581(.A1(new_n761), .A2(new_n782), .A3(new_n508), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n758), .A2(new_n519), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n783), .B1(new_n784), .B2(new_n782), .ZN(G1338gat));
  NOR3_X1   g584(.A1(new_n730), .A2(new_n439), .A3(G106gat), .ZN(new_n786));
  INV_X1    g585(.A(new_n786), .ZN(new_n787));
  AOI21_X1  g586(.A(new_n787), .B1(new_n753), .B2(new_n757), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(KEYINPUT107), .ZN(new_n789));
  INV_X1    g588(.A(KEYINPUT53), .ZN(new_n790));
  OAI211_X1 g589(.A(new_n438), .B(new_n760), .C1(new_n765), .C2(new_n766), .ZN(new_n791));
  XOR2_X1   g590(.A(KEYINPUT104), .B(G106gat), .Z(new_n792));
  NAND2_X1  g591(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n789), .A2(new_n790), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(KEYINPUT106), .ZN(new_n795));
  AOI21_X1  g594(.A(new_n748), .B1(new_n754), .B2(KEYINPUT100), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT51), .B1(new_n796), .B2(new_n756), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n751), .A2(new_n747), .A3(new_n752), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n786), .B1(new_n797), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n799), .A2(KEYINPUT105), .ZN(new_n800));
  INV_X1    g599(.A(KEYINPUT105), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n788), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n800), .A2(new_n802), .A3(new_n793), .ZN(new_n803));
  AOI21_X1  g602(.A(new_n795), .B1(new_n803), .B2(KEYINPUT53), .ZN(new_n804));
  OAI21_X1  g603(.A(new_n793), .B1(new_n788), .B2(new_n801), .ZN(new_n805));
  AOI211_X1 g604(.A(KEYINPUT105), .B(new_n787), .C1(new_n753), .C2(new_n757), .ZN(new_n806));
  OAI211_X1 g605(.A(new_n795), .B(KEYINPUT53), .C1(new_n805), .C2(new_n806), .ZN(new_n807));
  INV_X1    g606(.A(new_n807), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n794), .B1(new_n804), .B2(new_n808), .ZN(G1339gat));
  NAND2_X1  g608(.A1(new_n641), .A2(KEYINPUT95), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n626), .A2(new_n627), .A3(new_n628), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n633), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  OAI21_X1  g611(.A(KEYINPUT54), .B1(new_n641), .B2(new_n616), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT108), .B1(new_n812), .B2(new_n813), .ZN(new_n814));
  INV_X1    g613(.A(new_n813), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT108), .ZN(new_n816));
  NAND3_X1  g615(.A1(new_n631), .A2(new_n815), .A3(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(KEYINPUT54), .ZN(new_n818));
  AOI21_X1  g617(.A(new_n638), .B1(new_n643), .B2(new_n818), .ZN(new_n819));
  NAND4_X1  g618(.A1(new_n814), .A2(KEYINPUT55), .A3(new_n817), .A4(new_n819), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT109), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n820), .A2(new_n821), .A3(new_n639), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n814), .A2(new_n817), .A3(new_n819), .ZN(new_n823));
  INV_X1    g622(.A(KEYINPUT55), .ZN(new_n824));
  NAND2_X1  g623(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  AND2_X1   g624(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n820), .A2(new_n639), .ZN(new_n827));
  NAND2_X1  g626(.A1(new_n827), .A2(KEYINPUT109), .ZN(new_n828));
  NAND3_X1  g627(.A1(new_n826), .A2(new_n582), .A3(new_n828), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n560), .B1(new_n556), .B2(new_n559), .ZN(new_n830));
  AND2_X1   g629(.A1(new_n565), .A2(new_n567), .ZN(new_n831));
  OAI21_X1  g630(.A(new_n574), .B1(new_n830), .B2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n579), .A2(new_n832), .ZN(new_n833));
  INV_X1    g632(.A(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n646), .ZN(new_n835));
  AOI21_X1  g634(.A(new_n615), .B1(new_n829), .B2(new_n835), .ZN(new_n836));
  NAND4_X1  g635(.A1(new_n828), .A2(new_n615), .A3(new_n825), .A4(new_n822), .ZN(new_n837));
  NOR2_X1   g636(.A1(new_n837), .A2(new_n833), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n659), .B1(new_n836), .B2(new_n838), .ZN(new_n839));
  NOR2_X1   g638(.A1(new_n729), .A2(new_n646), .ZN(new_n840));
  INV_X1    g639(.A(new_n840), .ZN(new_n841));
  AND2_X1   g640(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n842), .A2(new_n438), .ZN(new_n843));
  NOR2_X1   g642(.A1(new_n448), .A2(new_n385), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n843), .A2(new_n519), .A3(new_n844), .ZN(new_n845));
  OAI21_X1  g644(.A(G113gat), .B1(new_n845), .B2(new_n583), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT110), .ZN(new_n847));
  AND2_X1   g646(.A1(new_n846), .A2(new_n847), .ZN(new_n848));
  NOR2_X1   g647(.A1(new_n846), .A2(new_n847), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n839), .A2(new_n841), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(new_n693), .ZN(new_n851));
  OR3_X1    g650(.A1(new_n851), .A2(new_n385), .A3(new_n510), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n582), .A2(new_n286), .ZN(new_n853));
  OAI22_X1  g652(.A1(new_n848), .A2(new_n849), .B1(new_n852), .B2(new_n853), .ZN(G1340gat));
  OAI21_X1  g653(.A(G120gat), .B1(new_n845), .B2(new_n730), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT111), .ZN(new_n856));
  AND2_X1   g655(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n855), .A2(new_n856), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n646), .A2(new_n287), .ZN(new_n859));
  OAI22_X1  g658(.A1(new_n857), .A2(new_n858), .B1(new_n852), .B2(new_n859), .ZN(G1341gat));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n659), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n658), .A2(new_n297), .ZN(new_n862));
  OAI22_X1  g661(.A1(new_n861), .A2(new_n297), .B1(new_n852), .B2(new_n862), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT112), .ZN(G1342gat));
  OR3_X1    g663(.A1(new_n852), .A2(G134gat), .A3(new_n678), .ZN(new_n865));
  OR2_X1    g664(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n866));
  OAI21_X1  g665(.A(G134gat), .B1(new_n845), .B2(new_n678), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n865), .A2(KEYINPUT56), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n866), .A2(new_n867), .A3(new_n868), .ZN(G1343gat));
  INV_X1    g668(.A(KEYINPUT58), .ZN(new_n870));
  AOI21_X1  g669(.A(KEYINPUT57), .B1(new_n850), .B2(new_n438), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT57), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n439), .A2(new_n872), .ZN(new_n873));
  INV_X1    g672(.A(new_n873), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT113), .ZN(new_n875));
  AND2_X1   g674(.A1(new_n823), .A2(new_n875), .ZN(new_n876));
  NOR2_X1   g675(.A1(new_n823), .A2(new_n875), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(KEYINPUT55), .ZN(new_n878));
  NAND4_X1  g677(.A1(new_n580), .A2(new_n581), .A3(new_n639), .A4(new_n820), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n835), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g679(.A1(new_n880), .A2(new_n678), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n881), .B1(new_n833), .B2(new_n837), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n882), .A2(new_n659), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n874), .B1(new_n883), .B2(new_n841), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n508), .B(new_n844), .C1(new_n871), .C2(new_n884), .ZN(new_n885));
  OAI21_X1  g684(.A(G141gat), .B1(new_n885), .B2(new_n583), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n870), .B1(new_n886), .B2(KEYINPUT115), .ZN(new_n887));
  OR2_X1    g686(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n851), .A2(KEYINPUT114), .ZN(new_n889));
  NAND2_X1  g688(.A1(new_n508), .A2(new_n438), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n385), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n888), .A2(new_n889), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n582), .A2(new_n306), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n886), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n887), .A2(new_n894), .ZN(new_n895));
  OAI221_X1 g694(.A(new_n886), .B1(KEYINPUT115), .B2(new_n870), .C1(new_n892), .C2(new_n893), .ZN(new_n896));
  NAND2_X1  g695(.A1(new_n895), .A2(new_n896), .ZN(G1344gat));
  INV_X1    g696(.A(new_n892), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n307), .A3(new_n646), .ZN(new_n899));
  INV_X1    g698(.A(new_n885), .ZN(new_n900));
  AOI211_X1 g699(.A(KEYINPUT59), .B(new_n307), .C1(new_n900), .C2(new_n646), .ZN(new_n901));
  INV_X1    g700(.A(KEYINPUT59), .ZN(new_n902));
  NAND2_X1  g701(.A1(new_n508), .A2(new_n844), .ZN(new_n903));
  XOR2_X1   g702(.A(new_n903), .B(KEYINPUT116), .Z(new_n904));
  INV_X1    g703(.A(KEYINPUT117), .ZN(new_n905));
  AOI21_X1  g704(.A(new_n833), .B1(new_n837), .B2(new_n905), .ZN(new_n906));
  NAND4_X1  g705(.A1(new_n826), .A2(KEYINPUT117), .A3(new_n615), .A4(new_n828), .ZN(new_n907));
  AOI22_X1  g706(.A1(new_n906), .A2(new_n907), .B1(new_n880), .B2(new_n678), .ZN(new_n908));
  OAI21_X1  g707(.A(new_n841), .B1(new_n908), .B2(new_n658), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT57), .B1(new_n909), .B2(new_n438), .ZN(new_n910));
  OAI22_X1  g709(.A1(new_n910), .A2(KEYINPUT118), .B1(new_n842), .B2(new_n874), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n837), .A2(new_n905), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n912), .A2(new_n907), .A3(new_n834), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n658), .B1(new_n913), .B2(new_n881), .ZN(new_n914));
  OAI21_X1  g713(.A(new_n438), .B1(new_n914), .B2(new_n840), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n872), .ZN(new_n916));
  INV_X1    g715(.A(KEYINPUT118), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  OAI211_X1 g717(.A(new_n646), .B(new_n904), .C1(new_n911), .C2(new_n918), .ZN(new_n919));
  AOI21_X1  g718(.A(new_n902), .B1(new_n919), .B2(G148gat), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n899), .B1(new_n901), .B2(new_n920), .ZN(G1345gat));
  AOI21_X1  g720(.A(new_n335), .B1(new_n898), .B2(new_n658), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n658), .A2(new_n335), .ZN(new_n923));
  XOR2_X1   g722(.A(new_n923), .B(KEYINPUT119), .Z(new_n924));
  AOI21_X1  g723(.A(new_n922), .B1(new_n900), .B2(new_n924), .ZN(G1346gat));
  OAI21_X1  g724(.A(G162gat), .B1(new_n885), .B2(new_n678), .ZN(new_n926));
  NAND2_X1  g725(.A1(new_n615), .A2(new_n304), .ZN(new_n927));
  OAI21_X1  g726(.A(new_n926), .B1(new_n892), .B2(new_n927), .ZN(G1347gat));
  NOR2_X1   g727(.A1(new_n693), .A2(new_n449), .ZN(new_n929));
  NAND4_X1  g728(.A1(new_n850), .A2(new_n519), .A3(new_n439), .A4(new_n929), .ZN(new_n930));
  NOR3_X1   g729(.A1(new_n930), .A2(new_n213), .A3(new_n583), .ZN(new_n931));
  NOR2_X1   g730(.A1(new_n510), .A2(new_n449), .ZN(new_n932));
  XOR2_X1   g731(.A(new_n932), .B(KEYINPUT120), .Z(new_n933));
  NOR3_X1   g732(.A1(new_n842), .A2(new_n693), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n934), .A2(new_n582), .ZN(new_n935));
  AOI21_X1  g734(.A(new_n931), .B1(new_n213), .B2(new_n935), .ZN(G1348gat));
  NAND3_X1  g735(.A1(new_n934), .A2(new_n214), .A3(new_n646), .ZN(new_n937));
  OAI21_X1  g736(.A(G176gat), .B1(new_n930), .B2(new_n730), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(G1349gat));
  OAI21_X1  g738(.A(G183gat), .B1(new_n930), .B2(new_n659), .ZN(new_n940));
  INV_X1    g739(.A(KEYINPUT121), .ZN(new_n941));
  NOR2_X1   g740(.A1(new_n659), .A2(new_n464), .ZN(new_n942));
  AND3_X1   g741(.A1(new_n934), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  AOI21_X1  g742(.A(new_n941), .B1(new_n934), .B2(new_n942), .ZN(new_n944));
  OAI21_X1  g743(.A(new_n940), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  XNOR2_X1  g744(.A(new_n945), .B(KEYINPUT60), .ZN(G1350gat));
  OAI21_X1  g745(.A(G190gat), .B1(new_n930), .B2(new_n678), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT122), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g748(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n950));
  NAND3_X1  g749(.A1(new_n934), .A2(new_n207), .A3(new_n615), .ZN(new_n951));
  NOR2_X1   g750(.A1(new_n947), .A2(new_n948), .ZN(new_n952));
  NAND2_X1  g751(.A1(new_n949), .A2(KEYINPUT61), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n950), .B(new_n951), .C1(new_n952), .C2(new_n953), .ZN(G1351gat));
  INV_X1    g753(.A(G197gat), .ZN(new_n955));
  NAND2_X1  g754(.A1(new_n508), .A2(new_n929), .ZN(new_n956));
  AOI21_X1  g755(.A(new_n874), .B1(new_n839), .B2(new_n841), .ZN(new_n957));
  AOI21_X1  g756(.A(new_n957), .B1(new_n916), .B2(new_n917), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n910), .A2(KEYINPUT118), .ZN(new_n959));
  AOI21_X1  g758(.A(new_n956), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  AOI21_X1  g759(.A(new_n955), .B1(new_n960), .B2(new_n582), .ZN(new_n961));
  NOR2_X1   g760(.A1(new_n890), .A2(new_n449), .ZN(new_n962));
  AND3_X1   g761(.A1(new_n850), .A2(new_n448), .A3(new_n962), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n963), .A2(new_n955), .A3(new_n582), .ZN(new_n964));
  XNOR2_X1  g763(.A(new_n964), .B(KEYINPUT123), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT124), .B1(new_n961), .B2(new_n965), .ZN(new_n966));
  INV_X1    g765(.A(new_n956), .ZN(new_n967));
  OAI21_X1  g766(.A(new_n967), .B1(new_n911), .B2(new_n918), .ZN(new_n968));
  OAI21_X1  g767(.A(G197gat), .B1(new_n968), .B2(new_n583), .ZN(new_n969));
  INV_X1    g768(.A(KEYINPUT124), .ZN(new_n970));
  INV_X1    g769(.A(KEYINPUT123), .ZN(new_n971));
  XNOR2_X1  g770(.A(new_n964), .B(new_n971), .ZN(new_n972));
  NAND3_X1  g771(.A1(new_n969), .A2(new_n970), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g772(.A1(new_n966), .A2(new_n973), .ZN(G1352gat));
  INV_X1    g773(.A(KEYINPUT125), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n968), .B2(new_n730), .ZN(new_n976));
  NAND3_X1  g775(.A1(new_n960), .A2(KEYINPUT125), .A3(new_n646), .ZN(new_n977));
  NAND3_X1  g776(.A1(new_n976), .A2(G204gat), .A3(new_n977), .ZN(new_n978));
  NAND3_X1  g777(.A1(new_n963), .A2(new_n637), .A3(new_n646), .ZN(new_n979));
  XOR2_X1   g778(.A(new_n979), .B(KEYINPUT62), .Z(new_n980));
  NAND2_X1  g779(.A1(new_n978), .A2(new_n980), .ZN(G1353gat));
  NAND3_X1  g780(.A1(new_n963), .A2(new_n257), .A3(new_n658), .ZN(new_n982));
  OAI211_X1 g781(.A(new_n658), .B(new_n967), .C1(new_n911), .C2(new_n918), .ZN(new_n983));
  AND3_X1   g782(.A1(new_n983), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n984));
  AOI21_X1  g783(.A(KEYINPUT63), .B1(new_n983), .B2(G211gat), .ZN(new_n985));
  OAI21_X1  g784(.A(new_n982), .B1(new_n984), .B2(new_n985), .ZN(G1354gat));
  NOR2_X1   g785(.A1(new_n678), .A2(new_n258), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n960), .A2(new_n987), .ZN(new_n988));
  NAND3_X1  g787(.A1(new_n850), .A2(new_n448), .A3(new_n962), .ZN(new_n989));
  OAI21_X1  g788(.A(new_n258), .B1(new_n989), .B2(new_n678), .ZN(new_n990));
  INV_X1    g789(.A(KEYINPUT126), .ZN(new_n991));
  XNOR2_X1  g790(.A(new_n990), .B(new_n991), .ZN(new_n992));
  NAND2_X1  g791(.A1(new_n988), .A2(new_n992), .ZN(new_n993));
  NAND2_X1  g792(.A1(new_n993), .A2(KEYINPUT127), .ZN(new_n994));
  INV_X1    g793(.A(KEYINPUT127), .ZN(new_n995));
  NAND3_X1  g794(.A1(new_n988), .A2(new_n992), .A3(new_n995), .ZN(new_n996));
  NAND2_X1  g795(.A1(new_n994), .A2(new_n996), .ZN(G1355gat));
endmodule


