//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 1 1 0 1 1 1 1 0 1 1 0 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 1 1 1 0 1 0 1 0 1 0 1 1 0 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:36 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n688, new_n689, new_n690,
    new_n691, new_n692, new_n693, new_n694, new_n695, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1085, new_n1086, new_n1087, new_n1088,
    new_n1089, new_n1090, new_n1091, new_n1092, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1240, new_n1241,
    new_n1242, new_n1243, new_n1244, new_n1245, new_n1246, new_n1247,
    new_n1248, new_n1249, new_n1250, new_n1251, new_n1252, new_n1253,
    new_n1254, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1268, new_n1269, new_n1270, new_n1271, new_n1273,
    new_n1274, new_n1275, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1359,
    new_n1360, new_n1361;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(KEYINPUT64), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT64), .ZN(new_n216));
  NAND3_X1  g0016(.A1(new_n216), .A2(G1), .A3(G13), .ZN(new_n217));
  NAND2_X1  g0017(.A1(new_n215), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g0018(.A1(new_n213), .A2(G20), .A3(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT65), .Z(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n222));
  AOI22_X1  g0022(.A1(G68), .A2(G238), .B1(G87), .B2(G250), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G97), .A2(G257), .B1(G107), .B2(G264), .ZN(new_n224));
  NAND3_X1  g0024(.A1(new_n222), .A2(new_n223), .A3(new_n224), .ZN(new_n225));
  OAI21_X1  g0025(.A(new_n208), .B1(new_n221), .B2(new_n225), .ZN(new_n226));
  OAI211_X1 g0026(.A(new_n211), .B(new_n219), .C1(KEYINPUT1), .C2(new_n226), .ZN(new_n227));
  AOI21_X1  g0027(.A(new_n227), .B1(KEYINPUT1), .B2(new_n226), .ZN(G361));
  XOR2_X1   g0028(.A(G238), .B(G244), .Z(new_n229));
  XNOR2_X1  g0029(.A(new_n229), .B(G232), .ZN(new_n230));
  XOR2_X1   g0030(.A(KEYINPUT2), .B(G226), .Z(new_n231));
  XNOR2_X1  g0031(.A(new_n230), .B(new_n231), .ZN(new_n232));
  XOR2_X1   g0032(.A(G264), .B(G270), .Z(new_n233));
  XNOR2_X1  g0033(.A(G250), .B(G257), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n232), .B(new_n235), .ZN(G358));
  XOR2_X1   g0036(.A(G87), .B(G97), .Z(new_n237));
  XNOR2_X1  g0037(.A(G107), .B(G116), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  INV_X1    g0039(.A(G50), .ZN(new_n240));
  NAND2_X1  g0040(.A1(new_n240), .A2(G68), .ZN(new_n241));
  INV_X1    g0041(.A(G68), .ZN(new_n242));
  NAND2_X1  g0042(.A1(new_n242), .A2(G50), .ZN(new_n243));
  NAND2_X1  g0043(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G58), .B(G77), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n239), .B(new_n246), .ZN(G351));
  INV_X1    g0047(.A(KEYINPUT13), .ZN(new_n248));
  INV_X1    g0048(.A(G41), .ZN(new_n249));
  INV_X1    g0049(.A(G45), .ZN(new_n250));
  AOI21_X1  g0050(.A(G1), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  NAND3_X1  g0052(.A1(new_n252), .A2(G1), .A3(G13), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n251), .A2(new_n253), .A3(G274), .ZN(new_n254));
  INV_X1    g0054(.A(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n253), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n256), .A2(new_n251), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n255), .B1(G238), .B2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G226), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1698), .ZN(new_n260));
  INV_X1    g0060(.A(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n261), .A2(KEYINPUT3), .ZN(new_n262));
  INV_X1    g0062(.A(KEYINPUT3), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n263), .A2(G33), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n260), .A2(new_n262), .A3(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT73), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n265), .A2(new_n266), .ZN(new_n267));
  XNOR2_X1  g0067(.A(KEYINPUT3), .B(G33), .ZN(new_n268));
  NAND3_X1  g0068(.A1(new_n268), .A2(KEYINPUT73), .A3(new_n260), .ZN(new_n269));
  NAND2_X1  g0069(.A1(new_n267), .A2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(KEYINPUT74), .ZN(new_n271));
  NAND4_X1  g0071(.A1(new_n262), .A2(new_n264), .A3(G232), .A4(G1698), .ZN(new_n272));
  NAND2_X1  g0072(.A1(G33), .A2(G97), .ZN(new_n273));
  AND2_X1   g0073(.A1(new_n272), .A2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n270), .A2(new_n271), .A3(new_n274), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n218), .A2(new_n252), .ZN(new_n276));
  INV_X1    g0076(.A(KEYINPUT67), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND3_X1  g0078(.A1(new_n218), .A2(KEYINPUT67), .A3(new_n252), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND2_X1  g0080(.A1(new_n275), .A2(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n271), .B1(new_n270), .B2(new_n274), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n248), .B(new_n258), .C1(new_n281), .C2(new_n282), .ZN(new_n283));
  INV_X1    g0083(.A(new_n283), .ZN(new_n284));
  AOI21_X1  g0084(.A(KEYINPUT73), .B1(new_n268), .B2(new_n260), .ZN(new_n285));
  AND4_X1   g0085(.A1(KEYINPUT73), .A2(new_n260), .A3(new_n262), .A4(new_n264), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n272), .A2(new_n273), .ZN(new_n288));
  OAI21_X1  g0088(.A(KEYINPUT74), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND3_X1  g0089(.A1(new_n289), .A2(new_n280), .A3(new_n275), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n248), .B1(new_n290), .B2(new_n258), .ZN(new_n291));
  OAI21_X1  g0091(.A(G200), .B1(new_n284), .B2(new_n291), .ZN(new_n292));
  INV_X1    g0092(.A(KEYINPUT75), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n292), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n258), .B1(new_n281), .B2(new_n282), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(KEYINPUT13), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n296), .A2(new_n283), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n297), .A2(KEYINPUT75), .A3(G200), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n294), .A2(new_n298), .ZN(new_n299));
  INV_X1    g0099(.A(G13), .ZN(new_n300));
  NOR3_X1   g0100(.A1(new_n300), .A2(new_n206), .A3(G1), .ZN(new_n301));
  INV_X1    g0101(.A(new_n301), .ZN(new_n302));
  NOR2_X1   g0102(.A1(new_n302), .A2(G68), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n303), .A2(KEYINPUT77), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT77), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n305), .B1(new_n302), .B2(G68), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(KEYINPUT12), .A3(new_n306), .ZN(new_n307));
  OR3_X1    g0107(.A1(new_n303), .A2(KEYINPUT77), .A3(KEYINPUT12), .ZN(new_n308));
  NAND3_X1  g0108(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n215), .A2(new_n217), .A3(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n301), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n205), .A2(G20), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n311), .A2(G68), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n307), .A2(new_n308), .A3(new_n313), .ZN(new_n314));
  INV_X1    g0114(.A(KEYINPUT78), .ZN(new_n315));
  OR2_X1    g0115(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n310), .A2(KEYINPUT68), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT68), .ZN(new_n318));
  NAND4_X1  g0118(.A1(new_n215), .A2(new_n217), .A3(new_n318), .A4(new_n309), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  NOR2_X1   g0120(.A1(G20), .A2(G33), .ZN(new_n321));
  AOI22_X1  g0121(.A1(new_n321), .A2(G50), .B1(G20), .B2(new_n242), .ZN(new_n322));
  INV_X1    g0122(.A(G77), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n206), .A2(G33), .ZN(new_n324));
  OAI21_X1  g0124(.A(new_n322), .B1(new_n323), .B2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g0126(.A(new_n326), .B(KEYINPUT11), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n314), .A2(new_n315), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n316), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  INV_X1    g0129(.A(KEYINPUT76), .ZN(new_n330));
  AOI211_X1 g0130(.A(new_n330), .B(new_n248), .C1(new_n290), .C2(new_n258), .ZN(new_n331));
  AOI21_X1  g0131(.A(KEYINPUT76), .B1(new_n295), .B2(KEYINPUT13), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G190), .ZN(new_n334));
  NOR2_X1   g0134(.A1(new_n284), .A2(new_n334), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n329), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  AND3_X1   g0136(.A1(new_n299), .A2(new_n336), .A3(KEYINPUT79), .ZN(new_n337));
  AOI21_X1  g0137(.A(KEYINPUT79), .B1(new_n299), .B2(new_n336), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n337), .A2(new_n338), .ZN(new_n339));
  INV_X1    g0139(.A(G179), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n284), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n333), .A2(new_n341), .ZN(new_n342));
  AOI21_X1  g0142(.A(KEYINPUT14), .B1(new_n297), .B2(G169), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT14), .ZN(new_n344));
  INV_X1    g0144(.A(G169), .ZN(new_n345));
  AOI211_X1 g0145(.A(new_n344), .B(new_n345), .C1(new_n296), .C2(new_n283), .ZN(new_n346));
  OAI21_X1  g0146(.A(new_n342), .B1(new_n343), .B2(new_n346), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n347), .A2(new_n329), .ZN(new_n348));
  INV_X1    g0148(.A(G1698), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n268), .A2(G222), .A3(new_n349), .ZN(new_n350));
  OAI21_X1  g0150(.A(new_n350), .B1(new_n323), .B2(new_n268), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n268), .A2(G1698), .ZN(new_n352));
  XNOR2_X1  g0152(.A(new_n352), .B(KEYINPUT66), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n351), .B1(new_n353), .B2(G223), .ZN(new_n354));
  AOI21_X1  g0154(.A(KEYINPUT67), .B1(new_n218), .B2(new_n252), .ZN(new_n355));
  AND2_X1   g0155(.A1(G33), .A2(G41), .ZN(new_n356));
  AOI211_X1 g0156(.A(new_n277), .B(new_n356), .C1(new_n215), .C2(new_n217), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n355), .A2(new_n357), .ZN(new_n358));
  NOR2_X1   g0158(.A1(new_n354), .A2(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(new_n257), .ZN(new_n360));
  OAI21_X1  g0160(.A(new_n254), .B1(new_n360), .B2(new_n259), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n359), .A2(new_n361), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n362), .A2(new_n340), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n363), .B1(new_n362), .B2(G169), .ZN(new_n364));
  XNOR2_X1  g0164(.A(KEYINPUT8), .B(G58), .ZN(new_n365));
  INV_X1    g0165(.A(G150), .ZN(new_n366));
  INV_X1    g0166(.A(new_n321), .ZN(new_n367));
  OAI22_X1  g0167(.A1(new_n365), .A2(new_n324), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(KEYINPUT69), .ZN(new_n369));
  AND2_X1   g0169(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G20), .B1(new_n202), .B2(G50), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(new_n368), .B2(new_n369), .ZN(new_n372));
  OAI21_X1  g0172(.A(new_n320), .B1(new_n370), .B2(new_n372), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT70), .ZN(new_n374));
  NAND3_X1  g0174(.A1(new_n317), .A2(new_n319), .A3(new_n302), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G50), .ZN(new_n376));
  AOI21_X1  g0176(.A(new_n301), .B1(G50), .B2(new_n312), .ZN(new_n377));
  INV_X1    g0177(.A(new_n377), .ZN(new_n378));
  AOI21_X1  g0178(.A(new_n374), .B1(new_n376), .B2(new_n378), .ZN(new_n379));
  AOI211_X1 g0179(.A(KEYINPUT70), .B(new_n377), .C1(new_n375), .C2(G50), .ZN(new_n380));
  OAI21_X1  g0180(.A(new_n373), .B1(new_n379), .B2(new_n380), .ZN(new_n381));
  INV_X1    g0181(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n364), .A2(new_n382), .ZN(new_n383));
  INV_X1    g0183(.A(G244), .ZN(new_n384));
  OAI21_X1  g0184(.A(new_n254), .B1(new_n360), .B2(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n268), .A2(G232), .A3(new_n349), .ZN(new_n387));
  INV_X1    g0187(.A(G107), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n387), .B1(new_n388), .B2(new_n268), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n389), .B1(new_n353), .B2(G238), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n386), .B1(new_n390), .B2(new_n358), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n391), .A2(G200), .ZN(new_n392));
  INV_X1    g0192(.A(new_n365), .ZN(new_n393));
  AOI22_X1  g0193(.A1(new_n393), .A2(new_n321), .B1(G20), .B2(G77), .ZN(new_n394));
  XNOR2_X1  g0194(.A(KEYINPUT15), .B(G87), .ZN(new_n395));
  OAI21_X1  g0195(.A(new_n394), .B1(new_n324), .B2(new_n395), .ZN(new_n396));
  AOI22_X1  g0196(.A1(new_n396), .A2(new_n310), .B1(new_n323), .B2(new_n301), .ZN(new_n397));
  INV_X1    g0197(.A(new_n312), .ZN(new_n398));
  NOR4_X1   g0198(.A1(new_n310), .A2(new_n301), .A3(new_n398), .A4(new_n323), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n397), .A2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(new_n401), .ZN(new_n402));
  OAI211_X1 g0202(.A(new_n392), .B(new_n402), .C1(new_n334), .C2(new_n391), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n391), .A2(new_n345), .ZN(new_n404));
  OAI211_X1 g0204(.A(new_n340), .B(new_n386), .C1(new_n390), .C2(new_n358), .ZN(new_n405));
  NAND3_X1  g0205(.A1(new_n404), .A2(new_n401), .A3(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n403), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g0207(.A1(new_n383), .A2(new_n407), .ZN(new_n408));
  INV_X1    g0208(.A(new_n375), .ZN(new_n409));
  NOR2_X1   g0209(.A1(new_n365), .A2(new_n398), .ZN(new_n410));
  AOI22_X1  g0210(.A1(new_n409), .A2(new_n410), .B1(new_n301), .B2(new_n365), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT81), .ZN(new_n412));
  OAI21_X1  g0212(.A(new_n412), .B1(new_n263), .B2(G33), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n261), .A2(KEYINPUT81), .A3(KEYINPUT3), .ZN(new_n414));
  NAND3_X1  g0214(.A1(new_n413), .A2(new_n264), .A3(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(KEYINPUT7), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n416), .A2(G20), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n415), .A2(KEYINPUT82), .A3(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n416), .B1(new_n268), .B2(G20), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  AOI21_X1  g0220(.A(KEYINPUT82), .B1(new_n415), .B2(new_n417), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(G58), .A2(G68), .ZN(new_n423));
  AOI21_X1  g0223(.A(new_n206), .B1(new_n202), .B2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(G159), .ZN(new_n425));
  NOR2_X1   g0225(.A1(new_n367), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT80), .B1(new_n424), .B2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(new_n423), .ZN(new_n428));
  OAI21_X1  g0228(.A(G20), .B1(new_n428), .B2(new_n201), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT80), .ZN(new_n430));
  OAI211_X1 g0230(.A(new_n429), .B(new_n430), .C1(new_n425), .C2(new_n367), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n427), .A2(new_n431), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI21_X1  g0233(.A(KEYINPUT16), .B1(new_n422), .B2(new_n433), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n262), .A2(new_n264), .ZN(new_n435));
  AOI21_X1  g0235(.A(KEYINPUT7), .B1(new_n435), .B2(new_n206), .ZN(new_n436));
  INV_X1    g0236(.A(new_n417), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n268), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(G68), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n439), .A2(KEYINPUT16), .A3(new_n431), .A4(new_n427), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n440), .A2(new_n310), .ZN(new_n441));
  OAI21_X1  g0241(.A(new_n411), .B1(new_n434), .B2(new_n441), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n259), .A2(G1698), .ZN(new_n443));
  OAI21_X1  g0243(.A(new_n443), .B1(G223), .B2(G1698), .ZN(new_n444));
  INV_X1    g0244(.A(G87), .ZN(new_n445));
  OAI22_X1  g0245(.A1(new_n444), .A2(new_n435), .B1(new_n261), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g0246(.A(new_n446), .B1(new_n355), .B2(new_n357), .ZN(new_n447));
  AOI21_X1  g0247(.A(new_n255), .B1(G232), .B2(new_n257), .ZN(new_n448));
  NAND3_X1  g0248(.A1(new_n447), .A2(new_n448), .A3(G179), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n448), .ZN(new_n450));
  OAI21_X1  g0250(.A(new_n449), .B1(new_n450), .B2(new_n345), .ZN(new_n451));
  AND3_X1   g0251(.A1(new_n442), .A2(KEYINPUT18), .A3(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(KEYINPUT18), .B1(new_n442), .B2(new_n451), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  NAND3_X1  g0254(.A1(new_n447), .A2(new_n448), .A3(new_n334), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(new_n450), .B2(G200), .ZN(new_n456));
  OAI211_X1 g0256(.A(new_n456), .B(new_n411), .C1(new_n434), .C2(new_n441), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT17), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  OR2_X1    g0259(.A1(new_n434), .A2(new_n441), .ZN(new_n460));
  NAND4_X1  g0260(.A1(new_n460), .A2(KEYINPUT17), .A3(new_n411), .A4(new_n456), .ZN(new_n461));
  NAND2_X1  g0261(.A1(new_n459), .A2(new_n461), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n454), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g0263(.A1(new_n348), .A2(new_n408), .A3(new_n463), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n339), .A2(new_n464), .ZN(new_n465));
  OAI21_X1  g0265(.A(G200), .B1(new_n359), .B2(new_n361), .ZN(new_n466));
  INV_X1    g0266(.A(new_n361), .ZN(new_n467));
  OAI211_X1 g0267(.A(G190), .B(new_n467), .C1(new_n354), .C2(new_n358), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT9), .ZN(new_n469));
  AOI21_X1  g0269(.A(new_n377), .B1(new_n375), .B2(G50), .ZN(new_n470));
  XNOR2_X1  g0270(.A(new_n470), .B(new_n374), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n469), .B1(new_n471), .B2(new_n373), .ZN(new_n472));
  OAI211_X1 g0272(.A(new_n469), .B(new_n373), .C1(new_n379), .C2(new_n380), .ZN(new_n473));
  INV_X1    g0273(.A(new_n473), .ZN(new_n474));
  OAI211_X1 g0274(.A(new_n466), .B(new_n468), .C1(new_n472), .C2(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT10), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT72), .ZN(new_n477));
  OAI21_X1  g0277(.A(KEYINPUT71), .B1(new_n472), .B2(new_n474), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n381), .A2(KEYINPUT9), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT71), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n479), .A2(new_n480), .A3(new_n473), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n478), .A2(new_n481), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT10), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n466), .A2(new_n483), .A3(new_n468), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n477), .B1(new_n482), .B2(new_n485), .ZN(new_n486));
  AOI211_X1 g0286(.A(KEYINPUT72), .B(new_n484), .C1(new_n478), .C2(new_n481), .ZN(new_n487));
  OAI21_X1  g0287(.A(new_n476), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n465), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g0289(.A(KEYINPUT25), .B1(new_n301), .B2(new_n388), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n490), .B(KEYINPUT89), .ZN(new_n491));
  NAND3_X1  g0291(.A1(new_n301), .A2(KEYINPUT25), .A3(new_n388), .ZN(new_n492));
  XNOR2_X1  g0292(.A(new_n492), .B(KEYINPUT88), .ZN(new_n493));
  NAND2_X1  g0293(.A1(new_n205), .A2(G33), .ZN(new_n494));
  NAND4_X1  g0294(.A1(new_n317), .A2(new_n319), .A3(new_n302), .A4(new_n494), .ZN(new_n495));
  OAI22_X1  g0295(.A1(new_n491), .A2(new_n493), .B1(new_n388), .B2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(new_n496), .ZN(new_n497));
  INV_X1    g0297(.A(KEYINPUT87), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n262), .A2(new_n264), .A3(new_n206), .A4(G87), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT22), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT22), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n268), .A2(new_n501), .A3(new_n206), .A4(G87), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT23), .ZN(new_n504));
  OAI21_X1  g0304(.A(new_n504), .B1(new_n206), .B2(G107), .ZN(new_n505));
  NAND3_X1  g0305(.A1(new_n388), .A2(KEYINPUT23), .A3(G20), .ZN(new_n506));
  INV_X1    g0306(.A(G116), .ZN(new_n507));
  NOR2_X1   g0307(.A1(new_n261), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g0308(.A1(new_n505), .A2(new_n506), .B1(new_n508), .B2(new_n206), .ZN(new_n509));
  NAND2_X1  g0309(.A1(new_n503), .A2(new_n509), .ZN(new_n510));
  XOR2_X1   g0310(.A(KEYINPUT86), .B(KEYINPUT24), .Z(new_n511));
  INV_X1    g0311(.A(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n503), .A2(new_n509), .A3(new_n511), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n513), .A2(new_n514), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n498), .B1(new_n515), .B2(new_n310), .ZN(new_n516));
  AND3_X1   g0316(.A1(new_n503), .A2(new_n509), .A3(new_n511), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n511), .B1(new_n503), .B2(new_n509), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n498), .B(new_n310), .C1(new_n517), .C2(new_n518), .ZN(new_n519));
  INV_X1    g0319(.A(new_n519), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n497), .B1(new_n516), .B2(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(G257), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G1698), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(G250), .B2(G1698), .ZN(new_n524));
  INV_X1    g0324(.A(G294), .ZN(new_n525));
  OAI22_X1  g0325(.A1(new_n524), .A2(new_n435), .B1(new_n261), .B2(new_n525), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n526), .B1(new_n355), .B2(new_n357), .ZN(new_n527));
  XNOR2_X1  g0327(.A(KEYINPUT5), .B(G41), .ZN(new_n528));
  NOR2_X1   g0328(.A1(new_n250), .A2(G1), .ZN(new_n529));
  NAND4_X1  g0329(.A1(new_n528), .A2(G274), .A3(new_n529), .A4(new_n253), .ZN(new_n530));
  AOI21_X1  g0330(.A(new_n256), .B1(new_n529), .B2(new_n528), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n531), .A2(G264), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n527), .A2(new_n530), .A3(new_n532), .ZN(new_n533));
  NAND2_X1  g0333(.A1(new_n533), .A2(new_n345), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(G179), .B2(new_n533), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n521), .A2(new_n536), .A3(KEYINPUT90), .ZN(new_n537));
  INV_X1    g0337(.A(KEYINPUT90), .ZN(new_n538));
  OAI21_X1  g0338(.A(new_n310), .B1(new_n517), .B2(new_n518), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(KEYINPUT87), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n496), .B1(new_n540), .B2(new_n519), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n535), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n537), .A2(new_n542), .ZN(new_n543));
  INV_X1    g0343(.A(G200), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n533), .A2(new_n544), .ZN(new_n545));
  OAI21_X1  g0345(.A(new_n545), .B1(G190), .B2(new_n533), .ZN(new_n546));
  OAI211_X1 g0346(.A(new_n546), .B(new_n497), .C1(new_n516), .C2(new_n520), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n262), .A2(new_n264), .A3(G238), .A4(new_n349), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(KEYINPUT84), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT84), .ZN(new_n550));
  NAND4_X1  g0350(.A1(new_n268), .A2(new_n550), .A3(G238), .A4(new_n349), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n549), .A2(new_n551), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(G1698), .ZN(new_n553));
  INV_X1    g0353(.A(new_n508), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n552), .A2(new_n556), .B1(new_n278), .B2(new_n279), .ZN(new_n557));
  INV_X1    g0357(.A(new_n529), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n558), .A2(G250), .A3(new_n253), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n253), .A2(G274), .A3(new_n529), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(G200), .B1(new_n557), .B2(new_n561), .ZN(new_n562));
  NOR3_X1   g0362(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n563));
  AND2_X1   g0363(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n564));
  NOR2_X1   g0364(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n565));
  OAI211_X1 g0365(.A(G33), .B(G97), .C1(new_n564), .C2(new_n565), .ZN(new_n566));
  AOI21_X1  g0366(.A(new_n563), .B1(new_n566), .B2(new_n206), .ZN(new_n567));
  OR2_X1    g0367(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n568));
  NAND2_X1  g0368(.A1(KEYINPUT85), .A2(KEYINPUT19), .ZN(new_n569));
  INV_X1    g0369(.A(G97), .ZN(new_n570));
  OAI211_X1 g0370(.A(new_n568), .B(new_n569), .C1(new_n324), .C2(new_n570), .ZN(new_n571));
  NAND4_X1  g0371(.A1(new_n262), .A2(new_n264), .A3(new_n206), .A4(G68), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n310), .B1(new_n567), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n395), .A2(new_n301), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g0376(.A1(new_n495), .A2(new_n445), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  INV_X1    g0378(.A(new_n561), .ZN(new_n579));
  AOI21_X1  g0379(.A(new_n555), .B1(new_n551), .B2(new_n549), .ZN(new_n580));
  OAI211_X1 g0380(.A(G190), .B(new_n579), .C1(new_n580), .C2(new_n358), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n562), .A2(new_n578), .A3(new_n581), .ZN(new_n582));
  OAI211_X1 g0382(.A(new_n574), .B(new_n575), .C1(new_n495), .C2(new_n395), .ZN(new_n583));
  OAI211_X1 g0383(.A(new_n340), .B(new_n579), .C1(new_n580), .C2(new_n358), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n552), .A2(new_n556), .ZN(new_n585));
  AOI21_X1  g0385(.A(new_n561), .B1(new_n585), .B2(new_n280), .ZN(new_n586));
  OAI211_X1 g0386(.A(new_n583), .B(new_n584), .C1(new_n586), .C2(G169), .ZN(new_n587));
  AND2_X1   g0387(.A1(new_n582), .A2(new_n587), .ZN(new_n588));
  NAND4_X1  g0388(.A1(new_n262), .A2(new_n264), .A3(G244), .A4(new_n349), .ZN(new_n589));
  INV_X1    g0389(.A(KEYINPUT4), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n589), .A2(new_n590), .ZN(new_n591));
  NAND4_X1  g0391(.A1(new_n268), .A2(KEYINPUT4), .A3(G244), .A4(new_n349), .ZN(new_n592));
  AND3_X1   g0392(.A1(KEYINPUT83), .A2(G33), .A3(G283), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT83), .B1(G33), .B2(G283), .ZN(new_n594));
  OR2_X1    g0394(.A1(new_n593), .A2(new_n594), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n268), .A2(G250), .A3(G1698), .ZN(new_n596));
  NAND4_X1  g0396(.A1(new_n591), .A2(new_n592), .A3(new_n595), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n280), .A2(new_n597), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n528), .A2(new_n529), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n599), .A2(new_n253), .ZN(new_n600));
  OAI21_X1  g0400(.A(new_n530), .B1(new_n600), .B2(new_n522), .ZN(new_n601));
  INV_X1    g0401(.A(new_n601), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n598), .A2(new_n602), .A3(new_n340), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n601), .B1(new_n280), .B2(new_n597), .ZN(new_n604));
  INV_X1    g0404(.A(new_n310), .ZN(new_n605));
  OAI21_X1  g0405(.A(G107), .B1(new_n420), .B2(new_n421), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n388), .A2(KEYINPUT6), .A3(G97), .ZN(new_n607));
  XOR2_X1   g0407(.A(G97), .B(G107), .Z(new_n608));
  OAI21_X1  g0408(.A(new_n607), .B1(new_n608), .B2(KEYINPUT6), .ZN(new_n609));
  AOI22_X1  g0409(.A1(new_n609), .A2(G20), .B1(G77), .B2(new_n321), .ZN(new_n610));
  AOI21_X1  g0410(.A(new_n605), .B1(new_n606), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n301), .A2(new_n570), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n612), .B1(new_n495), .B2(new_n570), .ZN(new_n613));
  OAI221_X1 g0413(.A(new_n603), .B1(new_n604), .B2(G169), .C1(new_n611), .C2(new_n613), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n611), .A2(new_n613), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n598), .A2(new_n602), .A3(new_n334), .ZN(new_n616));
  OAI21_X1  g0416(.A(new_n616), .B1(new_n604), .B2(G200), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n615), .A2(new_n617), .ZN(new_n618));
  NAND4_X1  g0418(.A1(new_n547), .A2(new_n588), .A3(new_n614), .A4(new_n618), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n599), .A2(G270), .A3(new_n253), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n620), .A2(new_n530), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n262), .A2(new_n264), .A3(G257), .A4(new_n349), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n262), .A2(new_n264), .A3(G264), .A4(G1698), .ZN(new_n623));
  INV_X1    g0423(.A(G303), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n622), .B(new_n623), .C1(new_n624), .C2(new_n268), .ZN(new_n625));
  OAI21_X1  g0425(.A(new_n625), .B1(new_n355), .B2(new_n357), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n345), .B1(new_n621), .B2(new_n626), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n507), .B1(new_n205), .B2(G33), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n300), .A2(G1), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n507), .A2(G20), .ZN(new_n630));
  INV_X1    g0430(.A(new_n630), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n311), .A2(new_n628), .B1(new_n629), .B2(new_n631), .ZN(new_n632));
  AOI21_X1  g0432(.A(G20), .B1(new_n261), .B2(G97), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n633), .B1(new_n593), .B2(new_n594), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n634), .A2(new_n310), .A3(new_n630), .ZN(new_n635));
  INV_X1    g0435(.A(KEYINPUT20), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  NOR2_X1   g0437(.A1(new_n635), .A2(new_n636), .ZN(new_n638));
  OAI21_X1  g0438(.A(new_n632), .B1(new_n637), .B2(new_n638), .ZN(new_n639));
  NAND3_X1  g0439(.A1(new_n627), .A2(new_n639), .A3(KEYINPUT21), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n620), .A2(new_n530), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n641), .B1(new_n280), .B2(new_n625), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n639), .A2(new_n642), .A3(G179), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n640), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT21), .B1(new_n627), .B2(new_n639), .ZN(new_n645));
  NOR2_X1   g0445(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g0446(.A1(new_n621), .A2(new_n626), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n639), .B1(G200), .B2(new_n647), .ZN(new_n648));
  OAI21_X1  g0448(.A(new_n648), .B1(new_n334), .B2(new_n647), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n646), .A2(new_n649), .ZN(new_n650));
  NOR4_X1   g0450(.A1(new_n489), .A2(new_n543), .A3(new_n619), .A4(new_n650), .ZN(G372));
  INV_X1    g0451(.A(new_n489), .ZN(new_n652));
  INV_X1    g0452(.A(KEYINPUT91), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n627), .A2(new_n639), .ZN(new_n654));
  INV_X1    g0454(.A(KEYINPUT21), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g0456(.A1(new_n656), .A2(new_n643), .A3(new_n640), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n657), .B1(new_n521), .B2(new_n536), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n653), .B1(new_n619), .B2(new_n658), .ZN(new_n659));
  AND4_X1   g0459(.A1(new_n614), .A2(new_n618), .A3(new_n587), .A4(new_n582), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n646), .B1(new_n541), .B2(new_n535), .ZN(new_n661));
  NAND4_X1  g0461(.A1(new_n660), .A2(new_n661), .A3(KEYINPUT91), .A4(new_n547), .ZN(new_n662));
  INV_X1    g0462(.A(new_n587), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n603), .B1(new_n604), .B2(G169), .ZN(new_n664));
  NOR2_X1   g0464(.A1(new_n615), .A2(new_n664), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n588), .A2(KEYINPUT26), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT26), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n582), .A2(new_n587), .ZN(new_n668));
  OAI21_X1  g0468(.A(new_n667), .B1(new_n614), .B2(new_n668), .ZN(new_n669));
  AOI21_X1  g0469(.A(new_n663), .B1(new_n666), .B2(new_n669), .ZN(new_n670));
  NAND3_X1  g0470(.A1(new_n659), .A2(new_n662), .A3(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n652), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n299), .A2(new_n336), .ZN(new_n673));
  INV_X1    g0473(.A(new_n406), .ZN(new_n674));
  AOI22_X1  g0474(.A1(new_n673), .A2(new_n674), .B1(new_n347), .B2(new_n329), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT92), .ZN(new_n676));
  NAND3_X1  g0476(.A1(new_n442), .A2(new_n676), .A3(new_n451), .ZN(new_n677));
  INV_X1    g0477(.A(new_n677), .ZN(new_n678));
  INV_X1    g0478(.A(KEYINPUT18), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n676), .B1(new_n442), .B2(new_n451), .ZN(new_n680));
  NOR3_X1   g0480(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  NAND2_X1  g0481(.A1(new_n442), .A2(new_n451), .ZN(new_n682));
  NAND2_X1  g0482(.A1(new_n682), .A2(KEYINPUT92), .ZN(new_n683));
  AOI21_X1  g0483(.A(KEYINPUT18), .B1(new_n683), .B2(new_n677), .ZN(new_n684));
  OAI22_X1  g0484(.A1(new_n675), .A2(new_n462), .B1(new_n681), .B2(new_n684), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n383), .B1(new_n685), .B2(new_n488), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n672), .A2(new_n686), .ZN(G369));
  AND2_X1   g0487(.A1(new_n537), .A2(new_n542), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n629), .A2(new_n206), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n689), .A2(KEYINPUT27), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(G213), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(G343), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  OAI211_X1 g0495(.A(new_n688), .B(new_n547), .C1(new_n541), .C2(new_n695), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n646), .A2(new_n694), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OR2_X1    g0498(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  NOR2_X1   g0499(.A1(new_n541), .A2(new_n535), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n700), .A2(new_n695), .ZN(new_n701));
  AND2_X1   g0501(.A1(new_n699), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n700), .A2(new_n694), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n696), .A2(new_n703), .ZN(new_n704));
  INV_X1    g0504(.A(KEYINPUT93), .ZN(new_n705));
  AND2_X1   g0505(.A1(new_n639), .A2(new_n694), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n657), .A2(new_n706), .ZN(new_n707));
  OAI211_X1 g0507(.A(new_n705), .B(new_n707), .C1(new_n650), .C2(new_n706), .ZN(new_n708));
  OAI21_X1  g0508(.A(new_n708), .B1(new_n705), .B2(new_n707), .ZN(new_n709));
  INV_X1    g0509(.A(G330), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n704), .A2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n702), .A2(new_n712), .ZN(G399));
  INV_X1    g0513(.A(new_n209), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n714), .A2(G41), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n563), .A2(new_n507), .ZN(new_n716));
  NOR3_X1   g0516(.A1(new_n715), .A2(new_n716), .A3(new_n205), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n213), .B2(new_n715), .ZN(new_n718));
  XOR2_X1   g0518(.A(new_n718), .B(KEYINPUT94), .Z(new_n719));
  XNOR2_X1  g0519(.A(new_n719), .B(KEYINPUT28), .ZN(new_n720));
  NOR2_X1   g0520(.A1(new_n619), .A2(new_n650), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n721), .A2(new_n688), .A3(new_n695), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n647), .A2(new_n340), .ZN(new_n723));
  AND2_X1   g0523(.A1(new_n527), .A2(new_n532), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n723), .A2(new_n724), .A3(new_n604), .A4(new_n586), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT30), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  AND2_X1   g0527(.A1(new_n604), .A2(new_n724), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n728), .A2(KEYINPUT30), .A3(new_n586), .A4(new_n723), .ZN(new_n729));
  NOR3_X1   g0529(.A1(new_n604), .A2(new_n642), .A3(G179), .ZN(new_n730));
  INV_X1    g0530(.A(new_n586), .ZN(new_n731));
  NAND3_X1  g0531(.A1(new_n730), .A2(new_n533), .A3(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n727), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  AND3_X1   g0533(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n734));
  AOI21_X1  g0534(.A(KEYINPUT31), .B1(new_n733), .B2(new_n694), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n734), .A2(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n710), .B1(new_n722), .B2(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n671), .A2(new_n695), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT29), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  OAI211_X1 g0540(.A(new_n547), .B(new_n660), .C1(new_n543), .C2(new_n657), .ZN(new_n741));
  NAND2_X1  g0541(.A1(new_n741), .A2(new_n670), .ZN(new_n742));
  NAND3_X1  g0542(.A1(new_n742), .A2(KEYINPUT29), .A3(new_n695), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n737), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  OAI21_X1  g0544(.A(new_n720), .B1(new_n744), .B2(G1), .ZN(G364));
  NOR2_X1   g0545(.A1(new_n300), .A2(G20), .ZN(new_n746));
  AOI21_X1  g0546(.A(new_n205), .B1(new_n746), .B2(G45), .ZN(new_n747));
  INV_X1    g0547(.A(new_n747), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n715), .A2(new_n748), .ZN(new_n749));
  OAI21_X1  g0549(.A(new_n218), .B1(new_n206), .B2(G169), .ZN(new_n750));
  INV_X1    g0550(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g0551(.A1(G13), .A2(G33), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(G20), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n714), .A2(new_n435), .ZN(new_n757));
  AOI22_X1  g0557(.A1(new_n757), .A2(G355), .B1(new_n507), .B2(new_n714), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n714), .A2(new_n268), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n759), .B1(G45), .B2(new_n212), .ZN(new_n760));
  NOR2_X1   g0560(.A1(new_n246), .A2(new_n250), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  INV_X1    g0562(.A(KEYINPUT95), .ZN(new_n763));
  AOI21_X1  g0563(.A(new_n756), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n764), .B1(new_n763), .B2(new_n762), .ZN(new_n765));
  NOR2_X1   g0565(.A1(new_n206), .A2(new_n340), .ZN(new_n766));
  NOR2_X1   g0566(.A1(G190), .A2(G200), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  INV_X1    g0568(.A(G58), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n334), .A2(G200), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n766), .A2(new_n770), .ZN(new_n771));
  OAI221_X1 g0571(.A(new_n268), .B1(new_n768), .B2(new_n323), .C1(new_n769), .C2(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n206), .A2(G179), .ZN(new_n773));
  NAND3_X1  g0573(.A1(new_n773), .A2(new_n334), .A3(G200), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n774), .A2(new_n388), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n766), .A2(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n334), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n775), .B1(G50), .B2(new_n777), .ZN(new_n778));
  NOR2_X1   g0578(.A1(new_n776), .A2(G190), .ZN(new_n779));
  INV_X1    g0579(.A(new_n779), .ZN(new_n780));
  NAND3_X1  g0580(.A1(new_n773), .A2(G190), .A3(G200), .ZN(new_n781));
  OAI221_X1 g0581(.A(new_n778), .B1(new_n242), .B2(new_n780), .C1(new_n445), .C2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n206), .B1(new_n770), .B2(new_n340), .ZN(new_n783));
  XOR2_X1   g0583(.A(new_n783), .B(KEYINPUT97), .Z(new_n784));
  AOI211_X1 g0584(.A(new_n772), .B(new_n782), .C1(G97), .C2(new_n784), .ZN(new_n785));
  AND2_X1   g0585(.A1(new_n773), .A2(new_n767), .ZN(new_n786));
  OR2_X1    g0586(.A1(new_n786), .A2(KEYINPUT96), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n786), .A2(KEYINPUT96), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n425), .ZN(new_n790));
  XNOR2_X1  g0590(.A(new_n790), .B(KEYINPUT32), .ZN(new_n791));
  INV_X1    g0591(.A(new_n789), .ZN(new_n792));
  AND2_X1   g0592(.A1(new_n792), .A2(G329), .ZN(new_n793));
  XOR2_X1   g0593(.A(new_n781), .B(KEYINPUT98), .Z(new_n794));
  INV_X1    g0594(.A(new_n794), .ZN(new_n795));
  NOR2_X1   g0595(.A1(new_n795), .A2(new_n624), .ZN(new_n796));
  INV_X1    g0596(.A(G311), .ZN(new_n797));
  OAI221_X1 g0597(.A(new_n435), .B1(new_n768), .B2(new_n797), .C1(new_n783), .C2(new_n525), .ZN(new_n798));
  INV_X1    g0598(.A(new_n777), .ZN(new_n799));
  INV_X1    g0599(.A(G326), .ZN(new_n800));
  INV_X1    g0600(.A(G283), .ZN(new_n801));
  OAI22_X1  g0601(.A1(new_n799), .A2(new_n800), .B1(new_n801), .B2(new_n774), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n793), .A2(new_n796), .A3(new_n798), .A4(new_n802), .ZN(new_n803));
  XOR2_X1   g0603(.A(KEYINPUT33), .B(G317), .Z(new_n804));
  INV_X1    g0604(.A(G322), .ZN(new_n805));
  OAI22_X1  g0605(.A1(new_n780), .A2(new_n804), .B1(new_n771), .B2(new_n805), .ZN(new_n806));
  XOR2_X1   g0606(.A(new_n806), .B(KEYINPUT99), .Z(new_n807));
  AOI22_X1  g0607(.A1(new_n785), .A2(new_n791), .B1(new_n803), .B2(new_n807), .ZN(new_n808));
  OAI211_X1 g0608(.A(new_n749), .B(new_n765), .C1(new_n808), .C2(new_n750), .ZN(new_n809));
  AOI21_X1  g0609(.A(new_n809), .B1(new_n709), .B2(new_n754), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n711), .A2(new_n749), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n709), .A2(new_n710), .ZN(new_n812));
  AOI21_X1  g0612(.A(new_n810), .B1(new_n811), .B2(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n813), .ZN(G396));
  INV_X1    g0614(.A(KEYINPUT100), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n674), .A2(new_n695), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n401), .A2(new_n694), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n403), .A2(new_n817), .ZN(new_n818));
  OAI21_X1  g0618(.A(new_n816), .B1(new_n818), .B2(new_n674), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n738), .A2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(new_n819), .ZN(new_n821));
  NAND3_X1  g0621(.A1(new_n671), .A2(new_n695), .A3(new_n821), .ZN(new_n822));
  NAND2_X1  g0622(.A1(new_n820), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g0623(.A1(new_n823), .A2(new_n737), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n722), .A2(new_n736), .ZN(new_n825));
  INV_X1    g0625(.A(new_n825), .ZN(new_n826));
  OAI211_X1 g0626(.A(new_n820), .B(new_n822), .C1(new_n710), .C2(new_n826), .ZN(new_n827));
  INV_X1    g0627(.A(new_n749), .ZN(new_n828));
  NAND3_X1  g0628(.A1(new_n824), .A2(new_n827), .A3(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n821), .A2(new_n753), .ZN(new_n830));
  INV_X1    g0630(.A(new_n771), .ZN(new_n831));
  INV_X1    g0631(.A(new_n768), .ZN(new_n832));
  AOI22_X1  g0632(.A1(G143), .A2(new_n831), .B1(new_n832), .B2(G159), .ZN(new_n833));
  INV_X1    g0633(.A(G137), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n833), .B1(new_n780), .B2(new_n366), .C1(new_n834), .C2(new_n799), .ZN(new_n835));
  XNOR2_X1  g0635(.A(new_n835), .B(KEYINPUT34), .ZN(new_n836));
  INV_X1    g0636(.A(new_n774), .ZN(new_n837));
  NAND2_X1  g0637(.A1(new_n837), .A2(G68), .ZN(new_n838));
  INV_X1    g0638(.A(new_n783), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n435), .B1(new_n839), .B2(G58), .ZN(new_n840));
  INV_X1    g0640(.A(G132), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n838), .B(new_n840), .C1(new_n789), .C2(new_n841), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(G50), .B2(new_n794), .ZN(new_n843));
  OAI221_X1 g0643(.A(new_n435), .B1(new_n768), .B2(new_n507), .C1(new_n525), .C2(new_n771), .ZN(new_n844));
  AOI22_X1  g0644(.A1(new_n779), .A2(G283), .B1(new_n837), .B2(G87), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n845), .B1(new_n624), .B2(new_n799), .ZN(new_n846));
  AOI211_X1 g0646(.A(new_n844), .B(new_n846), .C1(G311), .C2(new_n792), .ZN(new_n847));
  AOI22_X1  g0647(.A1(G97), .A2(new_n784), .B1(new_n794), .B2(G107), .ZN(new_n848));
  AOI22_X1  g0648(.A1(new_n836), .A2(new_n843), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  NOR2_X1   g0649(.A1(new_n751), .A2(new_n752), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  OAI22_X1  g0651(.A1(new_n849), .A2(new_n750), .B1(G77), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n749), .B1(new_n830), .B2(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n815), .B1(new_n829), .B2(new_n853), .ZN(new_n854));
  INV_X1    g0654(.A(new_n854), .ZN(new_n855));
  NAND3_X1  g0655(.A1(new_n829), .A2(new_n815), .A3(new_n853), .ZN(new_n856));
  NAND2_X1  g0656(.A1(new_n855), .A2(new_n856), .ZN(G384));
  XOR2_X1   g0657(.A(new_n609), .B(KEYINPUT101), .Z(new_n858));
  NAND2_X1  g0658(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n859));
  NAND4_X1  g0659(.A1(new_n859), .A2(G20), .A3(G116), .A4(new_n218), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n858), .A2(KEYINPUT35), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  XNOR2_X1  g0662(.A(KEYINPUT102), .B(KEYINPUT36), .ZN(new_n863));
  XNOR2_X1  g0663(.A(new_n862), .B(new_n863), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n213), .A2(G77), .A3(new_n423), .ZN(new_n865));
  AOI211_X1 g0665(.A(new_n205), .B(G13), .C1(new_n865), .C2(new_n241), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n864), .A2(new_n866), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n347), .A2(new_n329), .A3(new_n695), .ZN(new_n868));
  INV_X1    g0668(.A(KEYINPUT39), .ZN(new_n869));
  INV_X1    g0669(.A(new_n692), .ZN(new_n870));
  AOI21_X1  g0670(.A(KEYINPUT16), .B1(new_n433), .B2(new_n439), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n440), .A2(new_n320), .ZN(new_n872));
  NOR2_X1   g0672(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(new_n411), .ZN(new_n874));
  OAI21_X1  g0674(.A(new_n870), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  OAI21_X1  g0676(.A(new_n876), .B1(new_n454), .B2(new_n462), .ZN(new_n877));
  OAI22_X1  g0677(.A1(new_n873), .A2(new_n874), .B1(new_n451), .B2(new_n870), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n878), .A2(new_n457), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  INV_X1    g0680(.A(KEYINPUT104), .ZN(new_n881));
  AND3_X1   g0681(.A1(new_n442), .A2(new_n881), .A3(new_n870), .ZN(new_n882));
  AOI21_X1  g0682(.A(new_n881), .B1(new_n442), .B2(new_n870), .ZN(new_n883));
  NOR2_X1   g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(KEYINPUT37), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n682), .A2(new_n457), .A3(new_n885), .ZN(new_n886));
  OAI21_X1  g0686(.A(new_n880), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NAND3_X1  g0687(.A1(new_n877), .A2(new_n887), .A3(KEYINPUT38), .ZN(new_n888));
  NOR3_X1   g0688(.A1(new_n884), .A2(KEYINPUT106), .A3(new_n886), .ZN(new_n889));
  INV_X1    g0689(.A(KEYINPUT106), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n442), .A2(new_n870), .ZN(new_n891));
  NAND2_X1  g0691(.A1(new_n891), .A2(KEYINPUT104), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n442), .A2(new_n881), .A3(new_n870), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n892), .A2(new_n893), .ZN(new_n894));
  AND3_X1   g0694(.A1(new_n682), .A2(new_n457), .A3(new_n885), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n890), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  NOR2_X1   g0696(.A1(new_n889), .A2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n457), .B1(new_n678), .B2(new_n680), .ZN(new_n898));
  OAI21_X1  g0698(.A(KEYINPUT37), .B1(new_n898), .B2(new_n884), .ZN(new_n899));
  INV_X1    g0699(.A(new_n462), .ZN(new_n900));
  OAI21_X1  g0700(.A(new_n900), .B1(new_n681), .B2(new_n684), .ZN(new_n901));
  AOI22_X1  g0701(.A1(new_n897), .A2(new_n899), .B1(new_n884), .B2(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n869), .B(new_n888), .C1(new_n902), .C2(KEYINPUT38), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n888), .A2(KEYINPUT105), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT105), .ZN(new_n905));
  NAND4_X1  g0705(.A1(new_n877), .A2(new_n887), .A3(new_n905), .A4(KEYINPUT38), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n877), .A2(new_n887), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT38), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n907), .A2(new_n908), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n904), .A2(new_n906), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n910), .A2(KEYINPUT39), .ZN(new_n911));
  AOI21_X1  g0711(.A(new_n868), .B1(new_n903), .B2(new_n911), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n816), .B(KEYINPUT103), .ZN(new_n913));
  INV_X1    g0713(.A(new_n913), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n822), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n329), .A2(new_n694), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n348), .A2(new_n673), .A3(new_n916), .ZN(new_n917));
  INV_X1    g0717(.A(KEYINPUT79), .ZN(new_n918));
  AOI21_X1  g0718(.A(KEYINPUT75), .B1(new_n297), .B2(G200), .ZN(new_n919));
  AOI211_X1 g0719(.A(new_n293), .B(new_n544), .C1(new_n296), .C2(new_n283), .ZN(new_n920));
  NOR2_X1   g0720(.A1(new_n919), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g0721(.A1(new_n296), .A2(new_n330), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n291), .A2(KEYINPUT76), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n335), .A2(new_n922), .A3(new_n923), .ZN(new_n924));
  INV_X1    g0724(.A(new_n329), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n918), .B1(new_n921), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n299), .A2(new_n336), .A3(KEYINPUT79), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n347), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n917), .B1(new_n929), .B2(new_n916), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n910), .A2(new_n915), .A3(new_n930), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n681), .A2(new_n684), .A3(new_n870), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n912), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n740), .A2(new_n465), .A3(new_n743), .A4(new_n488), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n935), .A2(new_n686), .ZN(new_n936));
  XOR2_X1   g0736(.A(new_n934), .B(new_n936), .Z(new_n937));
  NOR4_X1   g0737(.A1(new_n543), .A2(new_n619), .A3(new_n650), .A4(new_n694), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n733), .A2(new_n694), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT31), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n939), .A2(new_n940), .ZN(new_n941));
  NAND3_X1  g0741(.A1(new_n733), .A2(KEYINPUT31), .A3(new_n694), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  OAI21_X1  g0743(.A(new_n821), .B1(new_n938), .B2(new_n943), .ZN(new_n944));
  INV_X1    g0744(.A(new_n347), .ZN(new_n945));
  OAI21_X1  g0745(.A(new_n945), .B1(new_n337), .B2(new_n338), .ZN(new_n946));
  INV_X1    g0746(.A(new_n916), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n944), .B1(new_n948), .B2(new_n917), .ZN(new_n949));
  OAI21_X1  g0749(.A(new_n888), .B1(new_n902), .B2(KEYINPUT38), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT40), .ZN(new_n951));
  INV_X1    g0751(.A(new_n951), .ZN(new_n952));
  AOI21_X1  g0752(.A(KEYINPUT40), .B1(new_n949), .B2(new_n910), .ZN(new_n953));
  OAI22_X1  g0753(.A1(new_n952), .A2(new_n953), .B1(new_n489), .B2(new_n826), .ZN(new_n954));
  AOI21_X1  g0754(.A(new_n819), .B1(new_n722), .B2(new_n736), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n910), .A2(new_n930), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND4_X1  g0758(.A1(new_n951), .A2(new_n958), .A3(new_n652), .A4(new_n825), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n954), .A2(G330), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n937), .A2(new_n960), .ZN(new_n961));
  OAI21_X1  g0761(.A(new_n961), .B1(new_n205), .B2(new_n746), .ZN(new_n962));
  NOR2_X1   g0762(.A1(new_n937), .A2(new_n960), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n867), .B1(new_n962), .B2(new_n963), .ZN(G367));
  INV_X1    g0764(.A(new_n759), .ZN(new_n965));
  NOR2_X1   g0765(.A1(new_n965), .A2(new_n235), .ZN(new_n966));
  OAI21_X1  g0766(.A(new_n755), .B1(new_n209), .B2(new_n395), .ZN(new_n967));
  OAI21_X1  g0767(.A(new_n749), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  XNOR2_X1  g0768(.A(new_n968), .B(KEYINPUT112), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n784), .A2(G68), .ZN(new_n970));
  AOI22_X1  g0770(.A1(new_n777), .A2(G143), .B1(new_n831), .B2(G150), .ZN(new_n971));
  NAND2_X1  g0771(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g0772(.A(new_n972), .B(KEYINPUT114), .Z(new_n973));
  OAI22_X1  g0773(.A1(new_n780), .A2(new_n425), .B1(new_n781), .B2(new_n769), .ZN(new_n974));
  OAI221_X1 g0774(.A(new_n268), .B1(new_n768), .B2(new_n240), .C1(new_n323), .C2(new_n774), .ZN(new_n975));
  NOR2_X1   g0775(.A1(new_n974), .A2(new_n975), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n973), .B(new_n976), .C1(new_n834), .C2(new_n789), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n435), .B1(new_n771), .B2(new_n624), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n780), .A2(new_n525), .B1(new_n799), .B2(new_n797), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(G97), .C2(new_n837), .ZN(new_n980));
  AOI22_X1  g0780(.A1(new_n839), .A2(G107), .B1(new_n832), .B2(G283), .ZN(new_n981));
  INV_X1    g0781(.A(new_n981), .ZN(new_n982));
  AND2_X1   g0782(.A1(KEYINPUT46), .A2(G116), .ZN(new_n983));
  AOI22_X1  g0783(.A1(new_n982), .A2(KEYINPUT113), .B1(new_n794), .B2(new_n983), .ZN(new_n984));
  INV_X1    g0784(.A(new_n781), .ZN(new_n985));
  AOI21_X1  g0785(.A(KEYINPUT46), .B1(new_n985), .B2(G116), .ZN(new_n986));
  AOI21_X1  g0786(.A(new_n986), .B1(new_n792), .B2(G317), .ZN(new_n987));
  OR2_X1    g0787(.A1(new_n982), .A2(KEYINPUT113), .ZN(new_n988));
  NAND4_X1  g0788(.A1(new_n980), .A2(new_n984), .A3(new_n987), .A4(new_n988), .ZN(new_n989));
  AOI21_X1  g0789(.A(KEYINPUT47), .B1(new_n977), .B2(new_n989), .ZN(new_n990));
  NOR2_X1   g0790(.A1(new_n990), .A2(new_n750), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n977), .A2(KEYINPUT47), .A3(new_n989), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n969), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  INV_X1    g0793(.A(new_n754), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n578), .A2(new_n695), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n663), .A2(new_n995), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n996), .B1(new_n668), .B2(new_n995), .ZN(new_n997));
  OAI21_X1  g0797(.A(new_n993), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n715), .B(KEYINPUT41), .Z(new_n999));
  OAI211_X1 g0799(.A(new_n614), .B(new_n618), .C1(new_n615), .C2(new_n695), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n665), .A2(new_n694), .ZN(new_n1001));
  NAND2_X1  g0801(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NOR2_X1   g0802(.A1(new_n702), .A2(new_n1002), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT44), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n702), .A2(new_n1002), .ZN(new_n1005));
  INV_X1    g0805(.A(KEYINPUT45), .ZN(new_n1006));
  XNOR2_X1  g0806(.A(new_n1005), .B(new_n1006), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1004), .A2(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n712), .ZN(new_n1009));
  NAND2_X1  g0809(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n1010), .A2(KEYINPUT111), .ZN(new_n1011));
  OAI21_X1  g0811(.A(new_n699), .B1(new_n704), .B2(new_n697), .ZN(new_n1012));
  XNOR2_X1  g0812(.A(new_n1012), .B(new_n711), .ZN(new_n1013));
  NAND2_X1  g0813(.A1(new_n1013), .A2(new_n744), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n1014), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1004), .A2(new_n1007), .A3(new_n712), .ZN(new_n1016));
  INV_X1    g0816(.A(KEYINPUT111), .ZN(new_n1017));
  NAND3_X1  g0817(.A1(new_n1008), .A2(new_n1017), .A3(new_n1009), .ZN(new_n1018));
  NAND4_X1  g0818(.A1(new_n1011), .A2(new_n1015), .A3(new_n1016), .A4(new_n1018), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n999), .B1(new_n1019), .B2(new_n744), .ZN(new_n1020));
  NOR2_X1   g0820(.A1(new_n1020), .A2(new_n748), .ZN(new_n1021));
  OR2_X1    g0821(.A1(new_n688), .A2(new_n1000), .ZN(new_n1022));
  AOI21_X1  g0822(.A(new_n694), .B1(new_n1022), .B2(new_n614), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n1002), .ZN(new_n1024));
  NOR2_X1   g0824(.A1(new_n699), .A2(new_n1024), .ZN(new_n1025));
  XNOR2_X1  g0825(.A(new_n1025), .B(KEYINPUT109), .ZN(new_n1026));
  AOI21_X1  g0826(.A(new_n1023), .B1(new_n1026), .B2(KEYINPUT42), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(KEYINPUT42), .B2(new_n1026), .ZN(new_n1028));
  NAND2_X1  g0828(.A1(new_n997), .A2(KEYINPUT43), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n1028), .A2(new_n1029), .ZN(new_n1030));
  OR2_X1    g0830(.A1(new_n997), .A2(KEYINPUT107), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n997), .A2(KEYINPUT107), .ZN(new_n1032));
  XOR2_X1   g0832(.A(KEYINPUT108), .B(KEYINPUT43), .Z(new_n1033));
  AND3_X1   g0833(.A1(new_n1031), .A2(new_n1032), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1030), .A2(new_n1034), .ZN(new_n1035));
  INV_X1    g0835(.A(new_n1034), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1028), .A2(new_n1036), .A3(new_n1029), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1035), .A2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g0838(.A1(new_n712), .A2(new_n1024), .ZN(new_n1039));
  NOR2_X1   g0839(.A1(new_n1039), .A2(KEYINPUT110), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n1038), .A2(new_n1040), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n1035), .A2(new_n1037), .B1(KEYINPUT110), .B2(new_n1039), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n1040), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n998), .B1(new_n1021), .B2(new_n1043), .ZN(G387));
  NAND3_X1  g0844(.A1(new_n696), .A2(new_n703), .A3(new_n754), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n757), .A2(new_n716), .ZN(new_n1046));
  OAI21_X1  g0846(.A(new_n1046), .B1(G107), .B2(new_n209), .ZN(new_n1047));
  OR2_X1    g0847(.A1(new_n232), .A2(new_n250), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n365), .A2(G50), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT50), .ZN(new_n1050));
  AOI211_X1 g0850(.A(G45), .B(new_n716), .C1(G68), .C2(G77), .ZN(new_n1051));
  AOI21_X1  g0851(.A(new_n965), .B1(new_n1050), .B2(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n1047), .B1(new_n1048), .B2(new_n1052), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n749), .B1(new_n1053), .B2(new_n756), .ZN(new_n1054));
  INV_X1    g0854(.A(new_n784), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1055), .A2(new_n395), .ZN(new_n1056));
  AOI22_X1  g0856(.A1(new_n985), .A2(G77), .B1(new_n837), .B2(G97), .ZN(new_n1057));
  AOI22_X1  g0857(.A1(G159), .A2(new_n777), .B1(new_n779), .B2(new_n393), .ZN(new_n1058));
  OAI221_X1 g0858(.A(new_n268), .B1(new_n768), .B2(new_n242), .C1(new_n240), .C2(new_n771), .ZN(new_n1059));
  XNOR2_X1  g0859(.A(KEYINPUT115), .B(G150), .ZN(new_n1060));
  AOI21_X1  g0860(.A(new_n1059), .B1(new_n792), .B2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1061), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n1062), .B(KEYINPUT116), .Z(new_n1063));
  AOI21_X1  g0863(.A(new_n268), .B1(new_n837), .B2(G116), .ZN(new_n1064));
  OAI22_X1  g0864(.A1(new_n783), .A2(new_n801), .B1(new_n781), .B2(new_n525), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G303), .A2(new_n832), .B1(new_n831), .B2(G317), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n780), .B2(new_n797), .C1(new_n805), .C2(new_n799), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  AOI21_X1  g0868(.A(new_n1065), .B1(new_n1067), .B2(new_n1068), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n1069), .B1(new_n1068), .B2(new_n1067), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT49), .ZN(new_n1071));
  OAI221_X1 g0871(.A(new_n1064), .B1(new_n800), .B2(new_n789), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1072));
  AND2_X1   g0872(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n1063), .B1(new_n1072), .B2(new_n1073), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n1054), .B1(new_n1074), .B2(new_n751), .ZN(new_n1075));
  AOI22_X1  g0875(.A1(new_n1013), .A2(new_n748), .B1(new_n1045), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1014), .A2(new_n715), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1013), .A2(new_n744), .ZN(new_n1078));
  OAI21_X1  g0878(.A(new_n1076), .B1(new_n1077), .B2(new_n1078), .ZN(G393));
  INV_X1    g0879(.A(new_n715), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1010), .A2(new_n1016), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n1080), .B1(new_n1081), .B2(new_n1014), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n1082), .A2(new_n1019), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1010), .A2(new_n748), .A3(new_n1016), .ZN(new_n1084));
  OAI221_X1 g0884(.A(new_n755), .B1(new_n570), .B2(new_n209), .C1(new_n965), .C2(new_n239), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT117), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n828), .B1(new_n1085), .B2(new_n1086), .ZN(new_n1087));
  OAI21_X1  g0887(.A(new_n1087), .B1(new_n1086), .B2(new_n1085), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n268), .B1(new_n768), .B2(new_n365), .ZN(new_n1089));
  OAI22_X1  g0889(.A1(new_n780), .A2(new_n240), .B1(new_n781), .B2(new_n242), .ZN(new_n1090));
  AOI211_X1 g0890(.A(new_n1089), .B(new_n1090), .C1(G87), .C2(new_n837), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n777), .A2(G150), .B1(new_n831), .B2(G159), .ZN(new_n1092));
  XOR2_X1   g0892(.A(new_n1092), .B(KEYINPUT51), .Z(new_n1093));
  NAND2_X1  g0893(.A1(new_n784), .A2(G77), .ZN(new_n1094));
  NAND2_X1  g0894(.A1(new_n792), .A2(G143), .ZN(new_n1095));
  NAND4_X1  g0895(.A1(new_n1091), .A2(new_n1093), .A3(new_n1094), .A4(new_n1095), .ZN(new_n1096));
  AOI22_X1  g0896(.A1(new_n777), .A2(G317), .B1(new_n831), .B2(G311), .ZN(new_n1097));
  XOR2_X1   g0897(.A(new_n1097), .B(KEYINPUT52), .Z(new_n1098));
  AOI211_X1 g0898(.A(new_n268), .B(new_n775), .C1(G283), .C2(new_n985), .ZN(new_n1099));
  OAI211_X1 g0899(.A(new_n1098), .B(new_n1099), .C1(new_n805), .C2(new_n789), .ZN(new_n1100));
  AOI22_X1  g0900(.A1(new_n839), .A2(G116), .B1(new_n832), .B2(G294), .ZN(new_n1101));
  OAI21_X1  g0901(.A(new_n1101), .B1(new_n624), .B2(new_n780), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT118), .Z(new_n1103));
  OAI21_X1  g0903(.A(new_n1096), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  AOI21_X1  g0904(.A(new_n1088), .B1(new_n1104), .B2(new_n751), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1105), .B1(new_n1002), .B2(new_n994), .ZN(new_n1106));
  AND2_X1   g0906(.A1(new_n1084), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1083), .A2(new_n1107), .ZN(G390));
  AOI22_X1  g0908(.A1(new_n948), .A2(new_n917), .B1(new_n822), .B2(new_n914), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n868), .ZN(new_n1110));
  OAI211_X1 g0910(.A(new_n911), .B(new_n903), .C1(new_n1109), .C2(new_n1110), .ZN(new_n1111));
  AOI211_X1 g0911(.A(new_n710), .B(new_n819), .C1(new_n722), .C2(new_n736), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n930), .A2(new_n1112), .ZN(new_n1113));
  AOI211_X1 g0913(.A(new_n694), .B(new_n819), .C1(new_n741), .C2(new_n670), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(new_n913), .ZN(new_n1115));
  INV_X1    g0915(.A(new_n930), .ZN(new_n1116));
  OAI211_X1 g0916(.A(new_n950), .B(new_n868), .C1(new_n1115), .C2(new_n1116), .ZN(new_n1117));
  AND3_X1   g0917(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1113), .B1(new_n1111), .B2(new_n1117), .ZN(new_n1119));
  NOR2_X1   g0919(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n903), .A2(new_n911), .A3(new_n752), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n749), .B1(new_n851), .B2(new_n393), .ZN(new_n1122));
  NOR2_X1   g0922(.A1(new_n789), .A2(new_n525), .ZN(new_n1123));
  OAI221_X1 g0923(.A(new_n435), .B1(new_n768), .B2(new_n570), .C1(new_n507), .C2(new_n771), .ZN(new_n1124));
  NOR2_X1   g0924(.A1(new_n1123), .A2(new_n1124), .ZN(new_n1125));
  AOI22_X1  g0925(.A1(new_n777), .A2(G283), .B1(new_n837), .B2(G68), .ZN(new_n1126));
  OAI211_X1 g0926(.A(new_n1125), .B(new_n1126), .C1(new_n388), .C2(new_n780), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n1094), .B1(new_n445), .B2(new_n795), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n985), .A2(new_n1060), .ZN(new_n1129));
  XOR2_X1   g0929(.A(new_n1129), .B(KEYINPUT53), .Z(new_n1130));
  NAND2_X1  g0930(.A1(new_n792), .A2(G125), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(KEYINPUT54), .B(G143), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n268), .B1(new_n768), .B2(new_n1132), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1133), .B1(G132), .B2(new_n831), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1130), .A2(new_n1131), .A3(new_n1134), .ZN(new_n1135));
  AOI22_X1  g0935(.A1(new_n779), .A2(G137), .B1(new_n837), .B2(G50), .ZN(new_n1136));
  INV_X1    g0936(.A(G128), .ZN(new_n1137));
  OAI221_X1 g0937(.A(new_n1136), .B1(new_n1137), .B2(new_n799), .C1(new_n1055), .C2(new_n425), .ZN(new_n1138));
  OAI22_X1  g0938(.A1(new_n1127), .A2(new_n1128), .B1(new_n1135), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g0939(.A(new_n1122), .B1(new_n1139), .B2(new_n751), .ZN(new_n1140));
  AOI22_X1  g0940(.A1(new_n1120), .A2(new_n748), .B1(new_n1121), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n465), .A2(new_n488), .A3(new_n737), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n935), .A2(new_n686), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(new_n1143), .ZN(new_n1144));
  OAI211_X1 g0944(.A(G330), .B(new_n821), .C1(new_n938), .C2(new_n943), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n948), .A2(new_n1145), .A3(new_n917), .ZN(new_n1146));
  AND3_X1   g0946(.A1(new_n1113), .A2(new_n1115), .A3(new_n1146), .ZN(new_n1147));
  AOI22_X1  g0947(.A1(new_n1113), .A2(new_n1146), .B1(new_n822), .B2(new_n914), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1144), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n1149), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1111), .A2(new_n1117), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1145), .B1(new_n948), .B2(new_n917), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1151), .A2(new_n1152), .ZN(new_n1153));
  NAND3_X1  g0953(.A1(new_n1111), .A2(new_n1113), .A3(new_n1117), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n930), .A2(new_n1112), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n915), .B1(new_n1155), .B2(new_n1152), .ZN(new_n1156));
  NAND3_X1  g0956(.A1(new_n1113), .A2(new_n1115), .A3(new_n1146), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1143), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n1153), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1159));
  NAND3_X1  g0959(.A1(new_n1150), .A2(new_n1159), .A3(new_n715), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1141), .A2(new_n1160), .ZN(G378));
  NOR2_X1   g0961(.A1(new_n382), .A2(new_n692), .ZN(new_n1162));
  AND3_X1   g0962(.A1(new_n479), .A2(new_n480), .A3(new_n473), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n480), .B1(new_n479), .B2(new_n473), .ZN(new_n1164));
  OAI21_X1  g0964(.A(new_n485), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1165), .A2(KEYINPUT72), .ZN(new_n1166));
  NAND3_X1  g0966(.A1(new_n482), .A2(new_n477), .A3(new_n485), .ZN(new_n1167));
  AOI22_X1  g0967(.A1(new_n1166), .A2(new_n1167), .B1(KEYINPUT10), .B2(new_n475), .ZN(new_n1168));
  OAI21_X1  g0968(.A(new_n1162), .B1(new_n1168), .B2(new_n383), .ZN(new_n1169));
  INV_X1    g0969(.A(new_n383), .ZN(new_n1170));
  INV_X1    g0970(.A(new_n1162), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n488), .A2(new_n1170), .A3(new_n1171), .ZN(new_n1172));
  XNOR2_X1  g0972(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1173));
  AND3_X1   g0973(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1173), .B1(new_n1169), .B2(new_n1172), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND3_X1  g0976(.A1(new_n930), .A2(KEYINPUT40), .A3(new_n955), .ZN(new_n1177));
  INV_X1    g0977(.A(new_n888), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n901), .A2(new_n884), .ZN(new_n1179));
  INV_X1    g0979(.A(new_n899), .ZN(new_n1180));
  OAI21_X1  g0980(.A(KEYINPUT106), .B1(new_n884), .B2(new_n886), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n894), .A2(new_n895), .A3(new_n890), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n1179), .B1(new_n1180), .B2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g0984(.A(new_n1178), .B1(new_n1184), .B2(new_n908), .ZN(new_n1185));
  OAI21_X1  g0985(.A(G330), .B1(new_n1177), .B2(new_n1185), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1176), .B1(new_n1186), .B2(new_n953), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1173), .ZN(new_n1188));
  NOR3_X1   g0988(.A1(new_n1168), .A2(new_n383), .A3(new_n1162), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1171), .B1(new_n488), .B2(new_n1170), .ZN(new_n1190));
  OAI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NAND3_X1  g0991(.A1(new_n1169), .A2(new_n1172), .A3(new_n1173), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n1191), .A2(new_n1192), .ZN(new_n1193));
  NAND4_X1  g0993(.A1(new_n1193), .A2(new_n951), .A3(new_n958), .A4(G330), .ZN(new_n1194));
  AND3_X1   g0994(.A1(new_n1187), .A2(new_n1194), .A3(new_n934), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n934), .B1(new_n1187), .B2(new_n1194), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NOR2_X1   g0997(.A1(new_n1193), .A2(new_n753), .ZN(new_n1198));
  NOR2_X1   g0998(.A1(new_n268), .A2(G41), .ZN(new_n1199));
  AOI211_X1 g0999(.A(G50), .B(new_n1199), .C1(new_n261), .C2(new_n249), .ZN(new_n1200));
  OAI211_X1 g1000(.A(new_n261), .B(new_n249), .C1(new_n774), .C2(new_n425), .ZN(new_n1201));
  OAI22_X1  g1001(.A1(new_n771), .A2(new_n1137), .B1(new_n768), .B2(new_n834), .ZN(new_n1202));
  AOI21_X1  g1002(.A(new_n1202), .B1(G132), .B2(new_n779), .ZN(new_n1203));
  INV_X1    g1003(.A(new_n1132), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n777), .A2(G125), .B1(new_n985), .B2(new_n1204), .ZN(new_n1205));
  OAI211_X1 g1005(.A(new_n1203), .B(new_n1205), .C1(new_n1055), .C2(new_n366), .ZN(new_n1206));
  AND2_X1   g1006(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1207));
  AOI211_X1 g1007(.A(new_n1201), .B(new_n1207), .C1(G124), .C2(new_n792), .ZN(new_n1208));
  OR2_X1    g1008(.A1(new_n1206), .A2(KEYINPUT59), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1200), .B1(new_n1208), .B2(new_n1209), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n970), .B1(new_n507), .B2(new_n799), .ZN(new_n1211));
  XOR2_X1   g1011(.A(new_n1211), .B(KEYINPUT120), .Z(new_n1212));
  NAND2_X1  g1012(.A1(new_n831), .A2(G107), .ZN(new_n1213));
  OAI221_X1 g1013(.A(new_n1213), .B1(new_n395), .B2(new_n768), .C1(new_n780), .C2(new_n570), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1214), .B1(G58), .B2(new_n837), .ZN(new_n1215));
  OAI21_X1  g1015(.A(new_n1215), .B1(new_n801), .B2(new_n789), .ZN(new_n1216));
  OAI21_X1  g1016(.A(new_n1199), .B1(new_n323), .B2(new_n781), .ZN(new_n1217));
  XNOR2_X1  g1017(.A(new_n1217), .B(KEYINPUT119), .ZN(new_n1218));
  NOR3_X1   g1018(.A1(new_n1212), .A2(new_n1216), .A3(new_n1218), .ZN(new_n1219));
  XOR2_X1   g1019(.A(KEYINPUT121), .B(KEYINPUT58), .Z(new_n1220));
  INV_X1    g1020(.A(new_n1220), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1210), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1219), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1223), .A2(new_n1220), .ZN(new_n1224));
  OAI21_X1  g1024(.A(new_n751), .B1(new_n1222), .B2(new_n1224), .ZN(new_n1225));
  OAI211_X1 g1025(.A(new_n1225), .B(new_n749), .C1(G50), .C2(new_n851), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n1197), .A2(new_n747), .B1(new_n1198), .B2(new_n1226), .ZN(new_n1227));
  INV_X1    g1027(.A(KEYINPUT57), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1187), .A2(new_n1194), .ZN(new_n1229));
  INV_X1    g1029(.A(new_n934), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1229), .A2(new_n1230), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1187), .A2(new_n1194), .A3(new_n934), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n1228), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1159), .A2(new_n1144), .ZN(new_n1234));
  AOI21_X1  g1034(.A(new_n1080), .B1(new_n1233), .B2(new_n1234), .ZN(new_n1235));
  AOI21_X1  g1035(.A(new_n1143), .B1(new_n1120), .B2(new_n1158), .ZN(new_n1236));
  OAI21_X1  g1036(.A(new_n1228), .B1(new_n1236), .B2(new_n1197), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1227), .B1(new_n1235), .B2(new_n1237), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(G375));
  AOI21_X1  g1039(.A(new_n747), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1116), .A2(new_n752), .ZN(new_n1241));
  NOR2_X1   g1041(.A1(new_n799), .A2(new_n841), .ZN(new_n1242));
  NOR2_X1   g1042(.A1(new_n789), .A2(new_n1137), .ZN(new_n1243));
  OAI22_X1  g1043(.A1(new_n780), .A2(new_n1132), .B1(new_n769), .B2(new_n774), .ZN(new_n1244));
  OAI221_X1 g1044(.A(new_n268), .B1(new_n768), .B2(new_n366), .C1(new_n834), .C2(new_n771), .ZN(new_n1245));
  OR4_X1    g1045(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1245), .ZN(new_n1246));
  OAI22_X1  g1046(.A1(new_n1055), .A2(new_n240), .B1(new_n795), .B2(new_n425), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1056), .B1(new_n570), .B2(new_n795), .ZN(new_n1248));
  NOR2_X1   g1048(.A1(new_n789), .A2(new_n624), .ZN(new_n1249));
  OAI221_X1 g1049(.A(new_n435), .B1(new_n768), .B2(new_n388), .C1(new_n801), .C2(new_n771), .ZN(new_n1250));
  NOR2_X1   g1050(.A1(new_n1249), .A2(new_n1250), .ZN(new_n1251));
  AOI22_X1  g1051(.A1(new_n777), .A2(G294), .B1(new_n837), .B2(G77), .ZN(new_n1252));
  OAI211_X1 g1052(.A(new_n1251), .B(new_n1252), .C1(new_n507), .C2(new_n780), .ZN(new_n1253));
  OAI22_X1  g1053(.A1(new_n1246), .A2(new_n1247), .B1(new_n1248), .B2(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(new_n1254), .A2(new_n751), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n850), .A2(new_n242), .ZN(new_n1256));
  NAND4_X1  g1056(.A1(new_n1241), .A2(new_n749), .A3(new_n1255), .A4(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(new_n1257), .ZN(new_n1258));
  OAI21_X1  g1058(.A(KEYINPUT122), .B1(new_n1240), .B2(new_n1258), .ZN(new_n1259));
  OAI21_X1  g1059(.A(new_n748), .B1(new_n1147), .B2(new_n1148), .ZN(new_n1260));
  INV_X1    g1060(.A(KEYINPUT122), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1260), .A2(new_n1261), .A3(new_n1257), .ZN(new_n1262));
  NAND2_X1  g1062(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n999), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1156), .A2(new_n1143), .A3(new_n1157), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1149), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1263), .A2(new_n1266), .ZN(G381));
  INV_X1    g1067(.A(G387), .ZN(new_n1268));
  INV_X1    g1068(.A(G378), .ZN(new_n1269));
  OR2_X1    g1069(.A1(G393), .A2(G396), .ZN(new_n1270));
  NOR4_X1   g1070(.A1(G390), .A2(G384), .A3(G381), .A4(new_n1270), .ZN(new_n1271));
  NAND4_X1  g1071(.A1(new_n1268), .A2(new_n1269), .A3(new_n1238), .A4(new_n1271), .ZN(G407));
  NAND2_X1  g1072(.A1(new_n693), .A2(G213), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  NAND3_X1  g1074(.A1(new_n1238), .A2(new_n1269), .A3(new_n1274), .ZN(new_n1275));
  NAND3_X1  g1075(.A1(G407), .A2(G213), .A3(new_n1275), .ZN(G409));
  INV_X1    g1076(.A(KEYINPUT127), .ZN(new_n1277));
  OAI221_X1 g1077(.A(new_n1041), .B1(new_n1042), .B2(new_n1040), .C1(new_n1020), .C2(new_n748), .ZN(new_n1278));
  XNOR2_X1  g1078(.A(G393), .B(new_n813), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(G390), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1279), .ZN(new_n1281));
  NAND3_X1  g1081(.A1(new_n1083), .A2(new_n1107), .A3(new_n1281), .ZN(new_n1282));
  NAND4_X1  g1082(.A1(new_n1278), .A2(new_n1280), .A3(new_n998), .A4(new_n1282), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1280), .A2(new_n1282), .ZN(new_n1284));
  NAND2_X1  g1084(.A1(G387), .A2(new_n1284), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1198), .A2(new_n1226), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n1287), .B1(new_n1288), .B2(new_n748), .ZN(new_n1289));
  OAI21_X1  g1089(.A(KEYINPUT57), .B1(new_n1195), .B2(new_n1196), .ZN(new_n1290));
  OAI21_X1  g1090(.A(new_n715), .B1(new_n1290), .B2(new_n1236), .ZN(new_n1291));
  AOI21_X1  g1091(.A(KEYINPUT57), .B1(new_n1288), .B2(new_n1234), .ZN(new_n1292));
  OAI211_X1 g1092(.A(G378), .B(new_n1289), .C1(new_n1291), .C2(new_n1292), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1288), .A2(new_n1234), .A3(new_n1264), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1289), .A2(new_n1294), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1295), .A2(new_n1269), .ZN(new_n1296));
  NAND2_X1  g1096(.A1(new_n1293), .A2(new_n1296), .ZN(new_n1297));
  INV_X1    g1097(.A(KEYINPUT123), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(G384), .A2(new_n1298), .ZN(new_n1299));
  INV_X1    g1099(.A(new_n856), .ZN(new_n1300));
  NOR2_X1   g1100(.A1(new_n1300), .A2(new_n854), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(KEYINPUT123), .ZN(new_n1302));
  AND2_X1   g1102(.A1(new_n1259), .A2(new_n1262), .ZN(new_n1303));
  NAND4_X1  g1103(.A1(new_n1156), .A2(new_n1143), .A3(KEYINPUT60), .A4(new_n1157), .ZN(new_n1304));
  NAND2_X1  g1104(.A1(new_n1304), .A2(new_n715), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1149), .A2(KEYINPUT60), .ZN(new_n1306));
  AOI21_X1  g1106(.A(new_n1305), .B1(new_n1306), .B2(new_n1265), .ZN(new_n1307));
  OAI211_X1 g1107(.A(new_n1299), .B(new_n1302), .C1(new_n1303), .C2(new_n1307), .ZN(new_n1308));
  INV_X1    g1108(.A(KEYINPUT60), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1265), .B1(new_n1158), .B2(new_n1309), .ZN(new_n1310));
  NAND3_X1  g1110(.A1(new_n1310), .A2(new_n715), .A3(new_n1304), .ZN(new_n1311));
  NAND4_X1  g1111(.A1(new_n1311), .A2(new_n1263), .A3(KEYINPUT123), .A4(new_n1301), .ZN(new_n1312));
  NAND2_X1  g1112(.A1(new_n1308), .A2(new_n1312), .ZN(new_n1313));
  XNOR2_X1  g1113(.A(KEYINPUT125), .B(KEYINPUT62), .ZN(new_n1314));
  AND4_X1   g1114(.A1(new_n1273), .A2(new_n1297), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1315));
  XNOR2_X1  g1115(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n1316));
  INV_X1    g1116(.A(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1274), .B1(new_n1293), .B2(new_n1296), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1274), .A2(G2897), .ZN(new_n1319));
  AND3_X1   g1119(.A1(new_n1308), .A2(new_n1312), .A3(new_n1319), .ZN(new_n1320));
  AOI21_X1  g1120(.A(new_n1319), .B1(new_n1308), .B2(new_n1312), .ZN(new_n1321));
  NOR2_X1   g1121(.A1(new_n1320), .A2(new_n1321), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1317), .B1(new_n1318), .B2(new_n1322), .ZN(new_n1323));
  NOR2_X1   g1123(.A1(new_n1315), .A2(new_n1323), .ZN(new_n1324));
  NAND3_X1  g1124(.A1(new_n1297), .A2(new_n1273), .A3(new_n1313), .ZN(new_n1325));
  INV_X1    g1125(.A(KEYINPUT62), .ZN(new_n1326));
  NOR2_X1   g1126(.A1(new_n1326), .A2(KEYINPUT125), .ZN(new_n1327));
  NAND2_X1  g1127(.A1(new_n1325), .A2(new_n1327), .ZN(new_n1328));
  AOI21_X1  g1128(.A(KEYINPUT126), .B1(new_n1324), .B2(new_n1328), .ZN(new_n1329));
  NAND2_X1  g1129(.A1(new_n1297), .A2(new_n1273), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1321), .ZN(new_n1331));
  NAND3_X1  g1131(.A1(new_n1308), .A2(new_n1312), .A3(new_n1319), .ZN(new_n1332));
  NAND2_X1  g1132(.A1(new_n1331), .A2(new_n1332), .ZN(new_n1333));
  AOI21_X1  g1133(.A(new_n1316), .B1(new_n1330), .B2(new_n1333), .ZN(new_n1334));
  NAND4_X1  g1134(.A1(new_n1297), .A2(new_n1273), .A3(new_n1313), .A4(new_n1314), .ZN(new_n1335));
  AND4_X1   g1135(.A1(KEYINPUT126), .A2(new_n1334), .A3(new_n1328), .A4(new_n1335), .ZN(new_n1336));
  OAI21_X1  g1136(.A(new_n1286), .B1(new_n1329), .B2(new_n1336), .ZN(new_n1337));
  INV_X1    g1137(.A(KEYINPUT61), .ZN(new_n1338));
  OAI21_X1  g1138(.A(new_n1338), .B1(new_n1318), .B2(new_n1322), .ZN(new_n1339));
  INV_X1    g1139(.A(new_n1325), .ZN(new_n1340));
  AOI21_X1  g1140(.A(new_n1339), .B1(new_n1340), .B2(KEYINPUT63), .ZN(new_n1341));
  OR2_X1    g1141(.A1(new_n1340), .A2(KEYINPUT63), .ZN(new_n1342));
  AOI21_X1  g1142(.A(new_n1286), .B1(new_n1341), .B2(new_n1342), .ZN(new_n1343));
  INV_X1    g1143(.A(new_n1343), .ZN(new_n1344));
  AOI21_X1  g1144(.A(new_n1277), .B1(new_n1337), .B2(new_n1344), .ZN(new_n1345));
  AND2_X1   g1145(.A1(new_n1283), .A2(new_n1285), .ZN(new_n1346));
  INV_X1    g1146(.A(KEYINPUT126), .ZN(new_n1347));
  AOI21_X1  g1147(.A(G378), .B1(new_n1289), .B2(new_n1294), .ZN(new_n1348));
  AOI21_X1  g1148(.A(new_n1348), .B1(new_n1238), .B2(G378), .ZN(new_n1349));
  OAI21_X1  g1149(.A(new_n1333), .B1(new_n1349), .B2(new_n1274), .ZN(new_n1350));
  NAND3_X1  g1150(.A1(new_n1350), .A2(new_n1335), .A3(new_n1317), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1327), .ZN(new_n1352));
  AOI21_X1  g1152(.A(new_n1352), .B1(new_n1318), .B2(new_n1313), .ZN(new_n1353));
  OAI21_X1  g1153(.A(new_n1347), .B1(new_n1351), .B2(new_n1353), .ZN(new_n1354));
  NAND4_X1  g1154(.A1(new_n1334), .A2(new_n1328), .A3(KEYINPUT126), .A4(new_n1335), .ZN(new_n1355));
  AOI21_X1  g1155(.A(new_n1346), .B1(new_n1354), .B2(new_n1355), .ZN(new_n1356));
  NOR3_X1   g1156(.A1(new_n1356), .A2(KEYINPUT127), .A3(new_n1343), .ZN(new_n1357));
  NOR2_X1   g1157(.A1(new_n1345), .A2(new_n1357), .ZN(G405));
  NAND2_X1  g1158(.A1(G375), .A2(new_n1269), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1359), .A2(new_n1293), .ZN(new_n1360));
  XNOR2_X1  g1160(.A(new_n1360), .B(new_n1313), .ZN(new_n1361));
  XNOR2_X1  g1161(.A(new_n1361), .B(new_n1286), .ZN(G402));
endmodule


