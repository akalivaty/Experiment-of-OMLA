

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333,
         n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344,
         n345, n346, n347, n348, n349, n350, n351, n352, n353, n354, n355,
         n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, n366,
         n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377,
         n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
         n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443,
         n444, n445, n446, n447, n448, n449, n450, n451, n452, n453, n454,
         n455, n456, n457, n458, n459, n460, n461, n462, n463, n464, n465,
         n466, n467, n468, n469, n470, n471, n472, n473, n474, n475, n476,
         n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, n487,
         n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
         n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509,
         n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584;

  XNOR2_X1 U322 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U323 ( .A(n456), .B(KEYINPUT38), .ZN(n476) );
  XOR2_X1 U324 ( .A(n550), .B(KEYINPUT28), .Z(n521) );
  XOR2_X1 U325 ( .A(G64GAT), .B(G92GAT), .Z(n290) );
  XOR2_X1 U326 ( .A(n420), .B(n419), .Z(n495) );
  INV_X1 U327 ( .A(KEYINPUT102), .ZN(n405) );
  XNOR2_X1 U328 ( .A(n545), .B(n421), .ZN(n443) );
  XNOR2_X1 U329 ( .A(n406), .B(n405), .ZN(n407) );
  INV_X1 U330 ( .A(KEYINPUT108), .ZN(n452) );
  XNOR2_X1 U331 ( .A(n408), .B(n407), .ZN(n409) );
  XNOR2_X1 U332 ( .A(n325), .B(n324), .ZN(n326) );
  XNOR2_X1 U333 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U334 ( .A(n327), .B(n326), .ZN(n574) );
  XNOR2_X1 U335 ( .A(n455), .B(n454), .ZN(n491) );
  XNOR2_X1 U336 ( .A(n414), .B(n413), .ZN(n420) );
  NOR2_X1 U337 ( .A1(n553), .A2(n552), .ZN(n565) );
  XNOR2_X1 U338 ( .A(n478), .B(KEYINPUT41), .ZN(n535) );
  INV_X1 U339 ( .A(G43GAT), .ZN(n457) );
  XNOR2_X1 U340 ( .A(n458), .B(n457), .ZN(n459) );
  XNOR2_X1 U341 ( .A(n460), .B(n459), .ZN(G1330GAT) );
  XOR2_X1 U342 ( .A(G127GAT), .B(KEYINPUT0), .Z(n292) );
  XNOR2_X1 U343 ( .A(G134GAT), .B(KEYINPUT88), .ZN(n291) );
  XNOR2_X1 U344 ( .A(n292), .B(n291), .ZN(n394) );
  XOR2_X1 U345 ( .A(n394), .B(G99GAT), .Z(n294) );
  NAND2_X1 U346 ( .A1(G227GAT), .A2(G233GAT), .ZN(n293) );
  XNOR2_X1 U347 ( .A(n294), .B(n293), .ZN(n298) );
  XOR2_X1 U348 ( .A(KEYINPUT91), .B(KEYINPUT20), .Z(n296) );
  XNOR2_X1 U349 ( .A(KEYINPUT90), .B(KEYINPUT89), .ZN(n295) );
  XNOR2_X1 U350 ( .A(n296), .B(n295), .ZN(n297) );
  XOR2_X1 U351 ( .A(n298), .B(n297), .Z(n304) );
  XNOR2_X1 U352 ( .A(KEYINPUT18), .B(KEYINPUT92), .ZN(n299) );
  XNOR2_X1 U353 ( .A(n299), .B(KEYINPUT17), .ZN(n300) );
  XOR2_X1 U354 ( .A(n300), .B(KEYINPUT19), .Z(n302) );
  XNOR2_X1 U355 ( .A(G183GAT), .B(G190GAT), .ZN(n301) );
  XNOR2_X1 U356 ( .A(n302), .B(n301), .ZN(n412) );
  XNOR2_X1 U357 ( .A(G43GAT), .B(n412), .ZN(n303) );
  XNOR2_X1 U358 ( .A(n304), .B(n303), .ZN(n312) );
  XOR2_X1 U359 ( .A(G176GAT), .B(G120GAT), .Z(n306) );
  XNOR2_X1 U360 ( .A(G169GAT), .B(KEYINPUT93), .ZN(n305) );
  XNOR2_X1 U361 ( .A(n306), .B(n305), .ZN(n310) );
  XOR2_X1 U362 ( .A(KEYINPUT65), .B(G71GAT), .Z(n308) );
  XNOR2_X1 U363 ( .A(G113GAT), .B(G15GAT), .ZN(n307) );
  XNOR2_X1 U364 ( .A(n308), .B(n307), .ZN(n309) );
  XOR2_X1 U365 ( .A(n310), .B(n309), .Z(n311) );
  XNOR2_X1 U366 ( .A(n312), .B(n311), .ZN(n553) );
  INV_X1 U367 ( .A(n553), .ZN(n518) );
  XOR2_X1 U368 ( .A(KEYINPUT75), .B(KEYINPUT78), .Z(n314) );
  NAND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n315) );
  XOR2_X1 U371 ( .A(n315), .B(KEYINPUT32), .Z(n319) );
  XNOR2_X1 U372 ( .A(G176GAT), .B(G204GAT), .ZN(n316) );
  XNOR2_X1 U373 ( .A(n290), .B(n316), .ZN(n408) );
  XNOR2_X1 U374 ( .A(G71GAT), .B(KEYINPUT13), .ZN(n317) );
  XNOR2_X1 U375 ( .A(n317), .B(KEYINPUT74), .ZN(n378) );
  XNOR2_X1 U376 ( .A(n408), .B(n378), .ZN(n318) );
  XNOR2_X1 U377 ( .A(n319), .B(n318), .ZN(n320) );
  XOR2_X1 U378 ( .A(n320), .B(KEYINPUT33), .Z(n327) );
  XOR2_X1 U379 ( .A(G78GAT), .B(G148GAT), .Z(n322) );
  XNOR2_X1 U380 ( .A(G106GAT), .B(KEYINPUT76), .ZN(n321) );
  XNOR2_X1 U381 ( .A(n322), .B(n321), .ZN(n431) );
  XNOR2_X1 U382 ( .A(G99GAT), .B(G85GAT), .ZN(n323) );
  XOR2_X1 U383 ( .A(n323), .B(KEYINPUT77), .Z(n358) );
  XNOR2_X1 U384 ( .A(n431), .B(n358), .ZN(n325) );
  XOR2_X1 U385 ( .A(G120GAT), .B(G57GAT), .Z(n388) );
  XNOR2_X1 U386 ( .A(n388), .B(KEYINPUT31), .ZN(n324) );
  INV_X1 U387 ( .A(n574), .ZN(n478) );
  XOR2_X1 U388 ( .A(KEYINPUT29), .B(KEYINPUT67), .Z(n329) );
  XNOR2_X1 U389 ( .A(KEYINPUT30), .B(KEYINPUT68), .ZN(n328) );
  XNOR2_X1 U390 ( .A(n329), .B(n328), .ZN(n340) );
  XOR2_X1 U391 ( .A(KEYINPUT72), .B(KEYINPUT69), .Z(n331) );
  XOR2_X1 U392 ( .A(G113GAT), .B(G1GAT), .Z(n389) );
  XOR2_X1 U393 ( .A(G169GAT), .B(G8GAT), .Z(n410) );
  XNOR2_X1 U394 ( .A(n389), .B(n410), .ZN(n330) );
  XNOR2_X1 U395 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U396 ( .A(n332), .B(G15GAT), .Z(n338) );
  XNOR2_X1 U397 ( .A(G50GAT), .B(G22GAT), .ZN(n333) );
  XNOR2_X1 U398 ( .A(n333), .B(G141GAT), .ZN(n434) );
  XOR2_X1 U399 ( .A(n434), .B(KEYINPUT70), .Z(n335) );
  NAND2_X1 U400 ( .A1(G229GAT), .A2(G233GAT), .ZN(n334) );
  XNOR2_X1 U401 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U402 ( .A(n336), .B(G197GAT), .ZN(n337) );
  XNOR2_X1 U403 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U404 ( .A(n340), .B(n339), .ZN(n345) );
  XOR2_X1 U405 ( .A(G29GAT), .B(KEYINPUT7), .Z(n342) );
  XNOR2_X1 U406 ( .A(G43GAT), .B(G36GAT), .ZN(n341) );
  XNOR2_X1 U407 ( .A(n342), .B(n341), .ZN(n344) );
  XOR2_X1 U408 ( .A(KEYINPUT71), .B(KEYINPUT8), .Z(n343) );
  XNOR2_X1 U409 ( .A(n344), .B(n343), .ZN(n347) );
  XOR2_X1 U410 ( .A(n345), .B(n347), .Z(n570) );
  INV_X1 U411 ( .A(n570), .ZN(n533) );
  XOR2_X1 U412 ( .A(KEYINPUT73), .B(n533), .Z(n554) );
  INV_X1 U413 ( .A(n554), .ZN(n510) );
  NOR2_X1 U414 ( .A1(n478), .A2(n510), .ZN(n346) );
  XNOR2_X1 U415 ( .A(n346), .B(KEYINPUT79), .ZN(n465) );
  INV_X1 U416 ( .A(n347), .ZN(n351) );
  XOR2_X1 U417 ( .A(KEYINPUT10), .B(KEYINPUT11), .Z(n349) );
  XNOR2_X1 U418 ( .A(G50GAT), .B(KEYINPUT9), .ZN(n348) );
  XNOR2_X1 U419 ( .A(n349), .B(n348), .ZN(n350) );
  XNOR2_X1 U420 ( .A(n351), .B(n350), .ZN(n365) );
  XOR2_X1 U421 ( .A(KEYINPUT82), .B(KEYINPUT81), .Z(n353) );
  XNOR2_X1 U422 ( .A(G134GAT), .B(KEYINPUT80), .ZN(n352) );
  XNOR2_X1 U423 ( .A(n353), .B(n352), .ZN(n357) );
  XOR2_X1 U424 ( .A(KEYINPUT66), .B(G92GAT), .Z(n355) );
  XNOR2_X1 U425 ( .A(G190GAT), .B(G106GAT), .ZN(n354) );
  XNOR2_X1 U426 ( .A(n355), .B(n354), .ZN(n356) );
  XOR2_X1 U427 ( .A(n357), .B(n356), .Z(n363) );
  XNOR2_X1 U428 ( .A(n358), .B(G162GAT), .ZN(n360) );
  NAND2_X1 U429 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U430 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U431 ( .A(G218GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U432 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U433 ( .A(n365), .B(n364), .ZN(n527) );
  XNOR2_X1 U434 ( .A(KEYINPUT36), .B(n527), .ZN(n581) );
  XOR2_X1 U435 ( .A(KEYINPUT84), .B(KEYINPUT12), .Z(n367) );
  XNOR2_X1 U436 ( .A(G64GAT), .B(KEYINPUT85), .ZN(n366) );
  XNOR2_X1 U437 ( .A(n367), .B(n366), .ZN(n371) );
  XOR2_X1 U438 ( .A(KEYINPUT86), .B(KEYINPUT14), .Z(n369) );
  XNOR2_X1 U439 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n368) );
  XNOR2_X1 U440 ( .A(n369), .B(n368), .ZN(n370) );
  XNOR2_X1 U441 ( .A(n371), .B(n370), .ZN(n385) );
  XOR2_X1 U442 ( .A(G155GAT), .B(G127GAT), .Z(n373) );
  XNOR2_X1 U443 ( .A(G22GAT), .B(G15GAT), .ZN(n372) );
  XNOR2_X1 U444 ( .A(n373), .B(n372), .ZN(n377) );
  XOR2_X1 U445 ( .A(G57GAT), .B(G183GAT), .Z(n375) );
  XNOR2_X1 U446 ( .A(G1GAT), .B(G8GAT), .ZN(n374) );
  XNOR2_X1 U447 ( .A(n375), .B(n374), .ZN(n376) );
  XOR2_X1 U448 ( .A(n377), .B(n376), .Z(n383) );
  XOR2_X1 U449 ( .A(n378), .B(G78GAT), .Z(n380) );
  NAND2_X1 U450 ( .A1(G231GAT), .A2(G233GAT), .ZN(n379) );
  XNOR2_X1 U451 ( .A(n380), .B(n379), .ZN(n381) );
  XNOR2_X1 U452 ( .A(G211GAT), .B(n381), .ZN(n382) );
  XNOR2_X1 U453 ( .A(n383), .B(n382), .ZN(n384) );
  XNOR2_X1 U454 ( .A(n385), .B(n384), .ZN(n578) );
  XOR2_X1 U455 ( .A(KEYINPUT100), .B(KEYINPUT4), .Z(n387) );
  XNOR2_X1 U456 ( .A(G141GAT), .B(G148GAT), .ZN(n386) );
  XNOR2_X1 U457 ( .A(n387), .B(n386), .ZN(n404) );
  XOR2_X1 U458 ( .A(G85GAT), .B(n388), .Z(n391) );
  XNOR2_X1 U459 ( .A(G29GAT), .B(n389), .ZN(n390) );
  XNOR2_X1 U460 ( .A(n391), .B(n390), .ZN(n400) );
  XOR2_X1 U461 ( .A(G155GAT), .B(KEYINPUT3), .Z(n393) );
  XNOR2_X1 U462 ( .A(G162GAT), .B(KEYINPUT2), .ZN(n392) );
  XNOR2_X1 U463 ( .A(n393), .B(n392), .ZN(n422) );
  XNOR2_X1 U464 ( .A(n394), .B(n422), .ZN(n398) );
  XOR2_X1 U465 ( .A(KEYINPUT1), .B(KEYINPUT5), .Z(n396) );
  XNOR2_X1 U466 ( .A(KEYINPUT99), .B(KEYINPUT6), .ZN(n395) );
  XNOR2_X1 U467 ( .A(n396), .B(n395), .ZN(n397) );
  XNOR2_X1 U468 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U469 ( .A(n400), .B(n399), .Z(n402) );
  NAND2_X1 U470 ( .A1(G225GAT), .A2(G233GAT), .ZN(n401) );
  XNOR2_X1 U471 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U472 ( .A(n404), .B(n403), .ZN(n447) );
  XNOR2_X1 U473 ( .A(KEYINPUT101), .B(n447), .ZN(n549) );
  NAND2_X1 U474 ( .A1(G226GAT), .A2(G233GAT), .ZN(n406) );
  XOR2_X1 U475 ( .A(n409), .B(KEYINPUT103), .Z(n414) );
  XNOR2_X1 U476 ( .A(G36GAT), .B(n410), .ZN(n411) );
  XNOR2_X1 U477 ( .A(G211GAT), .B(KEYINPUT96), .ZN(n415) );
  XNOR2_X1 U478 ( .A(n415), .B(KEYINPUT21), .ZN(n416) );
  XOR2_X1 U479 ( .A(n416), .B(KEYINPUT97), .Z(n418) );
  XNOR2_X1 U480 ( .A(G197GAT), .B(G218GAT), .ZN(n417) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n433) );
  INV_X1 U482 ( .A(n433), .ZN(n419) );
  INV_X1 U483 ( .A(n495), .ZN(n545) );
  XOR2_X1 U484 ( .A(KEYINPUT27), .B(KEYINPUT104), .Z(n421) );
  NAND2_X1 U485 ( .A1(n549), .A2(n443), .ZN(n516) );
  XOR2_X1 U486 ( .A(KEYINPUT22), .B(KEYINPUT24), .Z(n424) );
  XNOR2_X1 U487 ( .A(KEYINPUT23), .B(n422), .ZN(n423) );
  XNOR2_X1 U488 ( .A(n424), .B(n423), .ZN(n425) );
  XOR2_X1 U489 ( .A(n425), .B(KEYINPUT95), .Z(n430) );
  XOR2_X1 U490 ( .A(KEYINPUT94), .B(KEYINPUT98), .Z(n427) );
  NAND2_X1 U491 ( .A1(G228GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U492 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U493 ( .A(G204GAT), .B(n428), .ZN(n429) );
  XNOR2_X1 U494 ( .A(n430), .B(n429), .ZN(n432) );
  XOR2_X1 U495 ( .A(n432), .B(n431), .Z(n436) );
  XNOR2_X1 U496 ( .A(n434), .B(n433), .ZN(n435) );
  XNOR2_X1 U497 ( .A(n436), .B(n435), .ZN(n550) );
  NOR2_X1 U498 ( .A1(n516), .A2(n521), .ZN(n437) );
  NAND2_X1 U499 ( .A1(n437), .A2(n553), .ZN(n438) );
  XOR2_X1 U500 ( .A(KEYINPUT105), .B(n438), .Z(n450) );
  NAND2_X1 U501 ( .A1(n518), .A2(n495), .ZN(n439) );
  NAND2_X1 U502 ( .A1(n550), .A2(n439), .ZN(n440) );
  XOR2_X1 U503 ( .A(KEYINPUT25), .B(n440), .Z(n445) );
  XNOR2_X1 U504 ( .A(KEYINPUT106), .B(KEYINPUT26), .ZN(n442) );
  NOR2_X1 U505 ( .A1(n518), .A2(n550), .ZN(n441) );
  XNOR2_X1 U506 ( .A(n442), .B(n441), .ZN(n568) );
  NAND2_X1 U507 ( .A1(n443), .A2(n568), .ZN(n444) );
  NAND2_X1 U508 ( .A1(n445), .A2(n444), .ZN(n446) );
  XOR2_X1 U509 ( .A(KEYINPUT107), .B(n446), .Z(n448) );
  NAND2_X1 U510 ( .A1(n448), .A2(n447), .ZN(n449) );
  NAND2_X1 U511 ( .A1(n450), .A2(n449), .ZN(n463) );
  NAND2_X1 U512 ( .A1(n578), .A2(n463), .ZN(n451) );
  NOR2_X1 U513 ( .A1(n581), .A2(n451), .ZN(n455) );
  XNOR2_X1 U514 ( .A(KEYINPUT109), .B(KEYINPUT37), .ZN(n453) );
  NOR2_X1 U515 ( .A1(n465), .A2(n491), .ZN(n456) );
  NAND2_X1 U516 ( .A1(n518), .A2(n476), .ZN(n460) );
  XOR2_X1 U517 ( .A(KEYINPUT40), .B(KEYINPUT110), .Z(n458) );
  INV_X1 U518 ( .A(n578), .ZN(n562) );
  NAND2_X1 U519 ( .A1(n562), .A2(n527), .ZN(n461) );
  XNOR2_X1 U520 ( .A(n461), .B(KEYINPUT16), .ZN(n462) );
  XNOR2_X1 U521 ( .A(n462), .B(KEYINPUT87), .ZN(n464) );
  NAND2_X1 U522 ( .A1(n464), .A2(n463), .ZN(n479) );
  NOR2_X1 U523 ( .A1(n465), .A2(n479), .ZN(n471) );
  NAND2_X1 U524 ( .A1(n471), .A2(n549), .ZN(n466) );
  XNOR2_X1 U525 ( .A(n466), .B(KEYINPUT34), .ZN(n467) );
  XNOR2_X1 U526 ( .A(G1GAT), .B(n467), .ZN(G1324GAT) );
  NAND2_X1 U527 ( .A1(n471), .A2(n495), .ZN(n468) );
  XNOR2_X1 U528 ( .A(n468), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U529 ( .A(G15GAT), .B(KEYINPUT35), .Z(n470) );
  NAND2_X1 U530 ( .A1(n471), .A2(n518), .ZN(n469) );
  XNOR2_X1 U531 ( .A(n470), .B(n469), .ZN(G1326GAT) );
  NAND2_X1 U532 ( .A1(n471), .A2(n521), .ZN(n472) );
  XNOR2_X1 U533 ( .A(n472), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U534 ( .A(G29GAT), .B(KEYINPUT39), .Z(n474) );
  NAND2_X1 U535 ( .A1(n549), .A2(n476), .ZN(n473) );
  XNOR2_X1 U536 ( .A(n474), .B(n473), .ZN(G1328GAT) );
  NAND2_X1 U537 ( .A1(n476), .A2(n495), .ZN(n475) );
  XNOR2_X1 U538 ( .A(n475), .B(G36GAT), .ZN(G1329GAT) );
  NAND2_X1 U539 ( .A1(n476), .A2(n521), .ZN(n477) );
  XNOR2_X1 U540 ( .A(n477), .B(G50GAT), .ZN(G1331GAT) );
  XOR2_X1 U541 ( .A(KEYINPUT112), .B(KEYINPUT42), .Z(n481) );
  XNOR2_X1 U542 ( .A(KEYINPUT111), .B(n535), .ZN(n557) );
  NAND2_X1 U543 ( .A1(n570), .A2(n557), .ZN(n490) );
  NOR2_X1 U544 ( .A1(n490), .A2(n479), .ZN(n486) );
  NAND2_X1 U545 ( .A1(n486), .A2(n549), .ZN(n480) );
  XNOR2_X1 U546 ( .A(n481), .B(n480), .ZN(n482) );
  XOR2_X1 U547 ( .A(G57GAT), .B(n482), .Z(G1332GAT) );
  XOR2_X1 U548 ( .A(G64GAT), .B(KEYINPUT113), .Z(n484) );
  NAND2_X1 U549 ( .A1(n486), .A2(n495), .ZN(n483) );
  XNOR2_X1 U550 ( .A(n484), .B(n483), .ZN(G1333GAT) );
  NAND2_X1 U551 ( .A1(n486), .A2(n518), .ZN(n485) );
  XNOR2_X1 U552 ( .A(n485), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U553 ( .A(KEYINPUT43), .B(KEYINPUT114), .Z(n488) );
  NAND2_X1 U554 ( .A1(n486), .A2(n521), .ZN(n487) );
  XNOR2_X1 U555 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U556 ( .A(G78GAT), .B(n489), .ZN(G1335GAT) );
  XOR2_X1 U557 ( .A(KEYINPUT115), .B(KEYINPUT116), .Z(n493) );
  NOR2_X1 U558 ( .A1(n491), .A2(n490), .ZN(n499) );
  NAND2_X1 U559 ( .A1(n499), .A2(n549), .ZN(n492) );
  XNOR2_X1 U560 ( .A(n493), .B(n492), .ZN(n494) );
  XNOR2_X1 U561 ( .A(G85GAT), .B(n494), .ZN(G1336GAT) );
  XOR2_X1 U562 ( .A(G92GAT), .B(KEYINPUT117), .Z(n497) );
  NAND2_X1 U563 ( .A1(n499), .A2(n495), .ZN(n496) );
  XNOR2_X1 U564 ( .A(n497), .B(n496), .ZN(G1337GAT) );
  NAND2_X1 U565 ( .A1(n499), .A2(n518), .ZN(n498) );
  XNOR2_X1 U566 ( .A(n498), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U567 ( .A1(n499), .A2(n521), .ZN(n500) );
  XNOR2_X1 U568 ( .A(n500), .B(KEYINPUT44), .ZN(n501) );
  XNOR2_X1 U569 ( .A(G106GAT), .B(n501), .ZN(G1339GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT48), .B(KEYINPUT64), .Z(n515) );
  XOR2_X1 U571 ( .A(KEYINPUT47), .B(KEYINPUT118), .Z(n506) );
  NOR2_X1 U572 ( .A1(n570), .A2(n535), .ZN(n502) );
  XNOR2_X1 U573 ( .A(n502), .B(KEYINPUT46), .ZN(n503) );
  NOR2_X1 U574 ( .A1(n562), .A2(n503), .ZN(n504) );
  NAND2_X1 U575 ( .A1(n504), .A2(n527), .ZN(n505) );
  XNOR2_X1 U576 ( .A(n506), .B(n505), .ZN(n513) );
  NOR2_X1 U577 ( .A1(n578), .A2(n581), .ZN(n507) );
  XNOR2_X1 U578 ( .A(n507), .B(KEYINPUT45), .ZN(n508) );
  NAND2_X1 U579 ( .A1(n508), .A2(n574), .ZN(n509) );
  XNOR2_X1 U580 ( .A(KEYINPUT119), .B(n509), .ZN(n511) );
  NAND2_X1 U581 ( .A1(n511), .A2(n510), .ZN(n512) );
  NAND2_X1 U582 ( .A1(n513), .A2(n512), .ZN(n514) );
  XNOR2_X1 U583 ( .A(n515), .B(n514), .ZN(n544) );
  NOR2_X1 U584 ( .A1(n544), .A2(n516), .ZN(n517) );
  XNOR2_X1 U585 ( .A(KEYINPUT120), .B(n517), .ZN(n532) );
  AND2_X1 U586 ( .A1(n532), .A2(n518), .ZN(n519) );
  XNOR2_X1 U587 ( .A(n519), .B(KEYINPUT121), .ZN(n520) );
  NOR2_X1 U588 ( .A1(n521), .A2(n520), .ZN(n528) );
  NAND2_X1 U589 ( .A1(n554), .A2(n528), .ZN(n522) );
  XNOR2_X1 U590 ( .A(n522), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U591 ( .A(G120GAT), .B(KEYINPUT49), .Z(n524) );
  NAND2_X1 U592 ( .A1(n528), .A2(n557), .ZN(n523) );
  XNOR2_X1 U593 ( .A(n524), .B(n523), .ZN(G1341GAT) );
  NAND2_X1 U594 ( .A1(n562), .A2(n528), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n525), .B(KEYINPUT50), .ZN(n526) );
  XNOR2_X1 U596 ( .A(G127GAT), .B(n526), .ZN(G1342GAT) );
  XOR2_X1 U597 ( .A(KEYINPUT122), .B(KEYINPUT51), .Z(n530) );
  INV_X1 U598 ( .A(n527), .ZN(n564) );
  NAND2_X1 U599 ( .A1(n528), .A2(n564), .ZN(n529) );
  XNOR2_X1 U600 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U601 ( .A(G134GAT), .B(n531), .ZN(G1343GAT) );
  NAND2_X1 U602 ( .A1(n532), .A2(n568), .ZN(n536) );
  INV_X1 U603 ( .A(n536), .ZN(n542) );
  NAND2_X1 U604 ( .A1(n542), .A2(n533), .ZN(n534) );
  XNOR2_X1 U605 ( .A(G141GAT), .B(n534), .ZN(G1344GAT) );
  NOR2_X1 U606 ( .A1(n536), .A2(n535), .ZN(n540) );
  XOR2_X1 U607 ( .A(KEYINPUT123), .B(KEYINPUT52), .Z(n538) );
  XNOR2_X1 U608 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n537) );
  XNOR2_X1 U609 ( .A(n538), .B(n537), .ZN(n539) );
  XNOR2_X1 U610 ( .A(n540), .B(n539), .ZN(G1345GAT) );
  NAND2_X1 U611 ( .A1(n562), .A2(n542), .ZN(n541) );
  XNOR2_X1 U612 ( .A(n541), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U613 ( .A1(n564), .A2(n542), .ZN(n543) );
  XNOR2_X1 U614 ( .A(n543), .B(G162GAT), .ZN(G1347GAT) );
  XNOR2_X1 U615 ( .A(G169GAT), .B(KEYINPUT124), .ZN(n556) );
  INV_X1 U616 ( .A(n544), .ZN(n546) );
  NAND2_X1 U617 ( .A1(n546), .A2(n495), .ZN(n547) );
  XNOR2_X1 U618 ( .A(n547), .B(KEYINPUT54), .ZN(n548) );
  NOR2_X1 U619 ( .A1(n549), .A2(n548), .ZN(n569) );
  NAND2_X1 U620 ( .A1(n550), .A2(n569), .ZN(n551) );
  XOR2_X1 U621 ( .A(KEYINPUT55), .B(n551), .Z(n552) );
  NAND2_X1 U622 ( .A1(n565), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(G1348GAT) );
  XOR2_X1 U624 ( .A(G176GAT), .B(KEYINPUT125), .Z(n559) );
  NAND2_X1 U625 ( .A1(n557), .A2(n565), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(n561) );
  XOR2_X1 U627 ( .A(KEYINPUT56), .B(KEYINPUT57), .Z(n560) );
  XNOR2_X1 U628 ( .A(n561), .B(n560), .ZN(G1349GAT) );
  NAND2_X1 U629 ( .A1(n562), .A2(n565), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G183GAT), .ZN(G1350GAT) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(KEYINPUT58), .ZN(n567) );
  NAND2_X1 U632 ( .A1(n565), .A2(n564), .ZN(n566) );
  XNOR2_X1 U633 ( .A(n567), .B(n566), .ZN(G1351GAT) );
  NAND2_X1 U634 ( .A1(n569), .A2(n568), .ZN(n580) );
  NOR2_X1 U635 ( .A1(n570), .A2(n580), .ZN(n572) );
  XNOR2_X1 U636 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(n573) );
  XNOR2_X1 U638 ( .A(G197GAT), .B(n573), .ZN(G1352GAT) );
  NOR2_X1 U639 ( .A1(n574), .A2(n580), .ZN(n576) );
  XNOR2_X1 U640 ( .A(KEYINPUT126), .B(KEYINPUT61), .ZN(n575) );
  XNOR2_X1 U641 ( .A(n576), .B(n575), .ZN(n577) );
  XNOR2_X1 U642 ( .A(G204GAT), .B(n577), .ZN(G1353GAT) );
  NOR2_X1 U643 ( .A1(n578), .A2(n580), .ZN(n579) );
  XOR2_X1 U644 ( .A(G211GAT), .B(n579), .Z(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n583) );
  XNOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

