//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 0 1 0 1 1 1 0 0 0 1 0 1 0 1 0 0 1 0 0 1 0 0 0 1 0 1 0 1 1 1 1 1 0 1 1 1 0 1 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:37:16 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n234, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n243, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1044, new_n1045,
    new_n1046, new_n1047, new_n1048, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1071, new_n1072, new_n1073, new_n1074, new_n1075, new_n1076,
    new_n1077, new_n1078, new_n1079, new_n1080, new_n1081, new_n1082,
    new_n1083, new_n1084, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1235, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1291, new_n1292, new_n1293,
    new_n1294, new_n1295, new_n1296, new_n1297, new_n1298, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  XNOR2_X1  g0003(.A(new_n203), .B(KEYINPUT64), .ZN(new_n204));
  INV_X1    g0004(.A(G77), .ZN(new_n205));
  AND2_X1   g0005(.A1(new_n204), .A2(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  NOR2_X1   g0011(.A1(new_n211), .A2(G13), .ZN(new_n212));
  OAI211_X1 g0012(.A(new_n212), .B(G250), .C1(G257), .C2(G264), .ZN(new_n213));
  XOR2_X1   g0013(.A(new_n213), .B(KEYINPUT0), .Z(new_n214));
  NAND2_X1  g0014(.A1(G1), .A2(G13), .ZN(new_n215));
  INV_X1    g0015(.A(KEYINPUT65), .ZN(new_n216));
  NAND2_X1  g0016(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  NAND3_X1  g0017(.A1(KEYINPUT65), .A2(G1), .A3(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  INV_X1    g0019(.A(new_n219), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n220), .A2(new_n209), .ZN(new_n221));
  OAI21_X1  g0021(.A(G50), .B1(G58), .B2(G68), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  AOI21_X1  g0023(.A(new_n214), .B1(new_n221), .B2(new_n223), .ZN(new_n224));
  INV_X1    g0024(.A(G68), .ZN(new_n225));
  XNOR2_X1  g0025(.A(KEYINPUT67), .B(G238), .ZN(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT68), .B(G244), .ZN(new_n227));
  OAI22_X1  g0027(.A1(new_n225), .A2(new_n226), .B1(new_n227), .B2(new_n205), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G87), .A2(G250), .B1(G107), .B2(G264), .ZN(new_n229));
  AOI22_X1  g0029(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n230));
  AOI22_X1  g0030(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n231));
  NAND3_X1  g0031(.A1(new_n229), .A2(new_n230), .A3(new_n231), .ZN(new_n232));
  OAI21_X1  g0032(.A(new_n211), .B1(new_n228), .B2(new_n232), .ZN(new_n233));
  OAI21_X1  g0033(.A(new_n224), .B1(KEYINPUT1), .B2(new_n233), .ZN(new_n234));
  AOI21_X1  g0034(.A(new_n234), .B1(KEYINPUT1), .B2(new_n233), .ZN(G361));
  XNOR2_X1  g0035(.A(G238), .B(G244), .ZN(new_n236));
  INV_X1    g0036(.A(G232), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(KEYINPUT2), .B(G226), .ZN(new_n239));
  XOR2_X1   g0039(.A(new_n238), .B(new_n239), .Z(new_n240));
  XOR2_X1   g0040(.A(G264), .B(G270), .Z(new_n241));
  XNOR2_X1  g0041(.A(G250), .B(G257), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n241), .B(new_n242), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n240), .B(new_n243), .ZN(G358));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n245), .B(KEYINPUT69), .ZN(new_n246));
  XOR2_X1   g0046(.A(G107), .B(G116), .Z(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(G50), .B(G68), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n248), .B(new_n251), .Z(G351));
  INV_X1    g0052(.A(G33), .ZN(new_n253));
  OAI211_X1 g0053(.A(new_n217), .B(new_n218), .C1(new_n211), .C2(new_n253), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n204), .A2(new_n209), .ZN(new_n255));
  XOR2_X1   g0055(.A(KEYINPUT8), .B(G58), .Z(new_n256));
  INV_X1    g0056(.A(new_n256), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n209), .A2(G33), .ZN(new_n258));
  AND3_X1   g0058(.A1(new_n209), .A2(new_n253), .A3(KEYINPUT71), .ZN(new_n259));
  AOI21_X1  g0059(.A(KEYINPUT71), .B1(new_n209), .B2(new_n253), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n259), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(G150), .ZN(new_n262));
  OAI22_X1  g0062(.A1(new_n257), .A2(new_n258), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g0063(.A(new_n254), .B1(new_n255), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n254), .B1(new_n208), .B2(G20), .ZN(new_n265));
  NAND2_X1  g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  INV_X1    g0066(.A(G13), .ZN(new_n267));
  NOR3_X1   g0067(.A1(new_n267), .A2(new_n209), .A3(G1), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI211_X1 g0069(.A(new_n264), .B(new_n266), .C1(G50), .C2(new_n269), .ZN(new_n270));
  XNOR2_X1  g0070(.A(new_n270), .B(KEYINPUT9), .ZN(new_n271));
  OAI211_X1 g0071(.A(new_n208), .B(G274), .C1(G41), .C2(G45), .ZN(new_n272));
  XNOR2_X1  g0072(.A(new_n272), .B(KEYINPUT70), .ZN(new_n273));
  NAND2_X1  g0073(.A1(G33), .A2(G41), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(G1), .A3(G13), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n275), .A2(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g0078(.A(new_n273), .B1(G226), .B2(new_n278), .ZN(new_n279));
  XNOR2_X1  g0079(.A(KEYINPUT3), .B(G33), .ZN(new_n280));
  INV_X1    g0080(.A(G1698), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n280), .A2(G222), .A3(new_n281), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n280), .A2(G223), .A3(G1698), .ZN(new_n283));
  OAI211_X1 g0083(.A(new_n282), .B(new_n283), .C1(new_n205), .C2(new_n280), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n219), .A2(new_n274), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g0086(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n279), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g0088(.A1(new_n288), .A2(G200), .ZN(new_n289));
  INV_X1    g0089(.A(G190), .ZN(new_n290));
  OAI211_X1 g0090(.A(new_n271), .B(new_n289), .C1(new_n290), .C2(new_n288), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n291), .B(KEYINPUT10), .ZN(new_n292));
  INV_X1    g0092(.A(G169), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI211_X1 g0094(.A(new_n270), .B(new_n294), .C1(G179), .C2(new_n288), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n292), .A2(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(KEYINPUT17), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n300));
  XNOR2_X1  g0100(.A(KEYINPUT75), .B(G33), .ZN(new_n301));
  AOI21_X1  g0101(.A(new_n300), .B1(new_n301), .B2(KEYINPUT3), .ZN(new_n302));
  NAND2_X1  g0102(.A1(G226), .A2(G1698), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n281), .A2(G223), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n303), .B1(new_n304), .B2(KEYINPUT78), .ZN(new_n305));
  AOI22_X1  g0105(.A1(new_n302), .A2(new_n305), .B1(G33), .B2(G87), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n253), .A2(KEYINPUT75), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT75), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n308), .A2(G33), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n307), .A2(new_n309), .A3(KEYINPUT3), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT3), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(G33), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n310), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g0113(.A(KEYINPUT78), .B1(new_n313), .B2(new_n304), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n285), .B1(new_n306), .B2(new_n314), .ZN(new_n315));
  XOR2_X1   g0115(.A(new_n272), .B(KEYINPUT70), .Z(new_n316));
  OAI21_X1  g0116(.A(new_n316), .B1(new_n237), .B2(new_n277), .ZN(new_n317));
  OAI21_X1  g0117(.A(new_n299), .B1(new_n315), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(KEYINPUT78), .ZN(new_n319));
  INV_X1    g0119(.A(G223), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n320), .A2(G1698), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n319), .B1(new_n302), .B2(new_n321), .ZN(new_n322));
  AOI22_X1  g0122(.A1(new_n321), .A2(new_n319), .B1(G226), .B2(G1698), .ZN(new_n323));
  INV_X1    g0123(.A(G87), .ZN(new_n324));
  OAI22_X1  g0124(.A1(new_n313), .A2(new_n323), .B1(new_n253), .B2(new_n324), .ZN(new_n325));
  OAI21_X1  g0125(.A(new_n286), .B1(new_n322), .B2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n273), .B1(G232), .B2(new_n278), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n326), .A2(new_n290), .A3(new_n327), .ZN(new_n328));
  NAND3_X1  g0128(.A1(new_n318), .A2(new_n328), .A3(KEYINPUT79), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n315), .A2(new_n317), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT79), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n330), .A2(new_n331), .A3(new_n290), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n329), .A2(new_n332), .ZN(new_n333));
  NOR2_X1   g0133(.A1(new_n256), .A2(new_n268), .ZN(new_n334));
  INV_X1    g0134(.A(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n335), .B1(new_n265), .B2(new_n257), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n253), .A2(KEYINPUT3), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n337), .B1(new_n301), .B2(KEYINPUT3), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT7), .ZN(new_n339));
  NOR2_X1   g0139(.A1(new_n339), .A2(G20), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n338), .A2(new_n340), .ZN(new_n341));
  INV_X1    g0141(.A(KEYINPUT77), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n311), .A2(G33), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n209), .B1(new_n300), .B2(new_n343), .ZN(new_n344));
  AOI21_X1  g0144(.A(new_n342), .B1(new_n344), .B2(new_n339), .ZN(new_n345));
  AOI21_X1  g0145(.A(G20), .B1(new_n312), .B2(new_n337), .ZN(new_n346));
  NOR3_X1   g0146(.A1(new_n346), .A2(KEYINPUT77), .A3(KEYINPUT7), .ZN(new_n347));
  OAI21_X1  g0147(.A(new_n341), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n348), .A2(G68), .ZN(new_n349));
  INV_X1    g0149(.A(G58), .ZN(new_n350));
  NOR2_X1   g0150(.A1(new_n350), .A2(new_n225), .ZN(new_n351));
  OAI21_X1  g0151(.A(G20), .B1(new_n351), .B2(new_n201), .ZN(new_n352));
  INV_X1    g0152(.A(G159), .ZN(new_n353));
  OAI21_X1  g0153(.A(new_n352), .B1(new_n261), .B2(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT16), .B1(new_n349), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT76), .ZN(new_n357));
  OAI21_X1  g0157(.A(new_n209), .B1(new_n357), .B2(KEYINPUT7), .ZN(new_n358));
  INV_X1    g0158(.A(new_n358), .ZN(new_n359));
  NAND2_X1  g0159(.A1(new_n357), .A2(KEYINPUT7), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n313), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n361), .A2(G68), .ZN(new_n362));
  AOI21_X1  g0162(.A(new_n358), .B1(new_n310), .B2(new_n312), .ZN(new_n363));
  NOR2_X1   g0163(.A1(new_n363), .A2(new_n360), .ZN(new_n364));
  OAI211_X1 g0164(.A(KEYINPUT16), .B(new_n355), .C1(new_n362), .C2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n365), .A2(new_n254), .ZN(new_n366));
  OAI21_X1  g0166(.A(new_n336), .B1(new_n356), .B2(new_n366), .ZN(new_n367));
  OAI21_X1  g0167(.A(new_n298), .B1(new_n333), .B2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n293), .B1(new_n326), .B2(new_n327), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n369), .B1(G179), .B2(new_n330), .ZN(new_n370));
  INV_X1    g0170(.A(new_n336), .ZN(new_n371));
  AOI21_X1  g0171(.A(new_n219), .B1(G33), .B2(new_n210), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n225), .B1(new_n363), .B2(new_n360), .ZN(new_n373));
  OAI211_X1 g0173(.A(new_n357), .B(KEYINPUT7), .C1(new_n302), .C2(G20), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n354), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n372), .B1(new_n375), .B2(KEYINPUT16), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT16), .ZN(new_n377));
  OAI21_X1  g0177(.A(KEYINPUT77), .B1(new_n346), .B2(KEYINPUT7), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n342), .B(new_n339), .C1(new_n280), .C2(G20), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AOI21_X1  g0180(.A(new_n225), .B1(new_n380), .B2(new_n341), .ZN(new_n381));
  OAI21_X1  g0181(.A(new_n377), .B1(new_n381), .B2(new_n354), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n371), .B1(new_n376), .B2(new_n382), .ZN(new_n383));
  OAI21_X1  g0183(.A(KEYINPUT18), .B1(new_n370), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n330), .A2(G179), .ZN(new_n385));
  OAI21_X1  g0185(.A(new_n385), .B1(new_n293), .B2(new_n330), .ZN(new_n386));
  INV_X1    g0186(.A(KEYINPUT18), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n386), .A2(new_n367), .A3(new_n387), .ZN(new_n388));
  NAND4_X1  g0188(.A1(new_n383), .A2(KEYINPUT17), .A3(new_n332), .A4(new_n329), .ZN(new_n389));
  NAND4_X1  g0189(.A1(new_n368), .A2(new_n384), .A3(new_n388), .A4(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NOR2_X1   g0191(.A1(new_n261), .A2(new_n202), .ZN(new_n392));
  OAI22_X1  g0192(.A1(new_n258), .A2(new_n205), .B1(new_n209), .B2(G68), .ZN(new_n393));
  OAI21_X1  g0193(.A(new_n254), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  XNOR2_X1  g0194(.A(new_n394), .B(KEYINPUT11), .ZN(new_n395));
  NOR2_X1   g0195(.A1(new_n254), .A2(new_n268), .ZN(new_n396));
  AOI21_X1  g0196(.A(new_n225), .B1(new_n208), .B2(G20), .ZN(new_n397));
  INV_X1    g0197(.A(KEYINPUT74), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT12), .ZN(new_n399));
  OAI21_X1  g0199(.A(new_n225), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  OAI22_X1  g0200(.A1(new_n269), .A2(new_n400), .B1(KEYINPUT74), .B2(KEYINPUT12), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n268), .A2(new_n398), .A3(new_n399), .A4(new_n225), .ZN(new_n402));
  AOI22_X1  g0202(.A1(new_n396), .A2(new_n397), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  NAND2_X1  g0203(.A1(new_n395), .A2(new_n403), .ZN(new_n404));
  INV_X1    g0204(.A(G238), .ZN(new_n405));
  OAI21_X1  g0205(.A(new_n316), .B1(new_n405), .B2(new_n277), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n237), .A2(G1698), .ZN(new_n407));
  OAI211_X1 g0207(.A(new_n280), .B(new_n407), .C1(G226), .C2(G1698), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G97), .ZN(new_n409));
  INV_X1    g0209(.A(KEYINPUT73), .ZN(new_n410));
  XNOR2_X1  g0210(.A(new_n409), .B(new_n410), .ZN(new_n411));
  INV_X1    g0211(.A(new_n411), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n285), .B1(new_n408), .B2(new_n412), .ZN(new_n413));
  OR3_X1    g0213(.A1(new_n406), .A2(KEYINPUT13), .A3(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT13), .B1(new_n406), .B2(new_n413), .ZN(new_n415));
  AND2_X1   g0215(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n416), .A2(G179), .ZN(new_n417));
  INV_X1    g0217(.A(KEYINPUT14), .ZN(new_n418));
  AOI21_X1  g0218(.A(new_n293), .B1(new_n414), .B2(new_n415), .ZN(new_n419));
  OAI21_X1  g0219(.A(new_n417), .B1(new_n418), .B2(new_n419), .ZN(new_n420));
  AND2_X1   g0220(.A1(new_n419), .A2(new_n418), .ZN(new_n421));
  OAI21_X1  g0221(.A(new_n404), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  AOI21_X1  g0222(.A(new_n404), .B1(new_n416), .B2(G190), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(new_n299), .B2(new_n416), .ZN(new_n424));
  AND2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n265), .A2(G77), .ZN(new_n426));
  XNOR2_X1  g0226(.A(KEYINPUT15), .B(G87), .ZN(new_n427));
  OAI22_X1  g0227(.A1(new_n427), .A2(new_n258), .B1(new_n209), .B2(new_n205), .ZN(new_n428));
  OR2_X1    g0228(.A1(new_n259), .A2(new_n260), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n428), .B1(new_n429), .B2(new_n256), .ZN(new_n430));
  OAI221_X1 g0230(.A(new_n426), .B1(G77), .B2(new_n269), .C1(new_n372), .C2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT72), .B(G107), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n286), .B1(new_n280), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(new_n280), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n226), .A2(G1698), .ZN(new_n435));
  NAND2_X1  g0235(.A1(new_n237), .A2(new_n281), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n434), .B1(new_n435), .B2(new_n436), .ZN(new_n437));
  OAI221_X1 g0237(.A(new_n316), .B1(new_n227), .B2(new_n277), .C1(new_n433), .C2(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n431), .B1(G200), .B2(new_n438), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n439), .B1(new_n290), .B2(new_n438), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n438), .A2(new_n293), .ZN(new_n441));
  OAI211_X1 g0241(.A(new_n431), .B(new_n441), .C1(G179), .C2(new_n438), .ZN(new_n442));
  AND2_X1   g0242(.A1(new_n440), .A2(new_n442), .ZN(new_n443));
  NAND4_X1  g0243(.A1(new_n297), .A2(new_n391), .A3(new_n425), .A4(new_n443), .ZN(new_n444));
  NAND4_X1  g0244(.A1(new_n310), .A2(new_n209), .A3(G87), .A4(new_n312), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT22), .ZN(new_n446));
  NOR3_X1   g0246(.A1(new_n324), .A2(KEYINPUT22), .A3(G20), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n280), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n448), .A2(KEYINPUT86), .ZN(new_n449));
  INV_X1    g0249(.A(KEYINPUT86), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n280), .A2(new_n450), .A3(new_n447), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n446), .A2(new_n449), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT87), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n307), .A2(new_n309), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n454), .A2(G116), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT23), .ZN(new_n456));
  AOI21_X1  g0256(.A(G20), .B1(new_n455), .B2(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(G107), .ZN(new_n458));
  NAND3_X1  g0258(.A1(new_n456), .A2(new_n458), .A3(G20), .ZN(new_n459));
  INV_X1    g0259(.A(new_n432), .ZN(new_n460));
  OAI21_X1  g0260(.A(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n457), .A2(new_n461), .ZN(new_n462));
  NAND3_X1  g0262(.A1(new_n452), .A2(new_n453), .A3(new_n462), .ZN(new_n463));
  INV_X1    g0263(.A(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n453), .B1(new_n452), .B2(new_n462), .ZN(new_n465));
  OAI21_X1  g0265(.A(KEYINPUT24), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  INV_X1    g0266(.A(new_n465), .ZN(new_n467));
  INV_X1    g0267(.A(KEYINPUT24), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(new_n468), .A3(new_n463), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n466), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n254), .ZN(new_n471));
  MUX2_X1   g0271(.A(G250), .B(G257), .S(G1698), .Z(new_n472));
  AOI22_X1  g0272(.A1(new_n302), .A2(new_n472), .B1(G294), .B2(new_n454), .ZN(new_n473));
  INV_X1    g0273(.A(G264), .ZN(new_n474));
  XNOR2_X1  g0274(.A(KEYINPUT5), .B(G41), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n475), .A2(new_n208), .A3(G45), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n476), .A2(new_n275), .ZN(new_n477));
  OAI22_X1  g0277(.A1(new_n473), .A2(new_n285), .B1(new_n474), .B2(new_n477), .ZN(new_n478));
  INV_X1    g0278(.A(new_n478), .ZN(new_n479));
  INV_X1    g0279(.A(G274), .ZN(new_n480));
  INV_X1    g0280(.A(new_n275), .ZN(new_n481));
  OR3_X1    g0281(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g0283(.A(KEYINPUT89), .B1(new_n483), .B2(G190), .ZN(new_n484));
  NOR3_X1   g0284(.A1(new_n476), .A2(new_n480), .A3(new_n481), .ZN(new_n485));
  OR4_X1    g0285(.A1(KEYINPUT89), .A2(new_n478), .A3(G190), .A4(new_n485), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n483), .A2(new_n299), .ZN(new_n487));
  NAND3_X1  g0287(.A1(new_n484), .A2(new_n486), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g0288(.A1(new_n268), .A2(new_n458), .ZN(new_n489));
  INV_X1    g0289(.A(KEYINPUT25), .ZN(new_n490));
  XNOR2_X1  g0290(.A(new_n489), .B(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n208), .A2(G33), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n372), .A2(new_n269), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g0293(.A(new_n491), .B1(new_n493), .B2(new_n458), .ZN(new_n494));
  INV_X1    g0294(.A(new_n494), .ZN(new_n495));
  NAND3_X1  g0295(.A1(new_n471), .A2(new_n488), .A3(new_n495), .ZN(new_n496));
  NOR2_X1   g0296(.A1(new_n269), .A2(G97), .ZN(new_n497));
  INV_X1    g0297(.A(new_n493), .ZN(new_n498));
  AOI21_X1  g0298(.A(new_n497), .B1(new_n498), .B2(G97), .ZN(new_n499));
  XNOR2_X1  g0299(.A(G97), .B(G107), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT6), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(G97), .ZN(new_n503));
  NOR3_X1   g0303(.A1(new_n501), .A2(new_n503), .A3(G107), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n502), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n506), .A2(G20), .B1(new_n429), .B2(G77), .ZN(new_n507));
  AOI22_X1  g0307(.A1(new_n378), .A2(new_n379), .B1(new_n338), .B2(new_n340), .ZN(new_n508));
  OAI21_X1  g0308(.A(new_n507), .B1(new_n508), .B2(new_n460), .ZN(new_n509));
  AND3_X1   g0309(.A1(new_n509), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n510));
  AOI21_X1  g0310(.A(KEYINPUT80), .B1(new_n509), .B2(new_n254), .ZN(new_n511));
  OAI21_X1  g0311(.A(new_n499), .B1(new_n510), .B2(new_n511), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(KEYINPUT81), .ZN(new_n513));
  INV_X1    g0313(.A(KEYINPUT80), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n504), .B1(new_n501), .B2(new_n500), .ZN(new_n515));
  OAI22_X1  g0315(.A1(new_n515), .A2(new_n209), .B1(new_n205), .B2(new_n261), .ZN(new_n516));
  AOI21_X1  g0316(.A(new_n516), .B1(new_n348), .B2(new_n432), .ZN(new_n517));
  OAI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(new_n372), .ZN(new_n518));
  NAND3_X1  g0318(.A1(new_n509), .A2(KEYINPUT80), .A3(new_n254), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  INV_X1    g0320(.A(KEYINPUT81), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n520), .A2(new_n521), .A3(new_n499), .ZN(new_n522));
  INV_X1    g0322(.A(new_n477), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n485), .B1(G257), .B2(new_n523), .ZN(new_n524));
  INV_X1    g0324(.A(G244), .ZN(new_n525));
  NOR2_X1   g0325(.A1(new_n525), .A2(G1698), .ZN(new_n526));
  AOI21_X1  g0326(.A(KEYINPUT4), .B1(new_n302), .B2(new_n526), .ZN(new_n527));
  NAND4_X1  g0327(.A1(new_n280), .A2(KEYINPUT4), .A3(G244), .A4(new_n281), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n280), .A2(G250), .A3(G1698), .ZN(new_n529));
  NAND2_X1  g0329(.A1(G33), .A2(G283), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT82), .ZN(new_n531));
  XNOR2_X1  g0331(.A(new_n530), .B(new_n531), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n528), .A2(new_n529), .A3(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n286), .B1(new_n527), .B2(new_n533), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n524), .A2(new_n534), .ZN(new_n535));
  NOR2_X1   g0335(.A1(new_n535), .A2(new_n290), .ZN(new_n536));
  AOI21_X1  g0336(.A(new_n536), .B1(G200), .B2(new_n535), .ZN(new_n537));
  NAND3_X1  g0337(.A1(new_n513), .A2(new_n522), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n539), .A2(G179), .ZN(new_n540));
  NAND2_X1  g0340(.A1(new_n535), .A2(G169), .ZN(new_n541));
  NAND2_X1  g0341(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n512), .A2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(G238), .A2(G1698), .ZN(new_n544));
  AOI21_X1  g0344(.A(new_n544), .B1(new_n525), .B2(G1698), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n302), .A2(new_n545), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n546), .A2(new_n455), .ZN(new_n547));
  NAND2_X1  g0347(.A1(new_n547), .A2(new_n286), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n208), .A2(G45), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n275), .A2(G250), .A3(new_n549), .ZN(new_n550));
  NAND3_X1  g0350(.A1(new_n208), .A2(G45), .A3(G274), .ZN(new_n551));
  NAND2_X1  g0351(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n552), .A2(KEYINPUT83), .ZN(new_n553));
  INV_X1    g0353(.A(KEYINPUT83), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n550), .A2(new_n554), .A3(new_n551), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n553), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n548), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n302), .A2(new_n209), .A3(G68), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT19), .ZN(new_n560));
  OAI21_X1  g0360(.A(new_n560), .B1(new_n258), .B2(new_n503), .ZN(new_n561));
  AOI21_X1  g0361(.A(G20), .B1(new_n411), .B2(KEYINPUT19), .ZN(new_n562));
  NOR3_X1   g0362(.A1(new_n432), .A2(G87), .A3(G97), .ZN(new_n563));
  OAI211_X1 g0363(.A(new_n559), .B(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n254), .B1(new_n268), .B2(new_n427), .ZN(new_n565));
  OAI21_X1  g0365(.A(KEYINPUT84), .B1(new_n493), .B2(new_n324), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT84), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n396), .A2(new_n567), .A3(G87), .A4(new_n492), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n566), .A2(new_n568), .ZN(new_n569));
  NAND3_X1  g0369(.A1(new_n548), .A2(G190), .A3(new_n556), .ZN(new_n570));
  NAND4_X1  g0370(.A1(new_n558), .A2(new_n565), .A3(new_n569), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g0371(.A1(new_n564), .A2(new_n254), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n427), .A2(new_n268), .ZN(new_n573));
  INV_X1    g0373(.A(new_n427), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n498), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g0375(.A1(new_n572), .A2(new_n573), .A3(new_n575), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n557), .A2(new_n293), .ZN(new_n577));
  INV_X1    g0377(.A(G179), .ZN(new_n578));
  NAND3_X1  g0378(.A1(new_n548), .A2(new_n578), .A3(new_n556), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n576), .A2(new_n577), .A3(new_n579), .ZN(new_n580));
  AND2_X1   g0380(.A1(new_n571), .A2(new_n580), .ZN(new_n581));
  NAND4_X1  g0381(.A1(new_n496), .A2(new_n538), .A3(new_n543), .A4(new_n581), .ZN(new_n582));
  NOR2_X1   g0382(.A1(new_n483), .A2(G179), .ZN(new_n583));
  AOI21_X1  g0383(.A(new_n583), .B1(new_n293), .B2(new_n483), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n372), .B1(new_n466), .B2(new_n469), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n584), .B1(new_n585), .B2(new_n494), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n586), .A2(KEYINPUT88), .ZN(new_n587));
  OAI211_X1 g0387(.A(new_n532), .B(new_n209), .C1(G33), .C2(new_n503), .ZN(new_n588));
  INV_X1    g0388(.A(G116), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(G20), .ZN(new_n590));
  NAND4_X1  g0390(.A1(new_n588), .A2(KEYINPUT20), .A3(new_n254), .A4(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT85), .ZN(new_n592));
  AND2_X1   g0392(.A1(new_n254), .A2(new_n590), .ZN(new_n593));
  INV_X1    g0393(.A(KEYINPUT85), .ZN(new_n594));
  NAND4_X1  g0394(.A1(new_n593), .A2(new_n594), .A3(KEYINPUT20), .A4(new_n588), .ZN(new_n595));
  NAND3_X1  g0395(.A1(new_n588), .A2(new_n254), .A3(new_n590), .ZN(new_n596));
  INV_X1    g0396(.A(KEYINPUT20), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n596), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n592), .A2(new_n595), .A3(new_n598), .ZN(new_n599));
  NOR2_X1   g0399(.A1(new_n269), .A2(G116), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n600), .B1(new_n498), .B2(G116), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n599), .A2(new_n601), .ZN(new_n602));
  INV_X1    g0402(.A(G270), .ZN(new_n603));
  OAI21_X1  g0403(.A(new_n482), .B1(new_n603), .B2(new_n477), .ZN(new_n604));
  NOR2_X1   g0404(.A1(G257), .A2(G1698), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n605), .B1(new_n474), .B2(G1698), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n302), .A2(new_n606), .B1(G303), .B2(new_n434), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n607), .A2(new_n285), .ZN(new_n608));
  NOR3_X1   g0408(.A1(new_n604), .A2(new_n608), .A3(new_n578), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n602), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g0410(.A(G169), .B1(new_n604), .B2(new_n608), .ZN(new_n611));
  AOI21_X1  g0411(.A(new_n611), .B1(new_n599), .B2(new_n601), .ZN(new_n612));
  OAI21_X1  g0412(.A(new_n610), .B1(new_n612), .B2(KEYINPUT21), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n604), .A2(new_n608), .ZN(new_n614));
  NAND2_X1  g0414(.A1(new_n614), .A2(G190), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n615), .B1(new_n299), .B2(new_n614), .ZN(new_n616));
  NOR2_X1   g0416(.A1(new_n616), .A2(new_n602), .ZN(new_n617));
  INV_X1    g0417(.A(new_n611), .ZN(new_n618));
  NAND2_X1  g0418(.A1(new_n602), .A2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(KEYINPUT21), .ZN(new_n620));
  NOR2_X1   g0420(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  NOR3_X1   g0421(.A1(new_n613), .A2(new_n617), .A3(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT88), .ZN(new_n623));
  OAI211_X1 g0423(.A(new_n584), .B(new_n623), .C1(new_n585), .C2(new_n494), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n587), .A2(new_n622), .A3(new_n624), .ZN(new_n625));
  NOR3_X1   g0425(.A1(new_n444), .A2(new_n582), .A3(new_n625), .ZN(G372));
  NOR2_X1   g0426(.A1(new_n613), .A2(new_n621), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n582), .B1(new_n586), .B2(new_n627), .ZN(new_n628));
  INV_X1    g0428(.A(new_n543), .ZN(new_n629));
  NAND3_X1  g0429(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n581), .ZN(new_n630));
  INV_X1    g0430(.A(new_n542), .ZN(new_n631));
  AOI21_X1  g0431(.A(new_n631), .B1(new_n513), .B2(new_n522), .ZN(new_n632));
  AOI21_X1  g0432(.A(KEYINPUT26), .B1(new_n632), .B2(new_n581), .ZN(new_n633));
  INV_X1    g0433(.A(KEYINPUT90), .ZN(new_n634));
  OAI21_X1  g0434(.A(new_n630), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  AOI21_X1  g0435(.A(new_n521), .B1(new_n520), .B2(new_n499), .ZN(new_n636));
  INV_X1    g0436(.A(new_n499), .ZN(new_n637));
  AOI211_X1 g0437(.A(KEYINPUT81), .B(new_n637), .C1(new_n518), .C2(new_n519), .ZN(new_n638));
  OAI211_X1 g0438(.A(new_n542), .B(new_n581), .C1(new_n636), .C2(new_n638), .ZN(new_n639));
  INV_X1    g0439(.A(KEYINPUT26), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NOR2_X1   g0441(.A1(new_n641), .A2(KEYINPUT90), .ZN(new_n642));
  OAI21_X1  g0442(.A(new_n580), .B1(new_n635), .B2(new_n642), .ZN(new_n643));
  AOI21_X1  g0443(.A(new_n628), .B1(new_n643), .B2(KEYINPUT91), .ZN(new_n644));
  INV_X1    g0444(.A(new_n580), .ZN(new_n645));
  AND3_X1   g0445(.A1(new_n629), .A2(KEYINPUT26), .A3(new_n581), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n646), .B1(new_n641), .B2(KEYINPUT90), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n633), .A2(new_n634), .ZN(new_n648));
  AOI21_X1  g0448(.A(new_n645), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(KEYINPUT91), .ZN(new_n650));
  NAND2_X1  g0450(.A1(new_n649), .A2(new_n650), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n444), .B1(new_n644), .B2(new_n651), .ZN(new_n652));
  XNOR2_X1  g0452(.A(new_n652), .B(KEYINPUT92), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n422), .A2(new_n442), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n654), .A2(new_n424), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n368), .A2(new_n389), .ZN(new_n656));
  OAI211_X1 g0456(.A(new_n384), .B(new_n388), .C1(new_n655), .C2(new_n656), .ZN(new_n657));
  INV_X1    g0457(.A(KEYINPUT93), .ZN(new_n658));
  OR2_X1    g0458(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n657), .A2(new_n658), .ZN(new_n660));
  NAND3_X1  g0460(.A1(new_n659), .A2(new_n292), .A3(new_n660), .ZN(new_n661));
  AND2_X1   g0461(.A1(new_n661), .A2(new_n295), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n653), .A2(new_n662), .ZN(G369));
  INV_X1    g0463(.A(KEYINPUT95), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n665));
  OR2_X1    g0465(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(KEYINPUT27), .ZN(new_n667));
  NAND3_X1  g0467(.A1(new_n666), .A2(G213), .A3(new_n667), .ZN(new_n668));
  XNOR2_X1  g0468(.A(KEYINPUT94), .B(G343), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n668), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n602), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n622), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n627), .B2(new_n671), .ZN(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  OAI21_X1  g0474(.A(new_n670), .B1(new_n585), .B2(new_n494), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n587), .A2(new_n496), .A3(new_n624), .A4(new_n675), .ZN(new_n676));
  INV_X1    g0476(.A(new_n586), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n677), .A2(new_n670), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n676), .A2(new_n678), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n664), .B1(new_n674), .B2(new_n679), .ZN(new_n680));
  AND4_X1   g0480(.A1(new_n664), .A2(new_n679), .A3(G330), .A4(new_n673), .ZN(new_n681));
  NOR2_X1   g0481(.A1(new_n680), .A2(new_n681), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n627), .A2(new_n670), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n684), .A2(new_n496), .A3(new_n587), .A4(new_n624), .ZN(new_n685));
  INV_X1    g0485(.A(new_n670), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n677), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n685), .A2(new_n687), .ZN(new_n688));
  INV_X1    g0488(.A(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n683), .A2(new_n689), .ZN(G399));
  INV_X1    g0490(.A(new_n212), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(G41), .ZN(new_n692));
  INV_X1    g0492(.A(new_n692), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n563), .A2(new_n589), .ZN(new_n694));
  INV_X1    g0494(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g0495(.A1(new_n693), .A2(G1), .A3(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(new_n223), .ZN(new_n697));
  OAI21_X1  g0497(.A(new_n696), .B1(new_n697), .B2(new_n693), .ZN(new_n698));
  XNOR2_X1  g0498(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  XNOR2_X1  g0499(.A(new_n699), .B(KEYINPUT28), .ZN(new_n700));
  INV_X1    g0500(.A(new_n582), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n587), .A2(new_n624), .ZN(new_n702));
  INV_X1    g0502(.A(new_n627), .ZN(new_n703));
  OAI21_X1  g0503(.A(new_n701), .B1(new_n702), .B2(new_n703), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n629), .A2(new_n640), .A3(new_n581), .ZN(new_n705));
  XNOR2_X1  g0505(.A(new_n580), .B(KEYINPUT99), .ZN(new_n706));
  NAND2_X1  g0506(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  AOI21_X1  g0507(.A(new_n707), .B1(KEYINPUT26), .B2(new_n639), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n670), .B1(new_n704), .B2(new_n708), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT29), .ZN(new_n710));
  NOR2_X1   g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n670), .B1(new_n644), .B2(new_n651), .ZN(new_n712));
  AOI21_X1  g0512(.A(new_n711), .B1(new_n712), .B2(new_n710), .ZN(new_n713));
  AND3_X1   g0513(.A1(new_n587), .A2(new_n622), .A3(new_n624), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n714), .A2(new_n701), .A3(new_n686), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n557), .A2(new_n478), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n716), .A2(new_n539), .A3(new_n609), .ZN(new_n717));
  INV_X1    g0517(.A(KEYINPUT30), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n717), .A2(new_n718), .ZN(new_n719));
  NOR3_X1   g0519(.A1(new_n535), .A2(new_n557), .A3(new_n478), .ZN(new_n720));
  NAND3_X1  g0520(.A1(new_n720), .A2(KEYINPUT30), .A3(new_n609), .ZN(new_n721));
  INV_X1    g0521(.A(new_n614), .ZN(new_n722));
  AOI21_X1  g0522(.A(G179), .B1(new_n548), .B2(new_n556), .ZN(new_n723));
  NAND4_X1  g0523(.A1(new_n722), .A2(new_n535), .A3(new_n483), .A4(new_n723), .ZN(new_n724));
  NAND3_X1  g0524(.A1(new_n719), .A2(new_n721), .A3(new_n724), .ZN(new_n725));
  NAND3_X1  g0525(.A1(new_n725), .A2(KEYINPUT31), .A3(new_n670), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT97), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  NAND4_X1  g0528(.A1(new_n725), .A2(KEYINPUT97), .A3(KEYINPUT31), .A4(new_n670), .ZN(new_n729));
  NAND2_X1  g0529(.A1(new_n725), .A2(new_n670), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT31), .ZN(new_n731));
  NAND2_X1  g0531(.A1(new_n730), .A2(new_n731), .ZN(new_n732));
  NAND3_X1  g0532(.A1(new_n728), .A2(new_n729), .A3(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n733), .A2(KEYINPUT98), .ZN(new_n734));
  INV_X1    g0534(.A(KEYINPUT98), .ZN(new_n735));
  NAND4_X1  g0535(.A1(new_n728), .A2(new_n732), .A3(new_n735), .A4(new_n729), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n715), .A2(new_n734), .A3(new_n736), .ZN(new_n737));
  NAND2_X1  g0537(.A1(new_n737), .A2(G330), .ZN(new_n738));
  NAND2_X1  g0538(.A1(new_n713), .A2(new_n738), .ZN(new_n739));
  INV_X1    g0539(.A(new_n739), .ZN(new_n740));
  OAI21_X1  g0540(.A(new_n700), .B1(new_n740), .B2(G1), .ZN(G364));
  NOR2_X1   g0541(.A1(new_n267), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n208), .B1(new_n742), .B2(G45), .ZN(new_n743));
  INV_X1    g0543(.A(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n692), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g0545(.A1(new_n674), .A2(new_n745), .ZN(new_n746));
  OAI21_X1  g0546(.A(new_n746), .B1(G330), .B2(new_n673), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n220), .B1(G20), .B2(new_n293), .ZN(new_n748));
  NOR2_X1   g0548(.A1(G13), .A2(G33), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(G20), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n748), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g0552(.A1(new_n212), .A2(new_n280), .ZN(new_n753));
  INV_X1    g0553(.A(G355), .ZN(new_n754));
  OAI22_X1  g0554(.A1(new_n753), .A2(new_n754), .B1(G116), .B2(new_n212), .ZN(new_n755));
  XNOR2_X1  g0555(.A(new_n755), .B(KEYINPUT100), .ZN(new_n756));
  NAND2_X1  g0556(.A1(new_n251), .A2(G45), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n691), .A2(new_n302), .ZN(new_n758));
  OAI211_X1 g0558(.A(new_n757), .B(new_n758), .C1(G45), .C2(new_n697), .ZN(new_n759));
  NAND2_X1  g0559(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT101), .ZN(new_n761));
  OAI21_X1  g0561(.A(new_n752), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(new_n762), .B1(new_n761), .B2(new_n760), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n209), .A2(G190), .ZN(new_n764));
  NOR2_X1   g0564(.A1(G179), .A2(G200), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  OR3_X1    g0566(.A1(new_n766), .A2(KEYINPUT32), .A3(new_n353), .ZN(new_n767));
  OAI21_X1  g0567(.A(KEYINPUT32), .B1(new_n766), .B2(new_n353), .ZN(new_n768));
  AOI21_X1  g0568(.A(new_n209), .B1(new_n765), .B2(G190), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g0570(.A1(new_n770), .A2(G97), .ZN(new_n771));
  NAND3_X1  g0571(.A1(new_n767), .A2(new_n768), .A3(new_n771), .ZN(new_n772));
  NOR2_X1   g0572(.A1(new_n209), .A2(new_n290), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n578), .A2(new_n299), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n578), .A2(G200), .ZN(new_n777));
  NAND2_X1  g0577(.A1(new_n773), .A2(new_n777), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  AOI22_X1  g0579(.A1(G50), .A2(new_n776), .B1(new_n779), .B2(G58), .ZN(new_n780));
  NAND2_X1  g0580(.A1(new_n764), .A2(new_n777), .ZN(new_n781));
  OAI21_X1  g0581(.A(new_n780), .B1(new_n205), .B2(new_n781), .ZN(new_n782));
  AND3_X1   g0582(.A1(new_n774), .A2(KEYINPUT103), .A3(new_n764), .ZN(new_n783));
  AOI21_X1  g0583(.A(KEYINPUT103), .B1(new_n774), .B2(new_n764), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  AOI211_X1 g0586(.A(new_n772), .B(new_n782), .C1(G68), .C2(new_n786), .ZN(new_n787));
  NOR2_X1   g0587(.A1(new_n299), .A2(G179), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n764), .A2(new_n788), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n458), .ZN(new_n790));
  NAND2_X1  g0590(.A1(new_n773), .A2(new_n788), .ZN(new_n791));
  INV_X1    g0591(.A(new_n791), .ZN(new_n792));
  AOI211_X1 g0592(.A(new_n434), .B(new_n790), .C1(G87), .C2(new_n792), .ZN(new_n793));
  XNOR2_X1  g0593(.A(new_n793), .B(KEYINPUT102), .ZN(new_n794));
  INV_X1    g0594(.A(new_n766), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n776), .A2(G326), .B1(new_n795), .B2(G329), .ZN(new_n796));
  NAND2_X1  g0596(.A1(new_n770), .A2(G294), .ZN(new_n797));
  INV_X1    g0597(.A(new_n781), .ZN(new_n798));
  AOI21_X1  g0598(.A(new_n280), .B1(new_n798), .B2(G311), .ZN(new_n799));
  AND3_X1   g0599(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(G303), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n791), .A2(new_n801), .ZN(new_n802));
  INV_X1    g0602(.A(G322), .ZN(new_n803));
  INV_X1    g0603(.A(G283), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n778), .A2(new_n803), .B1(new_n789), .B2(new_n804), .ZN(new_n805));
  XNOR2_X1  g0605(.A(KEYINPUT33), .B(G317), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n802), .B(new_n805), .C1(new_n786), .C2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(new_n787), .A2(new_n794), .B1(new_n800), .B2(new_n807), .ZN(new_n808));
  INV_X1    g0608(.A(new_n748), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n745), .B1(new_n808), .B2(new_n809), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n763), .A2(new_n810), .ZN(new_n811));
  INV_X1    g0611(.A(new_n751), .ZN(new_n812));
  OAI21_X1  g0612(.A(new_n811), .B1(new_n673), .B2(new_n812), .ZN(new_n813));
  AND2_X1   g0613(.A1(new_n747), .A2(new_n813), .ZN(new_n814));
  INV_X1    g0614(.A(new_n814), .ZN(G396));
  NAND2_X1  g0615(.A1(new_n431), .A2(new_n670), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n440), .A2(new_n816), .ZN(new_n817));
  AND2_X1   g0617(.A1(new_n817), .A2(new_n442), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n442), .A2(new_n670), .ZN(new_n819));
  NOR2_X1   g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  XNOR2_X1  g0620(.A(new_n712), .B(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n745), .B1(new_n821), .B2(new_n738), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n822), .B1(new_n738), .B2(new_n821), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n775), .A2(new_n801), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n434), .B1(new_n781), .B2(new_n589), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n824), .B(new_n825), .C1(G311), .C2(new_n795), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n786), .A2(G283), .ZN(new_n827));
  NOR2_X1   g0627(.A1(new_n789), .A2(new_n324), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n791), .A2(new_n458), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n828), .B(new_n829), .C1(G294), .C2(new_n779), .ZN(new_n830));
  NAND4_X1  g0630(.A1(new_n826), .A2(new_n771), .A3(new_n827), .A4(new_n830), .ZN(new_n831));
  AOI22_X1  g0631(.A1(G137), .A2(new_n776), .B1(new_n779), .B2(G143), .ZN(new_n832));
  OAI221_X1 g0632(.A(new_n832), .B1(new_n353), .B2(new_n781), .C1(new_n785), .C2(new_n262), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n834), .A2(KEYINPUT34), .ZN(new_n835));
  INV_X1    g0635(.A(G132), .ZN(new_n836));
  OAI22_X1  g0636(.A1(new_n791), .A2(new_n202), .B1(new_n766), .B2(new_n836), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n302), .B1(new_n350), .B2(new_n769), .ZN(new_n838));
  INV_X1    g0638(.A(new_n789), .ZN(new_n839));
  AOI211_X1 g0639(.A(new_n837), .B(new_n838), .C1(G68), .C2(new_n839), .ZN(new_n840));
  INV_X1    g0640(.A(KEYINPUT34), .ZN(new_n841));
  OAI21_X1  g0641(.A(new_n840), .B1(new_n841), .B2(new_n833), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n831), .B1(new_n835), .B2(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n843), .A2(new_n748), .ZN(new_n844));
  INV_X1    g0644(.A(new_n745), .ZN(new_n845));
  NOR2_X1   g0645(.A1(new_n748), .A2(new_n749), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n845), .B1(new_n846), .B2(new_n205), .ZN(new_n847));
  OAI211_X1 g0647(.A(new_n844), .B(new_n847), .C1(new_n820), .C2(new_n750), .ZN(new_n848));
  NAND2_X1  g0648(.A1(new_n823), .A2(new_n848), .ZN(G384));
  OR2_X1    g0649(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n850));
  NAND2_X1  g0650(.A1(new_n506), .A2(KEYINPUT35), .ZN(new_n851));
  NAND4_X1  g0651(.A1(new_n850), .A2(G116), .A3(new_n221), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(new_n852), .B(KEYINPUT36), .Z(new_n853));
  OAI211_X1 g0653(.A(new_n223), .B(G77), .C1(new_n350), .C2(new_n225), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n202), .A2(G68), .ZN(new_n855));
  AOI211_X1 g0655(.A(new_n208), .B(G13), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n853), .A2(new_n856), .ZN(new_n857));
  INV_X1    g0657(.A(new_n668), .ZN(new_n858));
  AOI21_X1  g0658(.A(new_n858), .B1(new_n384), .B2(new_n388), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n375), .A2(KEYINPUT16), .ZN(new_n860));
  OAI21_X1  g0660(.A(new_n336), .B1(new_n366), .B2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n861), .A2(KEYINPUT104), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT104), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n863), .B(new_n336), .C1(new_n366), .C2(new_n860), .ZN(new_n864));
  NAND3_X1  g0664(.A1(new_n862), .A2(new_n858), .A3(new_n864), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n862), .A2(new_n386), .A3(new_n864), .ZN(new_n866));
  NAND3_X1  g0666(.A1(new_n383), .A2(new_n332), .A3(new_n329), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n865), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n868), .A2(KEYINPUT37), .ZN(new_n869));
  OAI21_X1  g0669(.A(KEYINPUT106), .B1(new_n383), .B2(new_n668), .ZN(new_n870));
  INV_X1    g0670(.A(KEYINPUT106), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n367), .A2(new_n871), .A3(new_n858), .ZN(new_n872));
  NAND2_X1  g0672(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT37), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n386), .A2(new_n367), .ZN(new_n875));
  NAND4_X1  g0675(.A1(new_n873), .A2(new_n874), .A3(new_n875), .A4(new_n867), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n869), .A2(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(KEYINPUT105), .ZN(new_n878));
  INV_X1    g0678(.A(new_n865), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n878), .B1(new_n390), .B2(new_n879), .ZN(new_n880));
  AND3_X1   g0680(.A1(new_n390), .A2(new_n878), .A3(new_n879), .ZN(new_n881));
  OAI211_X1 g0681(.A(new_n877), .B(KEYINPUT38), .C1(new_n880), .C2(new_n881), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n390), .A2(new_n879), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n884), .A2(KEYINPUT105), .ZN(new_n885));
  NAND3_X1  g0685(.A1(new_n390), .A2(new_n878), .A3(new_n879), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  AOI21_X1  g0687(.A(KEYINPUT38), .B1(new_n887), .B2(new_n877), .ZN(new_n888));
  OAI21_X1  g0688(.A(KEYINPUT39), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n889), .A2(KEYINPUT107), .ZN(new_n890));
  INV_X1    g0690(.A(KEYINPUT39), .ZN(new_n891));
  INV_X1    g0691(.A(KEYINPUT38), .ZN(new_n892));
  NAND3_X1  g0692(.A1(new_n873), .A2(new_n875), .A3(new_n867), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(KEYINPUT37), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT108), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n894), .A2(new_n895), .A3(new_n876), .ZN(new_n896));
  NAND3_X1  g0696(.A1(new_n390), .A2(new_n872), .A3(new_n870), .ZN(new_n897));
  NAND2_X1  g0697(.A1(new_n896), .A2(new_n897), .ZN(new_n898));
  AOI21_X1  g0698(.A(new_n895), .B1(new_n894), .B2(new_n876), .ZN(new_n899));
  OAI21_X1  g0699(.A(new_n892), .B1(new_n898), .B2(new_n899), .ZN(new_n900));
  AOI22_X1  g0700(.A1(new_n885), .A2(new_n886), .B1(new_n876), .B2(new_n869), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT109), .B1(new_n901), .B2(KEYINPUT38), .ZN(new_n902));
  INV_X1    g0702(.A(KEYINPUT109), .ZN(new_n903));
  NOR2_X1   g0703(.A1(new_n882), .A2(new_n903), .ZN(new_n904));
  OAI211_X1 g0704(.A(new_n891), .B(new_n900), .C1(new_n902), .C2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT107), .ZN(new_n906));
  OAI211_X1 g0706(.A(new_n906), .B(KEYINPUT39), .C1(new_n883), .C2(new_n888), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n890), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  OR2_X1    g0708(.A1(new_n422), .A2(new_n670), .ZN(new_n909));
  INV_X1    g0709(.A(new_n909), .ZN(new_n910));
  AOI21_X1  g0710(.A(new_n859), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n404), .A2(new_n670), .ZN(new_n912));
  NAND3_X1  g0712(.A1(new_n422), .A2(new_n424), .A3(new_n912), .ZN(new_n913));
  OAI211_X1 g0713(.A(new_n404), .B(new_n670), .C1(new_n420), .C2(new_n421), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g0715(.A(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n628), .ZN(new_n917));
  OAI21_X1  g0717(.A(new_n917), .B1(new_n649), .B2(new_n650), .ZN(new_n918));
  AOI211_X1 g0718(.A(KEYINPUT91), .B(new_n645), .C1(new_n647), .C2(new_n648), .ZN(new_n919));
  OAI211_X1 g0719(.A(new_n686), .B(new_n820), .C1(new_n918), .C2(new_n919), .ZN(new_n920));
  INV_X1    g0720(.A(new_n819), .ZN(new_n921));
  AOI21_X1  g0721(.A(new_n916), .B1(new_n920), .B2(new_n921), .ZN(new_n922));
  NOR2_X1   g0722(.A1(new_n883), .A2(new_n888), .ZN(new_n923));
  INV_X1    g0723(.A(new_n923), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n922), .A2(new_n924), .ZN(new_n925));
  AND2_X1   g0725(.A1(new_n911), .A2(new_n925), .ZN(new_n926));
  OAI211_X1 g0726(.A(new_n710), .B(new_n686), .C1(new_n918), .C2(new_n919), .ZN(new_n927));
  INV_X1    g0727(.A(new_n711), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n444), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n661), .A2(new_n295), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  XNOR2_X1  g0731(.A(new_n926), .B(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n900), .B1(new_n902), .B2(new_n904), .ZN(new_n933));
  NOR3_X1   g0733(.A1(new_n625), .A2(new_n582), .A3(new_n670), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n732), .A2(new_n726), .ZN(new_n935));
  OAI211_X1 g0735(.A(new_n820), .B(new_n915), .C1(new_n934), .C2(new_n935), .ZN(new_n936));
  INV_X1    g0736(.A(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n933), .A2(KEYINPUT40), .A3(new_n937), .ZN(new_n938));
  INV_X1    g0738(.A(KEYINPUT40), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n923), .B2(new_n936), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n938), .A2(new_n940), .ZN(new_n941));
  NOR2_X1   g0741(.A1(new_n934), .A2(new_n935), .ZN(new_n942));
  OAI21_X1  g0742(.A(new_n941), .B1(new_n444), .B2(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(new_n444), .ZN(new_n944));
  INV_X1    g0744(.A(new_n942), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n938), .A2(new_n944), .A3(new_n945), .A4(new_n940), .ZN(new_n946));
  NAND3_X1  g0746(.A1(new_n943), .A2(G330), .A3(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n932), .A2(new_n947), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n948), .B1(new_n208), .B2(new_n742), .ZN(new_n949));
  NOR2_X1   g0749(.A1(new_n932), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n857), .B1(new_n949), .B2(new_n950), .ZN(G367));
  INV_X1    g0751(.A(new_n758), .ZN(new_n952));
  OAI221_X1 g0752(.A(new_n752), .B1(new_n212), .B2(new_n427), .C1(new_n952), .C2(new_n243), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n953), .A2(new_n745), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n565), .A2(new_n569), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n955), .A2(new_n670), .ZN(new_n956));
  NAND2_X1  g0756(.A1(new_n581), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g0757(.A(new_n957), .B1(new_n580), .B2(new_n956), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n791), .A2(new_n350), .ZN(new_n959));
  OAI21_X1  g0759(.A(new_n280), .B1(new_n778), .B2(new_n262), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n959), .B(new_n960), .C1(G143), .C2(new_n776), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n770), .A2(G68), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n786), .A2(G159), .ZN(new_n963));
  OAI22_X1  g0763(.A1(new_n202), .A2(new_n781), .B1(new_n789), .B2(new_n205), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(G137), .B2(new_n795), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n961), .A2(new_n962), .A3(new_n963), .A4(new_n965), .ZN(new_n966));
  OAI211_X1 g0766(.A(new_n792), .B(G116), .C1(KEYINPUT112), .C2(KEYINPUT46), .ZN(new_n967));
  NAND2_X1  g0767(.A1(KEYINPUT112), .A2(KEYINPUT46), .ZN(new_n968));
  XOR2_X1   g0768(.A(new_n967), .B(new_n968), .Z(new_n969));
  NAND2_X1  g0769(.A1(new_n786), .A2(G294), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n779), .A2(G303), .ZN(new_n971));
  XOR2_X1   g0771(.A(KEYINPUT111), .B(G311), .Z(new_n972));
  AOI22_X1  g0772(.A1(new_n776), .A2(new_n972), .B1(new_n798), .B2(G283), .ZN(new_n973));
  NAND4_X1  g0773(.A1(new_n969), .A2(new_n970), .A3(new_n971), .A4(new_n973), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n789), .A2(new_n503), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G317), .B2(new_n795), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(new_n313), .C1(new_n460), .C2(new_n769), .ZN(new_n977));
  OAI21_X1  g0777(.A(new_n966), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  XOR2_X1   g0778(.A(new_n978), .B(KEYINPUT47), .Z(new_n979));
  OAI221_X1 g0779(.A(new_n954), .B1(new_n958), .B2(new_n812), .C1(new_n979), .C2(new_n809), .ZN(new_n980));
  INV_X1    g0780(.A(KEYINPUT110), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT45), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n670), .B1(new_n636), .B2(new_n638), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n983), .A2(new_n543), .A3(new_n538), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n632), .A2(new_n670), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(new_n986), .ZN(new_n987));
  NOR3_X1   g0787(.A1(new_n688), .A2(new_n982), .A3(new_n987), .ZN(new_n988));
  AOI21_X1  g0788(.A(KEYINPUT45), .B1(new_n689), .B2(new_n986), .ZN(new_n989));
  INV_X1    g0789(.A(KEYINPUT44), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n689), .A2(new_n990), .A3(new_n986), .ZN(new_n991));
  AOI21_X1  g0791(.A(KEYINPUT44), .B1(new_n688), .B2(new_n987), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n988), .A2(new_n989), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XNOR2_X1  g0793(.A(new_n683), .B(new_n993), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n685), .B1(new_n679), .B2(new_n684), .ZN(new_n995));
  XOR2_X1   g0795(.A(new_n995), .B(new_n674), .Z(new_n996));
  INV_X1    g0796(.A(new_n996), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n739), .B1(new_n994), .B2(new_n997), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n692), .B(KEYINPUT41), .Z(new_n999));
  OAI21_X1  g0799(.A(new_n981), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n993), .B(new_n682), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n740), .B1(new_n1001), .B2(new_n996), .ZN(new_n1002));
  INV_X1    g0802(.A(new_n999), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1002), .A2(KEYINPUT110), .A3(new_n1003), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n744), .B1(new_n1000), .B2(new_n1004), .ZN(new_n1005));
  AND2_X1   g0805(.A1(new_n986), .A2(new_n702), .ZN(new_n1006));
  OAI21_X1  g0806(.A(new_n686), .B1(new_n1006), .B2(new_n629), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n987), .A2(new_n685), .A3(KEYINPUT42), .ZN(new_n1008));
  OAI21_X1  g0808(.A(KEYINPUT42), .B1(new_n987), .B2(new_n685), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  NAND2_X1  g0810(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1011));
  NAND2_X1  g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g0812(.A1(new_n958), .A2(KEYINPUT43), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1012), .B(new_n1013), .Z(new_n1014));
  NOR2_X1   g0814(.A1(new_n683), .A2(new_n987), .ZN(new_n1015));
  XNOR2_X1  g0815(.A(new_n1014), .B(new_n1015), .ZN(new_n1016));
  OAI21_X1  g0816(.A(new_n980), .B1(new_n1005), .B2(new_n1016), .ZN(G387));
  NOR2_X1   g0817(.A1(new_n739), .A2(new_n996), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n1018), .ZN(new_n1019));
  NAND2_X1  g0819(.A1(new_n739), .A2(new_n996), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n1019), .A2(new_n692), .A3(new_n1020), .ZN(new_n1021));
  OR3_X1    g0821(.A1(new_n996), .A2(KEYINPUT113), .A3(new_n743), .ZN(new_n1022));
  OAI21_X1  g0822(.A(KEYINPUT113), .B1(new_n996), .B2(new_n743), .ZN(new_n1023));
  NAND3_X1  g0823(.A1(new_n676), .A2(new_n678), .A3(new_n751), .ZN(new_n1024));
  OAI22_X1  g0824(.A1(new_n695), .A2(new_n753), .B1(G107), .B2(new_n212), .ZN(new_n1025));
  INV_X1    g0825(.A(new_n240), .ZN(new_n1026));
  NAND2_X1  g0826(.A1(new_n1026), .A2(G45), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT114), .ZN(new_n1028));
  AOI211_X1 g0828(.A(G45), .B(new_n694), .C1(G68), .C2(G77), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n256), .A2(new_n202), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT50), .Z(new_n1031));
  AOI21_X1  g0831(.A(new_n952), .B1(new_n1029), .B2(new_n1031), .ZN(new_n1032));
  AOI21_X1  g0832(.A(new_n1025), .B1(new_n1028), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n752), .ZN(new_n1034));
  OAI21_X1  g0834(.A(new_n745), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n313), .B(new_n975), .C1(G77), .C2(new_n792), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n786), .A2(new_n256), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n770), .A2(new_n574), .ZN(new_n1038));
  OAI22_X1  g0838(.A1(new_n775), .A2(new_n353), .B1(new_n781), .B2(new_n225), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n778), .A2(new_n202), .B1(new_n766), .B2(new_n262), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND4_X1  g0841(.A1(new_n1036), .A2(new_n1037), .A3(new_n1038), .A4(new_n1041), .ZN(new_n1042));
  AOI22_X1  g0842(.A1(G322), .A2(new_n776), .B1(new_n779), .B2(G317), .ZN(new_n1043));
  OAI21_X1  g0843(.A(new_n1043), .B1(new_n801), .B2(new_n781), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1044), .B1(new_n786), .B2(new_n972), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT48), .ZN(new_n1046));
  INV_X1    g0846(.A(G294), .ZN(new_n1047));
  OAI22_X1  g0847(.A1(new_n791), .A2(new_n1047), .B1(new_n769), .B2(new_n804), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n1045), .B2(KEYINPUT48), .ZN(new_n1049));
  NAND3_X1  g0849(.A1(new_n1046), .A2(KEYINPUT49), .A3(new_n1049), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(G116), .A2(new_n839), .B1(new_n795), .B2(G326), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n313), .A3(new_n1051), .ZN(new_n1052));
  AOI21_X1  g0852(.A(KEYINPUT49), .B1(new_n1046), .B2(new_n1049), .ZN(new_n1053));
  OAI21_X1  g0853(.A(new_n1042), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g0854(.A(KEYINPUT115), .ZN(new_n1055));
  OR2_X1    g0855(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n809), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1057));
  AOI21_X1  g0857(.A(new_n1035), .B1(new_n1056), .B2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(new_n1022), .A2(new_n1023), .B1(new_n1024), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1021), .A2(new_n1059), .ZN(G393));
  NAND2_X1  g0860(.A1(new_n1019), .A2(new_n1001), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n693), .B1(new_n1018), .B2(new_n994), .ZN(new_n1062));
  AND2_X1   g0862(.A1(new_n1061), .A2(new_n1062), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n248), .A2(new_n952), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n752), .B1(new_n503), .B2(new_n212), .ZN(new_n1065));
  OAI21_X1  g0865(.A(new_n745), .B1(new_n1064), .B2(new_n1065), .ZN(new_n1066));
  OAI22_X1  g0866(.A1(new_n257), .A2(new_n781), .B1(new_n225), .B2(new_n791), .ZN(new_n1067));
  AOI211_X1 g0867(.A(new_n828), .B(new_n1067), .C1(G143), .C2(new_n795), .ZN(new_n1068));
  OAI22_X1  g0868(.A1(new_n775), .A2(new_n262), .B1(new_n778), .B2(new_n353), .ZN(new_n1069));
  XNOR2_X1  g0869(.A(new_n1069), .B(KEYINPUT51), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n786), .A2(G50), .ZN(new_n1071));
  AOI21_X1  g0871(.A(new_n313), .B1(G77), .B2(new_n770), .ZN(new_n1072));
  NAND4_X1  g0872(.A1(new_n1068), .A2(new_n1070), .A3(new_n1071), .A4(new_n1072), .ZN(new_n1073));
  AOI22_X1  g0873(.A1(G317), .A2(new_n776), .B1(new_n779), .B2(G311), .ZN(new_n1074));
  XNOR2_X1  g0874(.A(new_n1074), .B(KEYINPUT52), .ZN(new_n1075));
  AOI211_X1 g0875(.A(new_n280), .B(new_n790), .C1(G116), .C2(new_n770), .ZN(new_n1076));
  OAI22_X1  g0876(.A1(new_n791), .A2(new_n804), .B1(new_n766), .B2(new_n803), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n1077), .B1(G294), .B2(new_n798), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1076), .B(new_n1078), .C1(new_n801), .C2(new_n785), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1073), .B1(new_n1075), .B2(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1066), .B1(new_n1080), .B2(new_n748), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n1081), .B1(new_n986), .B2(new_n812), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1001), .B2(new_n743), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1063), .A2(new_n1083), .ZN(new_n1084));
  INV_X1    g0884(.A(new_n1084), .ZN(G390));
  AND3_X1   g0885(.A1(new_n890), .A2(new_n905), .A3(new_n907), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1086), .A2(new_n749), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n775), .A2(new_n804), .B1(new_n789), .B2(new_n225), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n280), .B(new_n1088), .C1(G87), .C2(new_n792), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n770), .A2(G77), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n786), .A2(new_n432), .ZN(new_n1091));
  OAI22_X1  g0891(.A1(new_n781), .A2(new_n503), .B1(new_n766), .B2(new_n1047), .ZN(new_n1092));
  AOI21_X1  g0892(.A(new_n1092), .B1(G116), .B2(new_n779), .ZN(new_n1093));
  NAND4_X1  g0893(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1093), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n769), .A2(new_n353), .ZN(new_n1095));
  AOI211_X1 g0895(.A(new_n434), .B(new_n1095), .C1(G125), .C2(new_n795), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n791), .A2(new_n262), .ZN(new_n1097));
  XNOR2_X1  g0897(.A(new_n1097), .B(KEYINPUT53), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n786), .A2(G137), .ZN(new_n1099));
  INV_X1    g0899(.A(G128), .ZN(new_n1100));
  OAI22_X1  g0900(.A1(new_n775), .A2(new_n1100), .B1(new_n778), .B2(new_n836), .ZN(new_n1101));
  XNOR2_X1  g0901(.A(KEYINPUT54), .B(G143), .ZN(new_n1102));
  OAI22_X1  g0902(.A1(new_n1102), .A2(new_n781), .B1(new_n789), .B2(new_n202), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n1101), .A2(new_n1103), .ZN(new_n1104));
  NAND4_X1  g0904(.A1(new_n1096), .A2(new_n1098), .A3(new_n1099), .A4(new_n1104), .ZN(new_n1105));
  AOI21_X1  g0905(.A(new_n809), .B1(new_n1094), .B2(new_n1105), .ZN(new_n1106));
  AOI211_X1 g0906(.A(new_n845), .B(new_n1106), .C1(new_n257), .C2(new_n846), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1087), .A2(new_n1107), .ZN(new_n1108));
  OAI21_X1  g0908(.A(new_n1086), .B1(new_n922), .B2(new_n910), .ZN(new_n1109));
  INV_X1    g0909(.A(new_n818), .ZN(new_n1110));
  AOI21_X1  g0910(.A(new_n819), .B1(new_n709), .B2(new_n1110), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1111), .A2(new_n916), .ZN(new_n1112));
  NAND3_X1  g0912(.A1(new_n1112), .A2(new_n909), .A3(new_n933), .ZN(new_n1113));
  NAND4_X1  g0913(.A1(new_n737), .A2(G330), .A3(new_n820), .A4(new_n915), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1109), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1115));
  AND3_X1   g0915(.A1(new_n1112), .A2(new_n909), .A3(new_n933), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n819), .B1(new_n712), .B2(new_n820), .ZN(new_n1117));
  OAI21_X1  g0917(.A(new_n909), .B1(new_n1117), .B2(new_n916), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n1116), .B1(new_n1118), .B2(new_n1086), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n937), .A2(G330), .ZN(new_n1120));
  OAI21_X1  g0920(.A(new_n1115), .B1(new_n1119), .B2(new_n1120), .ZN(new_n1121));
  OAI21_X1  g0921(.A(new_n1108), .B1(new_n1121), .B2(new_n743), .ZN(new_n1122));
  INV_X1    g0922(.A(G330), .ZN(new_n1123));
  NOR3_X1   g0923(.A1(new_n444), .A2(new_n942), .A3(new_n1123), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1124), .ZN(new_n1125));
  OAI211_X1 g0925(.A(new_n662), .B(new_n1125), .C1(new_n713), .C2(new_n444), .ZN(new_n1126));
  OAI211_X1 g0926(.A(G330), .B(new_n820), .C1(new_n934), .C2(new_n935), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1127), .A2(new_n916), .ZN(new_n1128));
  AND3_X1   g0928(.A1(new_n1114), .A2(new_n1128), .A3(new_n1111), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n920), .A2(new_n921), .ZN(new_n1130));
  NAND3_X1  g0930(.A1(new_n737), .A2(G330), .A3(new_n820), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n1131), .A2(new_n916), .ZN(new_n1132));
  NAND2_X1  g0932(.A1(new_n1132), .A2(new_n1120), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1129), .B1(new_n1130), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g0934(.A(KEYINPUT116), .ZN(new_n1135));
  NOR3_X1   g0935(.A1(new_n1126), .A2(new_n1134), .A3(new_n1135), .ZN(new_n1136));
  NOR3_X1   g0936(.A1(new_n929), .A2(new_n930), .A3(new_n1124), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n1130), .A2(new_n1133), .ZN(new_n1138));
  INV_X1    g0938(.A(new_n1129), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1138), .A2(new_n1139), .ZN(new_n1140));
  AOI21_X1  g0940(.A(KEYINPUT116), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NOR2_X1   g0941(.A1(new_n1136), .A2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n693), .B1(new_n1142), .B2(new_n1121), .ZN(new_n1143));
  AND3_X1   g0943(.A1(new_n1109), .A2(new_n1113), .A3(new_n1114), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1120), .B1(new_n1109), .B2(new_n1113), .ZN(new_n1145));
  NOR2_X1   g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1135), .B1(new_n1126), .B2(new_n1134), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1137), .A2(new_n1140), .A3(KEYINPUT116), .ZN(new_n1148));
  NAND2_X1  g0948(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  NAND2_X1  g0949(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n1122), .B1(new_n1143), .B2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(G378));
  NAND2_X1  g0952(.A1(new_n270), .A2(new_n858), .ZN(new_n1153));
  XNOR2_X1  g0953(.A(new_n296), .B(new_n1153), .ZN(new_n1154));
  XNOR2_X1  g0954(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1155));
  XNOR2_X1  g0955(.A(new_n1154), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g0956(.A(new_n1156), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n1157), .A2(new_n749), .ZN(new_n1158));
  AOI211_X1 g0958(.A(G33), .B(G41), .C1(new_n795), .C2(G124), .ZN(new_n1159));
  INV_X1    g0959(.A(new_n1102), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(G125), .A2(new_n776), .B1(new_n792), .B2(new_n1160), .ZN(new_n1161));
  OAI221_X1 g0961(.A(new_n1161), .B1(new_n1100), .B2(new_n778), .C1(new_n262), .C2(new_n769), .ZN(new_n1162));
  AOI22_X1  g0962(.A1(new_n786), .A2(G132), .B1(G137), .B2(new_n798), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT118), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(KEYINPUT118), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1162), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(KEYINPUT59), .ZN(new_n1167));
  OAI221_X1 g0967(.A(new_n1159), .B1(new_n353), .B2(new_n789), .C1(new_n1166), .C2(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1168), .B1(new_n1167), .B2(new_n1166), .ZN(new_n1169));
  OAI221_X1 g0969(.A(new_n962), .B1(new_n350), .B2(new_n789), .C1(new_n589), .C2(new_n775), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n795), .A2(G283), .ZN(new_n1171));
  OAI221_X1 g0971(.A(new_n1171), .B1(new_n458), .B2(new_n778), .C1(new_n427), .C2(new_n781), .ZN(new_n1172));
  AOI211_X1 g0972(.A(new_n1170), .B(new_n1172), .C1(G97), .C2(new_n786), .ZN(new_n1173));
  OR2_X1    g0973(.A1(new_n302), .A2(G41), .ZN(new_n1174));
  AOI21_X1  g0974(.A(new_n1174), .B1(G77), .B2(new_n792), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(KEYINPUT117), .ZN(new_n1176));
  OR2_X1    g0976(.A1(new_n1175), .A2(KEYINPUT117), .ZN(new_n1177));
  NAND3_X1  g0977(.A1(new_n1173), .A2(new_n1176), .A3(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT58), .ZN(new_n1179));
  OR2_X1    g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND2_X1  g0980(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1181));
  OAI211_X1 g0981(.A(new_n1174), .B(new_n202), .C1(G33), .C2(G41), .ZN(new_n1182));
  NAND3_X1  g0982(.A1(new_n1180), .A2(new_n1181), .A3(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n748), .B1(new_n1169), .B2(new_n1183), .ZN(new_n1184));
  XOR2_X1   g0984(.A(new_n1184), .B(KEYINPUT119), .Z(new_n1185));
  AOI211_X1 g0985(.A(new_n845), .B(new_n1185), .C1(new_n202), .C2(new_n846), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1158), .A2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(KEYINPUT120), .ZN(new_n1189));
  OAI21_X1  g0989(.A(new_n1157), .B1(new_n941), .B2(new_n1123), .ZN(new_n1190));
  NAND4_X1  g0990(.A1(new_n1156), .A2(new_n938), .A3(G330), .A4(new_n940), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n1189), .B1(new_n1190), .B2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n911), .A2(new_n925), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1192), .B(new_n1193), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1188), .B1(new_n1194), .B2(new_n744), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1126), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n926), .A2(new_n1191), .A3(new_n1190), .ZN(new_n1197));
  NAND2_X1  g0997(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1198), .A2(new_n1193), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1197), .A2(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1200), .A2(KEYINPUT57), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n692), .B1(new_n1196), .B2(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1137), .B1(new_n1142), .B2(new_n1121), .ZN(new_n1203));
  AOI21_X1  g1003(.A(KEYINPUT57), .B1(new_n1203), .B2(new_n1194), .ZN(new_n1204));
  OAI21_X1  g1004(.A(new_n1195), .B1(new_n1202), .B2(new_n1204), .ZN(G375));
  NAND2_X1  g1005(.A1(new_n916), .A2(new_n749), .ZN(new_n1206));
  XNOR2_X1  g1006(.A(new_n1206), .B(KEYINPUT121), .ZN(new_n1207));
  NOR3_X1   g1007(.A1(new_n748), .A2(G68), .A3(new_n749), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n302), .B1(new_n202), .B2(new_n769), .ZN(new_n1209));
  OAI22_X1  g1009(.A1(new_n350), .A2(new_n789), .B1(new_n781), .B2(new_n262), .ZN(new_n1210));
  OAI22_X1  g1010(.A1(new_n791), .A2(new_n353), .B1(new_n766), .B2(new_n1100), .ZN(new_n1211));
  NOR3_X1   g1011(.A1(new_n1209), .A2(new_n1210), .A3(new_n1211), .ZN(new_n1212));
  XOR2_X1   g1012(.A(new_n1212), .B(KEYINPUT123), .Z(new_n1213));
  AOI22_X1  g1013(.A1(G132), .A2(new_n776), .B1(new_n779), .B2(G137), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n785), .B2(new_n1102), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n280), .B1(new_n839), .B2(G77), .ZN(new_n1216));
  XNOR2_X1  g1016(.A(new_n1216), .B(KEYINPUT122), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n786), .A2(G116), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n503), .A2(new_n791), .B1(new_n778), .B2(new_n804), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1219), .B1(G303), .B2(new_n795), .ZN(new_n1220));
  AOI22_X1  g1020(.A1(G294), .A2(new_n776), .B1(new_n798), .B2(new_n432), .ZN(new_n1221));
  NAND4_X1  g1021(.A1(new_n1218), .A2(new_n1220), .A3(new_n1038), .A4(new_n1221), .ZN(new_n1222));
  OAI22_X1  g1022(.A1(new_n1213), .A2(new_n1215), .B1(new_n1217), .B2(new_n1222), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n845), .B(new_n1208), .C1(new_n1223), .C2(new_n748), .ZN(new_n1224));
  AOI22_X1  g1024(.A1(new_n1140), .A2(new_n744), .B1(new_n1207), .B2(new_n1224), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1126), .A2(new_n1134), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n1147), .A2(new_n1148), .A3(new_n1226), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1225), .B1(new_n1227), .B2(new_n999), .ZN(G381));
  OAI211_X1 g1028(.A(new_n1151), .B(new_n1195), .C1(new_n1202), .C2(new_n1204), .ZN(new_n1229));
  OAI211_X1 g1029(.A(new_n1084), .B(new_n980), .C1(new_n1005), .C2(new_n1016), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(G393), .A2(G396), .ZN(new_n1231));
  INV_X1    g1031(.A(G384), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1233));
  OR4_X1    g1033(.A1(G381), .A2(new_n1229), .A3(new_n1230), .A4(new_n1233), .ZN(G407));
  NAND2_X1  g1034(.A1(new_n669), .A2(G213), .ZN(new_n1235));
  OAI211_X1 g1035(.A(G407), .B(G213), .C1(new_n1229), .C2(new_n1235), .ZN(G409));
  NAND3_X1  g1036(.A1(new_n669), .A2(G213), .A3(G2897), .ZN(new_n1237));
  XOR2_X1   g1037(.A(new_n1237), .B(KEYINPUT125), .Z(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(KEYINPUT60), .ZN(new_n1240));
  AOI21_X1  g1040(.A(new_n693), .B1(new_n1226), .B2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(new_n1227), .ZN(new_n1242));
  OAI21_X1  g1042(.A(new_n1241), .B1(new_n1242), .B2(new_n1240), .ZN(new_n1243));
  NAND3_X1  g1043(.A1(new_n1243), .A2(G384), .A3(new_n1225), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(G384), .B1(new_n1243), .B2(new_n1225), .ZN(new_n1246));
  OAI21_X1  g1046(.A(new_n1239), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1246), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(new_n1244), .A3(new_n1238), .ZN(new_n1249));
  NAND2_X1  g1049(.A1(new_n1247), .A2(new_n1249), .ZN(new_n1250));
  NAND3_X1  g1050(.A1(new_n1203), .A2(new_n1003), .A3(new_n1194), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1188), .B1(new_n1200), .B2(new_n744), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1151), .A2(new_n1251), .A3(new_n1252), .ZN(new_n1253));
  XNOR2_X1  g1053(.A(new_n1192), .B(new_n926), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1187), .B1(new_n1254), .B2(new_n743), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT57), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n1256), .B1(new_n1196), .B2(new_n1254), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1197), .B2(new_n1199), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n693), .B1(new_n1203), .B2(new_n1258), .ZN(new_n1259));
  AOI21_X1  g1059(.A(new_n1255), .B1(new_n1257), .B2(new_n1259), .ZN(new_n1260));
  OAI211_X1 g1060(.A(new_n1235), .B(new_n1253), .C1(new_n1260), .C2(new_n1151), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT61), .B1(new_n1250), .B2(new_n1261), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1253), .A2(new_n1235), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(G375), .A2(G378), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1265));
  NAND3_X1  g1065(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1266), .A2(KEYINPUT62), .ZN(new_n1267));
  INV_X1    g1067(.A(KEYINPUT62), .ZN(new_n1268));
  NAND4_X1  g1068(.A1(new_n1263), .A2(new_n1264), .A3(new_n1265), .A4(new_n1268), .ZN(new_n1269));
  NAND3_X1  g1069(.A1(new_n1262), .A2(new_n1267), .A3(new_n1269), .ZN(new_n1270));
  NAND2_X1  g1070(.A1(G387), .A2(G390), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n814), .B1(new_n1021), .B2(new_n1059), .ZN(new_n1272));
  OAI21_X1  g1072(.A(KEYINPUT126), .B1(new_n1231), .B2(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1271), .A2(new_n1230), .A3(new_n1273), .ZN(new_n1274));
  NOR3_X1   g1074(.A1(new_n1231), .A2(KEYINPUT126), .A3(new_n1272), .ZN(new_n1275));
  NAND2_X1  g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  INV_X1    g1076(.A(new_n1275), .ZN(new_n1277));
  NAND4_X1  g1077(.A1(new_n1277), .A2(new_n1271), .A3(new_n1230), .A4(new_n1273), .ZN(new_n1278));
  NAND2_X1  g1078(.A1(new_n1276), .A2(new_n1278), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1270), .A2(new_n1279), .ZN(new_n1280));
  INV_X1    g1080(.A(KEYINPUT63), .ZN(new_n1281));
  OR2_X1    g1081(.A1(new_n1266), .A2(new_n1281), .ZN(new_n1282));
  NAND2_X1  g1082(.A1(new_n1261), .A2(KEYINPUT124), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT124), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1263), .A2(new_n1264), .A3(new_n1284), .ZN(new_n1285));
  NAND3_X1  g1085(.A1(new_n1283), .A2(new_n1250), .A3(new_n1285), .ZN(new_n1286));
  NOR2_X1   g1086(.A1(new_n1279), .A2(KEYINPUT61), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1266), .A2(new_n1281), .ZN(new_n1288));
  NAND4_X1  g1088(.A1(new_n1282), .A2(new_n1286), .A3(new_n1287), .A4(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1280), .A2(new_n1289), .ZN(G405));
  INV_X1    g1090(.A(KEYINPUT127), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1229), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1257), .A2(new_n1259), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1151), .B1(new_n1293), .B2(new_n1195), .ZN(new_n1294));
  OAI21_X1  g1094(.A(new_n1291), .B1(new_n1292), .B2(new_n1294), .ZN(new_n1295));
  INV_X1    g1095(.A(new_n1265), .ZN(new_n1296));
  NAND3_X1  g1096(.A1(new_n1264), .A2(KEYINPUT127), .A3(new_n1229), .ZN(new_n1297));
  AND3_X1   g1097(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1296), .B1(new_n1295), .B2(new_n1297), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1279), .B1(new_n1298), .B2(new_n1299), .ZN(new_n1300));
  INV_X1    g1100(.A(new_n1297), .ZN(new_n1301));
  AOI21_X1  g1101(.A(KEYINPUT127), .B1(new_n1264), .B2(new_n1229), .ZN(new_n1302));
  OAI21_X1  g1102(.A(new_n1265), .B1(new_n1301), .B2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1279), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1295), .A2(new_n1296), .A3(new_n1297), .ZN(new_n1305));
  NAND3_X1  g1105(.A1(new_n1303), .A2(new_n1304), .A3(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1300), .A2(new_n1306), .ZN(G402));
endmodule


