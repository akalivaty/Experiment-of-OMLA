

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X1 U549 ( .A1(n672), .A2(n671), .ZN(n635) );
  NOR2_X1 U550 ( .A1(n627), .A2(n626), .ZN(n628) );
  NOR2_X1 U551 ( .A1(n717), .A2(G1966), .ZN(n621) );
  NOR2_X1 U552 ( .A1(G2104), .A2(G2105), .ZN(n516) );
  NOR2_X1 U553 ( .A1(n717), .A2(n716), .ZN(n514) );
  XOR2_X2 U554 ( .A(KEYINPUT17), .B(n516), .Z(n895) );
  AND2_X1 U555 ( .A1(n711), .A2(n710), .ZN(n515) );
  XNOR2_X1 U556 ( .A(KEYINPUT30), .B(KEYINPUT100), .ZN(n623) );
  XNOR2_X1 U557 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U558 ( .A(KEYINPUT102), .B(KEYINPUT32), .ZN(n690) );
  XNOR2_X1 U559 ( .A(n691), .B(n690), .ZN(n721) );
  INV_X1 U560 ( .A(KEYINPUT13), .ZN(n641) );
  XNOR2_X1 U561 ( .A(n642), .B(n641), .ZN(n643) );
  AND2_X1 U562 ( .A1(n517), .A2(G2104), .ZN(n897) );
  NOR2_X1 U563 ( .A1(G651), .A2(G543), .ZN(n797) );
  NOR2_X1 U564 ( .A1(n517), .A2(G2104), .ZN(n892) );
  NOR2_X1 U565 ( .A1(G651), .A2(n588), .ZN(n794) );
  INV_X1 U566 ( .A(KEYINPUT65), .ZN(n533) );
  NAND2_X1 U567 ( .A1(n895), .A2(G138), .ZN(n520) );
  INV_X1 U568 ( .A(G2105), .ZN(n517) );
  NAND2_X1 U569 ( .A1(G102), .A2(n897), .ZN(n518) );
  XOR2_X1 U570 ( .A(KEYINPUT91), .B(n518), .Z(n519) );
  NAND2_X1 U571 ( .A1(n520), .A2(n519), .ZN(n524) );
  AND2_X1 U572 ( .A1(G2104), .A2(G2105), .ZN(n891) );
  NAND2_X1 U573 ( .A1(G114), .A2(n891), .ZN(n522) );
  NAND2_X1 U574 ( .A1(G126), .A2(n892), .ZN(n521) );
  NAND2_X1 U575 ( .A1(n522), .A2(n521), .ZN(n523) );
  NOR2_X1 U576 ( .A1(n524), .A2(n523), .ZN(G164) );
  NAND2_X1 U577 ( .A1(n897), .A2(G101), .ZN(n525) );
  XOR2_X1 U578 ( .A(KEYINPUT23), .B(n525), .Z(n527) );
  NAND2_X1 U579 ( .A1(n892), .A2(G125), .ZN(n526) );
  NAND2_X1 U580 ( .A1(n527), .A2(n526), .ZN(n528) );
  XNOR2_X1 U581 ( .A(n528), .B(KEYINPUT66), .ZN(n532) );
  NAND2_X1 U582 ( .A1(G137), .A2(n895), .ZN(n530) );
  NAND2_X1 U583 ( .A1(G113), .A2(n891), .ZN(n529) );
  NAND2_X1 U584 ( .A1(n530), .A2(n529), .ZN(n531) );
  NOR2_X1 U585 ( .A1(n532), .A2(n531), .ZN(n534) );
  XNOR2_X1 U586 ( .A(n534), .B(n533), .ZN(n615) );
  BUF_X1 U587 ( .A(n615), .Z(G160) );
  NAND2_X1 U588 ( .A1(G85), .A2(n797), .ZN(n536) );
  XOR2_X1 U589 ( .A(G543), .B(KEYINPUT0), .Z(n588) );
  INV_X1 U590 ( .A(G651), .ZN(n537) );
  NOR2_X1 U591 ( .A1(n588), .A2(n537), .ZN(n798) );
  NAND2_X1 U592 ( .A1(G72), .A2(n798), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n542) );
  NOR2_X1 U594 ( .A1(G543), .A2(n537), .ZN(n538) );
  XOR2_X1 U595 ( .A(KEYINPUT1), .B(n538), .Z(n793) );
  NAND2_X1 U596 ( .A1(G60), .A2(n793), .ZN(n540) );
  NAND2_X1 U597 ( .A1(G47), .A2(n794), .ZN(n539) );
  NAND2_X1 U598 ( .A1(n540), .A2(n539), .ZN(n541) );
  OR2_X1 U599 ( .A1(n542), .A2(n541), .ZN(G290) );
  NAND2_X1 U600 ( .A1(G64), .A2(n793), .ZN(n544) );
  NAND2_X1 U601 ( .A1(G52), .A2(n794), .ZN(n543) );
  NAND2_X1 U602 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U603 ( .A(KEYINPUT67), .B(n545), .Z(n551) );
  NAND2_X1 U604 ( .A1(n798), .A2(G77), .ZN(n546) );
  XNOR2_X1 U605 ( .A(n546), .B(KEYINPUT68), .ZN(n548) );
  NAND2_X1 U606 ( .A1(G90), .A2(n797), .ZN(n547) );
  NAND2_X1 U607 ( .A1(n548), .A2(n547), .ZN(n549) );
  XOR2_X1 U608 ( .A(KEYINPUT9), .B(n549), .Z(n550) );
  NOR2_X1 U609 ( .A1(n551), .A2(n550), .ZN(G171) );
  NAND2_X1 U610 ( .A1(G89), .A2(n797), .ZN(n552) );
  XNOR2_X1 U611 ( .A(n552), .B(KEYINPUT78), .ZN(n553) );
  XNOR2_X1 U612 ( .A(n553), .B(KEYINPUT4), .ZN(n555) );
  NAND2_X1 U613 ( .A1(G76), .A2(n798), .ZN(n554) );
  NAND2_X1 U614 ( .A1(n555), .A2(n554), .ZN(n556) );
  XNOR2_X1 U615 ( .A(KEYINPUT5), .B(n556), .ZN(n563) );
  XNOR2_X1 U616 ( .A(KEYINPUT6), .B(KEYINPUT80), .ZN(n561) );
  NAND2_X1 U617 ( .A1(n793), .A2(G63), .ZN(n559) );
  NAND2_X1 U618 ( .A1(n794), .A2(G51), .ZN(n557) );
  XOR2_X1 U619 ( .A(KEYINPUT79), .B(n557), .Z(n558) );
  NAND2_X1 U620 ( .A1(n559), .A2(n558), .ZN(n560) );
  XOR2_X1 U621 ( .A(n561), .B(n560), .Z(n562) );
  NAND2_X1 U622 ( .A1(n563), .A2(n562), .ZN(n564) );
  XNOR2_X1 U623 ( .A(KEYINPUT7), .B(n564), .ZN(G168) );
  NAND2_X1 U624 ( .A1(n797), .A2(G91), .ZN(n565) );
  XOR2_X1 U625 ( .A(KEYINPUT69), .B(n565), .Z(n567) );
  NAND2_X1 U626 ( .A1(n798), .A2(G78), .ZN(n566) );
  NAND2_X1 U627 ( .A1(n567), .A2(n566), .ZN(n568) );
  XOR2_X1 U628 ( .A(KEYINPUT70), .B(n568), .Z(n572) );
  NAND2_X1 U629 ( .A1(G65), .A2(n793), .ZN(n570) );
  NAND2_X1 U630 ( .A1(G53), .A2(n794), .ZN(n569) );
  AND2_X1 U631 ( .A1(n570), .A2(n569), .ZN(n571) );
  NAND2_X1 U632 ( .A1(n572), .A2(n571), .ZN(G299) );
  NAND2_X1 U633 ( .A1(G88), .A2(n797), .ZN(n574) );
  NAND2_X1 U634 ( .A1(G75), .A2(n798), .ZN(n573) );
  NAND2_X1 U635 ( .A1(n574), .A2(n573), .ZN(n577) );
  NAND2_X1 U636 ( .A1(n794), .A2(G50), .ZN(n575) );
  XOR2_X1 U637 ( .A(KEYINPUT86), .B(n575), .Z(n576) );
  NOR2_X1 U638 ( .A1(n577), .A2(n576), .ZN(n579) );
  NAND2_X1 U639 ( .A1(n793), .A2(G62), .ZN(n578) );
  NAND2_X1 U640 ( .A1(n579), .A2(n578), .ZN(G303) );
  XOR2_X1 U641 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U642 ( .A1(G73), .A2(n798), .ZN(n580) );
  XOR2_X1 U643 ( .A(KEYINPUT2), .B(n580), .Z(n585) );
  NAND2_X1 U644 ( .A1(G86), .A2(n797), .ZN(n582) );
  NAND2_X1 U645 ( .A1(G61), .A2(n793), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT85), .B(n583), .Z(n584) );
  NOR2_X1 U648 ( .A1(n585), .A2(n584), .ZN(n587) );
  NAND2_X1 U649 ( .A1(n794), .A2(G48), .ZN(n586) );
  NAND2_X1 U650 ( .A1(n587), .A2(n586), .ZN(G305) );
  NAND2_X1 U651 ( .A1(G74), .A2(G651), .ZN(n593) );
  NAND2_X1 U652 ( .A1(G49), .A2(n794), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G87), .A2(n588), .ZN(n589) );
  NAND2_X1 U654 ( .A1(n590), .A2(n589), .ZN(n591) );
  NOR2_X1 U655 ( .A1(n793), .A2(n591), .ZN(n592) );
  NAND2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n594) );
  XNOR2_X1 U657 ( .A(n594), .B(KEYINPUT84), .ZN(G288) );
  NOR2_X1 U658 ( .A1(G164), .A2(G1384), .ZN(n613) );
  NAND2_X1 U659 ( .A1(G160), .A2(G40), .ZN(n595) );
  NOR2_X1 U660 ( .A1(n613), .A2(n595), .ZN(n760) );
  NAND2_X1 U661 ( .A1(G105), .A2(n897), .ZN(n596) );
  XNOR2_X1 U662 ( .A(n596), .B(KEYINPUT38), .ZN(n603) );
  NAND2_X1 U663 ( .A1(G141), .A2(n895), .ZN(n598) );
  NAND2_X1 U664 ( .A1(G129), .A2(n892), .ZN(n597) );
  NAND2_X1 U665 ( .A1(n598), .A2(n597), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G117), .A2(n891), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT95), .B(n599), .ZN(n600) );
  NOR2_X1 U668 ( .A1(n601), .A2(n600), .ZN(n602) );
  NAND2_X1 U669 ( .A1(n603), .A2(n602), .ZN(n886) );
  NAND2_X1 U670 ( .A1(G1996), .A2(n886), .ZN(n611) );
  NAND2_X1 U671 ( .A1(G131), .A2(n895), .ZN(n605) );
  NAND2_X1 U672 ( .A1(G119), .A2(n892), .ZN(n604) );
  NAND2_X1 U673 ( .A1(n605), .A2(n604), .ZN(n609) );
  NAND2_X1 U674 ( .A1(G95), .A2(n897), .ZN(n607) );
  NAND2_X1 U675 ( .A1(G107), .A2(n891), .ZN(n606) );
  NAND2_X1 U676 ( .A1(n607), .A2(n606), .ZN(n608) );
  OR2_X1 U677 ( .A1(n609), .A2(n608), .ZN(n874) );
  NAND2_X1 U678 ( .A1(G1991), .A2(n874), .ZN(n610) );
  NAND2_X1 U679 ( .A1(n611), .A2(n610), .ZN(n930) );
  NAND2_X1 U680 ( .A1(n760), .A2(n930), .ZN(n752) );
  XNOR2_X1 U681 ( .A(G1986), .B(G290), .ZN(n976) );
  NAND2_X1 U682 ( .A1(n760), .A2(n976), .ZN(n612) );
  NAND2_X1 U683 ( .A1(n752), .A2(n612), .ZN(n735) );
  AND2_X1 U684 ( .A1(G40), .A2(n613), .ZN(n614) );
  NAND2_X1 U685 ( .A1(n615), .A2(n614), .ZN(n616) );
  XNOR2_X1 U686 ( .A(n616), .B(KEYINPUT64), .ZN(n620) );
  INV_X1 U687 ( .A(n620), .ZN(n617) );
  INV_X2 U688 ( .A(n617), .ZN(n680) );
  XNOR2_X1 U689 ( .A(G2078), .B(KEYINPUT25), .ZN(n950) );
  NOR2_X1 U690 ( .A1(n680), .A2(n950), .ZN(n619) );
  INV_X1 U691 ( .A(n680), .ZN(n663) );
  INV_X1 U692 ( .A(G1961), .ZN(n1017) );
  NOR2_X1 U693 ( .A1(n663), .A2(n1017), .ZN(n618) );
  NOR2_X1 U694 ( .A1(n619), .A2(n618), .ZN(n629) );
  NOR2_X1 U695 ( .A1(G171), .A2(n629), .ZN(n627) );
  NOR2_X1 U696 ( .A1(n680), .A2(G2084), .ZN(n697) );
  NAND2_X1 U697 ( .A1(n620), .A2(G8), .ZN(n717) );
  XNOR2_X1 U698 ( .A(n621), .B(KEYINPUT96), .ZN(n695) );
  NOR2_X1 U699 ( .A1(n697), .A2(n695), .ZN(n622) );
  NAND2_X1 U700 ( .A1(n622), .A2(G8), .ZN(n624) );
  NOR2_X1 U701 ( .A1(G168), .A2(n625), .ZN(n626) );
  XOR2_X1 U702 ( .A(KEYINPUT31), .B(n628), .Z(n692) );
  NAND2_X1 U703 ( .A1(G171), .A2(n629), .ZN(n679) );
  NAND2_X1 U704 ( .A1(G2072), .A2(n663), .ZN(n630) );
  XNOR2_X1 U705 ( .A(n630), .B(KEYINPUT27), .ZN(n632) );
  AND2_X1 U706 ( .A1(n680), .A2(G1956), .ZN(n631) );
  NOR2_X1 U707 ( .A1(n632), .A2(n631), .ZN(n672) );
  INV_X1 U708 ( .A(G299), .ZN(n671) );
  XNOR2_X1 U709 ( .A(KEYINPUT28), .B(KEYINPUT98), .ZN(n633) );
  XNOR2_X1 U710 ( .A(n633), .B(KEYINPUT97), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n635), .B(n634), .ZN(n676) );
  NAND2_X1 U712 ( .A1(n793), .A2(G56), .ZN(n636) );
  XOR2_X1 U713 ( .A(KEYINPUT14), .B(n636), .Z(n644) );
  NAND2_X1 U714 ( .A1(G81), .A2(n797), .ZN(n637) );
  XOR2_X1 U715 ( .A(KEYINPUT12), .B(n637), .Z(n638) );
  XNOR2_X1 U716 ( .A(n638), .B(KEYINPUT71), .ZN(n640) );
  NAND2_X1 U717 ( .A1(G68), .A2(n798), .ZN(n639) );
  NAND2_X1 U718 ( .A1(n640), .A2(n639), .ZN(n642) );
  NOR2_X1 U719 ( .A1(n644), .A2(n643), .ZN(n645) );
  XNOR2_X1 U720 ( .A(n645), .B(KEYINPUT72), .ZN(n647) );
  NAND2_X1 U721 ( .A1(G43), .A2(n794), .ZN(n646) );
  NAND2_X1 U722 ( .A1(n647), .A2(n646), .ZN(n648) );
  XOR2_X2 U723 ( .A(KEYINPUT73), .B(n648), .Z(n970) );
  XNOR2_X1 U724 ( .A(G1996), .B(KEYINPUT99), .ZN(n949) );
  NOR2_X1 U725 ( .A1(n680), .A2(n949), .ZN(n649) );
  XOR2_X1 U726 ( .A(n649), .B(KEYINPUT26), .Z(n651) );
  NAND2_X1 U727 ( .A1(n680), .A2(G1341), .ZN(n650) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U729 ( .A1(n970), .A2(n652), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n793), .A2(G66), .ZN(n653) );
  XOR2_X1 U731 ( .A(KEYINPUT75), .B(n653), .Z(n655) );
  NAND2_X1 U732 ( .A1(n797), .A2(G92), .ZN(n654) );
  NAND2_X1 U733 ( .A1(n655), .A2(n654), .ZN(n656) );
  XNOR2_X1 U734 ( .A(KEYINPUT76), .B(n656), .ZN(n660) );
  NAND2_X1 U735 ( .A1(G79), .A2(n798), .ZN(n658) );
  NAND2_X1 U736 ( .A1(G54), .A2(n794), .ZN(n657) );
  NAND2_X1 U737 ( .A1(n658), .A2(n657), .ZN(n659) );
  NOR2_X1 U738 ( .A1(n660), .A2(n659), .ZN(n661) );
  XOR2_X1 U739 ( .A(KEYINPUT15), .B(n661), .Z(n662) );
  XNOR2_X1 U740 ( .A(KEYINPUT77), .B(n662), .ZN(n768) );
  NAND2_X1 U741 ( .A1(G2067), .A2(n663), .ZN(n665) );
  NAND2_X1 U742 ( .A1(n680), .A2(G1348), .ZN(n664) );
  NAND2_X1 U743 ( .A1(n665), .A2(n664), .ZN(n668) );
  NOR2_X1 U744 ( .A1(n768), .A2(n668), .ZN(n666) );
  OR2_X1 U745 ( .A1(n667), .A2(n666), .ZN(n670) );
  NAND2_X1 U746 ( .A1(n768), .A2(n668), .ZN(n669) );
  NAND2_X1 U747 ( .A1(n670), .A2(n669), .ZN(n674) );
  NAND2_X1 U748 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U749 ( .A1(n674), .A2(n673), .ZN(n675) );
  NAND2_X1 U750 ( .A1(n676), .A2(n675), .ZN(n677) );
  XOR2_X1 U751 ( .A(KEYINPUT29), .B(n677), .Z(n678) );
  NAND2_X1 U752 ( .A1(n679), .A2(n678), .ZN(n693) );
  NOR2_X1 U753 ( .A1(n680), .A2(G2090), .ZN(n682) );
  NOR2_X1 U754 ( .A1(G1971), .A2(n717), .ZN(n681) );
  NOR2_X1 U755 ( .A1(n682), .A2(n681), .ZN(n683) );
  NAND2_X1 U756 ( .A1(n683), .A2(G303), .ZN(n685) );
  AND2_X1 U757 ( .A1(n693), .A2(n685), .ZN(n684) );
  NAND2_X1 U758 ( .A1(n692), .A2(n684), .ZN(n689) );
  INV_X1 U759 ( .A(n685), .ZN(n686) );
  OR2_X1 U760 ( .A1(n686), .A2(G286), .ZN(n687) );
  AND2_X1 U761 ( .A1(n687), .A2(G8), .ZN(n688) );
  NAND2_X1 U762 ( .A1(n689), .A2(n688), .ZN(n691) );
  NAND2_X1 U763 ( .A1(n693), .A2(n692), .ZN(n694) );
  XNOR2_X1 U764 ( .A(KEYINPUT101), .B(n694), .ZN(n696) );
  NOR2_X1 U765 ( .A1(n696), .A2(n695), .ZN(n699) );
  NAND2_X1 U766 ( .A1(n697), .A2(G8), .ZN(n698) );
  NAND2_X1 U767 ( .A1(n699), .A2(n698), .ZN(n719) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n700) );
  XOR2_X1 U769 ( .A(n700), .B(KEYINPUT24), .Z(n701) );
  NOR2_X1 U770 ( .A1(n717), .A2(n701), .ZN(n705) );
  OR2_X1 U771 ( .A1(n705), .A2(n717), .ZN(n703) );
  AND2_X1 U772 ( .A1(n719), .A2(n703), .ZN(n702) );
  NAND2_X1 U773 ( .A1(n721), .A2(n702), .ZN(n711) );
  INV_X1 U774 ( .A(n703), .ZN(n709) );
  NOR2_X1 U775 ( .A1(G2090), .A2(G303), .ZN(n704) );
  NAND2_X1 U776 ( .A1(G8), .A2(n704), .ZN(n707) );
  INV_X1 U777 ( .A(n705), .ZN(n706) );
  AND2_X1 U778 ( .A1(n707), .A2(n706), .ZN(n708) );
  OR2_X1 U779 ( .A1(n709), .A2(n708), .ZN(n710) );
  NAND2_X1 U780 ( .A1(G1976), .A2(G288), .ZN(n977) );
  INV_X1 U781 ( .A(n977), .ZN(n724) );
  NOR2_X1 U782 ( .A1(G1976), .A2(G288), .ZN(n979) );
  NAND2_X1 U783 ( .A1(n979), .A2(KEYINPUT33), .ZN(n712) );
  NOR2_X1 U784 ( .A1(n712), .A2(n717), .ZN(n714) );
  XOR2_X1 U785 ( .A(G1981), .B(G305), .Z(n986) );
  INV_X1 U786 ( .A(n986), .ZN(n713) );
  NOR2_X1 U787 ( .A1(n714), .A2(n713), .ZN(n715) );
  AND2_X1 U788 ( .A1(n715), .A2(KEYINPUT33), .ZN(n725) );
  INV_X1 U789 ( .A(n715), .ZN(n716) );
  NOR2_X1 U790 ( .A1(n725), .A2(n514), .ZN(n729) );
  NOR2_X1 U791 ( .A1(n724), .A2(n729), .ZN(n718) );
  AND2_X1 U792 ( .A1(n719), .A2(n718), .ZN(n720) );
  NAND2_X1 U793 ( .A1(n721), .A2(n720), .ZN(n731) );
  NOR2_X1 U794 ( .A1(G1971), .A2(G303), .ZN(n722) );
  NOR2_X1 U795 ( .A1(n979), .A2(n722), .ZN(n723) );
  OR2_X1 U796 ( .A1(n724), .A2(n723), .ZN(n727) );
  INV_X1 U797 ( .A(n725), .ZN(n726) );
  AND2_X1 U798 ( .A1(n727), .A2(n726), .ZN(n728) );
  OR2_X1 U799 ( .A1(n729), .A2(n728), .ZN(n730) );
  AND2_X1 U800 ( .A1(n731), .A2(n730), .ZN(n732) );
  NAND2_X1 U801 ( .A1(n515), .A2(n732), .ZN(n733) );
  XNOR2_X1 U802 ( .A(n733), .B(KEYINPUT103), .ZN(n734) );
  NOR2_X1 U803 ( .A1(n735), .A2(n734), .ZN(n748) );
  XNOR2_X1 U804 ( .A(KEYINPUT92), .B(KEYINPUT34), .ZN(n739) );
  NAND2_X1 U805 ( .A1(G104), .A2(n897), .ZN(n737) );
  NAND2_X1 U806 ( .A1(G140), .A2(n895), .ZN(n736) );
  NAND2_X1 U807 ( .A1(n737), .A2(n736), .ZN(n738) );
  XNOR2_X1 U808 ( .A(n739), .B(n738), .ZN(n745) );
  NAND2_X1 U809 ( .A1(n892), .A2(G128), .ZN(n740) );
  XOR2_X1 U810 ( .A(KEYINPUT93), .B(n740), .Z(n742) );
  NAND2_X1 U811 ( .A1(n891), .A2(G116), .ZN(n741) );
  NAND2_X1 U812 ( .A1(n742), .A2(n741), .ZN(n743) );
  XOR2_X1 U813 ( .A(KEYINPUT35), .B(n743), .Z(n744) );
  NOR2_X1 U814 ( .A1(n745), .A2(n744), .ZN(n746) );
  XNOR2_X1 U815 ( .A(KEYINPUT36), .B(n746), .ZN(n905) );
  XNOR2_X1 U816 ( .A(G2067), .B(KEYINPUT37), .ZN(n758) );
  NOR2_X1 U817 ( .A1(n905), .A2(n758), .ZN(n747) );
  XNOR2_X1 U818 ( .A(KEYINPUT94), .B(n747), .ZN(n943) );
  NAND2_X1 U819 ( .A1(n760), .A2(n943), .ZN(n757) );
  NAND2_X1 U820 ( .A1(n748), .A2(n757), .ZN(n749) );
  XNOR2_X1 U821 ( .A(n749), .B(KEYINPUT104), .ZN(n763) );
  NOR2_X1 U822 ( .A1(G1986), .A2(G290), .ZN(n750) );
  NOR2_X1 U823 ( .A1(G1991), .A2(n874), .ZN(n926) );
  NOR2_X1 U824 ( .A1(n750), .A2(n926), .ZN(n751) );
  XNOR2_X1 U825 ( .A(n751), .B(KEYINPUT105), .ZN(n753) );
  NAND2_X1 U826 ( .A1(n753), .A2(n752), .ZN(n754) );
  OR2_X1 U827 ( .A1(n886), .A2(G1996), .ZN(n931) );
  NAND2_X1 U828 ( .A1(n754), .A2(n931), .ZN(n755) );
  XOR2_X1 U829 ( .A(KEYINPUT39), .B(n755), .Z(n756) );
  NAND2_X1 U830 ( .A1(n757), .A2(n756), .ZN(n759) );
  NAND2_X1 U831 ( .A1(n905), .A2(n758), .ZN(n935) );
  NAND2_X1 U832 ( .A1(n759), .A2(n935), .ZN(n761) );
  NAND2_X1 U833 ( .A1(n761), .A2(n760), .ZN(n762) );
  NAND2_X1 U834 ( .A1(n763), .A2(n762), .ZN(n764) );
  XNOR2_X1 U835 ( .A(n764), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U836 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U837 ( .A(G57), .ZN(G237) );
  INV_X1 U838 ( .A(G69), .ZN(G235) );
  INV_X1 U839 ( .A(G108), .ZN(G238) );
  INV_X1 U840 ( .A(G120), .ZN(G236) );
  INV_X1 U841 ( .A(G132), .ZN(G219) );
  INV_X1 U842 ( .A(G82), .ZN(G220) );
  NAND2_X1 U843 ( .A1(G7), .A2(G661), .ZN(n765) );
  XNOR2_X1 U844 ( .A(n765), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U845 ( .A(G223), .ZN(n840) );
  NAND2_X1 U846 ( .A1(n840), .A2(G567), .ZN(n766) );
  XOR2_X1 U847 ( .A(KEYINPUT11), .B(n766), .Z(G234) );
  INV_X1 U848 ( .A(n970), .ZN(n767) );
  NAND2_X1 U849 ( .A1(n767), .A2(G860), .ZN(G153) );
  XOR2_X1 U850 ( .A(G171), .B(KEYINPUT74), .Z(G301) );
  NAND2_X1 U851 ( .A1(G868), .A2(G301), .ZN(n770) );
  BUF_X1 U852 ( .A(n768), .Z(n971) );
  INV_X1 U853 ( .A(G868), .ZN(n779) );
  NAND2_X1 U854 ( .A1(n971), .A2(n779), .ZN(n769) );
  NAND2_X1 U855 ( .A1(n770), .A2(n769), .ZN(G284) );
  NOR2_X1 U856 ( .A1(G286), .A2(n779), .ZN(n771) );
  XOR2_X1 U857 ( .A(KEYINPUT81), .B(n771), .Z(n773) );
  NOR2_X1 U858 ( .A1(G868), .A2(G299), .ZN(n772) );
  NOR2_X1 U859 ( .A1(n773), .A2(n772), .ZN(G297) );
  INV_X1 U860 ( .A(G559), .ZN(n777) );
  NOR2_X1 U861 ( .A1(G860), .A2(n777), .ZN(n774) );
  NOR2_X1 U862 ( .A1(n971), .A2(n774), .ZN(n775) );
  XOR2_X1 U863 ( .A(n775), .B(KEYINPUT82), .Z(n776) );
  XNOR2_X1 U864 ( .A(KEYINPUT16), .B(n776), .ZN(G148) );
  INV_X1 U865 ( .A(n971), .ZN(n909) );
  NAND2_X1 U866 ( .A1(n777), .A2(n909), .ZN(n778) );
  NAND2_X1 U867 ( .A1(n778), .A2(G868), .ZN(n781) );
  NAND2_X1 U868 ( .A1(n970), .A2(n779), .ZN(n780) );
  NAND2_X1 U869 ( .A1(n781), .A2(n780), .ZN(G282) );
  NAND2_X1 U870 ( .A1(G123), .A2(n892), .ZN(n782) );
  XOR2_X1 U871 ( .A(KEYINPUT83), .B(n782), .Z(n783) );
  XNOR2_X1 U872 ( .A(n783), .B(KEYINPUT18), .ZN(n785) );
  NAND2_X1 U873 ( .A1(G99), .A2(n897), .ZN(n784) );
  NAND2_X1 U874 ( .A1(n785), .A2(n784), .ZN(n789) );
  NAND2_X1 U875 ( .A1(G135), .A2(n895), .ZN(n787) );
  NAND2_X1 U876 ( .A1(G111), .A2(n891), .ZN(n786) );
  NAND2_X1 U877 ( .A1(n787), .A2(n786), .ZN(n788) );
  NOR2_X1 U878 ( .A1(n789), .A2(n788), .ZN(n925) );
  XNOR2_X1 U879 ( .A(n925), .B(G2096), .ZN(n791) );
  INV_X1 U880 ( .A(G2100), .ZN(n790) );
  NAND2_X1 U881 ( .A1(n791), .A2(n790), .ZN(G156) );
  NAND2_X1 U882 ( .A1(G559), .A2(n909), .ZN(n792) );
  XNOR2_X1 U883 ( .A(n792), .B(n970), .ZN(n811) );
  NOR2_X1 U884 ( .A1(n811), .A2(G860), .ZN(n803) );
  NAND2_X1 U885 ( .A1(G67), .A2(n793), .ZN(n796) );
  NAND2_X1 U886 ( .A1(G55), .A2(n794), .ZN(n795) );
  NAND2_X1 U887 ( .A1(n796), .A2(n795), .ZN(n802) );
  NAND2_X1 U888 ( .A1(G93), .A2(n797), .ZN(n800) );
  NAND2_X1 U889 ( .A1(G80), .A2(n798), .ZN(n799) );
  NAND2_X1 U890 ( .A1(n800), .A2(n799), .ZN(n801) );
  NOR2_X1 U891 ( .A1(n802), .A2(n801), .ZN(n805) );
  XNOR2_X1 U892 ( .A(n803), .B(n805), .ZN(G145) );
  NOR2_X1 U893 ( .A1(G868), .A2(n805), .ZN(n804) );
  XNOR2_X1 U894 ( .A(n804), .B(KEYINPUT87), .ZN(n814) );
  XNOR2_X1 U895 ( .A(n805), .B(G303), .ZN(n806) );
  XNOR2_X1 U896 ( .A(n806), .B(G305), .ZN(n807) );
  XNOR2_X1 U897 ( .A(KEYINPUT19), .B(n807), .ZN(n809) );
  XNOR2_X1 U898 ( .A(G290), .B(G288), .ZN(n808) );
  XNOR2_X1 U899 ( .A(n809), .B(n808), .ZN(n810) );
  XNOR2_X1 U900 ( .A(n810), .B(G299), .ZN(n910) );
  XNOR2_X1 U901 ( .A(n910), .B(n811), .ZN(n812) );
  NAND2_X1 U902 ( .A1(G868), .A2(n812), .ZN(n813) );
  NAND2_X1 U903 ( .A1(n814), .A2(n813), .ZN(n815) );
  XNOR2_X1 U904 ( .A(KEYINPUT88), .B(n815), .ZN(G295) );
  NAND2_X1 U905 ( .A1(G2078), .A2(G2084), .ZN(n816) );
  XOR2_X1 U906 ( .A(KEYINPUT20), .B(n816), .Z(n817) );
  NAND2_X1 U907 ( .A1(G2090), .A2(n817), .ZN(n818) );
  XNOR2_X1 U908 ( .A(KEYINPUT21), .B(n818), .ZN(n819) );
  NAND2_X1 U909 ( .A1(n819), .A2(G2072), .ZN(n820) );
  XOR2_X1 U910 ( .A(KEYINPUT89), .B(n820), .Z(G158) );
  XNOR2_X1 U911 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U912 ( .A1(G220), .A2(G219), .ZN(n821) );
  XOR2_X1 U913 ( .A(KEYINPUT22), .B(n821), .Z(n822) );
  NOR2_X1 U914 ( .A1(G218), .A2(n822), .ZN(n823) );
  NAND2_X1 U915 ( .A1(G96), .A2(n823), .ZN(n844) );
  NAND2_X1 U916 ( .A1(n844), .A2(G2106), .ZN(n828) );
  NOR2_X1 U917 ( .A1(G236), .A2(G238), .ZN(n825) );
  NOR2_X1 U918 ( .A1(G235), .A2(G237), .ZN(n824) );
  NAND2_X1 U919 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U920 ( .A(KEYINPUT90), .B(n826), .ZN(n845) );
  NAND2_X1 U921 ( .A1(n845), .A2(G567), .ZN(n827) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n846) );
  NAND2_X1 U923 ( .A1(G483), .A2(G661), .ZN(n829) );
  NOR2_X1 U924 ( .A1(n846), .A2(n829), .ZN(n843) );
  NAND2_X1 U925 ( .A1(n843), .A2(G36), .ZN(G176) );
  XNOR2_X1 U926 ( .A(G2430), .B(G2454), .ZN(n838) );
  XNOR2_X1 U927 ( .A(KEYINPUT106), .B(G2435), .ZN(n836) );
  XOR2_X1 U928 ( .A(G2451), .B(G2427), .Z(n831) );
  XNOR2_X1 U929 ( .A(G2438), .B(G2446), .ZN(n830) );
  XNOR2_X1 U930 ( .A(n831), .B(n830), .ZN(n832) );
  XOR2_X1 U931 ( .A(n832), .B(G2443), .Z(n834) );
  XNOR2_X1 U932 ( .A(G1341), .B(G1348), .ZN(n833) );
  XNOR2_X1 U933 ( .A(n834), .B(n833), .ZN(n835) );
  XNOR2_X1 U934 ( .A(n836), .B(n835), .ZN(n837) );
  XNOR2_X1 U935 ( .A(n838), .B(n837), .ZN(n839) );
  NAND2_X1 U936 ( .A1(n839), .A2(G14), .ZN(n915) );
  XNOR2_X1 U937 ( .A(KEYINPUT107), .B(n915), .ZN(G401) );
  NAND2_X1 U938 ( .A1(G2106), .A2(n840), .ZN(G217) );
  AND2_X1 U939 ( .A1(G15), .A2(G2), .ZN(n841) );
  NAND2_X1 U940 ( .A1(G661), .A2(n841), .ZN(G259) );
  NAND2_X1 U941 ( .A1(G3), .A2(G1), .ZN(n842) );
  NAND2_X1 U942 ( .A1(n843), .A2(n842), .ZN(G188) );
  NOR2_X1 U943 ( .A1(n845), .A2(n844), .ZN(G325) );
  XOR2_X1 U944 ( .A(KEYINPUT108), .B(G325), .Z(G261) );
  INV_X1 U946 ( .A(G96), .ZN(G221) );
  INV_X1 U947 ( .A(n846), .ZN(G319) );
  XNOR2_X1 U948 ( .A(G1996), .B(KEYINPUT41), .ZN(n856) );
  XOR2_X1 U949 ( .A(G1976), .B(G1956), .Z(n848) );
  XNOR2_X1 U950 ( .A(G1991), .B(G1961), .ZN(n847) );
  XNOR2_X1 U951 ( .A(n848), .B(n847), .ZN(n852) );
  XOR2_X1 U952 ( .A(G1981), .B(G1966), .Z(n850) );
  XNOR2_X1 U953 ( .A(G1986), .B(G1971), .ZN(n849) );
  XNOR2_X1 U954 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U955 ( .A(n852), .B(n851), .Z(n854) );
  XNOR2_X1 U956 ( .A(G2474), .B(KEYINPUT110), .ZN(n853) );
  XNOR2_X1 U957 ( .A(n854), .B(n853), .ZN(n855) );
  XNOR2_X1 U958 ( .A(n856), .B(n855), .ZN(G229) );
  XOR2_X1 U959 ( .A(G2678), .B(G2084), .Z(n858) );
  XNOR2_X1 U960 ( .A(G2078), .B(G2072), .ZN(n857) );
  XNOR2_X1 U961 ( .A(n858), .B(n857), .ZN(n859) );
  XOR2_X1 U962 ( .A(n859), .B(G2100), .Z(n861) );
  XNOR2_X1 U963 ( .A(G2067), .B(G2090), .ZN(n860) );
  XNOR2_X1 U964 ( .A(n861), .B(n860), .ZN(n865) );
  XOR2_X1 U965 ( .A(G2096), .B(KEYINPUT109), .Z(n863) );
  XNOR2_X1 U966 ( .A(KEYINPUT42), .B(KEYINPUT43), .ZN(n862) );
  XNOR2_X1 U967 ( .A(n863), .B(n862), .ZN(n864) );
  XOR2_X1 U968 ( .A(n865), .B(n864), .Z(G227) );
  NAND2_X1 U969 ( .A1(G100), .A2(n897), .ZN(n867) );
  NAND2_X1 U970 ( .A1(G112), .A2(n891), .ZN(n866) );
  NAND2_X1 U971 ( .A1(n867), .A2(n866), .ZN(n868) );
  XNOR2_X1 U972 ( .A(n868), .B(KEYINPUT111), .ZN(n870) );
  NAND2_X1 U973 ( .A1(G136), .A2(n895), .ZN(n869) );
  NAND2_X1 U974 ( .A1(n870), .A2(n869), .ZN(n873) );
  NAND2_X1 U975 ( .A1(n892), .A2(G124), .ZN(n871) );
  XOR2_X1 U976 ( .A(KEYINPUT44), .B(n871), .Z(n872) );
  NOR2_X1 U977 ( .A1(n873), .A2(n872), .ZN(G162) );
  XNOR2_X1 U978 ( .A(KEYINPUT46), .B(KEYINPUT48), .ZN(n876) );
  XNOR2_X1 U979 ( .A(n874), .B(KEYINPUT113), .ZN(n875) );
  XNOR2_X1 U980 ( .A(n876), .B(n875), .ZN(n877) );
  XNOR2_X1 U981 ( .A(G162), .B(n877), .ZN(n890) );
  NAND2_X1 U982 ( .A1(G103), .A2(n897), .ZN(n879) );
  NAND2_X1 U983 ( .A1(G139), .A2(n895), .ZN(n878) );
  NAND2_X1 U984 ( .A1(n879), .A2(n878), .ZN(n885) );
  NAND2_X1 U985 ( .A1(G115), .A2(n891), .ZN(n881) );
  NAND2_X1 U986 ( .A1(G127), .A2(n892), .ZN(n880) );
  NAND2_X1 U987 ( .A1(n881), .A2(n880), .ZN(n882) );
  XOR2_X1 U988 ( .A(KEYINPUT47), .B(n882), .Z(n883) );
  XNOR2_X1 U989 ( .A(KEYINPUT114), .B(n883), .ZN(n884) );
  NOR2_X1 U990 ( .A1(n885), .A2(n884), .ZN(n921) );
  XOR2_X1 U991 ( .A(n921), .B(n925), .Z(n888) );
  XOR2_X1 U992 ( .A(G164), .B(n886), .Z(n887) );
  XNOR2_X1 U993 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U994 ( .A(n890), .B(n889), .ZN(n904) );
  NAND2_X1 U995 ( .A1(G118), .A2(n891), .ZN(n894) );
  NAND2_X1 U996 ( .A1(G130), .A2(n892), .ZN(n893) );
  NAND2_X1 U997 ( .A1(n894), .A2(n893), .ZN(n902) );
  NAND2_X1 U998 ( .A1(n895), .A2(G142), .ZN(n896) );
  XNOR2_X1 U999 ( .A(n896), .B(KEYINPUT112), .ZN(n899) );
  NAND2_X1 U1000 ( .A1(G106), .A2(n897), .ZN(n898) );
  NAND2_X1 U1001 ( .A1(n899), .A2(n898), .ZN(n900) );
  XOR2_X1 U1002 ( .A(n900), .B(KEYINPUT45), .Z(n901) );
  NOR2_X1 U1003 ( .A1(n902), .A2(n901), .ZN(n903) );
  XOR2_X1 U1004 ( .A(n904), .B(n903), .Z(n907) );
  XNOR2_X1 U1005 ( .A(n905), .B(G160), .ZN(n906) );
  XNOR2_X1 U1006 ( .A(n907), .B(n906), .ZN(n908) );
  NOR2_X1 U1007 ( .A1(G37), .A2(n908), .ZN(G395) );
  XOR2_X1 U1008 ( .A(n910), .B(n909), .Z(n912) );
  XNOR2_X1 U1009 ( .A(G286), .B(G171), .ZN(n911) );
  XNOR2_X1 U1010 ( .A(n912), .B(n911), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(n913), .B(n970), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(G37), .A2(n914), .ZN(G397) );
  NAND2_X1 U1013 ( .A1(G319), .A2(n915), .ZN(n918) );
  NOR2_X1 U1014 ( .A1(G229), .A2(G227), .ZN(n916) );
  XNOR2_X1 U1015 ( .A(KEYINPUT49), .B(n916), .ZN(n917) );
  NOR2_X1 U1016 ( .A1(n918), .A2(n917), .ZN(n920) );
  NOR2_X1 U1017 ( .A1(G395), .A2(G397), .ZN(n919) );
  NAND2_X1 U1018 ( .A1(n920), .A2(n919), .ZN(G225) );
  INV_X1 U1019 ( .A(G225), .ZN(G308) );
  INV_X1 U1020 ( .A(G303), .ZN(G166) );
  XOR2_X1 U1021 ( .A(G2072), .B(n921), .Z(n923) );
  XOR2_X1 U1022 ( .A(G164), .B(G2078), .Z(n922) );
  NOR2_X1 U1023 ( .A1(n923), .A2(n922), .ZN(n924) );
  XNOR2_X1 U1024 ( .A(KEYINPUT50), .B(n924), .ZN(n928) );
  NOR2_X1 U1025 ( .A1(n926), .A2(n925), .ZN(n927) );
  NAND2_X1 U1026 ( .A1(n928), .A2(n927), .ZN(n929) );
  NOR2_X1 U1027 ( .A1(n930), .A2(n929), .ZN(n941) );
  XNOR2_X1 U1028 ( .A(G2090), .B(G162), .ZN(n932) );
  NAND2_X1 U1029 ( .A1(n932), .A2(n931), .ZN(n933) );
  XNOR2_X1 U1030 ( .A(n933), .B(KEYINPUT116), .ZN(n934) );
  XNOR2_X1 U1031 ( .A(n934), .B(KEYINPUT51), .ZN(n936) );
  NAND2_X1 U1032 ( .A1(n936), .A2(n935), .ZN(n939) );
  XNOR2_X1 U1033 ( .A(G2084), .B(G160), .ZN(n937) );
  XNOR2_X1 U1034 ( .A(KEYINPUT115), .B(n937), .ZN(n938) );
  NOR2_X1 U1035 ( .A1(n939), .A2(n938), .ZN(n940) );
  NAND2_X1 U1036 ( .A1(n941), .A2(n940), .ZN(n942) );
  NOR2_X1 U1037 ( .A1(n943), .A2(n942), .ZN(n944) );
  XOR2_X1 U1038 ( .A(KEYINPUT52), .B(n944), .Z(n945) );
  NOR2_X1 U1039 ( .A1(KEYINPUT55), .A2(n945), .ZN(n946) );
  XNOR2_X1 U1040 ( .A(KEYINPUT117), .B(n946), .ZN(n947) );
  NAND2_X1 U1041 ( .A1(n947), .A2(G29), .ZN(n1030) );
  XOR2_X1 U1042 ( .A(G1991), .B(G25), .Z(n948) );
  NAND2_X1 U1043 ( .A1(n948), .A2(G28), .ZN(n955) );
  XOR2_X1 U1044 ( .A(n949), .B(G32), .Z(n952) );
  XOR2_X1 U1045 ( .A(n950), .B(G27), .Z(n951) );
  NOR2_X1 U1046 ( .A1(n952), .A2(n951), .ZN(n953) );
  XOR2_X1 U1047 ( .A(KEYINPUT118), .B(n953), .Z(n954) );
  NOR2_X1 U1048 ( .A1(n955), .A2(n954), .ZN(n959) );
  XNOR2_X1 U1049 ( .A(G2067), .B(G26), .ZN(n957) );
  XNOR2_X1 U1050 ( .A(G33), .B(G2072), .ZN(n956) );
  NOR2_X1 U1051 ( .A1(n957), .A2(n956), .ZN(n958) );
  NAND2_X1 U1052 ( .A1(n959), .A2(n958), .ZN(n960) );
  XNOR2_X1 U1053 ( .A(n960), .B(KEYINPUT53), .ZN(n963) );
  XOR2_X1 U1054 ( .A(G2084), .B(G34), .Z(n961) );
  XNOR2_X1 U1055 ( .A(KEYINPUT54), .B(n961), .ZN(n962) );
  NAND2_X1 U1056 ( .A1(n963), .A2(n962), .ZN(n965) );
  XNOR2_X1 U1057 ( .A(G35), .B(G2090), .ZN(n964) );
  NOR2_X1 U1058 ( .A1(n965), .A2(n964), .ZN(n966) );
  XNOR2_X1 U1059 ( .A(KEYINPUT55), .B(n966), .ZN(n968) );
  INV_X1 U1060 ( .A(G29), .ZN(n967) );
  NAND2_X1 U1061 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1062 ( .A1(n969), .A2(G11), .ZN(n1028) );
  XNOR2_X1 U1063 ( .A(G16), .B(KEYINPUT56), .ZN(n994) );
  XNOR2_X1 U1064 ( .A(n970), .B(G1341), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n971), .B(G1348), .ZN(n972) );
  NOR2_X1 U1066 ( .A1(n973), .A2(n972), .ZN(n992) );
  XNOR2_X1 U1067 ( .A(G1971), .B(G166), .ZN(n974) );
  XNOR2_X1 U1068 ( .A(n974), .B(KEYINPUT120), .ZN(n985) );
  XNOR2_X1 U1069 ( .A(G1956), .B(G299), .ZN(n975) );
  NOR2_X1 U1070 ( .A1(n976), .A2(n975), .ZN(n978) );
  NAND2_X1 U1071 ( .A1(n978), .A2(n977), .ZN(n983) );
  XNOR2_X1 U1072 ( .A(n979), .B(KEYINPUT119), .ZN(n981) );
  XNOR2_X1 U1073 ( .A(G171), .B(G1961), .ZN(n980) );
  NAND2_X1 U1074 ( .A1(n981), .A2(n980), .ZN(n982) );
  NOR2_X1 U1075 ( .A1(n983), .A2(n982), .ZN(n984) );
  NAND2_X1 U1076 ( .A1(n985), .A2(n984), .ZN(n990) );
  XNOR2_X1 U1077 ( .A(G168), .B(G1966), .ZN(n987) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  XOR2_X1 U1079 ( .A(KEYINPUT57), .B(n988), .Z(n989) );
  NOR2_X1 U1080 ( .A1(n990), .A2(n989), .ZN(n991) );
  NAND2_X1 U1081 ( .A1(n992), .A2(n991), .ZN(n993) );
  NAND2_X1 U1082 ( .A1(n994), .A2(n993), .ZN(n1026) );
  INV_X1 U1083 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1084 ( .A(G1966), .B(G21), .Z(n1009) );
  XNOR2_X1 U1085 ( .A(KEYINPUT121), .B(G1956), .ZN(n995) );
  XNOR2_X1 U1086 ( .A(n995), .B(G20), .ZN(n1004) );
  XOR2_X1 U1087 ( .A(G1341), .B(G19), .Z(n999) );
  XOR2_X1 U1088 ( .A(KEYINPUT59), .B(KEYINPUT123), .Z(n996) );
  XNOR2_X1 U1089 ( .A(G4), .B(n996), .ZN(n997) );
  XNOR2_X1 U1090 ( .A(n997), .B(G1348), .ZN(n998) );
  NAND2_X1 U1091 ( .A1(n999), .A2(n998), .ZN(n1002) );
  XNOR2_X1 U1092 ( .A(KEYINPUT122), .B(G1981), .ZN(n1000) );
  XNOR2_X1 U1093 ( .A(G6), .B(n1000), .ZN(n1001) );
  NOR2_X1 U1094 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1007) );
  XNOR2_X1 U1096 ( .A(KEYINPUT124), .B(KEYINPUT125), .ZN(n1005) );
  XNOR2_X1 U1097 ( .A(n1005), .B(KEYINPUT60), .ZN(n1006) );
  XNOR2_X1 U1098 ( .A(n1007), .B(n1006), .ZN(n1008) );
  NAND2_X1 U1099 ( .A1(n1009), .A2(n1008), .ZN(n1021) );
  XOR2_X1 U1100 ( .A(G1986), .B(G24), .Z(n1012) );
  XOR2_X1 U1101 ( .A(G22), .B(KEYINPUT126), .Z(n1010) );
  XNOR2_X1 U1102 ( .A(n1010), .B(G1971), .ZN(n1011) );
  NAND2_X1 U1103 ( .A1(n1012), .A2(n1011), .ZN(n1015) );
  XOR2_X1 U1104 ( .A(KEYINPUT127), .B(G1976), .Z(n1013) );
  XNOR2_X1 U1105 ( .A(G23), .B(n1013), .ZN(n1014) );
  NOR2_X1 U1106 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1016), .ZN(n1019) );
  XNOR2_X1 U1108 ( .A(n1017), .B(G5), .ZN(n1018) );
  NAND2_X1 U1109 ( .A1(n1019), .A2(n1018), .ZN(n1020) );
  NOR2_X1 U1110 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1111 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1112 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1113 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  NOR2_X1 U1114 ( .A1(n1028), .A2(n1027), .ZN(n1029) );
  NAND2_X1 U1115 ( .A1(n1030), .A2(n1029), .ZN(n1031) );
  XOR2_X1 U1116 ( .A(KEYINPUT62), .B(n1031), .Z(G311) );
  INV_X1 U1117 ( .A(G311), .ZN(G150) );
endmodule

