

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583;

  XOR2_X1 U323 ( .A(n322), .B(KEYINPUT31), .Z(n291) );
  XNOR2_X1 U324 ( .A(n499), .B(KEYINPUT113), .ZN(n500) );
  XNOR2_X1 U325 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT119), .ZN(n542) );
  XNOR2_X1 U327 ( .A(n543), .B(n542), .ZN(n544) );
  XNOR2_X1 U328 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n511) );
  XNOR2_X1 U329 ( .A(n512), .B(n511), .ZN(n541) );
  XNOR2_X1 U330 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U331 ( .A(n332), .B(n331), .ZN(n473) );
  NOR2_X1 U332 ( .A1(n551), .A2(n550), .ZN(n562) );
  XNOR2_X1 U333 ( .A(n314), .B(n313), .ZN(n545) );
  XNOR2_X1 U334 ( .A(G1GAT), .B(KEYINPUT34), .ZN(n446) );
  XOR2_X1 U335 ( .A(KEYINPUT5), .B(G57GAT), .Z(n293) );
  XNOR2_X1 U336 ( .A(G1GAT), .B(G141GAT), .ZN(n292) );
  XNOR2_X1 U337 ( .A(n293), .B(n292), .ZN(n297) );
  XOR2_X1 U338 ( .A(G85GAT), .B(G148GAT), .Z(n295) );
  XNOR2_X1 U339 ( .A(G29GAT), .B(G120GAT), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n296) );
  XNOR2_X1 U341 ( .A(n297), .B(n296), .ZN(n314) );
  XOR2_X1 U342 ( .A(KEYINPUT92), .B(KEYINPUT4), .Z(n299) );
  XNOR2_X1 U343 ( .A(KEYINPUT94), .B(KEYINPUT90), .ZN(n298) );
  XNOR2_X1 U344 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U345 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n301) );
  XNOR2_X1 U346 ( .A(KEYINPUT93), .B(KEYINPUT91), .ZN(n300) );
  XNOR2_X1 U347 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U348 ( .A(n303), .B(n302), .Z(n312) );
  XOR2_X1 U349 ( .A(KEYINPUT3), .B(G162GAT), .Z(n305) );
  XNOR2_X1 U350 ( .A(KEYINPUT2), .B(G155GAT), .ZN(n304) );
  XNOR2_X1 U351 ( .A(n305), .B(n304), .ZN(n306) );
  XOR2_X1 U352 ( .A(KEYINPUT88), .B(n306), .Z(n430) );
  XOR2_X1 U353 ( .A(G134GAT), .B(KEYINPUT79), .Z(n350) );
  XNOR2_X1 U354 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n307) );
  XNOR2_X1 U355 ( .A(n307), .B(G127GAT), .ZN(n404) );
  XOR2_X1 U356 ( .A(n350), .B(n404), .Z(n309) );
  NAND2_X1 U357 ( .A1(G225GAT), .A2(G233GAT), .ZN(n308) );
  XNOR2_X1 U358 ( .A(n309), .B(n308), .ZN(n310) );
  XNOR2_X1 U359 ( .A(n430), .B(n310), .ZN(n311) );
  XNOR2_X1 U360 ( .A(n312), .B(n311), .ZN(n313) );
  XNOR2_X1 U361 ( .A(G176GAT), .B(G92GAT), .ZN(n315) );
  XNOR2_X1 U362 ( .A(n315), .B(G64GAT), .ZN(n389) );
  INV_X1 U363 ( .A(n389), .ZN(n316) );
  XOR2_X1 U364 ( .A(G120GAT), .B(G71GAT), .Z(n403) );
  NAND2_X1 U365 ( .A1(n316), .A2(n403), .ZN(n319) );
  INV_X1 U366 ( .A(n403), .ZN(n317) );
  NAND2_X1 U367 ( .A1(n389), .A2(n317), .ZN(n318) );
  NAND2_X1 U368 ( .A1(n319), .A2(n318), .ZN(n321) );
  NAND2_X1 U369 ( .A1(G230GAT), .A2(G233GAT), .ZN(n320) );
  XNOR2_X1 U370 ( .A(n321), .B(n320), .ZN(n322) );
  XNOR2_X1 U371 ( .A(G99GAT), .B(G85GAT), .ZN(n323) );
  XNOR2_X1 U372 ( .A(n323), .B(KEYINPUT74), .ZN(n349) );
  XNOR2_X1 U373 ( .A(n349), .B(KEYINPUT75), .ZN(n324) );
  XNOR2_X1 U374 ( .A(n291), .B(n324), .ZN(n332) );
  XNOR2_X1 U375 ( .A(G106GAT), .B(G78GAT), .ZN(n325) );
  XNOR2_X1 U376 ( .A(n325), .B(G148GAT), .ZN(n418) );
  XNOR2_X1 U377 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(KEYINPUT73), .ZN(n383) );
  XOR2_X1 U379 ( .A(n418), .B(n383), .Z(n330) );
  XOR2_X1 U380 ( .A(KEYINPUT32), .B(KEYINPUT76), .Z(n328) );
  XNOR2_X1 U381 ( .A(G204GAT), .B(KEYINPUT33), .ZN(n327) );
  XNOR2_X1 U382 ( .A(n328), .B(n327), .ZN(n329) );
  XNOR2_X1 U383 ( .A(G169GAT), .B(G36GAT), .ZN(n333) );
  XNOR2_X1 U384 ( .A(n333), .B(G8GAT), .ZN(n400) );
  XOR2_X1 U385 ( .A(n400), .B(G197GAT), .Z(n335) );
  XOR2_X1 U386 ( .A(G141GAT), .B(G22GAT), .Z(n419) );
  XNOR2_X1 U387 ( .A(G113GAT), .B(n419), .ZN(n334) );
  XNOR2_X1 U388 ( .A(n335), .B(n334), .ZN(n340) );
  XNOR2_X1 U389 ( .A(G15GAT), .B(G1GAT), .ZN(n336) );
  XNOR2_X1 U390 ( .A(n336), .B(KEYINPUT71), .ZN(n384) );
  XOR2_X1 U391 ( .A(n384), .B(KEYINPUT29), .Z(n338) );
  NAND2_X1 U392 ( .A1(G229GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n339) );
  XOR2_X1 U394 ( .A(n340), .B(n339), .Z(n348) );
  XOR2_X1 U395 ( .A(KEYINPUT7), .B(G50GAT), .Z(n342) );
  XNOR2_X1 U396 ( .A(G43GAT), .B(G29GAT), .ZN(n341) );
  XNOR2_X1 U397 ( .A(n342), .B(n341), .ZN(n343) );
  XOR2_X1 U398 ( .A(KEYINPUT8), .B(n343), .Z(n366) );
  XOR2_X1 U399 ( .A(KEYINPUT69), .B(KEYINPUT68), .Z(n345) );
  XNOR2_X1 U400 ( .A(KEYINPUT30), .B(KEYINPUT70), .ZN(n344) );
  XNOR2_X1 U401 ( .A(n345), .B(n344), .ZN(n346) );
  XNOR2_X1 U402 ( .A(n366), .B(n346), .ZN(n347) );
  XNOR2_X1 U403 ( .A(n348), .B(n347), .ZN(n568) );
  XNOR2_X1 U404 ( .A(n568), .B(KEYINPUT72), .ZN(n552) );
  NAND2_X1 U405 ( .A1(n473), .A2(n552), .ZN(n460) );
  XOR2_X1 U406 ( .A(KEYINPUT16), .B(KEYINPUT84), .Z(n388) );
  XOR2_X1 U407 ( .A(n350), .B(n349), .Z(n352) );
  XNOR2_X1 U408 ( .A(G36GAT), .B(G218GAT), .ZN(n351) );
  XNOR2_X1 U409 ( .A(n352), .B(n351), .ZN(n365) );
  XOR2_X1 U410 ( .A(KEYINPUT9), .B(KEYINPUT77), .Z(n354) );
  XNOR2_X1 U411 ( .A(G106GAT), .B(G92GAT), .ZN(n353) );
  XNOR2_X1 U412 ( .A(n354), .B(n353), .ZN(n358) );
  XOR2_X1 U413 ( .A(KEYINPUT67), .B(KEYINPUT10), .Z(n356) );
  XNOR2_X1 U414 ( .A(KEYINPUT11), .B(KEYINPUT78), .ZN(n355) );
  XNOR2_X1 U415 ( .A(n356), .B(n355), .ZN(n357) );
  XOR2_X1 U416 ( .A(n358), .B(n357), .Z(n363) );
  XOR2_X1 U417 ( .A(KEYINPUT80), .B(G162GAT), .Z(n360) );
  NAND2_X1 U418 ( .A1(G232GAT), .A2(G233GAT), .ZN(n359) );
  XNOR2_X1 U419 ( .A(n360), .B(n359), .ZN(n361) );
  XNOR2_X1 U420 ( .A(G190GAT), .B(n361), .ZN(n362) );
  XNOR2_X1 U421 ( .A(n363), .B(n362), .ZN(n364) );
  XNOR2_X1 U422 ( .A(n365), .B(n364), .ZN(n367) );
  XOR2_X1 U423 ( .A(n367), .B(n366), .Z(n454) );
  BUF_X1 U424 ( .A(n454), .Z(n561) );
  XOR2_X1 U425 ( .A(G78GAT), .B(G127GAT), .Z(n369) );
  XNOR2_X1 U426 ( .A(G183GAT), .B(G71GAT), .ZN(n368) );
  XNOR2_X1 U427 ( .A(n369), .B(n368), .ZN(n373) );
  XOR2_X1 U428 ( .A(G64GAT), .B(G211GAT), .Z(n371) );
  XNOR2_X1 U429 ( .A(G22GAT), .B(G155GAT), .ZN(n370) );
  XNOR2_X1 U430 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U431 ( .A(n373), .B(n372), .Z(n378) );
  XOR2_X1 U432 ( .A(KEYINPUT81), .B(KEYINPUT83), .Z(n375) );
  NAND2_X1 U433 ( .A1(G231GAT), .A2(G233GAT), .ZN(n374) );
  XNOR2_X1 U434 ( .A(n375), .B(n374), .ZN(n376) );
  XNOR2_X1 U435 ( .A(KEYINPUT82), .B(n376), .ZN(n377) );
  XNOR2_X1 U436 ( .A(n378), .B(n377), .ZN(n382) );
  XOR2_X1 U437 ( .A(KEYINPUT15), .B(KEYINPUT14), .Z(n380) );
  XNOR2_X1 U438 ( .A(G8GAT), .B(KEYINPUT12), .ZN(n379) );
  XNOR2_X1 U439 ( .A(n380), .B(n379), .ZN(n381) );
  XOR2_X1 U440 ( .A(n382), .B(n381), .Z(n386) );
  XNOR2_X1 U441 ( .A(n384), .B(n383), .ZN(n385) );
  XNOR2_X1 U442 ( .A(n386), .B(n385), .ZN(n521) );
  OR2_X1 U443 ( .A1(n561), .A2(n521), .ZN(n387) );
  XNOR2_X1 U444 ( .A(n388), .B(n387), .ZN(n444) );
  XOR2_X1 U445 ( .A(KEYINPUT95), .B(n389), .Z(n391) );
  NAND2_X1 U446 ( .A1(G226GAT), .A2(G233GAT), .ZN(n390) );
  XNOR2_X1 U447 ( .A(n391), .B(n390), .ZN(n396) );
  XNOR2_X1 U448 ( .A(G211GAT), .B(G218GAT), .ZN(n392) );
  XNOR2_X1 U449 ( .A(n392), .B(KEYINPUT87), .ZN(n393) );
  XOR2_X1 U450 ( .A(n393), .B(KEYINPUT21), .Z(n395) );
  XNOR2_X1 U451 ( .A(G197GAT), .B(G204GAT), .ZN(n394) );
  XNOR2_X1 U452 ( .A(n395), .B(n394), .ZN(n426) );
  XOR2_X1 U453 ( .A(n396), .B(n426), .Z(n402) );
  XOR2_X1 U454 ( .A(KEYINPUT17), .B(G190GAT), .Z(n398) );
  XNOR2_X1 U455 ( .A(KEYINPUT19), .B(G183GAT), .ZN(n397) );
  XNOR2_X1 U456 ( .A(n398), .B(n397), .ZN(n399) );
  XOR2_X1 U457 ( .A(KEYINPUT18), .B(n399), .Z(n417) );
  XNOR2_X1 U458 ( .A(n400), .B(n417), .ZN(n401) );
  XOR2_X1 U459 ( .A(n402), .B(n401), .Z(n539) );
  XOR2_X1 U460 ( .A(n404), .B(n403), .Z(n406) );
  XNOR2_X1 U461 ( .A(G43GAT), .B(G99GAT), .ZN(n405) );
  XNOR2_X1 U462 ( .A(n406), .B(n405), .ZN(n410) );
  XOR2_X1 U463 ( .A(G176GAT), .B(KEYINPUT86), .Z(n408) );
  NAND2_X1 U464 ( .A1(G227GAT), .A2(G233GAT), .ZN(n407) );
  XNOR2_X1 U465 ( .A(n408), .B(n407), .ZN(n409) );
  XOR2_X1 U466 ( .A(n410), .B(n409), .Z(n415) );
  XOR2_X1 U467 ( .A(KEYINPUT85), .B(KEYINPUT20), .Z(n412) );
  XNOR2_X1 U468 ( .A(G15GAT), .B(G134GAT), .ZN(n411) );
  XNOR2_X1 U469 ( .A(n412), .B(n411), .ZN(n413) );
  XNOR2_X1 U470 ( .A(G169GAT), .B(n413), .ZN(n414) );
  XNOR2_X1 U471 ( .A(n415), .B(n414), .ZN(n416) );
  XNOR2_X1 U472 ( .A(n417), .B(n416), .ZN(n550) );
  INV_X1 U473 ( .A(n550), .ZN(n513) );
  NAND2_X1 U474 ( .A1(n539), .A2(n513), .ZN(n431) );
  XOR2_X1 U475 ( .A(KEYINPUT89), .B(n418), .Z(n421) );
  XNOR2_X1 U476 ( .A(G50GAT), .B(n419), .ZN(n420) );
  XNOR2_X1 U477 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U478 ( .A(KEYINPUT24), .B(KEYINPUT23), .Z(n423) );
  NAND2_X1 U479 ( .A1(G228GAT), .A2(G233GAT), .ZN(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U481 ( .A(n425), .B(n424), .Z(n428) );
  XNOR2_X1 U482 ( .A(n426), .B(KEYINPUT22), .ZN(n427) );
  XNOR2_X1 U483 ( .A(n428), .B(n427), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n547) );
  NAND2_X1 U485 ( .A1(n431), .A2(n547), .ZN(n432) );
  XNOR2_X1 U486 ( .A(n432), .B(KEYINPUT97), .ZN(n433) );
  XOR2_X1 U487 ( .A(n433), .B(KEYINPUT25), .Z(n436) );
  XNOR2_X1 U488 ( .A(n539), .B(KEYINPUT27), .ZN(n438) );
  NOR2_X1 U489 ( .A1(n547), .A2(n513), .ZN(n434) );
  XNOR2_X1 U490 ( .A(n434), .B(KEYINPUT26), .ZN(n566) );
  NAND2_X1 U491 ( .A1(n438), .A2(n566), .ZN(n529) );
  XOR2_X1 U492 ( .A(n529), .B(KEYINPUT96), .Z(n435) );
  NOR2_X1 U493 ( .A1(n436), .A2(n435), .ZN(n437) );
  NOR2_X1 U494 ( .A1(n545), .A2(n437), .ZN(n442) );
  INV_X1 U495 ( .A(n438), .ZN(n439) );
  XOR2_X1 U496 ( .A(KEYINPUT28), .B(n547), .Z(n494) );
  NOR2_X1 U497 ( .A1(n439), .A2(n494), .ZN(n440) );
  NAND2_X1 U498 ( .A1(n545), .A2(n440), .ZN(n515) );
  NOR2_X1 U499 ( .A1(n513), .A2(n515), .ZN(n441) );
  NOR2_X1 U500 ( .A1(n442), .A2(n441), .ZN(n456) );
  INV_X1 U501 ( .A(n456), .ZN(n443) );
  NAND2_X1 U502 ( .A1(n444), .A2(n443), .ZN(n475) );
  NOR2_X1 U503 ( .A1(n460), .A2(n475), .ZN(n452) );
  NAND2_X1 U504 ( .A1(n545), .A2(n452), .ZN(n445) );
  XNOR2_X1 U505 ( .A(n446), .B(n445), .ZN(G1324GAT) );
  NAND2_X1 U506 ( .A1(n539), .A2(n452), .ZN(n447) );
  XNOR2_X1 U507 ( .A(n447), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U508 ( .A(KEYINPUT35), .B(KEYINPUT99), .Z(n449) );
  NAND2_X1 U509 ( .A1(n452), .A2(n513), .ZN(n448) );
  XNOR2_X1 U510 ( .A(n449), .B(n448), .ZN(n451) );
  XOR2_X1 U511 ( .A(G15GAT), .B(KEYINPUT98), .Z(n450) );
  XNOR2_X1 U512 ( .A(n451), .B(n450), .ZN(G1326GAT) );
  NAND2_X1 U513 ( .A1(n494), .A2(n452), .ZN(n453) );
  XNOR2_X1 U514 ( .A(n453), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U515 ( .A(KEYINPUT39), .B(KEYINPUT102), .Z(n463) );
  XNOR2_X1 U516 ( .A(KEYINPUT101), .B(KEYINPUT37), .ZN(n459) );
  XOR2_X1 U517 ( .A(n454), .B(KEYINPUT100), .Z(n455) );
  XNOR2_X1 U518 ( .A(n455), .B(KEYINPUT36), .ZN(n580) );
  NOR2_X1 U519 ( .A1(n580), .A2(n456), .ZN(n457) );
  NAND2_X1 U520 ( .A1(n521), .A2(n457), .ZN(n458) );
  XNOR2_X1 U521 ( .A(n459), .B(n458), .ZN(n487) );
  NOR2_X1 U522 ( .A1(n460), .A2(n487), .ZN(n461) );
  XNOR2_X1 U523 ( .A(n461), .B(KEYINPUT38), .ZN(n470) );
  NAND2_X1 U524 ( .A1(n545), .A2(n470), .ZN(n462) );
  XNOR2_X1 U525 ( .A(n463), .B(n462), .ZN(n464) );
  XNOR2_X1 U526 ( .A(G29GAT), .B(n464), .ZN(G1328GAT) );
  XOR2_X1 U527 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n466) );
  NAND2_X1 U528 ( .A1(n470), .A2(n539), .ZN(n465) );
  XNOR2_X1 U529 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U530 ( .A(G36GAT), .B(n467), .ZN(G1329GAT) );
  NAND2_X1 U531 ( .A1(n470), .A2(n513), .ZN(n468) );
  XNOR2_X1 U532 ( .A(n468), .B(KEYINPUT40), .ZN(n469) );
  XNOR2_X1 U533 ( .A(G43GAT), .B(n469), .ZN(G1330GAT) );
  XOR2_X1 U534 ( .A(G50GAT), .B(KEYINPUT105), .Z(n472) );
  NAND2_X1 U535 ( .A1(n470), .A2(n494), .ZN(n471) );
  XNOR2_X1 U536 ( .A(n472), .B(n471), .ZN(G1331GAT) );
  INV_X1 U537 ( .A(n568), .ZN(n474) );
  XNOR2_X1 U538 ( .A(n473), .B(KEYINPUT41), .ZN(n557) );
  NAND2_X1 U539 ( .A1(n474), .A2(n557), .ZN(n488) );
  NOR2_X1 U540 ( .A1(n488), .A2(n475), .ZN(n476) );
  XNOR2_X1 U541 ( .A(KEYINPUT106), .B(n476), .ZN(n482) );
  NAND2_X1 U542 ( .A1(n482), .A2(n545), .ZN(n479) );
  XOR2_X1 U543 ( .A(G57GAT), .B(KEYINPUT42), .Z(n477) );
  XNOR2_X1 U544 ( .A(KEYINPUT107), .B(n477), .ZN(n478) );
  XNOR2_X1 U545 ( .A(n479), .B(n478), .ZN(G1332GAT) );
  NAND2_X1 U546 ( .A1(n482), .A2(n539), .ZN(n480) );
  XNOR2_X1 U547 ( .A(n480), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U548 ( .A1(n482), .A2(n513), .ZN(n481) );
  XNOR2_X1 U549 ( .A(n481), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U550 ( .A(KEYINPUT109), .B(KEYINPUT43), .Z(n484) );
  NAND2_X1 U551 ( .A1(n482), .A2(n494), .ZN(n483) );
  XNOR2_X1 U552 ( .A(n484), .B(n483), .ZN(n486) );
  XOR2_X1 U553 ( .A(G78GAT), .B(KEYINPUT108), .Z(n485) );
  XNOR2_X1 U554 ( .A(n486), .B(n485), .ZN(G1335GAT) );
  NOR2_X1 U555 ( .A1(n488), .A2(n487), .ZN(n489) );
  XNOR2_X1 U556 ( .A(n489), .B(KEYINPUT110), .ZN(n495) );
  NAND2_X1 U557 ( .A1(n545), .A2(n495), .ZN(n490) );
  XNOR2_X1 U558 ( .A(G85GAT), .B(n490), .ZN(G1336GAT) );
  XOR2_X1 U559 ( .A(G92GAT), .B(KEYINPUT111), .Z(n492) );
  NAND2_X1 U560 ( .A1(n495), .A2(n539), .ZN(n491) );
  XNOR2_X1 U561 ( .A(n492), .B(n491), .ZN(G1337GAT) );
  NAND2_X1 U562 ( .A1(n495), .A2(n513), .ZN(n493) );
  XNOR2_X1 U563 ( .A(n493), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U564 ( .A(KEYINPUT44), .B(KEYINPUT112), .Z(n497) );
  NAND2_X1 U565 ( .A1(n495), .A2(n494), .ZN(n496) );
  XNOR2_X1 U566 ( .A(n497), .B(n496), .ZN(n498) );
  XOR2_X1 U567 ( .A(G106GAT), .B(n498), .Z(G1339GAT) );
  AND2_X1 U568 ( .A1(n557), .A2(n568), .ZN(n501) );
  INV_X1 U569 ( .A(KEYINPUT46), .ZN(n499) );
  NOR2_X1 U570 ( .A1(n561), .A2(n502), .ZN(n503) );
  NAND2_X1 U571 ( .A1(n521), .A2(n503), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n504), .B(KEYINPUT47), .ZN(n510) );
  NOR2_X1 U573 ( .A1(n580), .A2(n521), .ZN(n505) );
  XNOR2_X1 U574 ( .A(n505), .B(KEYINPUT45), .ZN(n506) );
  XNOR2_X1 U575 ( .A(n506), .B(KEYINPUT66), .ZN(n507) );
  NAND2_X1 U576 ( .A1(n507), .A2(n473), .ZN(n508) );
  NOR2_X1 U577 ( .A1(n552), .A2(n508), .ZN(n509) );
  NOR2_X1 U578 ( .A1(n510), .A2(n509), .ZN(n512) );
  INV_X1 U579 ( .A(n541), .ZN(n527) );
  NAND2_X1 U580 ( .A1(n513), .A2(n527), .ZN(n514) );
  NOR2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n524) );
  NAND2_X1 U582 ( .A1(n524), .A2(n552), .ZN(n516) );
  XNOR2_X1 U583 ( .A(G113GAT), .B(n516), .ZN(G1340GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT49), .B(KEYINPUT115), .Z(n518) );
  NAND2_X1 U585 ( .A1(n524), .A2(n557), .ZN(n517) );
  XNOR2_X1 U586 ( .A(n518), .B(n517), .ZN(n520) );
  XOR2_X1 U587 ( .A(G120GAT), .B(KEYINPUT114), .Z(n519) );
  XNOR2_X1 U588 ( .A(n520), .B(n519), .ZN(G1341GAT) );
  INV_X1 U589 ( .A(n521), .ZN(n577) );
  NAND2_X1 U590 ( .A1(n577), .A2(n524), .ZN(n522) );
  XNOR2_X1 U591 ( .A(n522), .B(KEYINPUT50), .ZN(n523) );
  XNOR2_X1 U592 ( .A(G127GAT), .B(n523), .ZN(G1342GAT) );
  XOR2_X1 U593 ( .A(G134GAT), .B(KEYINPUT51), .Z(n526) );
  NAND2_X1 U594 ( .A1(n524), .A2(n561), .ZN(n525) );
  XNOR2_X1 U595 ( .A(n526), .B(n525), .ZN(G1343GAT) );
  NAND2_X1 U596 ( .A1(n545), .A2(n527), .ZN(n528) );
  NOR2_X1 U597 ( .A1(n529), .A2(n528), .ZN(n537) );
  NAND2_X1 U598 ( .A1(n537), .A2(n568), .ZN(n530) );
  XNOR2_X1 U599 ( .A(n530), .B(G141GAT), .ZN(G1344GAT) );
  XNOR2_X1 U600 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n534) );
  XOR2_X1 U601 ( .A(KEYINPUT116), .B(KEYINPUT52), .Z(n532) );
  NAND2_X1 U602 ( .A1(n537), .A2(n557), .ZN(n531) );
  XNOR2_X1 U603 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U604 ( .A(n534), .B(n533), .ZN(G1345GAT) );
  XOR2_X1 U605 ( .A(G155GAT), .B(KEYINPUT117), .Z(n536) );
  NAND2_X1 U606 ( .A1(n537), .A2(n577), .ZN(n535) );
  XNOR2_X1 U607 ( .A(n536), .B(n535), .ZN(G1346GAT) );
  NAND2_X1 U608 ( .A1(n561), .A2(n537), .ZN(n538) );
  XNOR2_X1 U609 ( .A(n538), .B(G162GAT), .ZN(G1347GAT) );
  XOR2_X1 U610 ( .A(n539), .B(KEYINPUT118), .Z(n540) );
  NOR2_X1 U611 ( .A1(n541), .A2(n540), .ZN(n543) );
  NOR2_X1 U612 ( .A1(n545), .A2(n544), .ZN(n546) );
  XOR2_X1 U613 ( .A(KEYINPUT65), .B(n546), .Z(n567) );
  NAND2_X1 U614 ( .A1(n567), .A2(n547), .ZN(n549) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(KEYINPUT55), .Z(n548) );
  XNOR2_X1 U616 ( .A(n549), .B(n548), .ZN(n551) );
  NAND2_X1 U617 ( .A1(n562), .A2(n552), .ZN(n553) );
  XNOR2_X1 U618 ( .A(G169GAT), .B(n553), .ZN(G1348GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT57), .B(KEYINPUT122), .Z(n555) );
  XNOR2_X1 U620 ( .A(G176GAT), .B(KEYINPUT121), .ZN(n554) );
  XNOR2_X1 U621 ( .A(n555), .B(n554), .ZN(n556) );
  XOR2_X1 U622 ( .A(KEYINPUT56), .B(n556), .Z(n559) );
  NAND2_X1 U623 ( .A1(n562), .A2(n557), .ZN(n558) );
  XNOR2_X1 U624 ( .A(n559), .B(n558), .ZN(G1349GAT) );
  NAND2_X1 U625 ( .A1(n577), .A2(n562), .ZN(n560) );
  XNOR2_X1 U626 ( .A(n560), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n562), .A2(n561), .ZN(n564) );
  XOR2_X1 U628 ( .A(KEYINPUT123), .B(KEYINPUT58), .Z(n563) );
  XNOR2_X1 U629 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U630 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT124), .ZN(n572) );
  XOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT59), .Z(n570) );
  NAND2_X1 U633 ( .A1(n567), .A2(n566), .ZN(n579) );
  INV_X1 U634 ( .A(n579), .ZN(n576) );
  NAND2_X1 U635 ( .A1(n576), .A2(n568), .ZN(n569) );
  XNOR2_X1 U636 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U637 ( .A(n572), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U638 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n574) );
  OR2_X1 U639 ( .A1(n579), .A2(n473), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(G204GAT), .B(n575), .Z(G1353GAT) );
  NAND2_X1 U642 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U643 ( .A(n578), .B(G211GAT), .ZN(G1354GAT) );
  NOR2_X1 U644 ( .A1(n580), .A2(n579), .ZN(n582) );
  XNOR2_X1 U645 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n581) );
  XNOR2_X1 U646 ( .A(n582), .B(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(G218GAT), .B(n583), .Z(G1355GAT) );
endmodule

