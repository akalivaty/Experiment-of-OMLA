//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 1 0 0 1 1 1 1 0 1 1 1 1 0 1 0 1 0 1 1 1 0 0 0 0 0 0 0 1 0 1 0 0 1 0 1 1 1 1 0 0 1 0 1 0 0 1 1 0 0 0 1 0 1 1 1 0 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:25 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n677, new_n678, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n687, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n694, new_n695, new_n696, new_n697, new_n698, new_n699,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n741, new_n742, new_n743, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n897, new_n898,
    new_n899, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n934, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978;
  INV_X1    g000(.A(KEYINPUT64), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT11), .ZN(new_n188));
  INV_X1    g002(.A(G134), .ZN(new_n189));
  OAI22_X1  g003(.A1(new_n187), .A2(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n190));
  INV_X1    g004(.A(G137), .ZN(new_n191));
  NAND4_X1  g005(.A1(new_n191), .A2(KEYINPUT64), .A3(KEYINPUT11), .A4(G134), .ZN(new_n192));
  AND2_X1   g006(.A1(new_n190), .A2(new_n192), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT65), .ZN(new_n194));
  INV_X1    g008(.A(G131), .ZN(new_n195));
  AOI22_X1  g009(.A1(new_n187), .A2(new_n188), .B1(new_n189), .B2(G137), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n193), .A2(new_n194), .A3(new_n195), .A4(new_n196), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n196), .A2(new_n190), .A3(new_n195), .A4(new_n192), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n193), .A2(new_n196), .ZN(new_n200));
  AOI22_X1  g014(.A1(new_n197), .A2(new_n199), .B1(new_n200), .B2(G131), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT84), .ZN(new_n202));
  NOR2_X1   g016(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G101), .ZN(new_n204));
  INV_X1    g018(.A(G107), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G104), .ZN(new_n206));
  INV_X1    g020(.A(G104), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n207), .A2(G107), .ZN(new_n208));
  AOI21_X1  g022(.A(new_n204), .B1(new_n206), .B2(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G146), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(G143), .ZN(new_n211));
  INV_X1    g025(.A(G143), .ZN(new_n212));
  NAND2_X1  g026(.A1(new_n212), .A2(G146), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT1), .ZN(new_n215));
  AOI21_X1  g029(.A(new_n215), .B1(G143), .B2(new_n210), .ZN(new_n216));
  INV_X1    g030(.A(G128), .ZN(new_n217));
  OAI21_X1  g031(.A(new_n214), .B1(new_n216), .B2(new_n217), .ZN(new_n218));
  XNOR2_X1  g032(.A(G143), .B(G146), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n219), .A2(new_n215), .A3(G128), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n209), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  OAI21_X1  g035(.A(KEYINPUT3), .B1(new_n207), .B2(G107), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n223));
  NAND3_X1  g037(.A1(new_n223), .A2(new_n205), .A3(G104), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(new_n224), .A3(new_n204), .A4(new_n208), .ZN(new_n225));
  AND2_X1   g039(.A1(new_n225), .A2(KEYINPUT82), .ZN(new_n226));
  NOR2_X1   g040(.A1(new_n225), .A2(KEYINPUT82), .ZN(new_n227));
  OAI21_X1  g041(.A(new_n221), .B1(new_n226), .B2(new_n227), .ZN(new_n228));
  OR2_X1    g042(.A1(new_n225), .A2(KEYINPUT82), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n225), .A2(KEYINPUT82), .ZN(new_n230));
  AOI21_X1  g044(.A(new_n209), .B1(new_n229), .B2(new_n230), .ZN(new_n231));
  XNOR2_X1  g045(.A(KEYINPUT68), .B(G128), .ZN(new_n232));
  OAI21_X1  g046(.A(new_n214), .B1(new_n232), .B2(new_n216), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n233), .A2(new_n220), .ZN(new_n234));
  OAI21_X1  g048(.A(new_n228), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n203), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT12), .ZN(new_n237));
  XNOR2_X1  g051(.A(new_n236), .B(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(KEYINPUT10), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n228), .A2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT4), .ZN(new_n241));
  NAND3_X1  g055(.A1(new_n222), .A2(new_n224), .A3(new_n208), .ZN(new_n242));
  AOI21_X1  g056(.A(new_n241), .B1(new_n242), .B2(G101), .ZN(new_n243));
  OAI21_X1  g057(.A(new_n243), .B1(new_n226), .B2(new_n227), .ZN(new_n244));
  AND3_X1   g058(.A1(new_n242), .A2(new_n241), .A3(G101), .ZN(new_n245));
  OR2_X1    g059(.A1(KEYINPUT0), .A2(G128), .ZN(new_n246));
  NAND2_X1  g060(.A1(KEYINPUT0), .A2(G128), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n214), .A2(new_n246), .A3(new_n247), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n219), .A2(KEYINPUT0), .A3(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  NOR2_X1   g064(.A1(new_n245), .A2(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n244), .A2(new_n251), .ZN(new_n252));
  XNOR2_X1  g066(.A(new_n225), .B(KEYINPUT82), .ZN(new_n253));
  INV_X1    g067(.A(new_n209), .ZN(new_n254));
  AOI21_X1  g068(.A(new_n239), .B1(new_n233), .B2(new_n220), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n253), .A2(new_n254), .A3(new_n255), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n240), .A2(new_n252), .A3(new_n201), .A4(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT83), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  AOI22_X1  g073(.A1(new_n239), .A2(new_n228), .B1(new_n244), .B2(new_n251), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n260), .A2(KEYINPUT83), .A3(new_n201), .A4(new_n256), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(G953), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT71), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT71), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G953), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n264), .A2(new_n266), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n267), .A2(G227), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G140), .ZN(new_n269));
  XNOR2_X1  g083(.A(new_n268), .B(new_n269), .ZN(new_n270));
  AOI21_X1  g084(.A(KEYINPUT86), .B1(new_n262), .B2(new_n270), .ZN(new_n271));
  INV_X1    g085(.A(KEYINPUT86), .ZN(new_n272));
  INV_X1    g086(.A(new_n270), .ZN(new_n273));
  AOI211_X1 g087(.A(new_n272), .B(new_n273), .C1(new_n259), .C2(new_n261), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n238), .B1(new_n271), .B2(new_n274), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n275), .A2(KEYINPUT87), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n201), .B1(new_n260), .B2(new_n256), .ZN(new_n277));
  INV_X1    g091(.A(KEYINPUT85), .ZN(new_n278));
  XNOR2_X1  g092(.A(new_n277), .B(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n262), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n280), .A2(new_n273), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT87), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n282), .B(new_n238), .C1(new_n271), .C2(new_n274), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n276), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  NAND2_X1  g101(.A1(new_n238), .A2(new_n262), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n273), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n279), .A2(new_n262), .A3(new_n270), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  INV_X1    g105(.A(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G469), .B1(new_n292), .B2(G902), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n287), .A2(new_n293), .ZN(new_n294));
  XOR2_X1   g108(.A(KEYINPUT9), .B(G234), .Z(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G221), .B1(new_n296), .B2(G902), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n294), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n298), .A2(KEYINPUT88), .ZN(new_n299));
  INV_X1    g113(.A(KEYINPUT88), .ZN(new_n300));
  NAND3_X1  g114(.A1(new_n294), .A2(new_n300), .A3(new_n297), .ZN(new_n301));
  NAND2_X1  g115(.A1(new_n299), .A2(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT32), .ZN(new_n303));
  NOR2_X1   g117(.A1(G472), .A2(G902), .ZN(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT2), .B(G113), .ZN(new_n306));
  INV_X1    g120(.A(G119), .ZN(new_n307));
  OR2_X1    g121(.A1(KEYINPUT69), .A2(G116), .ZN(new_n308));
  NAND2_X1  g122(.A1(KEYINPUT69), .A2(G116), .ZN(new_n309));
  AOI21_X1  g123(.A(new_n307), .B1(new_n308), .B2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(G116), .ZN(new_n311));
  NOR2_X1   g125(.A1(new_n311), .A2(G119), .ZN(new_n312));
  OAI21_X1  g126(.A(new_n306), .B1(new_n310), .B2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(new_n306), .ZN(new_n314));
  INV_X1    g128(.A(new_n309), .ZN(new_n315));
  NOR2_X1   g129(.A1(KEYINPUT69), .A2(G116), .ZN(new_n316));
  OAI21_X1  g130(.A(G119), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  INV_X1    g131(.A(new_n312), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n314), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n313), .A2(new_n319), .ZN(new_n320));
  INV_X1    g134(.A(KEYINPUT67), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n321), .B1(new_n191), .B2(G134), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n189), .A2(KEYINPUT67), .A3(G137), .ZN(new_n323));
  OAI211_X1 g137(.A(new_n322), .B(new_n323), .C1(new_n189), .C2(G137), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n324), .A2(G131), .ZN(new_n325));
  AND2_X1   g139(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n326));
  NOR2_X1   g140(.A1(new_n198), .A2(KEYINPUT65), .ZN(new_n327));
  OAI211_X1 g141(.A(new_n325), .B(new_n234), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  OAI211_X1 g142(.A(new_n328), .B(KEYINPUT30), .C1(new_n201), .C2(new_n250), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT70), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g145(.A(new_n329), .ZN(new_n332));
  OAI21_X1  g146(.A(KEYINPUT66), .B1(new_n201), .B2(new_n250), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n200), .A2(G131), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n334), .B1(new_n326), .B2(new_n327), .ZN(new_n335));
  INV_X1    g149(.A(KEYINPUT66), .ZN(new_n336));
  INV_X1    g150(.A(new_n250), .ZN(new_n337));
  NAND3_X1  g151(.A1(new_n335), .A2(new_n336), .A3(new_n337), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n333), .A2(new_n338), .A3(new_n328), .ZN(new_n339));
  INV_X1    g153(.A(KEYINPUT30), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n332), .B1(new_n339), .B2(new_n340), .ZN(new_n341));
  OAI211_X1 g155(.A(new_n320), .B(new_n331), .C1(new_n341), .C2(new_n330), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n335), .A2(new_n337), .ZN(new_n343));
  INV_X1    g157(.A(new_n320), .ZN(new_n344));
  NAND3_X1  g158(.A1(new_n343), .A2(new_n344), .A3(new_n328), .ZN(new_n345));
  INV_X1    g159(.A(G237), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n267), .A2(G210), .A3(new_n346), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n347), .B(new_n204), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n349));
  XOR2_X1   g163(.A(new_n348), .B(new_n349), .Z(new_n350));
  NAND3_X1  g164(.A1(new_n342), .A2(new_n345), .A3(new_n350), .ZN(new_n351));
  INV_X1    g165(.A(new_n350), .ZN(new_n352));
  INV_X1    g166(.A(new_n345), .ZN(new_n353));
  OR2_X1    g167(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n339), .A2(new_n320), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n353), .A2(KEYINPUT28), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n354), .A2(new_n355), .A3(new_n356), .ZN(new_n357));
  AOI22_X1  g171(.A1(new_n351), .A2(KEYINPUT31), .B1(new_n352), .B2(new_n357), .ZN(new_n358));
  INV_X1    g172(.A(KEYINPUT31), .ZN(new_n359));
  NAND4_X1  g173(.A1(new_n342), .A2(new_n359), .A3(new_n345), .A4(new_n350), .ZN(new_n360));
  AOI211_X1 g174(.A(new_n303), .B(new_n305), .C1(new_n358), .C2(new_n360), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n351), .A2(KEYINPUT31), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n357), .A2(new_n352), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n362), .A2(new_n360), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g178(.A(KEYINPUT32), .B1(new_n364), .B2(new_n304), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n361), .A2(new_n365), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n350), .B1(new_n342), .B2(new_n345), .ZN(new_n367));
  NOR2_X1   g181(.A1(new_n357), .A2(new_n352), .ZN(new_n368));
  NOR3_X1   g182(.A1(new_n367), .A2(new_n368), .A3(KEYINPUT29), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n343), .A2(new_n328), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n370), .A2(new_n320), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(KEYINPUT72), .A3(new_n345), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT72), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n370), .A2(new_n373), .A3(new_n320), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n372), .A2(KEYINPUT28), .A3(new_n374), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n375), .A2(new_n354), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n350), .A2(KEYINPUT29), .ZN(new_n377));
  OAI21_X1  g191(.A(new_n286), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OAI21_X1  g192(.A(G472), .B1(new_n369), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(KEYINPUT16), .ZN(new_n380));
  NOR2_X1   g194(.A1(KEYINPUT74), .A2(G125), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  NAND2_X1  g196(.A1(KEYINPUT74), .A2(G125), .ZN(new_n383));
  NAND3_X1  g197(.A1(new_n382), .A2(G140), .A3(new_n383), .ZN(new_n384));
  NOR2_X1   g198(.A1(G125), .A2(G140), .ZN(new_n385));
  INV_X1    g199(.A(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n380), .B1(new_n384), .B2(new_n386), .ZN(new_n387));
  XNOR2_X1  g201(.A(KEYINPUT74), .B(G125), .ZN(new_n388));
  NOR3_X1   g202(.A1(new_n388), .A2(KEYINPUT16), .A3(G140), .ZN(new_n389));
  OAI21_X1  g203(.A(new_n210), .B1(new_n387), .B2(new_n389), .ZN(new_n390));
  AND2_X1   g204(.A1(KEYINPUT74), .A2(G125), .ZN(new_n391));
  NOR2_X1   g205(.A1(new_n391), .A2(new_n381), .ZN(new_n392));
  INV_X1    g206(.A(G140), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n392), .A2(new_n380), .A3(new_n393), .ZN(new_n394));
  AOI21_X1  g208(.A(new_n385), .B1(new_n392), .B2(G140), .ZN(new_n395));
  OAI211_X1 g209(.A(G146), .B(new_n394), .C1(new_n395), .C2(new_n380), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n390), .A2(new_n396), .A3(KEYINPUT75), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n232), .A2(G119), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n307), .A2(G128), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  XNOR2_X1  g214(.A(KEYINPUT24), .B(G110), .ZN(new_n401));
  OR2_X1    g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT23), .ZN(new_n403));
  OAI21_X1  g217(.A(new_n403), .B1(new_n307), .B2(G128), .ZN(new_n404));
  OAI211_X1 g218(.A(new_n399), .B(new_n404), .C1(new_n398), .C2(new_n403), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(G110), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT75), .ZN(new_n407));
  OAI211_X1 g221(.A(new_n407), .B(new_n210), .C1(new_n387), .C2(new_n389), .ZN(new_n408));
  NAND4_X1  g222(.A1(new_n397), .A2(new_n402), .A3(new_n406), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n400), .A2(new_n401), .ZN(new_n410));
  OAI21_X1  g224(.A(new_n410), .B1(new_n405), .B2(G110), .ZN(new_n411));
  XNOR2_X1  g225(.A(G125), .B(G140), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n210), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n411), .A2(new_n396), .A3(new_n413), .ZN(new_n414));
  AND3_X1   g228(.A1(new_n409), .A2(KEYINPUT78), .A3(new_n414), .ZN(new_n415));
  AOI21_X1  g229(.A(KEYINPUT78), .B1(new_n409), .B2(new_n414), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n267), .A2(G221), .A3(G234), .ZN(new_n417));
  XNOR2_X1  g231(.A(KEYINPUT76), .B(KEYINPUT77), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n417), .B(new_n418), .ZN(new_n419));
  XOR2_X1   g233(.A(KEYINPUT22), .B(G137), .Z(new_n420));
  XNOR2_X1  g234(.A(new_n419), .B(new_n420), .ZN(new_n421));
  NOR3_X1   g235(.A1(new_n415), .A2(new_n416), .A3(new_n421), .ZN(new_n422));
  AND4_X1   g236(.A1(KEYINPUT78), .A2(new_n421), .A3(new_n409), .A4(new_n414), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n286), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n424), .A2(KEYINPUT25), .ZN(new_n425));
  INV_X1    g239(.A(KEYINPUT25), .ZN(new_n426));
  OAI211_X1 g240(.A(new_n426), .B(new_n286), .C1(new_n422), .C2(new_n423), .ZN(new_n427));
  INV_X1    g241(.A(G217), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n428), .B1(G234), .B2(new_n286), .ZN(new_n429));
  XNOR2_X1  g243(.A(new_n429), .B(KEYINPUT73), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n425), .A2(new_n427), .A3(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT79), .ZN(new_n432));
  OR3_X1    g246(.A1(new_n415), .A2(new_n416), .A3(new_n421), .ZN(new_n433));
  INV_X1    g247(.A(new_n423), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NOR2_X1   g249(.A1(new_n429), .A2(G902), .ZN(new_n436));
  AND3_X1   g250(.A1(new_n435), .A2(KEYINPUT80), .A3(new_n436), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT80), .B1(new_n435), .B2(new_n436), .ZN(new_n438));
  NOR2_X1   g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT79), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n425), .A2(new_n440), .A3(new_n427), .A4(new_n430), .ZN(new_n441));
  NAND3_X1  g255(.A1(new_n432), .A2(new_n439), .A3(new_n441), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n442), .A2(KEYINPUT81), .ZN(new_n443));
  INV_X1    g257(.A(KEYINPUT81), .ZN(new_n444));
  NAND4_X1  g258(.A1(new_n432), .A2(new_n439), .A3(new_n444), .A4(new_n441), .ZN(new_n445));
  AOI22_X1  g259(.A1(new_n366), .A2(new_n379), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  OAI21_X1  g260(.A(G214), .B1(G237), .B2(G902), .ZN(new_n447));
  INV_X1    g261(.A(G952), .ZN(new_n448));
  AOI211_X1 g262(.A(G953), .B(new_n448), .C1(G234), .C2(G237), .ZN(new_n449));
  INV_X1    g263(.A(new_n449), .ZN(new_n450));
  AOI211_X1 g264(.A(new_n286), .B(new_n267), .C1(G234), .C2(G237), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  XOR2_X1   g266(.A(KEYINPUT21), .B(G898), .Z(new_n453));
  OAI21_X1  g267(.A(new_n450), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n242), .A2(G101), .ZN(new_n455));
  AOI22_X1  g269(.A1(new_n455), .A2(new_n241), .B1(new_n313), .B2(new_n319), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(new_n244), .ZN(new_n457));
  NAND3_X1  g271(.A1(new_n317), .A2(KEYINPUT5), .A3(new_n318), .ZN(new_n458));
  INV_X1    g272(.A(G113), .ZN(new_n459));
  INV_X1    g273(.A(KEYINPUT5), .ZN(new_n460));
  AOI21_X1  g274(.A(new_n459), .B1(new_n312), .B2(new_n460), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n458), .A2(new_n461), .ZN(new_n462));
  NAND4_X1  g276(.A1(new_n253), .A2(new_n319), .A3(new_n254), .A4(new_n462), .ZN(new_n463));
  XNOR2_X1  g277(.A(G110), .B(G122), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n457), .A2(new_n463), .A3(new_n464), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT90), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND4_X1  g281(.A1(new_n457), .A2(new_n463), .A3(KEYINPUT90), .A4(new_n464), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  INV_X1    g283(.A(KEYINPUT91), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT6), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n457), .A2(new_n463), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n464), .B(KEYINPUT89), .ZN(new_n473));
  AOI21_X1  g287(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND3_X1   g288(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g289(.A(new_n470), .B1(new_n469), .B2(new_n474), .ZN(new_n476));
  NAND3_X1  g290(.A1(new_n472), .A2(new_n471), .A3(new_n473), .ZN(new_n477));
  INV_X1    g291(.A(new_n477), .ZN(new_n478));
  NOR3_X1   g292(.A1(new_n475), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n250), .A2(new_n392), .ZN(new_n480));
  OAI21_X1  g294(.A(new_n480), .B1(new_n234), .B2(new_n392), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n263), .A2(G224), .ZN(new_n482));
  XOR2_X1   g296(.A(new_n481), .B(new_n482), .Z(new_n483));
  NAND3_X1  g297(.A1(new_n479), .A2(KEYINPUT92), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n469), .A2(new_n474), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(KEYINPUT91), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n469), .A2(new_n470), .A3(new_n474), .ZN(new_n487));
  NAND4_X1  g301(.A1(new_n486), .A2(new_n477), .A3(new_n487), .A4(new_n483), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT92), .ZN(new_n489));
  NAND2_X1  g303(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n484), .A2(new_n490), .ZN(new_n491));
  OAI21_X1  g305(.A(G210), .B1(G237), .B2(G902), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n458), .A2(KEYINPUT93), .ZN(new_n493));
  INV_X1    g307(.A(KEYINPUT93), .ZN(new_n494));
  NAND4_X1  g308(.A1(new_n317), .A2(new_n494), .A3(KEYINPUT5), .A4(new_n318), .ZN(new_n495));
  NAND3_X1  g309(.A1(new_n493), .A2(new_n461), .A3(new_n495), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n231), .A2(new_n496), .A3(new_n319), .ZN(new_n497));
  INV_X1    g311(.A(KEYINPUT94), .ZN(new_n498));
  NAND2_X1  g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  AND2_X1   g313(.A1(new_n462), .A2(new_n319), .ZN(new_n500));
  OR2_X1    g314(.A1(new_n500), .A2(new_n231), .ZN(new_n501));
  NAND4_X1  g315(.A1(new_n231), .A2(new_n496), .A3(KEYINPUT94), .A4(new_n319), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n499), .A2(new_n501), .A3(new_n502), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n464), .B(KEYINPUT8), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n482), .A2(KEYINPUT7), .ZN(new_n506));
  XNOR2_X1  g320(.A(new_n481), .B(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n505), .A2(new_n469), .A3(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT95), .ZN(new_n510));
  AND3_X1   g324(.A1(new_n509), .A2(new_n510), .A3(new_n286), .ZN(new_n511));
  AOI21_X1  g325(.A(new_n510), .B1(new_n509), .B2(new_n286), .ZN(new_n512));
  OR2_X1    g326(.A1(new_n511), .A2(new_n512), .ZN(new_n513));
  AND3_X1   g327(.A1(new_n491), .A2(new_n492), .A3(new_n513), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n492), .B1(new_n491), .B2(new_n513), .ZN(new_n515));
  OAI211_X1 g329(.A(new_n447), .B(new_n454), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G122), .B1(new_n315), .B2(new_n316), .ZN(new_n517));
  OAI21_X1  g331(.A(new_n517), .B1(new_n311), .B2(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(G107), .ZN(new_n519));
  AND2_X1   g333(.A1(new_n232), .A2(G143), .ZN(new_n520));
  OAI21_X1  g334(.A(G134), .B1(new_n520), .B2(KEYINPUT13), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n232), .A2(G143), .ZN(new_n522));
  INV_X1    g336(.A(KEYINPUT99), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n523), .B1(new_n217), .B2(G143), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n212), .A2(KEYINPUT99), .A3(G128), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n522), .A2(new_n524), .A3(new_n525), .ZN(new_n526));
  AND2_X1   g340(.A1(new_n521), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g341(.A1(new_n521), .A2(new_n526), .ZN(new_n528));
  OAI21_X1  g342(.A(new_n519), .B1(new_n527), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT100), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n529), .A2(new_n530), .ZN(new_n531));
  OAI211_X1 g345(.A(KEYINPUT100), .B(new_n519), .C1(new_n527), .C2(new_n528), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n526), .B(G134), .ZN(new_n534));
  OR2_X1    g348(.A1(new_n518), .A2(G107), .ZN(new_n535));
  OAI211_X1 g349(.A(KEYINPUT14), .B(G122), .C1(new_n315), .C2(new_n316), .ZN(new_n536));
  OAI211_X1 g350(.A(G107), .B(new_n536), .C1(new_n518), .C2(KEYINPUT14), .ZN(new_n537));
  NAND3_X1  g351(.A1(new_n534), .A2(new_n535), .A3(new_n537), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n538), .A2(KEYINPUT101), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT101), .ZN(new_n540));
  NAND4_X1  g354(.A1(new_n534), .A2(new_n540), .A3(new_n535), .A4(new_n537), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n539), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  NOR3_X1   g357(.A1(new_n296), .A2(new_n428), .A3(G953), .ZN(new_n544));
  INV_X1    g358(.A(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n543), .A2(new_n545), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n533), .A2(new_n542), .A3(new_n544), .ZN(new_n547));
  AOI21_X1  g361(.A(G902), .B1(new_n546), .B2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(G478), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n548), .B1(KEYINPUT15), .B2(new_n549), .ZN(new_n550));
  INV_X1    g364(.A(new_n547), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n544), .B1(new_n533), .B2(new_n542), .ZN(new_n552));
  OAI21_X1  g366(.A(new_n286), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NOR2_X1   g367(.A1(new_n549), .A2(KEYINPUT15), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n553), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n550), .A2(new_n555), .ZN(new_n556));
  INV_X1    g370(.A(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n267), .A2(G214), .A3(new_n346), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n212), .ZN(new_n559));
  NAND4_X1  g373(.A1(new_n267), .A2(G143), .A3(G214), .A4(new_n346), .ZN(new_n560));
  INV_X1    g374(.A(KEYINPUT18), .ZN(new_n561));
  OAI211_X1 g375(.A(new_n559), .B(new_n560), .C1(new_n561), .C2(new_n195), .ZN(new_n562));
  INV_X1    g376(.A(new_n395), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n413), .B1(new_n563), .B2(new_n210), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n559), .A2(new_n560), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(G131), .ZN(new_n566));
  OAI211_X1 g380(.A(new_n562), .B(new_n564), .C1(new_n566), .C2(new_n561), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT17), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n195), .A3(new_n560), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n565), .A2(KEYINPUT17), .A3(G131), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n570), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g386(.A1(new_n397), .A2(new_n408), .ZN(new_n573));
  OAI21_X1  g387(.A(new_n567), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  XNOR2_X1  g388(.A(G113), .B(G122), .ZN(new_n575));
  XNOR2_X1  g389(.A(KEYINPUT96), .B(G104), .ZN(new_n576));
  XNOR2_X1  g390(.A(new_n575), .B(new_n576), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n574), .A2(new_n577), .ZN(new_n578));
  INV_X1    g392(.A(new_n577), .ZN(new_n579));
  OAI211_X1 g393(.A(new_n579), .B(new_n567), .C1(new_n572), .C2(new_n573), .ZN(new_n580));
  AOI21_X1  g394(.A(G902), .B1(new_n578), .B2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(KEYINPUT98), .B(G475), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n566), .A2(new_n569), .ZN(new_n584));
  MUX2_X1   g398(.A(new_n412), .B(new_n395), .S(KEYINPUT19), .Z(new_n585));
  OAI21_X1  g399(.A(new_n396), .B1(new_n585), .B2(G146), .ZN(new_n586));
  OAI21_X1  g400(.A(new_n567), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n577), .ZN(new_n588));
  AOI21_X1  g402(.A(G475), .B1(new_n580), .B2(new_n588), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT20), .ZN(new_n590));
  NAND3_X1  g404(.A1(new_n589), .A2(new_n590), .A3(new_n286), .ZN(new_n591));
  AOI21_X1  g405(.A(new_n590), .B1(new_n589), .B2(new_n286), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n591), .B1(new_n592), .B2(KEYINPUT97), .ZN(new_n593));
  INV_X1    g407(.A(KEYINPUT97), .ZN(new_n594));
  NAND4_X1  g408(.A1(new_n589), .A2(new_n594), .A3(new_n590), .A4(new_n286), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n583), .B1(new_n593), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n557), .A2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n516), .A2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n302), .A2(new_n446), .A3(new_n598), .ZN(new_n599));
  XNOR2_X1  g413(.A(new_n599), .B(G101), .ZN(G3));
  NAND2_X1  g414(.A1(new_n443), .A2(new_n445), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n364), .A2(new_n286), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(G472), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n364), .A2(new_n304), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  INV_X1    g419(.A(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n302), .A2(new_n601), .A3(new_n606), .ZN(new_n607));
  INV_X1    g421(.A(new_n607), .ZN(new_n608));
  INV_X1    g422(.A(new_n596), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT102), .B1(new_n548), .B2(G478), .ZN(new_n610));
  INV_X1    g424(.A(KEYINPUT102), .ZN(new_n611));
  NAND3_X1  g425(.A1(new_n553), .A2(new_n611), .A3(new_n549), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n610), .A2(new_n612), .ZN(new_n613));
  INV_X1    g427(.A(KEYINPUT33), .ZN(new_n614));
  OAI21_X1  g428(.A(new_n614), .B1(new_n551), .B2(new_n552), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n546), .A2(KEYINPUT33), .A3(new_n547), .ZN(new_n616));
  NAND4_X1  g430(.A1(new_n615), .A2(new_n616), .A3(G478), .A4(new_n286), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n613), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n609), .A2(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n516), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n608), .A2(new_n620), .ZN(new_n621));
  XNOR2_X1  g435(.A(new_n621), .B(G104), .ZN(new_n622));
  XOR2_X1   g436(.A(KEYINPUT103), .B(KEYINPUT34), .Z(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n592), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n591), .ZN(new_n626));
  XNOR2_X1  g440(.A(new_n626), .B(KEYINPUT104), .ZN(new_n627));
  INV_X1    g441(.A(new_n583), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n627), .A2(new_n556), .A3(new_n628), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n516), .A2(new_n629), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n608), .A2(new_n630), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n631), .B(KEYINPUT105), .ZN(new_n632));
  XNOR2_X1  g446(.A(KEYINPUT35), .B(G107), .ZN(new_n633));
  XNOR2_X1  g447(.A(new_n632), .B(new_n633), .ZN(G9));
  NOR2_X1   g448(.A1(new_n421), .A2(KEYINPUT36), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n409), .A2(new_n414), .ZN(new_n636));
  XNOR2_X1  g450(.A(new_n635), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n637), .A2(new_n436), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n432), .A2(new_n441), .A3(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n302), .A2(new_n598), .A3(new_n606), .A4(new_n639), .ZN(new_n640));
  XOR2_X1   g454(.A(KEYINPUT37), .B(G110), .Z(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  XNOR2_X1  g456(.A(KEYINPUT106), .B(G900), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n449), .B1(new_n451), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND4_X1  g459(.A1(new_n627), .A2(new_n556), .A3(new_n628), .A4(new_n645), .ZN(new_n646));
  AOI21_X1  g460(.A(new_n646), .B1(new_n299), .B2(new_n301), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n604), .A2(new_n303), .ZN(new_n648));
  NAND3_X1  g462(.A1(new_n364), .A2(KEYINPUT32), .A3(new_n304), .ZN(new_n649));
  NAND3_X1  g463(.A1(new_n648), .A2(new_n379), .A3(new_n649), .ZN(new_n650));
  INV_X1    g464(.A(new_n447), .ZN(new_n651));
  AOI21_X1  g465(.A(KEYINPUT92), .B1(new_n479), .B2(new_n483), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n488), .A2(new_n489), .ZN(new_n653));
  OAI21_X1  g467(.A(new_n513), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n492), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n654), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n491), .A2(new_n492), .A3(new_n513), .ZN(new_n657));
  AOI21_X1  g471(.A(new_n651), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND3_X1   g472(.A1(new_n650), .A2(new_n658), .A3(new_n639), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n647), .A2(new_n659), .ZN(new_n660));
  XNOR2_X1  g474(.A(new_n660), .B(G128), .ZN(G30));
  XOR2_X1   g475(.A(new_n644), .B(KEYINPUT39), .Z(new_n662));
  NAND2_X1  g476(.A1(new_n302), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(KEYINPUT40), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n372), .A2(new_n352), .A3(new_n374), .ZN(new_n665));
  AND2_X1   g479(.A1(new_n351), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g480(.A(G472), .B1(new_n666), .B2(G902), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n639), .B1(new_n366), .B2(new_n667), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n664), .A2(new_n447), .A3(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n557), .A2(new_n596), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n656), .A2(new_n657), .ZN(new_n671));
  XNOR2_X1  g485(.A(KEYINPUT107), .B(KEYINPUT38), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n671), .B(new_n672), .ZN(new_n673));
  OAI211_X1 g487(.A(new_n670), .B(new_n673), .C1(new_n663), .C2(KEYINPUT40), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n669), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(new_n212), .ZN(G45));
  NOR2_X1   g490(.A1(new_n619), .A2(new_n644), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n302), .A2(new_n659), .A3(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G146), .ZN(G48));
  AND3_X1   g493(.A1(new_n284), .A2(new_n285), .A3(new_n286), .ZN(new_n680));
  AOI21_X1  g494(.A(new_n285), .B1(new_n284), .B2(new_n286), .ZN(new_n681));
  INV_X1    g495(.A(new_n297), .ZN(new_n682));
  NOR3_X1   g496(.A1(new_n680), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND3_X1  g497(.A1(new_n620), .A2(new_n446), .A3(new_n683), .ZN(new_n684));
  XNOR2_X1  g498(.A(KEYINPUT41), .B(G113), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n684), .B(new_n685), .ZN(G15));
  NAND3_X1  g500(.A1(new_n630), .A2(new_n446), .A3(new_n683), .ZN(new_n687));
  XNOR2_X1  g501(.A(new_n687), .B(G116), .ZN(G18));
  OAI21_X1  g502(.A(new_n447), .B1(new_n514), .B2(new_n515), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n284), .A2(new_n286), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n690), .A2(G469), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n691), .A2(new_n297), .A3(new_n287), .ZN(new_n692));
  OAI21_X1  g506(.A(KEYINPUT108), .B1(new_n689), .B2(new_n692), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT108), .ZN(new_n694));
  NAND3_X1  g508(.A1(new_n683), .A2(new_n658), .A3(new_n694), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n693), .A2(new_n695), .ZN(new_n696));
  INV_X1    g510(.A(new_n597), .ZN(new_n697));
  AND3_X1   g511(.A1(new_n650), .A2(new_n454), .A3(new_n639), .ZN(new_n698));
  NAND3_X1  g512(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  XNOR2_X1  g513(.A(new_n699), .B(G119), .ZN(G21));
  INV_X1    g514(.A(KEYINPUT109), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n376), .A2(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n375), .A2(KEYINPUT109), .A3(new_n354), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n702), .A2(new_n352), .A3(new_n703), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n704), .A2(KEYINPUT110), .A3(new_n362), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n705), .A2(new_n360), .ZN(new_n706));
  AOI21_X1  g520(.A(KEYINPUT110), .B1(new_n704), .B2(new_n362), .ZN(new_n707));
  OAI21_X1  g521(.A(new_n304), .B1(new_n706), .B2(new_n707), .ZN(new_n708));
  INV_X1    g522(.A(new_n442), .ZN(new_n709));
  AND3_X1   g523(.A1(new_n708), .A2(new_n709), .A3(new_n603), .ZN(new_n710));
  INV_X1    g524(.A(new_n516), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n710), .A2(new_n711), .A3(new_n670), .A4(new_n683), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  AND4_X1   g527(.A1(new_n603), .A2(new_n677), .A3(new_n639), .A4(new_n708), .ZN(new_n714));
  NAND2_X1  g528(.A1(new_n696), .A2(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(G125), .ZN(G27));
  NAND2_X1  g530(.A1(G469), .A2(G902), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n289), .A2(KEYINPUT111), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT111), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n288), .A2(new_n719), .A3(new_n273), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n718), .A2(G469), .A3(new_n290), .A4(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n287), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(KEYINPUT112), .ZN(new_n723));
  AND3_X1   g537(.A1(new_n722), .A2(new_n723), .A3(new_n297), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n723), .B1(new_n722), .B2(new_n297), .ZN(new_n725));
  NOR2_X1   g539(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  INV_X1    g540(.A(new_n677), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n656), .A2(new_n447), .A3(new_n657), .ZN(new_n728));
  NOR2_X1   g542(.A1(new_n727), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g543(.A(KEYINPUT113), .B1(new_n650), .B2(new_n709), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n650), .A2(KEYINPUT113), .A3(new_n709), .ZN(new_n731));
  OAI211_X1 g545(.A(new_n726), .B(new_n729), .C1(new_n730), .C2(new_n731), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n722), .A2(new_n297), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n733), .A2(KEYINPUT112), .ZN(new_n734));
  INV_X1    g548(.A(new_n728), .ZN(new_n735));
  NAND3_X1  g549(.A1(new_n722), .A2(new_n723), .A3(new_n297), .ZN(new_n736));
  AND4_X1   g550(.A1(new_n446), .A2(new_n734), .A3(new_n735), .A4(new_n736), .ZN(new_n737));
  NOR2_X1   g551(.A1(new_n727), .A2(KEYINPUT42), .ZN(new_n738));
  AOI22_X1  g552(.A1(new_n732), .A2(KEYINPUT42), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  XNOR2_X1  g553(.A(new_n739), .B(G131), .ZN(G33));
  INV_X1    g554(.A(new_n646), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n737), .A2(new_n741), .ZN(new_n742));
  XOR2_X1   g556(.A(KEYINPUT114), .B(G134), .Z(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G36));
  OR2_X1    g558(.A1(new_n609), .A2(KEYINPUT117), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n609), .A2(KEYINPUT117), .ZN(new_n746));
  NAND3_X1  g560(.A1(new_n745), .A2(new_n618), .A3(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n747), .A2(KEYINPUT43), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  NAND3_X1  g563(.A1(new_n618), .A2(new_n749), .A3(new_n596), .ZN(new_n750));
  AND2_X1   g564(.A1(new_n605), .A2(new_n639), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n748), .A2(new_n750), .A3(new_n751), .ZN(new_n752));
  INV_X1    g566(.A(KEYINPUT44), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n752), .A2(new_n753), .ZN(new_n754));
  NAND4_X1  g568(.A1(new_n748), .A2(KEYINPUT44), .A3(new_n750), .A4(new_n751), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n754), .A2(new_n735), .A3(new_n755), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT118), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND4_X1  g572(.A1(new_n718), .A2(KEYINPUT45), .A3(new_n290), .A4(new_n720), .ZN(new_n759));
  INV_X1    g573(.A(KEYINPUT45), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n291), .A2(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n759), .A2(G469), .A3(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n717), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT46), .ZN(new_n764));
  NAND2_X1  g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n765), .A2(KEYINPUT115), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n762), .A2(KEYINPUT46), .A3(new_n717), .ZN(new_n767));
  AND2_X1   g581(.A1(new_n767), .A2(new_n287), .ZN(new_n768));
  INV_X1    g582(.A(KEYINPUT115), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n763), .A2(new_n769), .A3(new_n764), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n766), .A2(new_n768), .A3(new_n770), .ZN(new_n771));
  NAND3_X1  g585(.A1(new_n771), .A2(new_n297), .A3(new_n662), .ZN(new_n772));
  XNOR2_X1  g586(.A(new_n772), .B(KEYINPUT116), .ZN(new_n773));
  NAND4_X1  g587(.A1(new_n754), .A2(KEYINPUT118), .A3(new_n735), .A4(new_n755), .ZN(new_n774));
  NAND3_X1  g588(.A1(new_n758), .A2(new_n773), .A3(new_n774), .ZN(new_n775));
  XNOR2_X1  g589(.A(new_n775), .B(G137), .ZN(G39));
  NAND2_X1  g590(.A1(KEYINPUT119), .A2(KEYINPUT47), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n771), .B2(new_n297), .ZN(new_n778));
  AOI21_X1  g592(.A(new_n769), .B1(new_n763), .B2(new_n764), .ZN(new_n779));
  AOI211_X1 g593(.A(KEYINPUT115), .B(KEYINPUT46), .C1(new_n762), .C2(new_n717), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n767), .A2(new_n287), .ZN(new_n781));
  NOR3_X1   g595(.A1(new_n779), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  OAI22_X1  g596(.A1(new_n782), .A2(new_n682), .B1(KEYINPUT119), .B2(KEYINPUT47), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n778), .B1(new_n783), .B2(new_n777), .ZN(new_n784));
  NOR3_X1   g598(.A1(new_n727), .A2(new_n601), .A3(new_n728), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n784), .A2(new_n366), .A3(new_n379), .A4(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  NAND3_X1  g601(.A1(new_n748), .A2(new_n449), .A3(new_n750), .ZN(new_n788));
  NOR3_X1   g602(.A1(new_n788), .A2(new_n692), .A3(new_n728), .ZN(new_n789));
  OR2_X1    g603(.A1(new_n731), .A2(new_n730), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT123), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  OR2_X1    g607(.A1(new_n793), .A2(KEYINPUT48), .ZN(new_n794));
  NOR2_X1   g608(.A1(new_n448), .A2(G953), .ZN(new_n795));
  INV_X1    g609(.A(new_n710), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n788), .A2(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n797), .A2(new_n696), .ZN(new_n798));
  NAND3_X1  g612(.A1(new_n789), .A2(KEYINPUT123), .A3(new_n790), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n793), .A2(KEYINPUT48), .A3(new_n799), .ZN(new_n800));
  NAND4_X1  g614(.A1(new_n794), .A2(new_n795), .A3(new_n798), .A4(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n691), .A2(new_n287), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n297), .ZN(new_n803));
  OAI211_X1 g617(.A(new_n735), .B(new_n797), .C1(new_n784), .C2(new_n803), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n673), .A2(new_n447), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n797), .A2(new_n683), .A3(new_n805), .ZN(new_n806));
  XOR2_X1   g620(.A(KEYINPUT122), .B(KEYINPUT50), .Z(new_n807));
  NAND2_X1  g621(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g622(.A1(new_n366), .A2(new_n667), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n450), .ZN(new_n810));
  NAND4_X1  g624(.A1(new_n810), .A2(new_n601), .A3(new_n683), .A4(new_n735), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n811), .A2(new_n609), .A3(new_n618), .ZN(new_n812));
  AND3_X1   g626(.A1(new_n804), .A2(new_n808), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n814));
  AND2_X1   g628(.A1(new_n708), .A2(new_n603), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n789), .A2(new_n639), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(KEYINPUT122), .A2(KEYINPUT50), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n797), .A2(new_n683), .A3(new_n817), .A4(new_n805), .ZN(new_n818));
  NAND4_X1  g632(.A1(new_n813), .A2(new_n814), .A3(new_n816), .A4(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n804), .A2(new_n818), .A3(new_n808), .A4(new_n812), .ZN(new_n820));
  INV_X1    g634(.A(new_n816), .ZN(new_n821));
  OAI21_X1  g635(.A(KEYINPUT51), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n801), .B1(new_n819), .B2(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n671), .A2(new_n447), .A3(new_n670), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n824), .A2(new_n733), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n825), .A2(new_n645), .A3(new_n668), .ZN(new_n826));
  NAND4_X1  g640(.A1(new_n715), .A2(new_n660), .A3(new_n678), .A4(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT121), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI22_X1  g645(.A1(new_n696), .A2(new_n714), .B1(new_n647), .B2(new_n659), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .A3(new_n678), .A4(new_n826), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n827), .A2(KEYINPUT121), .A3(new_n828), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n831), .A2(new_n833), .A3(new_n834), .ZN(new_n835));
  AND2_X1   g649(.A1(new_n650), .A2(new_n639), .ZN(new_n836));
  NAND3_X1  g650(.A1(new_n627), .A2(new_n628), .A3(new_n645), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n728), .A2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n302), .A2(new_n557), .A3(new_n836), .A4(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT120), .ZN(new_n840));
  AOI22_X1  g654(.A1(new_n741), .A2(new_n737), .B1(new_n839), .B2(new_n840), .ZN(new_n841));
  OR2_X1    g655(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n739), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n596), .B1(new_n613), .B2(new_n617), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n596), .A2(new_n556), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  NOR2_X1   g660(.A1(new_n516), .A2(new_n846), .ZN(new_n847));
  NAND4_X1  g661(.A1(new_n302), .A2(new_n601), .A3(new_n606), .A4(new_n847), .ZN(new_n848));
  AND3_X1   g662(.A1(new_n640), .A2(new_n848), .A3(new_n599), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n714), .A2(new_n726), .A3(new_n735), .ZN(new_n850));
  AND3_X1   g664(.A1(new_n712), .A2(new_n684), .A3(new_n687), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n699), .A3(new_n850), .A4(new_n851), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n843), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n835), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n739), .A2(new_n841), .A3(new_n842), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n699), .A2(new_n640), .A3(new_n848), .A4(new_n599), .ZN(new_n856));
  INV_X1    g670(.A(new_n850), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n712), .A2(new_n684), .A3(new_n687), .ZN(new_n858));
  NOR3_X1   g672(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n829), .A2(new_n833), .ZN(new_n860));
  AND4_X1   g674(.A1(KEYINPUT53), .A2(new_n855), .A3(new_n859), .A4(new_n860), .ZN(new_n861));
  OAI21_X1  g675(.A(KEYINPUT54), .B1(new_n854), .B2(new_n861), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n835), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n863));
  NAND3_X1  g677(.A1(new_n855), .A2(new_n859), .A3(new_n860), .ZN(new_n864));
  INV_X1    g678(.A(KEYINPUT53), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  INV_X1    g680(.A(KEYINPUT54), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n868));
  NAND3_X1  g682(.A1(new_n823), .A2(new_n862), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n811), .A2(new_n619), .ZN(new_n870));
  OAI22_X1  g684(.A1(new_n869), .A2(new_n870), .B1(G952), .B2(G953), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n673), .A2(new_n651), .A3(new_n747), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n802), .B(KEYINPUT49), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n873), .A2(new_n809), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n872), .A2(new_n874), .A3(new_n709), .A4(new_n297), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n871), .A2(new_n875), .ZN(G75));
  XOR2_X1   g690(.A(new_n479), .B(new_n483), .Z(new_n877));
  XOR2_X1   g691(.A(new_n877), .B(KEYINPUT55), .Z(new_n878));
  INV_X1    g692(.A(G210), .ZN(new_n879));
  AOI211_X1 g693(.A(new_n879), .B(new_n286), .C1(new_n863), .C2(new_n866), .ZN(new_n880));
  OAI21_X1  g694(.A(new_n878), .B1(new_n880), .B2(KEYINPUT56), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n267), .A2(G952), .ZN(new_n882));
  INV_X1    g696(.A(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT56), .ZN(new_n884));
  INV_X1    g698(.A(new_n878), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n863), .A2(new_n866), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n886), .A2(G902), .ZN(new_n887));
  OAI211_X1 g701(.A(new_n884), .B(new_n885), .C1(new_n887), .C2(new_n879), .ZN(new_n888));
  AND3_X1   g702(.A1(new_n881), .A2(new_n883), .A3(new_n888), .ZN(G51));
  XOR2_X1   g703(.A(new_n717), .B(KEYINPUT57), .Z(new_n890));
  AND3_X1   g704(.A1(new_n863), .A2(new_n866), .A3(new_n867), .ZN(new_n891));
  AOI21_X1  g705(.A(new_n867), .B1(new_n863), .B2(new_n866), .ZN(new_n892));
  OAI21_X1  g706(.A(new_n890), .B1(new_n891), .B2(new_n892), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n893), .A2(new_n284), .ZN(new_n894));
  OR2_X1    g708(.A1(new_n887), .A2(new_n762), .ZN(new_n895));
  AOI21_X1  g709(.A(new_n882), .B1(new_n894), .B2(new_n895), .ZN(G54));
  NAND2_X1  g710(.A1(KEYINPUT58), .A2(G475), .ZN(new_n897));
  INV_X1    g711(.A(new_n897), .ZN(new_n898));
  NAND3_X1  g712(.A1(new_n886), .A2(G902), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n580), .A2(new_n588), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n883), .B1(new_n899), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g716(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n903), .A2(KEYINPUT124), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT124), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n899), .A2(new_n905), .A3(new_n901), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n902), .B1(new_n904), .B2(new_n906), .ZN(G60));
  NAND2_X1  g721(.A1(G478), .A2(G902), .ZN(new_n908));
  XOR2_X1   g722(.A(new_n908), .B(KEYINPUT59), .Z(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n862), .B2(new_n868), .ZN(new_n910));
  AND2_X1   g724(.A1(new_n615), .A2(new_n616), .ZN(new_n911));
  OAI21_X1  g725(.A(new_n883), .B1(new_n910), .B2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n909), .ZN(new_n913));
  OAI211_X1 g727(.A(new_n911), .B(new_n913), .C1(new_n891), .C2(new_n892), .ZN(new_n914));
  INV_X1    g728(.A(new_n914), .ZN(new_n915));
  NOR2_X1   g729(.A1(new_n912), .A2(new_n915), .ZN(G63));
  XNOR2_X1  g730(.A(KEYINPUT126), .B(KEYINPUT61), .ZN(new_n917));
  INV_X1    g731(.A(new_n917), .ZN(new_n918));
  XNOR2_X1  g732(.A(KEYINPUT125), .B(KEYINPUT60), .ZN(new_n919));
  NOR2_X1   g733(.A1(new_n428), .A2(new_n286), .ZN(new_n920));
  XNOR2_X1  g734(.A(new_n919), .B(new_n920), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n886), .A2(new_n637), .A3(new_n921), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(new_n883), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n435), .B1(new_n886), .B2(new_n921), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n918), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  INV_X1    g739(.A(new_n924), .ZN(new_n926));
  NAND4_X1  g740(.A1(new_n926), .A2(new_n883), .A3(new_n922), .A4(new_n917), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n925), .A2(new_n927), .ZN(G66));
  NOR2_X1   g742(.A1(new_n856), .A2(new_n858), .ZN(new_n929));
  INV_X1    g743(.A(new_n267), .ZN(new_n930));
  AND2_X1   g744(.A1(new_n453), .A2(G224), .ZN(new_n931));
  OAI22_X1  g745(.A1(new_n929), .A2(new_n930), .B1(new_n263), .B2(new_n931), .ZN(new_n932));
  INV_X1    g746(.A(new_n479), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n933), .B1(G898), .B2(new_n267), .ZN(new_n934));
  XNOR2_X1  g748(.A(new_n932), .B(new_n934), .ZN(G69));
  OAI21_X1  g749(.A(new_n331), .B1(new_n341), .B2(new_n330), .ZN(new_n936));
  XNOR2_X1  g750(.A(new_n936), .B(new_n585), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n930), .A2(G900), .ZN(new_n938));
  NAND2_X1  g752(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g753(.A(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n832), .A2(new_n678), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n775), .A2(new_n742), .A3(new_n786), .A4(new_n942), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n773), .A2(new_n790), .ZN(new_n944));
  OAI21_X1  g758(.A(new_n739), .B1(new_n944), .B2(new_n824), .ZN(new_n945));
  OR2_X1    g759(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n940), .B1(new_n946), .B2(new_n930), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n267), .B1(G227), .B2(G900), .ZN(new_n948));
  AND2_X1   g762(.A1(new_n775), .A2(new_n786), .ZN(new_n949));
  INV_X1    g763(.A(KEYINPUT62), .ZN(new_n950));
  OAI21_X1  g764(.A(new_n950), .B1(new_n675), .B2(new_n941), .ZN(new_n951));
  OAI211_X1 g765(.A(new_n942), .B(KEYINPUT62), .C1(new_n674), .C2(new_n669), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n446), .ZN(new_n954));
  OR4_X1    g768(.A1(new_n954), .A2(new_n663), .A3(new_n728), .A4(new_n846), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n949), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  AND2_X1   g770(.A1(new_n956), .A2(new_n267), .ZN(new_n957));
  OAI211_X1 g771(.A(new_n947), .B(new_n948), .C1(new_n957), .C2(new_n937), .ZN(new_n958));
  INV_X1    g772(.A(new_n948), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n937), .B1(new_n956), .B2(new_n267), .ZN(new_n960));
  NOR2_X1   g774(.A1(new_n943), .A2(new_n945), .ZN(new_n961));
  AOI21_X1  g775(.A(new_n939), .B1(new_n961), .B2(new_n267), .ZN(new_n962));
  OAI21_X1  g776(.A(new_n959), .B1(new_n960), .B2(new_n962), .ZN(new_n963));
  AND2_X1   g777(.A1(new_n958), .A2(new_n963), .ZN(G72));
  NAND2_X1  g778(.A1(new_n342), .A2(new_n345), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n965), .B(KEYINPUT127), .ZN(new_n966));
  NOR2_X1   g780(.A1(new_n966), .A2(new_n352), .ZN(new_n967));
  NAND4_X1  g781(.A1(new_n949), .A2(new_n953), .A3(new_n955), .A4(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n966), .A2(new_n352), .ZN(new_n969));
  OAI21_X1  g783(.A(new_n968), .B1(new_n946), .B2(new_n969), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n882), .B1(new_n970), .B2(new_n929), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  INV_X1    g787(.A(new_n973), .ZN(new_n974));
  INV_X1    g788(.A(new_n969), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n974), .B1(new_n975), .B2(new_n967), .ZN(new_n976));
  INV_X1    g790(.A(new_n351), .ZN(new_n977));
  OAI221_X1 g791(.A(new_n973), .B1(new_n977), .B2(new_n367), .C1(new_n854), .C2(new_n861), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n971), .A2(new_n976), .A3(new_n978), .ZN(G57));
endmodule


