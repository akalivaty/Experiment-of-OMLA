//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1 1 1 1 0 1 1 0 0 1 0 0 1 0 0 0 1 1 1 0 0 1 0 0 1 0 0 1 1 1 0 0 0 0 0 1 0 1 0 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:28:26 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n455,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n513, new_n514, new_n515, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n538, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n546, new_n548, new_n549, new_n551, new_n552,
    new_n553, new_n554, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n606, new_n607, new_n610, new_n612,
    new_n613, new_n614, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n823, new_n824,
    new_n825, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1161, new_n1162;
  BUF_X1    g000(.A(G452), .Z(G350));
  XOR2_X1   g001(.A(KEYINPUT64), .B(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  INV_X1    g015(.A(G57), .ZN(G237));
  INV_X1    g016(.A(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  INV_X1    g027(.A(new_n452), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n453), .A2(new_n455), .ZN(G325));
  INV_X1    g031(.A(G325), .ZN(G261));
  AOI22_X1  g032(.A1(new_n453), .A2(G2106), .B1(G567), .B2(new_n455), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n460), .A2(G125), .ZN(new_n461));
  NAND2_X1  g036(.A1(G113), .A2(G2104), .ZN(new_n462));
  AOI21_X1  g037(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n460), .A2(G137), .ZN(new_n464));
  NAND2_X1  g039(.A1(G101), .A2(G2104), .ZN(new_n465));
  AOI21_X1  g040(.A(G2105), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NOR2_X1   g041(.A1(new_n463), .A2(new_n466), .ZN(G160));
  INV_X1    g042(.A(KEYINPUT66), .ZN(new_n468));
  INV_X1    g043(.A(G2104), .ZN(new_n469));
  NAND2_X1  g044(.A1(new_n469), .A2(KEYINPUT3), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT3), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n471), .A2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n470), .A2(new_n472), .ZN(new_n473));
  OAI21_X1  g048(.A(new_n468), .B1(new_n473), .B2(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n460), .A2(KEYINPUT66), .A3(new_n459), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n474), .A2(new_n475), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n459), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n460), .A2(G2105), .ZN(new_n481));
  INV_X1    g056(.A(G124), .ZN(new_n482));
  OAI21_X1  g057(.A(KEYINPUT67), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  OR3_X1    g058(.A1(new_n481), .A2(KEYINPUT67), .A3(new_n482), .ZN(new_n484));
  AND4_X1   g059(.A1(new_n478), .A2(new_n480), .A3(new_n483), .A4(new_n484), .ZN(G162));
  NAND3_X1  g060(.A1(new_n470), .A2(new_n472), .A3(G126), .ZN(new_n486));
  NAND2_X1  g061(.A1(G114), .A2(G2104), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G2105), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n469), .A2(G2105), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n490), .A2(G102), .ZN(new_n491));
  NAND4_X1  g066(.A1(new_n470), .A2(new_n472), .A3(G138), .A4(new_n459), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NAND4_X1  g069(.A1(new_n460), .A2(KEYINPUT4), .A3(G138), .A4(new_n459), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n489), .A2(new_n491), .A3(new_n494), .A4(new_n495), .ZN(new_n496));
  INV_X1    g071(.A(new_n496), .ZN(G164));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  INV_X1    g073(.A(G651), .ZN(new_n499));
  OAI21_X1  g074(.A(new_n498), .B1(new_n499), .B2(KEYINPUT68), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT68), .ZN(new_n501));
  NAND3_X1  g076(.A1(new_n501), .A2(KEYINPUT6), .A3(G651), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n503), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  XNOR2_X1  g081(.A(KEYINPUT5), .B(G543), .ZN(new_n507));
  NAND3_X1  g082(.A1(new_n507), .A2(G62), .A3(G651), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n503), .A2(new_n507), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  OAI21_X1  g085(.A(new_n508), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n506), .A2(new_n511), .ZN(G166));
  NAND3_X1  g087(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n513));
  XNOR2_X1  g088(.A(new_n513), .B(KEYINPUT7), .ZN(new_n514));
  INV_X1    g089(.A(G89), .ZN(new_n515));
  INV_X1    g090(.A(KEYINPUT69), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n503), .A2(new_n516), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n500), .A2(KEYINPUT69), .A3(new_n502), .ZN(new_n518));
  NAND3_X1  g093(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G51), .ZN(new_n520));
  INV_X1    g095(.A(G63), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT5), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G543), .ZN(new_n524));
  NAND3_X1  g099(.A1(new_n522), .A2(new_n524), .A3(G651), .ZN(new_n525));
  OAI22_X1  g100(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n525), .ZN(new_n526));
  AND2_X1   g101(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n526), .A2(KEYINPUT70), .ZN(new_n528));
  OAI221_X1 g103(.A(new_n514), .B1(new_n515), .B2(new_n509), .C1(new_n527), .C2(new_n528), .ZN(G286));
  INV_X1    g104(.A(G286), .ZN(G168));
  AND3_X1   g105(.A1(new_n517), .A2(G543), .A3(new_n518), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G52), .ZN(new_n532));
  AOI22_X1  g107(.A1(new_n507), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n533));
  OR2_X1    g108(.A1(new_n533), .A2(new_n499), .ZN(new_n534));
  INV_X1    g109(.A(new_n509), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n535), .A2(G90), .ZN(new_n536));
  AND3_X1   g111(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(G171));
  INV_X1    g112(.A(G43), .ZN(new_n538));
  INV_X1    g113(.A(G81), .ZN(new_n539));
  OAI22_X1  g114(.A1(new_n519), .A2(new_n538), .B1(new_n539), .B2(new_n509), .ZN(new_n540));
  XNOR2_X1  g115(.A(new_n540), .B(KEYINPUT71), .ZN(new_n541));
  AOI22_X1  g116(.A1(new_n507), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(new_n499), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n541), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n544), .A2(G860), .ZN(G153));
  AND3_X1   g120(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G36), .ZN(G176));
  NAND2_X1  g122(.A1(G1), .A2(G3), .ZN(new_n548));
  XNOR2_X1  g123(.A(new_n548), .B(KEYINPUT8), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n546), .A2(new_n549), .ZN(G188));
  NAND3_X1  g125(.A1(new_n531), .A2(KEYINPUT9), .A3(G53), .ZN(new_n551));
  INV_X1    g126(.A(KEYINPUT9), .ZN(new_n552));
  INV_X1    g127(.A(G53), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n552), .B1(new_n519), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(G78), .A2(G543), .ZN(new_n555));
  XOR2_X1   g130(.A(KEYINPUT72), .B(G65), .Z(new_n556));
  NAND2_X1  g131(.A1(new_n522), .A2(new_n524), .ZN(new_n557));
  OAI21_X1  g132(.A(new_n555), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n535), .A2(G91), .B1(new_n558), .B2(G651), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n551), .A2(new_n554), .A3(new_n559), .ZN(new_n560));
  OR2_X1    g135(.A1(new_n560), .A2(KEYINPUT73), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n560), .A2(KEYINPUT73), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n561), .A2(new_n562), .ZN(G299));
  NAND3_X1  g138(.A1(new_n532), .A2(new_n534), .A3(new_n536), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT74), .ZN(G301));
  OAI221_X1 g140(.A(new_n508), .B1(new_n509), .B2(new_n510), .C1(new_n504), .C2(new_n505), .ZN(G303));
  NAND4_X1  g141(.A1(new_n517), .A2(G49), .A3(G543), .A4(new_n518), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  OAI211_X1 g143(.A(new_n568), .B(G651), .C1(new_n507), .C2(G74), .ZN(new_n569));
  NAND2_X1  g144(.A1(G74), .A2(G651), .ZN(new_n570));
  NAND3_X1  g145(.A1(new_n525), .A2(KEYINPUT75), .A3(new_n570), .ZN(new_n571));
  NAND2_X1  g146(.A1(new_n569), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n503), .A2(G87), .A3(new_n507), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n567), .A2(new_n572), .A3(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(KEYINPUT76), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g151(.A1(new_n567), .A2(new_n572), .A3(KEYINPUT76), .A4(new_n573), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n576), .A2(new_n577), .ZN(G288));
  NAND3_X1  g153(.A1(new_n522), .A2(new_n524), .A3(G61), .ZN(new_n579));
  NAND2_X1  g154(.A1(G73), .A2(G543), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n499), .B1(new_n579), .B2(new_n580), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(new_n582));
  NAND3_X1  g157(.A1(new_n522), .A2(new_n524), .A3(G86), .ZN(new_n583));
  NAND2_X1  g158(.A1(G48), .A2(G543), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n583), .A2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(new_n503), .ZN(new_n586));
  NAND2_X1  g161(.A1(new_n582), .A2(new_n586), .ZN(G305));
  AND2_X1   g162(.A1(new_n531), .A2(G47), .ZN(new_n588));
  AOI22_X1  g163(.A1(new_n507), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n589));
  INV_X1    g164(.A(G85), .ZN(new_n590));
  OAI22_X1  g165(.A1(new_n589), .A2(new_n499), .B1(new_n509), .B2(new_n590), .ZN(new_n591));
  NOR2_X1   g166(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(new_n535), .A2(G92), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  INV_X1    g170(.A(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n507), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OAI22_X1  g172(.A1(new_n519), .A2(new_n596), .B1(new_n499), .B2(new_n597), .ZN(new_n598));
  NOR2_X1   g173(.A1(new_n595), .A2(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  INV_X1    g175(.A(G868), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(new_n602));
  XNOR2_X1  g177(.A(G171), .B(KEYINPUT74), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G284));
  OAI21_X1  g179(.A(new_n602), .B1(new_n603), .B2(new_n601), .ZN(G321));
  NAND2_X1  g180(.A1(G286), .A2(G868), .ZN(new_n606));
  XOR2_X1   g181(.A(G299), .B(KEYINPUT77), .Z(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(G868), .ZN(G297));
  XNOR2_X1  g183(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g184(.A(G559), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n599), .B1(new_n610), .B2(G860), .ZN(G148));
  NAND2_X1  g186(.A1(new_n599), .A2(new_n610), .ZN(new_n612));
  XOR2_X1   g187(.A(new_n612), .B(KEYINPUT79), .Z(new_n613));
  NAND2_X1  g188(.A1(new_n613), .A2(G868), .ZN(new_n614));
  OAI21_X1  g189(.A(new_n614), .B1(G868), .B2(new_n544), .ZN(G323));
  XNOR2_X1  g190(.A(G323), .B(KEYINPUT11), .ZN(G282));
  INV_X1    g191(.A(new_n481), .ZN(new_n617));
  AOI22_X1  g192(.A1(new_n477), .A2(G135), .B1(G123), .B2(new_n617), .ZN(new_n618));
  OR2_X1    g193(.A1(G99), .A2(G2105), .ZN(new_n619));
  OAI211_X1 g194(.A(new_n619), .B(G2104), .C1(G111), .C2(new_n459), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(G2096), .Z(new_n622));
  NAND2_X1  g197(.A1(new_n460), .A2(new_n490), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT12), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT13), .ZN(new_n625));
  XNOR2_X1  g200(.A(new_n625), .B(G2100), .ZN(new_n626));
  NAND2_X1  g201(.A1(new_n622), .A2(new_n626), .ZN(G156));
  XOR2_X1   g202(.A(KEYINPUT15), .B(G2435), .Z(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2438), .ZN(new_n629));
  XNOR2_X1  g204(.A(G2427), .B(G2430), .ZN(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(KEYINPUT81), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n629), .B(new_n631), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n632), .A2(KEYINPUT14), .ZN(new_n633));
  XNOR2_X1  g208(.A(KEYINPUT80), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n633), .B(new_n634), .ZN(new_n635));
  XNOR2_X1  g210(.A(G2443), .B(G2446), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(G2451), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2454), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n635), .B(new_n638), .ZN(new_n639));
  XOR2_X1   g214(.A(G1341), .B(G1348), .Z(new_n640));
  NOR2_X1   g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(new_n641), .B(KEYINPUT82), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n639), .A2(new_n640), .ZN(new_n643));
  AND3_X1   g218(.A1(new_n642), .A2(G14), .A3(new_n643), .ZN(G401));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  XOR2_X1   g220(.A(new_n645), .B(KEYINPUT85), .Z(new_n646));
  XNOR2_X1  g221(.A(new_n646), .B(KEYINPUT17), .ZN(new_n647));
  XOR2_X1   g222(.A(G2067), .B(G2678), .Z(new_n648));
  XOR2_X1   g223(.A(new_n648), .B(KEYINPUT84), .Z(new_n649));
  XNOR2_X1  g224(.A(G2084), .B(G2090), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT83), .ZN(new_n651));
  OAI21_X1  g226(.A(new_n647), .B1(new_n649), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g227(.A1(new_n649), .A2(new_n651), .ZN(new_n653));
  OR3_X1    g228(.A1(new_n649), .A2(new_n645), .A3(new_n651), .ZN(new_n654));
  NAND3_X1  g229(.A1(new_n652), .A2(new_n653), .A3(new_n654), .ZN(new_n655));
  NAND3_X1  g230(.A1(new_n649), .A2(new_n645), .A3(new_n651), .ZN(new_n656));
  XOR2_X1   g231(.A(new_n656), .B(KEYINPUT18), .Z(new_n657));
  NAND2_X1  g232(.A1(new_n655), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g233(.A(new_n658), .B(KEYINPUT86), .Z(new_n659));
  XOR2_X1   g234(.A(G2096), .B(G2100), .Z(new_n660));
  XOR2_X1   g235(.A(new_n659), .B(new_n660), .Z(new_n661));
  INV_X1    g236(.A(new_n661), .ZN(G227));
  XOR2_X1   g237(.A(G1956), .B(G2474), .Z(new_n663));
  XOR2_X1   g238(.A(G1961), .B(G1966), .Z(new_n664));
  NOR2_X1   g239(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n665), .ZN(new_n666));
  XNOR2_X1  g241(.A(G1971), .B(G1976), .ZN(new_n667));
  XNOR2_X1  g242(.A(new_n667), .B(KEYINPUT19), .ZN(new_n668));
  NOR2_X1   g243(.A1(new_n666), .A2(new_n668), .ZN(new_n669));
  XOR2_X1   g244(.A(new_n669), .B(KEYINPUT88), .Z(new_n670));
  NAND2_X1  g245(.A1(new_n663), .A2(new_n664), .ZN(new_n671));
  NOR2_X1   g246(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(KEYINPUT87), .B(KEYINPUT20), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n666), .A2(new_n668), .A3(new_n671), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n670), .A2(new_n674), .A3(new_n675), .ZN(new_n676));
  XNOR2_X1  g251(.A(KEYINPUT21), .B(G1986), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1991), .B(G1996), .Z(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT89), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  XOR2_X1   g256(.A(KEYINPUT22), .B(G1981), .Z(new_n682));
  XNOR2_X1  g257(.A(new_n681), .B(new_n682), .ZN(G229));
  XOR2_X1   g258(.A(KEYINPUT31), .B(G11), .Z(new_n684));
  INV_X1    g259(.A(G16), .ZN(new_n685));
  AND3_X1   g260(.A1(new_n685), .A2(KEYINPUT23), .A3(G20), .ZN(new_n686));
  AOI21_X1  g261(.A(KEYINPUT23), .B1(new_n685), .B2(G20), .ZN(new_n687));
  AOI211_X1 g262(.A(new_n686), .B(new_n687), .C1(G299), .C2(G16), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(G1956), .ZN(new_n689));
  INV_X1    g264(.A(G2090), .ZN(new_n690));
  INV_X1    g265(.A(G29), .ZN(new_n691));
  NAND2_X1  g266(.A1(new_n691), .A2(G35), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(G162), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(new_n693), .B(KEYINPUT29), .Z(new_n694));
  OAI21_X1  g269(.A(new_n689), .B1(new_n690), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g270(.A(new_n684), .B1(new_n695), .B2(KEYINPUT100), .ZN(new_n696));
  AOI22_X1  g271(.A1(new_n477), .A2(G140), .B1(G128), .B2(new_n617), .ZN(new_n697));
  OR2_X1    g272(.A1(G104), .A2(G2105), .ZN(new_n698));
  OAI211_X1 g273(.A(new_n698), .B(G2104), .C1(G116), .C2(new_n459), .ZN(new_n699));
  XOR2_X1   g274(.A(new_n699), .B(KEYINPUT94), .Z(new_n700));
  NAND2_X1  g275(.A1(new_n697), .A2(new_n700), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT95), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g278(.A1(new_n697), .A2(KEYINPUT95), .A3(new_n700), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n703), .A2(new_n704), .ZN(new_n705));
  INV_X1    g280(.A(new_n705), .ZN(new_n706));
  NOR2_X1   g281(.A1(new_n706), .A2(new_n691), .ZN(new_n707));
  AND2_X1   g282(.A1(new_n691), .A2(G26), .ZN(new_n708));
  OAI21_X1  g283(.A(KEYINPUT28), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(KEYINPUT28), .B2(new_n708), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n710), .B(G2067), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n685), .A2(G19), .ZN(new_n712));
  OAI21_X1  g287(.A(new_n712), .B1(new_n544), .B2(new_n685), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(G1341), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n711), .A2(new_n714), .ZN(new_n715));
  NOR2_X1   g290(.A1(G16), .A2(G22), .ZN(new_n716));
  AOI21_X1  g291(.A(new_n716), .B1(G166), .B2(G16), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT93), .ZN(new_n718));
  INV_X1    g293(.A(G1971), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n718), .B(new_n719), .ZN(new_n720));
  NOR2_X1   g295(.A1(G16), .A2(G23), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n574), .A2(KEYINPUT92), .ZN(new_n722));
  INV_X1    g297(.A(KEYINPUT92), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n567), .A2(new_n572), .A3(new_n723), .A4(new_n573), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n722), .A2(new_n724), .ZN(new_n725));
  AOI21_X1  g300(.A(new_n721), .B1(new_n725), .B2(G16), .ZN(new_n726));
  XNOR2_X1  g301(.A(KEYINPUT33), .B(G1976), .ZN(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  MUX2_X1   g303(.A(G6), .B(G305), .S(G16), .Z(new_n729));
  XOR2_X1   g304(.A(KEYINPUT32), .B(G1981), .Z(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  NAND3_X1  g306(.A1(new_n720), .A2(new_n728), .A3(new_n731), .ZN(new_n732));
  XOR2_X1   g307(.A(new_n732), .B(KEYINPUT34), .Z(new_n733));
  NOR2_X1   g308(.A1(new_n592), .A2(new_n685), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n734), .B1(new_n685), .B2(G24), .ZN(new_n735));
  INV_X1    g310(.A(G1986), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n735), .A2(new_n736), .ZN(new_n738));
  AOI22_X1  g313(.A1(new_n477), .A2(G131), .B1(G119), .B2(new_n617), .ZN(new_n739));
  OR2_X1    g314(.A1(G95), .A2(G2105), .ZN(new_n740));
  OAI211_X1 g315(.A(new_n740), .B(G2104), .C1(G107), .C2(new_n459), .ZN(new_n741));
  NAND2_X1  g316(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  MUX2_X1   g317(.A(G25), .B(new_n742), .S(G29), .Z(new_n743));
  XNOR2_X1  g318(.A(KEYINPUT90), .B(KEYINPUT91), .ZN(new_n744));
  XNOR2_X1  g319(.A(KEYINPUT35), .B(G1991), .ZN(new_n745));
  XNOR2_X1  g320(.A(new_n744), .B(new_n745), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n743), .B(new_n746), .ZN(new_n747));
  NAND4_X1  g322(.A1(new_n733), .A2(new_n737), .A3(new_n738), .A4(new_n747), .ZN(new_n748));
  AND2_X1   g323(.A1(new_n748), .A2(KEYINPUT36), .ZN(new_n749));
  NOR2_X1   g324(.A1(new_n748), .A2(KEYINPUT36), .ZN(new_n750));
  OAI211_X1 g325(.A(new_n696), .B(new_n715), .C1(new_n749), .C2(new_n750), .ZN(new_n751));
  NOR2_X1   g326(.A1(G29), .A2(G32), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n477), .A2(G141), .ZN(new_n753));
  XOR2_X1   g328(.A(new_n753), .B(KEYINPUT97), .Z(new_n754));
  AOI22_X1  g329(.A1(new_n617), .A2(G129), .B1(G105), .B2(new_n490), .ZN(new_n755));
  AND2_X1   g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT98), .ZN(new_n758));
  XNOR2_X1  g333(.A(new_n758), .B(KEYINPUT26), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n756), .A2(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(new_n760), .ZN(new_n761));
  AOI21_X1  g336(.A(new_n752), .B1(new_n761), .B2(G29), .ZN(new_n762));
  XNOR2_X1  g337(.A(KEYINPUT27), .B(G1996), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g339(.A(G2072), .ZN(new_n765));
  OR2_X1    g340(.A1(G29), .A2(G33), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n490), .A2(G103), .ZN(new_n767));
  XOR2_X1   g342(.A(new_n767), .B(KEYINPUT25), .Z(new_n768));
  AOI22_X1  g343(.A1(new_n460), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n769));
  INV_X1    g344(.A(G139), .ZN(new_n770));
  OAI221_X1 g345(.A(new_n768), .B1(new_n459), .B2(new_n769), .C1(new_n476), .C2(new_n770), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n766), .B1(new_n771), .B2(new_n691), .ZN(new_n772));
  OAI21_X1  g347(.A(new_n764), .B1(new_n765), .B2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(G171), .A2(G16), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G5), .B2(G16), .ZN(new_n775));
  INV_X1    g350(.A(G1961), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(KEYINPUT30), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(G28), .ZN(new_n779));
  NAND2_X1  g354(.A1(new_n778), .A2(G28), .ZN(new_n780));
  NAND3_X1  g355(.A1(new_n779), .A2(new_n780), .A3(new_n691), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n621), .B2(new_n691), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n694), .A2(new_n690), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n772), .A2(new_n765), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n775), .A2(new_n776), .ZN(new_n785));
  NAND3_X1  g360(.A1(new_n783), .A2(new_n784), .A3(new_n785), .ZN(new_n786));
  NOR4_X1   g361(.A1(new_n773), .A2(new_n777), .A3(new_n782), .A4(new_n786), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n695), .A2(KEYINPUT100), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n685), .A2(G21), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n789), .B1(G168), .B2(new_n685), .ZN(new_n790));
  INV_X1    g365(.A(G1966), .ZN(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n685), .A2(G4), .ZN(new_n793));
  OAI21_X1  g368(.A(new_n793), .B1(new_n599), .B2(new_n685), .ZN(new_n794));
  INV_X1    g369(.A(G1348), .ZN(new_n795));
  XNOR2_X1  g370(.A(new_n794), .B(new_n795), .ZN(new_n796));
  NAND4_X1  g371(.A1(new_n787), .A2(new_n788), .A3(new_n792), .A4(new_n796), .ZN(new_n797));
  OR2_X1    g372(.A1(KEYINPUT24), .A2(G34), .ZN(new_n798));
  NAND2_X1  g373(.A1(KEYINPUT24), .A2(G34), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n798), .A2(new_n691), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g375(.A(new_n800), .B1(G160), .B2(new_n691), .ZN(new_n801));
  XNOR2_X1  g376(.A(KEYINPUT96), .B(G2084), .ZN(new_n802));
  XNOR2_X1  g377(.A(new_n801), .B(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n691), .A2(G27), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G164), .B2(new_n691), .ZN(new_n805));
  XNOR2_X1  g380(.A(KEYINPUT99), .B(G2078), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  NOR4_X1   g382(.A1(new_n751), .A2(new_n797), .A3(new_n803), .A4(new_n807), .ZN(G311));
  INV_X1    g383(.A(G311), .ZN(G150));
  NAND2_X1  g384(.A1(new_n531), .A2(G55), .ZN(new_n810));
  AOI22_X1  g385(.A1(new_n507), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT101), .B(G93), .Z(new_n812));
  OAI221_X1 g387(.A(new_n810), .B1(new_n499), .B2(new_n811), .C1(new_n509), .C2(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n813), .A2(G860), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT37), .Z(new_n815));
  NAND2_X1  g390(.A1(new_n541), .A2(new_n543), .ZN(new_n816));
  XNOR2_X1  g391(.A(new_n816), .B(new_n813), .ZN(new_n817));
  XNOR2_X1  g392(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(new_n600), .A2(new_n610), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n819), .B(new_n820), .ZN(new_n821));
  OAI21_X1  g396(.A(new_n815), .B1(new_n821), .B2(G860), .ZN(G145));
  INV_X1    g397(.A(G160), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n621), .B(new_n823), .ZN(new_n824));
  XNOR2_X1  g399(.A(new_n824), .B(G162), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n705), .B(new_n771), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  AOI22_X1  g402(.A1(new_n477), .A2(G142), .B1(G130), .B2(new_n617), .ZN(new_n828));
  NOR2_X1   g403(.A1(G106), .A2(G2105), .ZN(new_n829));
  OAI21_X1  g404(.A(G2104), .B1(new_n459), .B2(G118), .ZN(new_n830));
  OAI21_X1  g405(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  XOR2_X1   g406(.A(new_n831), .B(new_n742), .Z(new_n832));
  XNOR2_X1  g407(.A(new_n760), .B(new_n832), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n827), .B(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n496), .B(new_n624), .ZN(new_n835));
  OR2_X1    g410(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  INV_X1    g411(.A(G37), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n834), .A2(new_n835), .ZN(new_n838));
  NAND3_X1  g413(.A1(new_n836), .A2(new_n837), .A3(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g415(.A(new_n544), .B(new_n813), .ZN(new_n841));
  XNOR2_X1  g416(.A(new_n613), .B(new_n841), .ZN(new_n842));
  INV_X1    g417(.A(KEYINPUT41), .ZN(new_n843));
  NOR2_X1   g418(.A1(G299), .A2(new_n600), .ZN(new_n844));
  AOI21_X1  g419(.A(new_n599), .B1(new_n561), .B2(new_n562), .ZN(new_n845));
  OAI21_X1  g420(.A(new_n843), .B1(new_n844), .B2(new_n845), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n844), .A2(new_n845), .ZN(new_n847));
  NAND2_X1  g422(.A1(new_n847), .A2(KEYINPUT41), .ZN(new_n848));
  NAND3_X1  g423(.A1(new_n842), .A2(new_n846), .A3(new_n848), .ZN(new_n849));
  INV_X1    g424(.A(new_n847), .ZN(new_n850));
  OAI21_X1  g425(.A(new_n849), .B1(new_n842), .B2(new_n850), .ZN(new_n851));
  INV_X1    g426(.A(KEYINPUT104), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  XOR2_X1   g428(.A(new_n725), .B(KEYINPUT102), .Z(new_n854));
  NAND2_X1  g429(.A1(new_n854), .A2(new_n592), .ZN(new_n855));
  XNOR2_X1  g430(.A(new_n725), .B(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(new_n856), .A2(G290), .ZN(new_n857));
  XNOR2_X1  g432(.A(G303), .B(G305), .ZN(new_n858));
  AND3_X1   g433(.A1(new_n855), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g434(.A(new_n858), .B1(new_n855), .B2(new_n857), .ZN(new_n860));
  NOR2_X1   g435(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  XNOR2_X1  g436(.A(KEYINPUT103), .B(KEYINPUT42), .ZN(new_n862));
  XNOR2_X1  g437(.A(new_n861), .B(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n853), .A2(new_n863), .ZN(new_n864));
  NOR2_X1   g439(.A1(new_n864), .A2(new_n601), .ZN(new_n865));
  OR2_X1    g440(.A1(new_n851), .A2(new_n852), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n866), .A2(new_n853), .A3(new_n863), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT105), .ZN(new_n869));
  AOI22_X1  g444(.A1(new_n865), .A2(new_n867), .B1(new_n601), .B2(new_n813), .ZN(new_n870));
  OAI21_X1  g445(.A(new_n869), .B1(new_n870), .B2(KEYINPUT105), .ZN(G295));
  OAI21_X1  g446(.A(new_n869), .B1(new_n870), .B2(KEYINPUT105), .ZN(G331));
  OAI21_X1  g447(.A(KEYINPUT106), .B1(new_n603), .B2(G286), .ZN(new_n873));
  NAND2_X1  g448(.A1(G286), .A2(G171), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n527), .A2(new_n528), .ZN(new_n875));
  NOR2_X1   g450(.A1(new_n509), .A2(new_n515), .ZN(new_n876));
  NOR2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  INV_X1    g452(.A(KEYINPUT106), .ZN(new_n878));
  NAND4_X1  g453(.A1(new_n877), .A2(G301), .A3(new_n878), .A4(new_n514), .ZN(new_n879));
  NAND3_X1  g454(.A1(new_n873), .A2(new_n874), .A3(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n880), .A2(new_n841), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n817), .A2(new_n873), .A3(new_n874), .A4(new_n879), .ZN(new_n882));
  NAND3_X1  g457(.A1(new_n881), .A2(new_n850), .A3(new_n882), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  AOI22_X1  g459(.A1(new_n881), .A2(new_n882), .B1(new_n848), .B2(new_n846), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n861), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  INV_X1    g461(.A(new_n861), .ZN(new_n887));
  AND2_X1   g462(.A1(new_n881), .A2(new_n882), .ZN(new_n888));
  AND2_X1   g463(.A1(new_n848), .A2(new_n846), .ZN(new_n889));
  OAI211_X1 g464(.A(new_n887), .B(new_n883), .C1(new_n888), .C2(new_n889), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n886), .A2(new_n890), .A3(new_n837), .ZN(new_n891));
  INV_X1    g466(.A(KEYINPUT43), .ZN(new_n892));
  NOR2_X1   g467(.A1(new_n892), .A2(KEYINPUT108), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(new_n893), .ZN(new_n895));
  NAND4_X1  g470(.A1(new_n886), .A2(new_n890), .A3(new_n837), .A4(new_n895), .ZN(new_n896));
  AND3_X1   g471(.A1(new_n894), .A2(KEYINPUT44), .A3(new_n896), .ZN(new_n897));
  OR2_X1    g472(.A1(new_n897), .A2(KEYINPUT109), .ZN(new_n898));
  AND2_X1   g473(.A1(new_n886), .A2(new_n890), .ZN(new_n899));
  NAND4_X1  g474(.A1(new_n899), .A2(KEYINPUT107), .A3(new_n892), .A4(new_n837), .ZN(new_n900));
  INV_X1    g475(.A(KEYINPUT107), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n901), .B1(new_n891), .B2(KEYINPUT43), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n891), .A2(KEYINPUT43), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n900), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT44), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n897), .B1(new_n904), .B2(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(KEYINPUT109), .ZN(new_n907));
  OAI21_X1  g482(.A(new_n898), .B1(new_n906), .B2(new_n907), .ZN(G397));
  AND2_X1   g483(.A1(new_n494), .A2(new_n495), .ZN(new_n909));
  AOI22_X1  g484(.A1(new_n488), .A2(G2105), .B1(G102), .B2(new_n490), .ZN(new_n910));
  AOI21_X1  g485(.A(G1384), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  NOR2_X1   g486(.A1(new_n911), .A2(KEYINPUT45), .ZN(new_n912));
  INV_X1    g487(.A(new_n912), .ZN(new_n913));
  NAND2_X1  g488(.A1(G160), .A2(G40), .ZN(new_n914));
  NOR2_X1   g489(.A1(new_n913), .A2(new_n914), .ZN(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  NAND3_X1  g491(.A1(new_n760), .A2(G1996), .A3(new_n915), .ZN(new_n917));
  XNOR2_X1  g492(.A(new_n917), .B(KEYINPUT110), .ZN(new_n918));
  INV_X1    g493(.A(G2067), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n705), .B(new_n919), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n920), .B1(G1996), .B2(new_n760), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n918), .B1(new_n915), .B2(new_n921), .ZN(new_n922));
  INV_X1    g497(.A(new_n745), .ZN(new_n923));
  NAND4_X1  g498(.A1(new_n922), .A2(new_n739), .A3(new_n741), .A4(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n706), .A2(new_n919), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n916), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  XNOR2_X1  g501(.A(new_n742), .B(new_n923), .ZN(new_n927));
  OAI21_X1  g502(.A(new_n922), .B1(new_n916), .B2(new_n927), .ZN(new_n928));
  NOR2_X1   g503(.A1(G290), .A2(G1986), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(new_n915), .ZN(new_n930));
  XNOR2_X1  g505(.A(new_n930), .B(KEYINPUT127), .ZN(new_n931));
  XOR2_X1   g506(.A(new_n931), .B(KEYINPUT48), .Z(new_n932));
  NOR2_X1   g507(.A1(new_n928), .A2(new_n932), .ZN(new_n933));
  AOI21_X1  g508(.A(new_n916), .B1(new_n761), .B2(new_n920), .ZN(new_n934));
  OAI21_X1  g509(.A(KEYINPUT46), .B1(new_n916), .B2(G1996), .ZN(new_n935));
  OR3_X1    g510(.A1(new_n916), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n936));
  AOI21_X1  g511(.A(new_n934), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  XOR2_X1   g512(.A(KEYINPUT126), .B(KEYINPUT47), .Z(new_n938));
  XNOR2_X1  g513(.A(new_n937), .B(new_n938), .ZN(new_n939));
  NOR3_X1   g514(.A1(new_n926), .A2(new_n933), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(KEYINPUT125), .ZN(new_n941));
  INV_X1    g516(.A(new_n929), .ZN(new_n942));
  NAND2_X1  g517(.A1(G290), .A2(G1986), .ZN(new_n943));
  AOI21_X1  g518(.A(new_n916), .B1(new_n942), .B2(new_n943), .ZN(new_n944));
  OR2_X1    g519(.A1(new_n928), .A2(new_n944), .ZN(new_n945));
  INV_X1    g520(.A(KEYINPUT120), .ZN(new_n946));
  INV_X1    g521(.A(KEYINPUT57), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n560), .A2(new_n947), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n551), .A2(new_n554), .A3(new_n559), .A4(KEYINPUT57), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n948), .A2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G1384), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n496), .A2(KEYINPUT45), .A3(new_n951), .ZN(new_n952));
  INV_X1    g527(.A(G40), .ZN(new_n953));
  NOR3_X1   g528(.A1(new_n463), .A2(new_n466), .A3(new_n953), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n952), .A2(new_n954), .ZN(new_n955));
  NOR2_X1   g530(.A1(new_n955), .A2(new_n912), .ZN(new_n956));
  XNOR2_X1  g531(.A(KEYINPUT56), .B(G2072), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  INV_X1    g533(.A(new_n487), .ZN(new_n959));
  AOI21_X1  g534(.A(new_n959), .B1(new_n460), .B2(G126), .ZN(new_n960));
  OAI21_X1  g535(.A(new_n491), .B1(new_n960), .B2(new_n459), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n494), .A2(new_n495), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n951), .B1(new_n961), .B2(new_n962), .ZN(new_n963));
  INV_X1    g538(.A(KEYINPUT111), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  OAI211_X1 g540(.A(KEYINPUT111), .B(new_n951), .C1(new_n961), .C2(new_n962), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n965), .A2(KEYINPUT50), .A3(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(KEYINPUT50), .ZN(new_n968));
  AOI21_X1  g543(.A(new_n914), .B1(new_n968), .B2(new_n911), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g545(.A(new_n950), .B(new_n958), .C1(new_n970), .C2(G1956), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n948), .A2(new_n949), .ZN(new_n972));
  AOI21_X1  g547(.A(G1956), .B1(new_n967), .B2(new_n969), .ZN(new_n973));
  INV_X1    g548(.A(new_n957), .ZN(new_n974));
  NOR3_X1   g549(.A1(new_n955), .A2(new_n912), .A3(new_n974), .ZN(new_n975));
  OAI21_X1  g550(.A(new_n972), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n971), .A2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(KEYINPUT61), .ZN(new_n978));
  AOI21_X1  g553(.A(KEYINPUT119), .B1(new_n977), .B2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT119), .ZN(new_n980));
  AOI211_X1 g555(.A(new_n980), .B(KEYINPUT61), .C1(new_n971), .C2(new_n976), .ZN(new_n981));
  NOR2_X1   g556(.A1(new_n979), .A2(new_n981), .ZN(new_n982));
  NOR2_X1   g557(.A1(new_n950), .A2(KEYINPUT118), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT118), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n984), .B1(new_n948), .B2(new_n949), .ZN(new_n985));
  OAI22_X1  g560(.A1(new_n983), .A2(new_n985), .B1(new_n973), .B2(new_n975), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n986), .A2(new_n971), .A3(KEYINPUT61), .ZN(new_n987));
  NOR3_X1   g562(.A1(new_n955), .A2(new_n912), .A3(G1996), .ZN(new_n988));
  XNOR2_X1  g563(.A(KEYINPUT58), .B(G1341), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n965), .A2(new_n966), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n989), .B1(new_n990), .B2(new_n954), .ZN(new_n991));
  OAI21_X1  g566(.A(new_n544), .B1(new_n988), .B2(new_n991), .ZN(new_n992));
  NAND2_X1  g567(.A1(new_n992), .A2(KEYINPUT59), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT59), .ZN(new_n994));
  OAI211_X1 g569(.A(new_n544), .B(new_n994), .C1(new_n988), .C2(new_n991), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n993), .A2(new_n995), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n987), .A2(new_n996), .ZN(new_n997));
  OAI21_X1  g572(.A(new_n946), .B1(new_n982), .B2(new_n997), .ZN(new_n998));
  AND2_X1   g573(.A1(new_n987), .A2(new_n996), .ZN(new_n999));
  OAI211_X1 g574(.A(new_n999), .B(KEYINPUT120), .C1(new_n979), .C2(new_n981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1001));
  AOI21_X1  g576(.A(KEYINPUT50), .B1(new_n965), .B2(new_n966), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n954), .B1(new_n911), .B2(new_n968), .ZN(new_n1003));
  NOR2_X1   g578(.A1(new_n1002), .A2(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(KEYINPUT117), .ZN(new_n1005));
  NAND2_X1  g580(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  OAI21_X1  g581(.A(KEYINPUT117), .B1(new_n1002), .B2(new_n1003), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n1006), .A2(new_n795), .A3(new_n1007), .ZN(new_n1008));
  NAND3_X1  g583(.A1(new_n990), .A2(new_n919), .A3(new_n954), .ZN(new_n1009));
  AND2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  OR2_X1    g585(.A1(new_n599), .A2(KEYINPUT60), .ZN(new_n1011));
  AOI21_X1  g586(.A(new_n1001), .B1(new_n1010), .B2(new_n1011), .ZN(new_n1012));
  AND4_X1   g587(.A1(new_n1009), .A2(new_n1008), .A3(new_n1011), .A4(new_n1001), .ZN(new_n1013));
  NOR2_X1   g588(.A1(new_n1012), .A2(new_n1013), .ZN(new_n1014));
  NAND3_X1  g589(.A1(new_n998), .A2(new_n1000), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(new_n986), .ZN(new_n1016));
  INV_X1    g591(.A(new_n971), .ZN(new_n1017));
  NOR2_X1   g592(.A1(new_n1010), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1016), .B1(new_n1018), .B2(new_n599), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1015), .A2(new_n1019), .ZN(new_n1020));
  INV_X1    g595(.A(G2084), .ZN(new_n1021));
  INV_X1    g596(.A(new_n955), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n1022), .B1(new_n990), .B2(KEYINPUT45), .ZN(new_n1023));
  AOI22_X1  g598(.A1(new_n1021), .A2(new_n1004), .B1(new_n1023), .B2(new_n791), .ZN(new_n1024));
  OAI21_X1  g599(.A(KEYINPUT51), .B1(new_n1024), .B2(G168), .ZN(new_n1025));
  INV_X1    g600(.A(G8), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n1026), .B1(new_n1024), .B2(G168), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1025), .A2(new_n1027), .ZN(new_n1028));
  INV_X1    g603(.A(KEYINPUT51), .ZN(new_n1029));
  OAI21_X1  g604(.A(new_n1028), .B1(new_n1029), .B2(new_n1027), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT55), .B1(G166), .B2(new_n1026), .ZN(new_n1031));
  INV_X1    g606(.A(KEYINPUT55), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n1032), .B(G8), .C1(new_n506), .C2(new_n511), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1031), .A2(new_n1033), .ZN(new_n1034));
  NAND3_X1  g609(.A1(new_n967), .A2(new_n969), .A3(new_n690), .ZN(new_n1035));
  OAI21_X1  g610(.A(new_n719), .B1(new_n955), .B2(new_n912), .ZN(new_n1036));
  AND2_X1   g611(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1034), .B1(new_n1037), .B2(new_n1026), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n725), .A2(G1976), .ZN(new_n1039));
  INV_X1    g614(.A(new_n966), .ZN(new_n1040));
  AOI21_X1  g615(.A(KEYINPUT111), .B1(new_n496), .B2(new_n951), .ZN(new_n1041));
  OAI21_X1  g616(.A(new_n954), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1039), .A2(new_n1042), .A3(G8), .ZN(new_n1043));
  XOR2_X1   g618(.A(KEYINPUT113), .B(G1976), .Z(new_n1044));
  NAND2_X1  g619(.A1(G288), .A2(new_n1044), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT52), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1045), .A2(new_n1046), .ZN(new_n1047));
  NOR2_X1   g622(.A1(new_n1043), .A2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g623(.A(new_n1026), .B1(new_n990), .B2(new_n954), .ZN(new_n1049));
  AOI21_X1  g624(.A(new_n1046), .B1(new_n1049), .B2(new_n1039), .ZN(new_n1050));
  NOR2_X1   g625(.A1(new_n1048), .A2(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1032), .B1(G303), .B2(G8), .ZN(new_n1052));
  INV_X1    g627(.A(new_n1033), .ZN(new_n1053));
  OAI21_X1  g628(.A(KEYINPUT112), .B1(new_n1052), .B2(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT112), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n1031), .A2(new_n1055), .A3(new_n1033), .ZN(new_n1056));
  NAND2_X1  g631(.A1(new_n1054), .A2(new_n1056), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n968), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1058));
  INV_X1    g633(.A(new_n1003), .ZN(new_n1059));
  NAND3_X1  g634(.A1(new_n1058), .A2(new_n1059), .A3(new_n690), .ZN(new_n1060));
  INV_X1    g635(.A(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1036), .ZN(new_n1062));
  OAI211_X1 g637(.A(G8), .B(new_n1057), .C1(new_n1061), .C2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(G1981), .ZN(new_n1064));
  NAND3_X1  g639(.A1(new_n582), .A2(new_n586), .A3(new_n1064), .ZN(new_n1065));
  AOI22_X1  g640(.A1(new_n583), .A2(new_n584), .B1(new_n500), .B2(new_n502), .ZN(new_n1066));
  OAI21_X1  g641(.A(G1981), .B1(new_n1066), .B2(new_n581), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n1065), .A2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g643(.A1(new_n1068), .A2(KEYINPUT49), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT49), .ZN(new_n1070));
  NAND3_X1  g645(.A1(new_n1065), .A2(new_n1067), .A3(new_n1070), .ZN(new_n1071));
  NAND2_X1  g646(.A1(new_n1069), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1042), .A2(new_n1072), .A3(G8), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT114), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1073), .A2(new_n1074), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1049), .A2(KEYINPUT114), .A3(new_n1072), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1075), .A2(new_n1076), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1038), .A2(new_n1051), .A3(new_n1063), .A4(new_n1077), .ZN(new_n1078));
  INV_X1    g653(.A(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1030), .A2(new_n1079), .ZN(new_n1080));
  XNOR2_X1  g655(.A(KEYINPUT121), .B(G1961), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1006), .A2(new_n1007), .A3(new_n1081), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT53), .ZN(new_n1083));
  INV_X1    g658(.A(new_n956), .ZN(new_n1084));
  OAI21_X1  g659(.A(new_n1083), .B1(new_n1084), .B2(G2078), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n913), .A2(KEYINPUT122), .A3(new_n954), .ZN(new_n1086));
  NOR2_X1   g661(.A1(new_n1083), .A2(G2078), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT122), .ZN(new_n1088));
  OAI21_X1  g663(.A(new_n1088), .B1(new_n912), .B2(new_n914), .ZN(new_n1089));
  NAND4_X1  g664(.A1(new_n1086), .A2(new_n952), .A3(new_n1087), .A4(new_n1089), .ZN(new_n1090));
  NAND3_X1  g665(.A1(new_n1082), .A2(new_n1085), .A3(new_n1090), .ZN(new_n1091));
  NAND2_X1  g666(.A1(new_n1091), .A2(G171), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1092), .A2(KEYINPUT123), .ZN(new_n1093));
  OAI211_X1 g668(.A(new_n1022), .B(new_n1087), .C1(new_n990), .C2(KEYINPUT45), .ZN(new_n1094));
  NAND3_X1  g669(.A1(new_n1082), .A2(new_n1094), .A3(new_n1085), .ZN(new_n1095));
  OR2_X1    g670(.A1(new_n1095), .A2(new_n603), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT123), .ZN(new_n1097));
  NAND3_X1  g672(.A1(new_n1091), .A2(new_n1097), .A3(G171), .ZN(new_n1098));
  NAND3_X1  g673(.A1(new_n1093), .A2(new_n1096), .A3(new_n1098), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(KEYINPUT54), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1095), .A2(new_n603), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT54), .ZN(new_n1102));
  OAI211_X1 g677(.A(new_n1101), .B(new_n1102), .C1(new_n603), .C2(new_n1091), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1080), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1101), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1105), .B1(new_n1030), .B2(KEYINPUT62), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1004), .A2(new_n1021), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1023), .A2(new_n791), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1107), .A2(new_n1108), .A3(G168), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1029), .B1(new_n1109), .B2(G8), .ZN(new_n1110));
  AOI21_X1  g685(.A(new_n1110), .B1(new_n1027), .B2(new_n1025), .ZN(new_n1111));
  INV_X1    g686(.A(KEYINPUT62), .ZN(new_n1112));
  OAI21_X1  g687(.A(new_n1079), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  OAI21_X1  g688(.A(KEYINPUT124), .B1(new_n1106), .B2(new_n1113), .ZN(new_n1114));
  AOI21_X1  g689(.A(new_n1078), .B1(new_n1030), .B2(KEYINPUT62), .ZN(new_n1115));
  INV_X1    g690(.A(KEYINPUT124), .ZN(new_n1116));
  AOI21_X1  g691(.A(new_n1101), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1117));
  NAND3_X1  g692(.A1(new_n1115), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  AOI22_X1  g693(.A1(new_n1020), .A2(new_n1104), .B1(new_n1114), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(KEYINPUT115), .ZN(new_n1120));
  NAND3_X1  g695(.A1(new_n1109), .A2(G8), .A3(G168), .ZN(new_n1121));
  OAI21_X1  g696(.A(new_n1120), .B1(new_n1078), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1049), .A2(new_n1046), .A3(new_n1039), .A4(new_n1045), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1043), .A2(KEYINPUT52), .ZN(new_n1124));
  AOI21_X1  g699(.A(KEYINPUT114), .B1(new_n1049), .B2(new_n1072), .ZN(new_n1125));
  AND4_X1   g700(.A1(KEYINPUT114), .A2(new_n1042), .A3(G8), .A4(new_n1072), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1123), .B(new_n1124), .C1(new_n1125), .C2(new_n1126), .ZN(new_n1127));
  AOI221_X4 g702(.A(new_n1026), .B1(new_n1054), .B2(new_n1056), .C1(new_n1060), .C2(new_n1036), .ZN(new_n1128));
  NOR2_X1   g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NOR3_X1   g704(.A1(new_n1024), .A2(new_n1026), .A3(G286), .ZN(new_n1130));
  NAND4_X1  g705(.A1(new_n1129), .A2(KEYINPUT115), .A3(new_n1038), .A4(new_n1130), .ZN(new_n1131));
  INV_X1    g706(.A(KEYINPUT63), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1122), .A2(new_n1131), .A3(new_n1132), .ZN(new_n1133));
  OAI21_X1  g708(.A(G8), .B1(new_n1061), .B2(new_n1062), .ZN(new_n1134));
  AOI21_X1  g709(.A(new_n1132), .B1(new_n1134), .B2(new_n1034), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1129), .A2(new_n1130), .A3(new_n1135), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1133), .A2(new_n1136), .ZN(new_n1137));
  NOR2_X1   g712(.A1(G305), .A2(G1981), .ZN(new_n1138));
  NOR2_X1   g713(.A1(G288), .A2(G1976), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1138), .B1(new_n1077), .B2(new_n1139), .ZN(new_n1140));
  INV_X1    g715(.A(new_n1049), .ZN(new_n1141));
  NOR2_X1   g716(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1127), .A2(new_n1063), .ZN(new_n1143));
  OR2_X1    g718(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  INV_X1    g719(.A(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(KEYINPUT116), .B1(new_n1137), .B2(new_n1145), .ZN(new_n1146));
  INV_X1    g721(.A(KEYINPUT116), .ZN(new_n1147));
  AOI211_X1 g722(.A(new_n1147), .B(new_n1144), .C1(new_n1133), .C2(new_n1136), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1146), .A2(new_n1148), .ZN(new_n1149));
  AOI211_X1 g724(.A(new_n941), .B(new_n945), .C1(new_n1119), .C2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1020), .A2(new_n1104), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1137), .A2(new_n1145), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1152), .A2(new_n1147), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1137), .A2(KEYINPUT116), .A3(new_n1145), .ZN(new_n1155));
  NAND4_X1  g730(.A1(new_n1151), .A2(new_n1153), .A3(new_n1154), .A4(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(new_n945), .ZN(new_n1157));
  AOI21_X1  g732(.A(KEYINPUT125), .B1(new_n1156), .B2(new_n1157), .ZN(new_n1158));
  OAI21_X1  g733(.A(new_n940), .B1(new_n1150), .B2(new_n1158), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g734(.A1(G401), .A2(G229), .ZN(new_n1161));
  AND2_X1   g735(.A1(new_n839), .A2(new_n1161), .ZN(new_n1162));
  NAND4_X1  g736(.A1(new_n1162), .A2(G319), .A3(new_n661), .A4(new_n904), .ZN(G225));
  INV_X1    g737(.A(G225), .ZN(G308));
endmodule


