//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n544, new_n545, new_n546, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n568, new_n569, new_n571, new_n572, new_n573, new_n574,
    new_n575, new_n576, new_n577, new_n578, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n593, new_n594, new_n595, new_n596, new_n597, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n624, new_n625, new_n628, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n696, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1199, new_n1200, new_n1201;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(new_n451), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n455), .A2(G2106), .ZN(new_n456));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  OR2_X1    g032(.A1(new_n452), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n456), .A2(new_n458), .ZN(new_n459));
  INV_X1    g034(.A(new_n459), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(G125), .ZN(new_n462));
  OR2_X1    g037(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n463));
  NAND2_X1  g038(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OAI21_X1  g040(.A(new_n461), .B1(new_n465), .B2(KEYINPUT68), .ZN(new_n466));
  AND2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NOR2_X1   g042(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n468));
  OAI211_X1 g043(.A(KEYINPUT68), .B(G125), .C1(new_n467), .C2(new_n468), .ZN(new_n469));
  INV_X1    g044(.A(new_n469), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n466), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n467), .A2(new_n468), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n474), .A2(G101), .A3(G2104), .ZN(new_n475));
  OR2_X1    g050(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n475), .A2(KEYINPUT69), .ZN(new_n477));
  AOI22_X1  g052(.A1(new_n473), .A2(G137), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  XNOR2_X1  g054(.A(new_n479), .B(KEYINPUT70), .ZN(G160));
  NOR2_X1   g055(.A1(new_n472), .A2(KEYINPUT71), .ZN(new_n481));
  AND3_X1   g056(.A1(new_n463), .A2(KEYINPUT71), .A3(new_n464), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n483), .A2(G2105), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G136), .ZN(new_n485));
  OAI21_X1  g060(.A(G2105), .B1(new_n481), .B2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(G124), .ZN(new_n488));
  NOR2_X1   g063(.A1(new_n474), .A2(G112), .ZN(new_n489));
  OAI21_X1  g064(.A(G2104), .B1(G100), .B2(G2105), .ZN(new_n490));
  OAI211_X1 g065(.A(new_n485), .B(new_n488), .C1(new_n489), .C2(new_n490), .ZN(new_n491));
  XOR2_X1   g066(.A(new_n491), .B(KEYINPUT72), .Z(G162));
  INV_X1    g067(.A(G138), .ZN(new_n493));
  NOR2_X1   g068(.A1(new_n493), .A2(G2105), .ZN(new_n494));
  OAI211_X1 g069(.A(new_n494), .B(KEYINPUT75), .C1(new_n468), .C2(new_n467), .ZN(new_n495));
  INV_X1    g070(.A(KEYINPUT4), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT73), .ZN(new_n498));
  OAI21_X1  g073(.A(new_n498), .B1(new_n474), .B2(G114), .ZN(new_n499));
  INV_X1    g074(.A(G114), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n501));
  OR2_X1    g076(.A1(G102), .A2(G2105), .ZN(new_n502));
  NAND4_X1  g077(.A1(new_n499), .A2(new_n501), .A3(new_n502), .A4(G2104), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n463), .A2(new_n464), .ZN(new_n504));
  NAND3_X1  g079(.A1(new_n504), .A2(G126), .A3(G2105), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n497), .A2(new_n503), .A3(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT74), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n474), .A2(G138), .ZN(new_n508));
  AOI21_X1  g083(.A(new_n508), .B1(new_n463), .B2(new_n464), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(KEYINPUT4), .ZN(new_n510));
  AOI22_X1  g085(.A1(new_n507), .A2(new_n495), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  NOR2_X1   g086(.A1(new_n506), .A2(new_n511), .ZN(G164));
  INV_X1    g087(.A(KEYINPUT77), .ZN(new_n513));
  AND3_X1   g088(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT5), .B1(KEYINPUT76), .B2(G543), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n514), .A2(new_n515), .ZN(new_n516));
  AND2_X1   g091(.A1(KEYINPUT6), .A2(G651), .ZN(new_n517));
  NOR2_X1   g092(.A1(KEYINPUT6), .A2(G651), .ZN(new_n518));
  NOR2_X1   g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  OAI21_X1  g094(.A(new_n513), .B1(new_n516), .B2(new_n519), .ZN(new_n520));
  OAI221_X1 g095(.A(KEYINPUT77), .B1(new_n517), .B2(new_n518), .C1(new_n514), .C2(new_n515), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(new_n522), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(G88), .ZN(new_n524));
  NAND2_X1  g099(.A1(G75), .A2(G543), .ZN(new_n525));
  INV_X1    g100(.A(G62), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n516), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g102(.A(G543), .B1(new_n517), .B2(new_n518), .ZN(new_n528));
  INV_X1    g103(.A(new_n528), .ZN(new_n529));
  AOI22_X1  g104(.A1(new_n527), .A2(G651), .B1(G50), .B2(new_n529), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n524), .A2(new_n530), .ZN(G303));
  INV_X1    g106(.A(G303), .ZN(G166));
  INV_X1    g107(.A(KEYINPUT78), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n516), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g109(.A1(KEYINPUT76), .A2(G543), .ZN(new_n535));
  INV_X1    g110(.A(KEYINPUT5), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n535), .A2(new_n536), .ZN(new_n537));
  NAND3_X1  g112(.A1(KEYINPUT76), .A2(KEYINPUT5), .A3(G543), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g114(.A1(new_n539), .A2(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n534), .A2(new_n540), .A3(G63), .A4(G651), .ZN(new_n541));
  NAND3_X1  g116(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n543));
  OR2_X1    g118(.A1(new_n542), .A2(KEYINPUT7), .ZN(new_n544));
  AOI22_X1  g119(.A1(new_n529), .A2(G51), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G89), .ZN(new_n546));
  OAI211_X1 g121(.A(new_n541), .B(new_n545), .C1(new_n522), .C2(new_n546), .ZN(G286));
  INV_X1    g122(.A(G286), .ZN(G168));
  INV_X1    g123(.A(G651), .ZN(new_n549));
  AND2_X1   g124(.A1(new_n534), .A2(new_n540), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G64), .ZN(new_n551));
  NAND2_X1  g126(.A1(G77), .A2(G543), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n549), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n529), .A2(G52), .ZN(new_n554));
  INV_X1    g129(.A(G90), .ZN(new_n555));
  OAI21_X1  g130(.A(new_n554), .B1(new_n522), .B2(new_n555), .ZN(new_n556));
  NOR2_X1   g131(.A1(new_n553), .A2(new_n556), .ZN(G171));
  NAND2_X1  g132(.A1(new_n529), .A2(G43), .ZN(new_n558));
  INV_X1    g133(.A(G81), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n558), .B1(new_n522), .B2(new_n559), .ZN(new_n560));
  NAND3_X1  g135(.A1(new_n534), .A2(new_n540), .A3(G56), .ZN(new_n561));
  NAND2_X1  g136(.A1(G68), .A2(G543), .ZN(new_n562));
  AOI21_X1  g137(.A(new_n549), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  NOR2_X1   g138(.A1(new_n560), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n564), .A2(G860), .ZN(new_n565));
  XOR2_X1   g140(.A(new_n565), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g141(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g142(.A1(G1), .A2(G3), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT8), .ZN(new_n569));
  NAND4_X1  g144(.A1(G319), .A2(G483), .A3(G661), .A4(new_n569), .ZN(G188));
  NAND2_X1  g145(.A1(new_n523), .A2(G91), .ZN(new_n571));
  OAI211_X1 g146(.A(G53), .B(G543), .C1(new_n517), .C2(new_n518), .ZN(new_n572));
  OR2_X1    g147(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n572), .A2(KEYINPUT9), .ZN(new_n574));
  NAND2_X1  g149(.A1(G78), .A2(G543), .ZN(new_n575));
  INV_X1    g150(.A(G65), .ZN(new_n576));
  OAI21_X1  g151(.A(new_n575), .B1(new_n516), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g152(.A1(new_n573), .A2(new_n574), .B1(new_n577), .B2(G651), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n571), .A2(new_n578), .ZN(G299));
  INV_X1    g154(.A(G171), .ZN(G301));
  NAND2_X1  g155(.A1(new_n534), .A2(new_n540), .ZN(new_n581));
  INV_X1    g156(.A(G74), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  AOI22_X1  g158(.A1(new_n583), .A2(G651), .B1(G49), .B2(new_n529), .ZN(new_n584));
  INV_X1    g159(.A(G87), .ZN(new_n585));
  OAI21_X1  g160(.A(new_n584), .B1(new_n585), .B2(new_n522), .ZN(G288));
  NAND2_X1  g161(.A1(G73), .A2(G543), .ZN(new_n587));
  INV_X1    g162(.A(G61), .ZN(new_n588));
  OAI21_X1  g163(.A(new_n587), .B1(new_n516), .B2(new_n588), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n589), .A2(G651), .ZN(new_n590));
  INV_X1    g165(.A(KEYINPUT80), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n539), .A2(G61), .ZN(new_n593));
  AOI21_X1  g168(.A(new_n549), .B1(new_n593), .B2(new_n587), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n594), .A2(KEYINPUT80), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n520), .A2(new_n521), .A3(G86), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n529), .A2(G48), .ZN(new_n597));
  NAND4_X1  g172(.A1(new_n592), .A2(new_n595), .A3(new_n596), .A4(new_n597), .ZN(G305));
  NAND2_X1  g173(.A1(new_n550), .A2(G60), .ZN(new_n599));
  NAND2_X1  g174(.A1(G72), .A2(G543), .ZN(new_n600));
  AOI21_X1  g175(.A(new_n549), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n529), .A2(G47), .ZN(new_n602));
  INV_X1    g177(.A(G85), .ZN(new_n603));
  OAI21_X1  g178(.A(new_n602), .B1(new_n522), .B2(new_n603), .ZN(new_n604));
  NOR2_X1   g179(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  INV_X1    g180(.A(new_n605), .ZN(G290));
  NAND2_X1  g181(.A1(G301), .A2(G868), .ZN(new_n607));
  NAND2_X1  g182(.A1(G79), .A2(G543), .ZN(new_n608));
  INV_X1    g183(.A(G66), .ZN(new_n609));
  OAI21_X1  g184(.A(new_n608), .B1(new_n516), .B2(new_n609), .ZN(new_n610));
  AOI22_X1  g185(.A1(new_n610), .A2(G651), .B1(G54), .B2(new_n529), .ZN(new_n611));
  INV_X1    g186(.A(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(G92), .ZN(new_n613));
  OAI21_X1  g188(.A(KEYINPUT81), .B1(new_n522), .B2(new_n613), .ZN(new_n614));
  INV_X1    g189(.A(KEYINPUT81), .ZN(new_n615));
  NAND4_X1  g190(.A1(new_n520), .A2(new_n521), .A3(new_n615), .A4(G92), .ZN(new_n616));
  NAND2_X1  g191(.A1(new_n614), .A2(new_n616), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n617), .A2(KEYINPUT10), .ZN(new_n618));
  INV_X1    g193(.A(KEYINPUT10), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n614), .A2(new_n619), .A3(new_n616), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n612), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g196(.A(new_n607), .B1(new_n621), .B2(G868), .ZN(G284));
  OAI21_X1  g197(.A(new_n607), .B1(new_n621), .B2(G868), .ZN(G321));
  NAND2_X1  g198(.A1(G286), .A2(G868), .ZN(new_n624));
  INV_X1    g199(.A(G299), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G297));
  OAI21_X1  g201(.A(new_n624), .B1(new_n625), .B2(G868), .ZN(G280));
  INV_X1    g202(.A(G559), .ZN(new_n628));
  OAI21_X1  g203(.A(new_n621), .B1(new_n628), .B2(G860), .ZN(G148));
  NAND2_X1  g204(.A1(new_n621), .A2(new_n628), .ZN(new_n630));
  INV_X1    g205(.A(new_n630), .ZN(new_n631));
  INV_X1    g206(.A(G868), .ZN(new_n632));
  OR3_X1    g207(.A1(new_n631), .A2(KEYINPUT82), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g208(.A(KEYINPUT82), .B1(new_n631), .B2(new_n632), .ZN(new_n634));
  OAI211_X1 g209(.A(new_n633), .B(new_n634), .C1(G868), .C2(new_n564), .ZN(G323));
  XNOR2_X1  g210(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g211(.A1(new_n473), .A2(G2104), .ZN(new_n637));
  XNOR2_X1  g212(.A(KEYINPUT83), .B(KEYINPUT12), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(new_n639), .B(KEYINPUT13), .ZN(new_n640));
  XOR2_X1   g215(.A(new_n640), .B(G2100), .Z(new_n641));
  NAND2_X1  g216(.A1(new_n484), .A2(G135), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n487), .A2(G123), .ZN(new_n643));
  NOR2_X1   g218(.A1(new_n474), .A2(G111), .ZN(new_n644));
  OAI21_X1  g219(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n645));
  OAI211_X1 g220(.A(new_n642), .B(new_n643), .C1(new_n644), .C2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(KEYINPUT84), .B(G2096), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  NAND2_X1  g223(.A1(new_n641), .A2(new_n648), .ZN(G156));
  XNOR2_X1  g224(.A(G2451), .B(G2454), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT16), .ZN(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT86), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n658), .ZN(new_n661));
  NAND2_X1  g236(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XOR2_X1   g237(.A(G2443), .B(G2446), .Z(new_n663));
  NAND2_X1  g238(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  XNOR2_X1  g239(.A(G1341), .B(G1348), .ZN(new_n665));
  XOR2_X1   g240(.A(new_n665), .B(KEYINPUT87), .Z(new_n666));
  INV_X1    g241(.A(new_n663), .ZN(new_n667));
  NAND3_X1  g242(.A1(new_n660), .A2(new_n661), .A3(new_n667), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n664), .A2(new_n666), .A3(new_n668), .ZN(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n666), .B1(new_n664), .B2(new_n668), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n652), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n673), .A2(new_n651), .A3(new_n669), .ZN(new_n674));
  NAND3_X1  g249(.A1(new_n672), .A2(new_n674), .A3(G14), .ZN(new_n675));
  INV_X1    g250(.A(KEYINPUT88), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  NAND4_X1  g252(.A1(new_n672), .A2(new_n674), .A3(KEYINPUT88), .A4(G14), .ZN(new_n678));
  AND2_X1   g253(.A1(new_n677), .A2(new_n678), .ZN(G401));
  XOR2_X1   g254(.A(G2084), .B(G2090), .Z(new_n680));
  XNOR2_X1  g255(.A(G2067), .B(G2678), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT90), .ZN(new_n682));
  XNOR2_X1  g257(.A(G2072), .B(G2078), .ZN(new_n683));
  INV_X1    g258(.A(new_n683), .ZN(new_n684));
  AOI21_X1  g259(.A(new_n680), .B1(new_n682), .B2(new_n684), .ZN(new_n685));
  XOR2_X1   g260(.A(new_n683), .B(KEYINPUT17), .Z(new_n686));
  OAI21_X1  g261(.A(new_n685), .B1(new_n682), .B2(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT91), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n686), .A2(new_n682), .A3(new_n680), .ZN(new_n689));
  NAND3_X1  g264(.A1(new_n680), .A2(new_n681), .A3(new_n683), .ZN(new_n690));
  XOR2_X1   g265(.A(KEYINPUT89), .B(KEYINPUT18), .Z(new_n691));
  XNOR2_X1  g266(.A(new_n690), .B(new_n691), .ZN(new_n692));
  NAND3_X1  g267(.A1(new_n688), .A2(new_n689), .A3(new_n692), .ZN(new_n693));
  XOR2_X1   g268(.A(G2096), .B(G2100), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(G227));
  XNOR2_X1  g270(.A(G1971), .B(G1976), .ZN(new_n696));
  INV_X1    g271(.A(KEYINPUT19), .ZN(new_n697));
  XNOR2_X1  g272(.A(new_n696), .B(new_n697), .ZN(new_n698));
  XOR2_X1   g273(.A(G1956), .B(G2474), .Z(new_n699));
  XOR2_X1   g274(.A(G1961), .B(G1966), .Z(new_n700));
  AND2_X1   g275(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n698), .A2(new_n701), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n702), .B(KEYINPUT20), .ZN(new_n703));
  NOR2_X1   g278(.A1(new_n699), .A2(new_n700), .ZN(new_n704));
  NOR3_X1   g279(.A1(new_n698), .A2(new_n701), .A3(new_n704), .ZN(new_n705));
  AOI21_X1  g280(.A(new_n705), .B1(new_n698), .B2(new_n704), .ZN(new_n706));
  AND2_X1   g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n707), .B(new_n708), .ZN(new_n709));
  XNOR2_X1  g284(.A(G1991), .B(G1996), .ZN(new_n710));
  XNOR2_X1  g285(.A(new_n709), .B(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(G1981), .B(G1986), .ZN(new_n712));
  AND2_X1   g287(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  NOR2_X1   g288(.A1(new_n711), .A2(new_n712), .ZN(new_n714));
  NOR2_X1   g289(.A1(new_n713), .A2(new_n714), .ZN(G229));
  MUX2_X1   g290(.A(G6), .B(G305), .S(G16), .Z(new_n716));
  XOR2_X1   g291(.A(KEYINPUT32), .B(G1981), .Z(new_n717));
  XNOR2_X1  g292(.A(new_n716), .B(new_n717), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n718), .A2(KEYINPUT93), .ZN(new_n720));
  INV_X1    g295(.A(G16), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n721), .A2(G23), .ZN(new_n722));
  INV_X1    g297(.A(G288), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n722), .B1(new_n723), .B2(new_n721), .ZN(new_n724));
  XOR2_X1   g299(.A(KEYINPUT33), .B(G1976), .Z(new_n725));
  NAND2_X1  g300(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n721), .A2(G22), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(G166), .B2(new_n721), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(G1971), .ZN(new_n729));
  INV_X1    g304(.A(new_n725), .ZN(new_n730));
  OAI211_X1 g305(.A(new_n722), .B(new_n730), .C1(new_n723), .C2(new_n721), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n728), .A2(G1971), .ZN(new_n732));
  AND4_X1   g307(.A1(new_n726), .A2(new_n729), .A3(new_n731), .A4(new_n732), .ZN(new_n733));
  NAND3_X1  g308(.A1(new_n719), .A2(new_n720), .A3(new_n733), .ZN(new_n734));
  OR2_X1    g309(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n735));
  NAND2_X1  g310(.A1(new_n734), .A2(KEYINPUT34), .ZN(new_n736));
  NOR2_X1   g311(.A1(G16), .A2(G24), .ZN(new_n737));
  XNOR2_X1  g312(.A(new_n605), .B(KEYINPUT92), .ZN(new_n738));
  AOI21_X1  g313(.A(new_n737), .B1(new_n738), .B2(G16), .ZN(new_n739));
  INV_X1    g314(.A(G1986), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  INV_X1    g316(.A(G29), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n742), .A2(G25), .ZN(new_n743));
  OR2_X1    g318(.A1(new_n474), .A2(G107), .ZN(new_n744));
  OAI21_X1  g319(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n745));
  INV_X1    g320(.A(new_n745), .ZN(new_n746));
  AOI22_X1  g321(.A1(new_n487), .A2(G119), .B1(new_n744), .B2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n484), .A2(G131), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g324(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n743), .B1(new_n750), .B2(new_n742), .ZN(new_n751));
  XOR2_X1   g326(.A(KEYINPUT35), .B(G1991), .Z(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND4_X1  g328(.A1(new_n735), .A2(new_n736), .A3(new_n741), .A4(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n755));
  OR2_X1    g330(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  OR2_X1    g331(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n754), .A2(new_n755), .A3(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n742), .A2(G35), .ZN(new_n759));
  XOR2_X1   g334(.A(new_n759), .B(KEYINPUT101), .Z(new_n760));
  OAI21_X1  g335(.A(new_n760), .B1(G162), .B2(new_n742), .ZN(new_n761));
  INV_X1    g336(.A(KEYINPUT29), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n761), .B(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(G2090), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g340(.A1(new_n721), .A2(G21), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(G168), .B2(new_n721), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n767), .B(G1966), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n484), .A2(G141), .ZN(new_n769));
  NAND2_X1  g344(.A1(new_n487), .A2(G129), .ZN(new_n770));
  NAND3_X1  g345(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n771));
  INV_X1    g346(.A(KEYINPUT26), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n771), .A2(new_n772), .ZN(new_n774));
  AND2_X1   g349(.A1(new_n474), .A2(G2104), .ZN(new_n775));
  AOI22_X1  g350(.A1(new_n773), .A2(new_n774), .B1(G105), .B2(new_n775), .ZN(new_n776));
  NAND3_X1  g351(.A1(new_n769), .A2(new_n770), .A3(new_n776), .ZN(new_n777));
  INV_X1    g352(.A(new_n777), .ZN(new_n778));
  NOR2_X1   g353(.A1(new_n778), .A2(new_n742), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n742), .B2(G32), .ZN(new_n780));
  XNOR2_X1  g355(.A(KEYINPUT27), .B(G1996), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n768), .B1(new_n780), .B2(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n742), .A2(G33), .ZN(new_n783));
  NAND3_X1  g358(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT25), .Z(new_n785));
  AOI22_X1  g360(.A1(new_n504), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n785), .B1(new_n786), .B2(new_n474), .ZN(new_n787));
  AOI21_X1  g362(.A(new_n787), .B1(new_n484), .B2(G139), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n783), .B1(new_n788), .B2(new_n742), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2072), .ZN(new_n790));
  NOR2_X1   g365(.A1(new_n780), .A2(new_n781), .ZN(new_n791));
  NOR2_X1   g366(.A1(G5), .A2(G16), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n792), .B1(G171), .B2(G16), .ZN(new_n793));
  XNOR2_X1  g368(.A(KEYINPUT99), .B(G1961), .ZN(new_n794));
  AOI211_X1 g369(.A(new_n790), .B(new_n791), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  NOR2_X1   g370(.A1(new_n793), .A2(new_n794), .ZN(new_n796));
  INV_X1    g371(.A(KEYINPUT100), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n742), .A2(G27), .ZN(new_n798));
  OAI21_X1  g373(.A(new_n798), .B1(G164), .B2(new_n742), .ZN(new_n799));
  INV_X1    g374(.A(G2078), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n799), .B(new_n800), .ZN(new_n801));
  AOI21_X1  g376(.A(new_n796), .B1(new_n797), .B2(new_n801), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n765), .A2(new_n782), .A3(new_n795), .A4(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n621), .A2(G16), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(G4), .B2(G16), .ZN(new_n805));
  XOR2_X1   g380(.A(KEYINPUT95), .B(G1348), .Z(new_n806));
  NAND2_X1  g381(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  OR2_X1    g382(.A1(new_n805), .A2(new_n806), .ZN(new_n808));
  OAI211_X1 g383(.A(new_n807), .B(new_n808), .C1(new_n763), .C2(new_n764), .ZN(new_n809));
  NOR2_X1   g384(.A1(new_n801), .A2(new_n797), .ZN(new_n810));
  NAND2_X1  g385(.A1(new_n721), .A2(G20), .ZN(new_n811));
  XOR2_X1   g386(.A(new_n811), .B(KEYINPUT23), .Z(new_n812));
  AOI21_X1  g387(.A(new_n812), .B1(G299), .B2(G16), .ZN(new_n813));
  INV_X1    g388(.A(G1956), .ZN(new_n814));
  XNOR2_X1  g389(.A(new_n813), .B(new_n814), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n721), .A2(G19), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n564), .B2(new_n721), .ZN(new_n817));
  AOI211_X1 g392(.A(new_n810), .B(new_n815), .C1(G1341), .C2(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n742), .A2(G26), .ZN(new_n819));
  XOR2_X1   g394(.A(new_n819), .B(KEYINPUT28), .Z(new_n820));
  NAND3_X1  g395(.A1(new_n487), .A2(KEYINPUT96), .A3(G128), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT96), .ZN(new_n822));
  INV_X1    g397(.A(G128), .ZN(new_n823));
  OAI21_X1  g398(.A(new_n822), .B1(new_n486), .B2(new_n823), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n821), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n826));
  INV_X1    g401(.A(G116), .ZN(new_n827));
  AOI21_X1  g402(.A(new_n826), .B1(new_n827), .B2(G2105), .ZN(new_n828));
  OR2_X1    g403(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n829));
  NAND2_X1  g404(.A1(new_n828), .A2(KEYINPUT97), .ZN(new_n830));
  AOI22_X1  g405(.A1(new_n484), .A2(G140), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n825), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g407(.A(new_n820), .B1(new_n832), .B2(G29), .ZN(new_n833));
  INV_X1    g408(.A(G2067), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n833), .B(new_n834), .ZN(new_n835));
  XNOR2_X1  g410(.A(KEYINPUT30), .B(G28), .ZN(new_n836));
  OR2_X1    g411(.A1(KEYINPUT31), .A2(G11), .ZN(new_n837));
  NAND2_X1  g412(.A1(KEYINPUT31), .A2(G11), .ZN(new_n838));
  AOI22_X1  g413(.A1(new_n836), .A2(new_n742), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n646), .B2(new_n742), .ZN(new_n840));
  XNOR2_X1  g415(.A(new_n840), .B(KEYINPUT98), .ZN(new_n841));
  NOR2_X1   g416(.A1(new_n817), .A2(G1341), .ZN(new_n842));
  NOR3_X1   g417(.A1(new_n835), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  INV_X1    g418(.A(G34), .ZN(new_n844));
  AND2_X1   g419(.A1(new_n844), .A2(KEYINPUT24), .ZN(new_n845));
  NOR2_X1   g420(.A1(new_n844), .A2(KEYINPUT24), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n742), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n847), .B1(G160), .B2(new_n742), .ZN(new_n848));
  INV_X1    g423(.A(G2084), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n818), .A2(new_n843), .A3(new_n850), .ZN(new_n851));
  NOR3_X1   g426(.A1(new_n803), .A2(new_n809), .A3(new_n851), .ZN(new_n852));
  AND3_X1   g427(.A1(new_n756), .A2(new_n758), .A3(new_n852), .ZN(G311));
  NAND3_X1  g428(.A1(new_n756), .A2(new_n758), .A3(new_n852), .ZN(G150));
  NAND3_X1  g429(.A1(new_n534), .A2(new_n540), .A3(G67), .ZN(new_n855));
  INV_X1    g430(.A(KEYINPUT102), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n856), .B1(new_n855), .B2(new_n857), .ZN(new_n859));
  NOR3_X1   g434(.A1(new_n858), .A2(new_n859), .A3(new_n549), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n529), .A2(G55), .ZN(new_n861));
  INV_X1    g436(.A(G93), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n861), .B1(new_n522), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  INV_X1    g439(.A(G860), .ZN(new_n865));
  NOR2_X1   g440(.A1(new_n864), .A2(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT37), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n621), .A2(G559), .ZN(new_n868));
  XNOR2_X1  g443(.A(new_n868), .B(KEYINPUT103), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT38), .ZN(new_n870));
  INV_X1    g445(.A(new_n564), .ZN(new_n871));
  OAI21_X1  g446(.A(new_n871), .B1(new_n860), .B2(new_n863), .ZN(new_n872));
  INV_X1    g447(.A(new_n859), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n855), .A2(new_n856), .A3(new_n857), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n873), .A2(G651), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(new_n863), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n564), .A3(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n872), .A2(new_n877), .ZN(new_n878));
  XNOR2_X1  g453(.A(new_n870), .B(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT39), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n881), .A2(new_n865), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n879), .A2(new_n880), .ZN(new_n883));
  OAI21_X1  g458(.A(new_n867), .B1(new_n882), .B2(new_n883), .ZN(G145));
  XNOR2_X1  g459(.A(KEYINPUT106), .B(G37), .ZN(new_n885));
  INV_X1    g460(.A(new_n885), .ZN(new_n886));
  XNOR2_X1  g461(.A(G160), .B(new_n646), .ZN(new_n887));
  XOR2_X1   g462(.A(new_n887), .B(G162), .Z(new_n888));
  NAND3_X1  g463(.A1(new_n825), .A2(G164), .A3(new_n831), .ZN(new_n889));
  INV_X1    g464(.A(new_n889), .ZN(new_n890));
  AOI21_X1  g465(.A(G164), .B1(new_n825), .B2(new_n831), .ZN(new_n891));
  OAI21_X1  g466(.A(new_n778), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  INV_X1    g467(.A(new_n891), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n893), .A2(new_n777), .A3(new_n889), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n788), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n895), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g472(.A1(new_n749), .A2(new_n639), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n484), .A2(G142), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n487), .A2(G130), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n474), .A2(KEYINPUT104), .A3(G118), .ZN(new_n902));
  OAI21_X1  g477(.A(KEYINPUT104), .B1(new_n474), .B2(G118), .ZN(new_n903));
  OR2_X1    g478(.A1(G106), .A2(G2105), .ZN(new_n904));
  NAND4_X1  g479(.A1(new_n902), .A2(G2104), .A3(new_n903), .A4(new_n904), .ZN(new_n905));
  NAND3_X1  g480(.A1(new_n900), .A2(new_n901), .A3(new_n905), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n749), .A2(new_n639), .ZN(new_n908));
  AND3_X1   g483(.A1(new_n899), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  AOI21_X1  g484(.A(new_n907), .B1(new_n899), .B2(new_n908), .ZN(new_n910));
  NOR2_X1   g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n892), .A2(new_n894), .A3(new_n788), .ZN(new_n912));
  NAND3_X1  g487(.A1(new_n897), .A2(new_n911), .A3(new_n912), .ZN(new_n913));
  INV_X1    g488(.A(new_n913), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  AOI21_X1  g490(.A(new_n888), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n897), .A2(new_n912), .ZN(new_n917));
  OR2_X1    g492(.A1(new_n909), .A2(new_n910), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n919), .A2(KEYINPUT105), .A3(new_n913), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n886), .B1(new_n916), .B2(new_n920), .ZN(new_n921));
  NAND3_X1  g496(.A1(new_n919), .A2(new_n913), .A3(new_n888), .ZN(new_n922));
  AND2_X1   g497(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n923));
  NOR2_X1   g498(.A1(new_n922), .A2(KEYINPUT107), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n921), .B1(new_n923), .B2(new_n924), .ZN(new_n925));
  XNOR2_X1  g500(.A(new_n925), .B(KEYINPUT40), .ZN(G395));
  INV_X1    g501(.A(KEYINPUT109), .ZN(new_n927));
  XNOR2_X1  g502(.A(new_n630), .B(new_n878), .ZN(new_n928));
  INV_X1    g503(.A(new_n620), .ZN(new_n929));
  AOI21_X1  g504(.A(new_n619), .B1(new_n614), .B2(new_n616), .ZN(new_n930));
  OAI21_X1  g505(.A(new_n611), .B1(new_n929), .B2(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n625), .ZN(new_n932));
  OAI211_X1 g507(.A(G299), .B(new_n611), .C1(new_n929), .C2(new_n930), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n928), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g510(.A(KEYINPUT108), .B1(new_n621), .B2(G299), .ZN(new_n936));
  INV_X1    g511(.A(KEYINPUT108), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n931), .A2(new_n937), .A3(new_n625), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n936), .A2(new_n938), .A3(new_n933), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT41), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n940), .B1(new_n621), .B2(G299), .ZN(new_n941));
  AOI22_X1  g516(.A1(new_n939), .A2(new_n940), .B1(new_n932), .B2(new_n941), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n935), .B1(new_n942), .B2(new_n928), .ZN(new_n943));
  NAND2_X1  g518(.A1(new_n943), .A2(KEYINPUT42), .ZN(new_n944));
  INV_X1    g519(.A(KEYINPUT42), .ZN(new_n945));
  OAI211_X1 g520(.A(new_n935), .B(new_n945), .C1(new_n942), .C2(new_n928), .ZN(new_n946));
  NAND2_X1  g521(.A1(new_n944), .A2(new_n946), .ZN(new_n947));
  XOR2_X1   g522(.A(new_n605), .B(G305), .Z(new_n948));
  XNOR2_X1  g523(.A(G166), .B(G288), .ZN(new_n949));
  XOR2_X1   g524(.A(new_n948), .B(new_n949), .Z(new_n950));
  NAND2_X1  g525(.A1(new_n947), .A2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(new_n950), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n944), .A2(new_n952), .A3(new_n946), .ZN(new_n953));
  AND4_X1   g528(.A1(new_n927), .A2(new_n951), .A3(G868), .A4(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(KEYINPUT109), .B1(new_n864), .B2(G868), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n632), .B1(new_n947), .B2(new_n950), .ZN(new_n956));
  AOI21_X1  g531(.A(new_n955), .B1(new_n956), .B2(new_n953), .ZN(new_n957));
  NOR2_X1   g532(.A1(new_n954), .A2(new_n957), .ZN(G295));
  NOR2_X1   g533(.A1(new_n954), .A2(new_n957), .ZN(G331));
  AOI21_X1  g534(.A(G286), .B1(G171), .B2(KEYINPUT110), .ZN(new_n960));
  INV_X1    g535(.A(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(KEYINPUT110), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n962), .B1(new_n553), .B2(new_n556), .ZN(new_n963));
  NAND3_X1  g538(.A1(new_n872), .A2(new_n877), .A3(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  AOI21_X1  g540(.A(new_n963), .B1(new_n872), .B2(new_n877), .ZN(new_n966));
  OAI21_X1  g541(.A(new_n961), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g542(.A(new_n963), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n878), .A2(new_n968), .ZN(new_n969));
  NAND3_X1  g544(.A1(new_n969), .A2(new_n964), .A3(new_n960), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n967), .A2(new_n970), .A3(new_n934), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n967), .A2(new_n970), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n934), .A2(new_n940), .ZN(new_n973));
  NAND3_X1  g548(.A1(new_n936), .A2(new_n941), .A3(new_n938), .ZN(new_n974));
  NAND2_X1  g549(.A1(new_n973), .A2(new_n974), .ZN(new_n975));
  AOI22_X1  g550(.A1(new_n971), .A2(KEYINPUT111), .B1(new_n972), .B2(new_n975), .ZN(new_n976));
  OR2_X1    g551(.A1(new_n971), .A2(KEYINPUT111), .ZN(new_n977));
  AOI21_X1  g552(.A(new_n950), .B1(new_n976), .B2(new_n977), .ZN(new_n978));
  AND2_X1   g553(.A1(new_n967), .A2(new_n970), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n950), .B(new_n971), .C1(new_n979), .C2(new_n942), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n980), .A2(new_n885), .ZN(new_n981));
  INV_X1    g556(.A(KEYINPUT43), .ZN(new_n982));
  NOR3_X1   g557(.A1(new_n978), .A2(new_n981), .A3(new_n982), .ZN(new_n983));
  OAI21_X1  g558(.A(new_n971), .B1(new_n979), .B2(new_n942), .ZN(new_n984));
  AOI21_X1  g559(.A(G37), .B1(new_n984), .B2(new_n952), .ZN(new_n985));
  AOI21_X1  g560(.A(KEYINPUT43), .B1(new_n985), .B2(new_n980), .ZN(new_n986));
  OAI21_X1  g561(.A(KEYINPUT44), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  INV_X1    g562(.A(KEYINPUT44), .ZN(new_n988));
  NOR3_X1   g563(.A1(new_n978), .A2(new_n981), .A3(KEYINPUT43), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n982), .B1(new_n985), .B2(new_n980), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n988), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g566(.A1(new_n987), .A2(new_n991), .ZN(G397));
  OAI21_X1  g567(.A(G125), .B1(new_n467), .B2(new_n468), .ZN(new_n993));
  INV_X1    g568(.A(KEYINPUT68), .ZN(new_n994));
  AOI22_X1  g569(.A1(new_n993), .A2(new_n994), .B1(G113), .B2(G2104), .ZN(new_n995));
  AOI21_X1  g570(.A(new_n474), .B1(new_n995), .B2(new_n469), .ZN(new_n996));
  XNOR2_X1  g571(.A(new_n475), .B(KEYINPUT69), .ZN(new_n997));
  INV_X1    g572(.A(G137), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n504), .A2(new_n474), .ZN(new_n999));
  OAI21_X1  g574(.A(new_n997), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(G40), .ZN(new_n1001));
  NOR3_X1   g576(.A1(new_n996), .A2(new_n1000), .A3(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT45), .ZN(new_n1003));
  INV_X1    g578(.A(G1384), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1004), .B1(new_n506), .B2(new_n511), .ZN(new_n1005));
  NAND3_X1  g580(.A1(new_n1002), .A2(new_n1003), .A3(new_n1005), .ZN(new_n1006));
  OR2_X1    g581(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1006), .A2(KEYINPUT112), .ZN(new_n1008));
  AND2_X1   g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  XNOR2_X1  g584(.A(new_n832), .B(new_n834), .ZN(new_n1010));
  INV_X1    g585(.A(G1996), .ZN(new_n1011));
  XNOR2_X1  g586(.A(new_n777), .B(new_n1011), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n750), .A2(new_n752), .ZN(new_n1013));
  OR2_X1    g588(.A1(new_n750), .A2(new_n752), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .A4(new_n1014), .ZN(new_n1015));
  XNOR2_X1  g590(.A(new_n605), .B(new_n740), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1009), .B1(new_n1015), .B2(new_n1016), .ZN(new_n1017));
  XOR2_X1   g592(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1018));
  INV_X1    g593(.A(G8), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n1005), .A2(new_n1003), .ZN(new_n1020));
  OAI211_X1 g595(.A(KEYINPUT45), .B(new_n1004), .C1(new_n506), .C2(new_n511), .ZN(new_n1021));
  NAND3_X1  g596(.A1(new_n1020), .A2(new_n1002), .A3(new_n1021), .ZN(new_n1022));
  INV_X1    g597(.A(G1966), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1005), .A2(KEYINPUT50), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT50), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1026), .B(new_n1004), .C1(new_n506), .C2(new_n511), .ZN(new_n1027));
  NAND4_X1  g602(.A1(new_n1025), .A2(new_n849), .A3(new_n1002), .A4(new_n1027), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1019), .B1(new_n1024), .B2(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT121), .ZN(new_n1030));
  AOI21_X1  g605(.A(new_n1030), .B1(G286), .B2(G8), .ZN(new_n1031));
  INV_X1    g606(.A(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(G286), .A2(new_n1030), .A3(G8), .ZN(new_n1033));
  NAND2_X1  g608(.A1(new_n1032), .A2(new_n1033), .ZN(new_n1034));
  OAI21_X1  g609(.A(new_n1018), .B1(new_n1029), .B2(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(KEYINPUT51), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1032), .A2(new_n1036), .A3(new_n1033), .ZN(new_n1037));
  OAI21_X1  g612(.A(KEYINPUT123), .B1(new_n1029), .B2(new_n1037), .ZN(new_n1038));
  INV_X1    g613(.A(KEYINPUT123), .ZN(new_n1039));
  INV_X1    g614(.A(new_n1037), .ZN(new_n1040));
  AND3_X1   g615(.A1(new_n1025), .A2(new_n1002), .A3(new_n1027), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1041), .A2(new_n849), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1042));
  OAI211_X1 g617(.A(new_n1039), .B(new_n1040), .C1(new_n1042), .C2(new_n1019), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1035), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  INV_X1    g619(.A(new_n1042), .ZN(new_n1045));
  NAND2_X1  g620(.A1(new_n1045), .A2(new_n1034), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g622(.A1(new_n1047), .A2(KEYINPUT62), .ZN(new_n1048));
  INV_X1    g623(.A(G1971), .ZN(new_n1049));
  NAND2_X1  g624(.A1(new_n1022), .A2(new_n1049), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1025), .A2(new_n1002), .A3(new_n1027), .ZN(new_n1051));
  OAI21_X1  g626(.A(new_n1050), .B1(G2090), .B2(new_n1051), .ZN(new_n1052));
  INV_X1    g627(.A(KEYINPUT55), .ZN(new_n1053));
  OAI21_X1  g628(.A(new_n1053), .B1(G166), .B2(new_n1019), .ZN(new_n1054));
  NAND3_X1  g629(.A1(G303), .A2(KEYINPUT55), .A3(G8), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  AND3_X1   g631(.A1(new_n1052), .A2(G8), .A3(new_n1056), .ZN(new_n1057));
  AOI21_X1  g632(.A(new_n1056), .B1(new_n1052), .B2(G8), .ZN(new_n1058));
  NOR2_X1   g633(.A1(new_n1057), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G1981), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n596), .A2(new_n597), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n594), .B1(new_n1061), .B2(KEYINPUT114), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT114), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n596), .A2(new_n1063), .A3(new_n597), .ZN(new_n1064));
  AOI21_X1  g639(.A(new_n1060), .B1(new_n1062), .B2(new_n1064), .ZN(new_n1065));
  NOR2_X1   g640(.A1(G305), .A2(G1981), .ZN(new_n1066));
  OAI21_X1  g641(.A(KEYINPUT115), .B1(new_n1065), .B2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT115), .ZN(new_n1068));
  INV_X1    g643(.A(new_n1061), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n1069), .A2(new_n1060), .A3(new_n592), .A4(new_n595), .ZN(new_n1070));
  AND3_X1   g645(.A1(new_n596), .A2(new_n1063), .A3(new_n597), .ZN(new_n1071));
  AOI21_X1  g646(.A(new_n1063), .B1(new_n596), .B2(new_n597), .ZN(new_n1072));
  NOR3_X1   g647(.A1(new_n1071), .A2(new_n1072), .A3(new_n594), .ZN(new_n1073));
  OAI211_X1 g648(.A(new_n1068), .B(new_n1070), .C1(new_n1073), .C2(new_n1060), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT116), .ZN(new_n1075));
  INV_X1    g650(.A(KEYINPUT49), .ZN(new_n1076));
  NAND4_X1  g651(.A1(new_n1067), .A2(new_n1074), .A3(new_n1075), .A4(new_n1076), .ZN(new_n1077));
  NAND3_X1  g652(.A1(new_n471), .A2(G40), .A3(new_n478), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1078), .A2(new_n1005), .ZN(new_n1079));
  NOR2_X1   g654(.A1(new_n1079), .A2(new_n1019), .ZN(new_n1080));
  AND3_X1   g655(.A1(new_n1067), .A2(new_n1076), .A3(new_n1074), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1065), .A2(new_n1066), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT116), .B1(new_n1082), .B2(KEYINPUT49), .ZN(new_n1083));
  OAI211_X1 g658(.A(new_n1077), .B(new_n1080), .C1(new_n1081), .C2(new_n1083), .ZN(new_n1084));
  INV_X1    g659(.A(G1976), .ZN(new_n1085));
  OAI21_X1  g660(.A(new_n1080), .B1(new_n1085), .B2(G288), .ZN(new_n1086));
  AND2_X1   g661(.A1(new_n1086), .A2(KEYINPUT52), .ZN(new_n1087));
  INV_X1    g662(.A(new_n1086), .ZN(new_n1088));
  XOR2_X1   g663(.A(KEYINPUT113), .B(G1976), .Z(new_n1089));
  AOI21_X1  g664(.A(KEYINPUT52), .B1(G288), .B2(new_n1089), .ZN(new_n1090));
  AOI21_X1  g665(.A(new_n1087), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1091));
  AND3_X1   g666(.A1(new_n1059), .A2(new_n1084), .A3(new_n1091), .ZN(new_n1092));
  INV_X1    g667(.A(KEYINPUT62), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n1044), .A2(new_n1093), .A3(new_n1046), .ZN(new_n1094));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n1095));
  NAND4_X1  g670(.A1(new_n1020), .A2(new_n800), .A3(new_n1002), .A4(new_n1021), .ZN(new_n1096));
  XNOR2_X1  g671(.A(KEYINPUT125), .B(G1961), .ZN(new_n1097));
  AOI22_X1  g672(.A1(new_n1095), .A2(new_n1096), .B1(new_n1051), .B2(new_n1097), .ZN(new_n1098));
  OR2_X1    g673(.A1(new_n1096), .A2(new_n1095), .ZN(new_n1099));
  AOI21_X1  g674(.A(G301), .B1(new_n1098), .B2(new_n1099), .ZN(new_n1100));
  NAND4_X1  g675(.A1(new_n1048), .A2(new_n1092), .A3(new_n1094), .A4(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT127), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  NOR3_X1   g678(.A1(new_n1042), .A2(new_n1019), .A3(G286), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1059), .A2(new_n1084), .A3(new_n1091), .A4(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1105), .B(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1103), .A2(new_n1107), .ZN(new_n1108));
  INV_X1    g683(.A(new_n1100), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1109), .B1(new_n1047), .B2(KEYINPUT62), .ZN(new_n1110));
  NAND4_X1  g685(.A1(new_n1110), .A2(KEYINPUT127), .A3(new_n1092), .A4(new_n1094), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  XNOR2_X1  g687(.A(new_n1112), .B(KEYINPUT117), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1020), .A2(new_n1002), .A3(new_n1021), .A4(new_n1113), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1115), .A2(KEYINPUT118), .B1(new_n814), .B2(new_n1051), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT57), .ZN(new_n1117));
  AND3_X1   g692(.A1(new_n571), .A2(new_n1117), .A3(new_n578), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1117), .B1(new_n571), .B2(new_n578), .ZN(new_n1119));
  NOR2_X1   g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT118), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1114), .A2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1116), .A2(KEYINPUT119), .A3(new_n1120), .A4(new_n1122), .ZN(new_n1123));
  AOI21_X1  g698(.A(new_n1078), .B1(new_n1003), .B2(new_n1005), .ZN(new_n1124));
  NAND4_X1  g699(.A1(new_n1124), .A2(KEYINPUT118), .A3(new_n1021), .A4(new_n1113), .ZN(new_n1125));
  NAND2_X1  g700(.A1(new_n1051), .A2(new_n814), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1125), .A2(new_n1122), .A3(new_n1120), .A4(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT119), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1123), .A2(new_n1129), .ZN(new_n1130));
  INV_X1    g705(.A(G1348), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1051), .A2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1079), .A2(new_n834), .ZN(new_n1133));
  AOI21_X1  g708(.A(new_n931), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  NAND3_X1  g709(.A1(new_n1125), .A2(new_n1122), .A3(new_n1126), .ZN(new_n1135));
  INV_X1    g710(.A(new_n1120), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  INV_X1    g712(.A(new_n1137), .ZN(new_n1138));
  OAI21_X1  g713(.A(new_n1130), .B1(new_n1134), .B2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(KEYINPUT61), .B1(new_n1130), .B2(new_n1137), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT60), .ZN(new_n1141));
  AND4_X1   g716(.A1(new_n1141), .A2(new_n621), .A3(new_n1132), .A4(new_n1133), .ZN(new_n1142));
  XOR2_X1   g717(.A(KEYINPUT58), .B(G1341), .Z(new_n1143));
  OAI21_X1  g718(.A(new_n1143), .B1(new_n1078), .B2(new_n1005), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1144), .B1(new_n1022), .B2(G1996), .ZN(new_n1145));
  NOR2_X1   g720(.A1(new_n871), .A2(KEYINPUT120), .ZN(new_n1146));
  NAND2_X1  g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1147), .A2(KEYINPUT59), .ZN(new_n1148));
  INV_X1    g723(.A(KEYINPUT59), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1145), .A2(new_n1149), .A3(new_n1146), .ZN(new_n1150));
  AOI21_X1  g725(.A(new_n1142), .B1(new_n1148), .B2(new_n1150), .ZN(new_n1151));
  NAND3_X1  g726(.A1(new_n1137), .A2(KEYINPUT61), .A3(new_n1127), .ZN(new_n1152));
  AND3_X1   g727(.A1(new_n931), .A2(new_n1132), .A3(new_n1133), .ZN(new_n1153));
  OAI21_X1  g728(.A(KEYINPUT60), .B1(new_n1153), .B2(new_n1134), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1151), .A2(new_n1152), .A3(new_n1154), .ZN(new_n1155));
  OAI21_X1  g730(.A(new_n1139), .B1(new_n1140), .B2(new_n1155), .ZN(new_n1156));
  XNOR2_X1  g731(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1096), .A2(new_n1095), .ZN(new_n1158));
  NAND2_X1  g733(.A1(new_n1051), .A2(new_n1097), .ZN(new_n1159));
  OR2_X1    g734(.A1(KEYINPUT126), .A2(G2078), .ZN(new_n1160));
  NAND2_X1  g735(.A1(KEYINPUT126), .A2(G2078), .ZN(new_n1161));
  AOI21_X1  g736(.A(new_n1095), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1124), .A2(new_n1021), .A3(new_n1162), .ZN(new_n1163));
  AND4_X1   g738(.A1(G301), .A2(new_n1158), .A3(new_n1159), .A4(new_n1163), .ZN(new_n1164));
  OAI21_X1  g739(.A(new_n1157), .B1(new_n1100), .B2(new_n1164), .ZN(new_n1165));
  NAND3_X1  g740(.A1(new_n1158), .A2(new_n1163), .A3(new_n1159), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1166), .A2(G171), .ZN(new_n1167));
  NAND3_X1  g742(.A1(new_n1098), .A2(new_n1099), .A3(G301), .ZN(new_n1168));
  NAND3_X1  g743(.A1(new_n1167), .A2(new_n1168), .A3(KEYINPUT54), .ZN(new_n1169));
  NAND2_X1  g744(.A1(new_n1165), .A2(new_n1169), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1170), .B1(new_n1046), .B2(new_n1044), .ZN(new_n1171));
  NAND3_X1  g746(.A1(new_n1156), .A2(new_n1171), .A3(new_n1092), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1084), .A2(new_n1085), .A3(new_n723), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1173), .A2(new_n1070), .ZN(new_n1174));
  AND2_X1   g749(.A1(new_n1084), .A2(new_n1091), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1174), .A2(new_n1080), .B1(new_n1175), .B2(new_n1057), .ZN(new_n1176));
  NAND3_X1  g751(.A1(new_n1111), .A2(new_n1172), .A3(new_n1176), .ZN(new_n1177));
  OAI21_X1  g752(.A(new_n1017), .B1(new_n1108), .B2(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1179));
  OAI22_X1  g754(.A1(new_n1179), .A2(new_n1013), .B1(G2067), .B2(new_n832), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(new_n1009), .ZN(new_n1181));
  NAND2_X1  g756(.A1(new_n1015), .A2(new_n1009), .ZN(new_n1182));
  INV_X1    g757(.A(KEYINPUT48), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1009), .A2(new_n740), .A3(new_n605), .ZN(new_n1184));
  OAI21_X1  g759(.A(new_n1182), .B1(new_n1183), .B2(new_n1184), .ZN(new_n1185));
  INV_X1    g760(.A(new_n1184), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n1186), .A2(KEYINPUT48), .ZN(new_n1187));
  OAI21_X1  g762(.A(new_n1181), .B1(new_n1185), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1189));
  XNOR2_X1  g764(.A(new_n1189), .B(KEYINPUT46), .ZN(new_n1190));
  INV_X1    g765(.A(new_n1010), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1009), .B1(new_n1191), .B2(new_n777), .ZN(new_n1192));
  NAND2_X1  g767(.A1(new_n1190), .A2(new_n1192), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1193), .A2(KEYINPUT47), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(KEYINPUT47), .ZN(new_n1195));
  AOI21_X1  g770(.A(new_n1188), .B1(new_n1194), .B2(new_n1195), .ZN(new_n1196));
  NAND2_X1  g771(.A1(new_n1178), .A2(new_n1196), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g772(.A1(G227), .A2(new_n459), .ZN(new_n1199));
  OAI21_X1  g773(.A(new_n1199), .B1(new_n713), .B2(new_n714), .ZN(new_n1200));
  AOI21_X1  g774(.A(new_n1200), .B1(new_n677), .B2(new_n678), .ZN(new_n1201));
  OAI211_X1 g775(.A(new_n925), .B(new_n1201), .C1(new_n989), .C2(new_n990), .ZN(G225));
  INV_X1    g776(.A(G225), .ZN(G308));
endmodule


