//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 0 1 1 1 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 0 1 1 1 0 0 0 1 0 0 1 1 0 0 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:09 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n719, new_n720,
    new_n721, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n737, new_n738, new_n739, new_n740, new_n741, new_n742, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n946, new_n947,
    new_n948, new_n950, new_n951, new_n952, new_n953, new_n954, new_n955,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n980, new_n981, new_n982, new_n983, new_n984, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1026, new_n1027, new_n1028, new_n1029, new_n1030;
  OR2_X1    g000(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n187));
  INV_X1    g001(.A(G107), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G104), .ZN(new_n189));
  AND2_X1   g003(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n187), .B1(new_n189), .B2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G101), .ZN(new_n192));
  NOR2_X1   g006(.A1(new_n188), .A2(G104), .ZN(new_n193));
  INV_X1    g007(.A(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT80), .A2(KEYINPUT3), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  NAND4_X1  g012(.A1(new_n191), .A2(new_n192), .A3(new_n194), .A4(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G146), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G143), .ZN(new_n201));
  INV_X1    g015(.A(G143), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G146), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  OAI211_X1 g018(.A(new_n201), .B(new_n203), .C1(KEYINPUT1), .C2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT81), .ZN(new_n206));
  OAI21_X1  g020(.A(new_n206), .B1(new_n188), .B2(G104), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n195), .A2(KEYINPUT81), .A3(G107), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n207), .A2(new_n189), .A3(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G101), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n201), .A2(new_n203), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n201), .A2(KEYINPUT1), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n211), .A2(new_n212), .A3(G128), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n199), .A2(new_n205), .A3(new_n210), .A4(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT10), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n216), .A2(KEYINPUT82), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT82), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n218), .A3(new_n215), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n217), .A2(new_n219), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT11), .ZN(new_n221));
  INV_X1    g035(.A(G134), .ZN(new_n222));
  OAI21_X1  g036(.A(new_n221), .B1(new_n222), .B2(G137), .ZN(new_n223));
  INV_X1    g037(.A(G137), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n224), .A2(KEYINPUT11), .A3(G134), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n222), .A2(G137), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n223), .A2(new_n225), .A3(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(G131), .ZN(new_n228));
  INV_X1    g042(.A(G131), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n223), .A2(new_n225), .A3(new_n229), .A4(new_n226), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n228), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n193), .B1(new_n197), .B2(new_n196), .ZN(new_n233));
  AOI21_X1  g047(.A(new_n192), .B1(new_n233), .B2(new_n191), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  NOR2_X1   g050(.A1(KEYINPUT0), .A2(G128), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT64), .ZN(new_n238));
  AOI22_X1  g052(.A1(new_n201), .A2(new_n203), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  OAI21_X1  g053(.A(KEYINPUT64), .B1(KEYINPUT0), .B2(G128), .ZN(new_n240));
  NAND2_X1  g054(.A1(KEYINPUT0), .A2(G128), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  XNOR2_X1  g056(.A(G143), .B(G146), .ZN(new_n243));
  INV_X1    g057(.A(new_n241), .ZN(new_n244));
  AOI22_X1  g058(.A1(new_n239), .A2(new_n242), .B1(new_n243), .B2(new_n244), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n199), .A2(KEYINPUT4), .ZN(new_n246));
  OAI211_X1 g060(.A(new_n236), .B(new_n245), .C1(new_n234), .C2(new_n246), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n199), .A2(new_n210), .ZN(new_n248));
  NAND2_X1  g062(.A1(new_n213), .A2(new_n205), .ZN(new_n249));
  INV_X1    g063(.A(new_n249), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n248), .A2(KEYINPUT83), .A3(KEYINPUT10), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT83), .ZN(new_n252));
  OAI21_X1  g066(.A(new_n252), .B1(new_n214), .B2(new_n215), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n251), .A2(new_n253), .ZN(new_n254));
  NAND4_X1  g068(.A1(new_n220), .A2(new_n232), .A3(new_n247), .A4(new_n254), .ZN(new_n255));
  INV_X1    g069(.A(G953), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n256), .A2(G227), .ZN(new_n257));
  XNOR2_X1  g071(.A(new_n257), .B(KEYINPUT79), .ZN(new_n258));
  XNOR2_X1  g072(.A(G110), .B(G140), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n258), .B(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n220), .A2(new_n254), .A3(new_n247), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(new_n231), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n263), .A2(KEYINPUT84), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT84), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n262), .A2(new_n265), .A3(new_n231), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n261), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n248), .A2(new_n250), .ZN(new_n268));
  INV_X1    g082(.A(new_n214), .ZN(new_n269));
  OAI21_X1  g083(.A(new_n231), .B1(new_n268), .B2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  XNOR2_X1  g085(.A(new_n270), .B(new_n271), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n260), .B1(new_n272), .B2(new_n255), .ZN(new_n273));
  OAI21_X1  g087(.A(KEYINPUT85), .B1(new_n267), .B2(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(new_n261), .ZN(new_n275));
  AND3_X1   g089(.A1(new_n262), .A2(new_n265), .A3(new_n231), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n265), .B1(new_n262), .B2(new_n231), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n275), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n272), .A2(new_n255), .ZN(new_n279));
  INV_X1    g093(.A(new_n260), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  INV_X1    g095(.A(KEYINPUT85), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n278), .A2(new_n281), .A3(new_n282), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n274), .A2(G469), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(G469), .ZN(new_n285));
  INV_X1    g099(.A(G902), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n264), .A2(new_n266), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n260), .B1(new_n287), .B2(new_n255), .ZN(new_n288));
  AND3_X1   g102(.A1(new_n272), .A2(new_n260), .A3(new_n255), .ZN(new_n289));
  OAI211_X1 g103(.A(new_n285), .B(new_n286), .C1(new_n288), .C2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(G469), .A2(G902), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n284), .A2(new_n290), .A3(new_n291), .ZN(new_n292));
  OAI21_X1  g106(.A(G214), .B1(G237), .B2(G902), .ZN(new_n293));
  INV_X1    g107(.A(new_n293), .ZN(new_n294));
  OAI21_X1  g108(.A(G210), .B1(G237), .B2(G902), .ZN(new_n295));
  INV_X1    g109(.A(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(G119), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n297), .A2(KEYINPUT66), .A3(G116), .ZN(new_n298));
  INV_X1    g112(.A(G116), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n299), .A2(G119), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  XOR2_X1   g115(.A(KEYINPUT2), .B(G113), .Z(new_n302));
  INV_X1    g116(.A(KEYINPUT67), .ZN(new_n303));
  INV_X1    g117(.A(KEYINPUT66), .ZN(new_n304));
  OAI21_X1  g118(.A(new_n304), .B1(new_n299), .B2(G119), .ZN(new_n305));
  NAND4_X1  g119(.A1(new_n301), .A2(new_n302), .A3(new_n303), .A4(new_n305), .ZN(new_n306));
  NAND3_X1  g120(.A1(new_n305), .A2(new_n298), .A3(new_n300), .ZN(new_n307));
  XNOR2_X1  g121(.A(KEYINPUT2), .B(G113), .ZN(new_n308));
  OAI21_X1  g122(.A(KEYINPUT67), .B1(new_n307), .B2(new_n308), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n306), .A2(new_n309), .ZN(new_n310));
  INV_X1    g124(.A(KEYINPUT5), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n311), .A2(new_n297), .A3(G116), .ZN(new_n312));
  OAI211_X1 g126(.A(G113), .B(new_n312), .C1(new_n307), .C2(new_n311), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n248), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n236), .B1(new_n246), .B2(new_n234), .ZN(new_n315));
  AOI22_X1  g129(.A1(new_n306), .A2(new_n309), .B1(new_n308), .B2(new_n307), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n314), .B1(new_n315), .B2(new_n316), .ZN(new_n317));
  XNOR2_X1  g131(.A(G110), .B(G122), .ZN(new_n318));
  INV_X1    g132(.A(new_n318), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n317), .A2(new_n319), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n314), .B(new_n318), .C1(new_n315), .C2(new_n316), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n320), .A2(KEYINPUT6), .A3(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G125), .ZN(new_n323));
  NOR2_X1   g137(.A1(new_n245), .A2(new_n323), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n324), .B1(new_n323), .B2(new_n249), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n256), .A2(G224), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n325), .B(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT6), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n317), .A2(new_n328), .A3(new_n319), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n322), .A2(new_n327), .A3(new_n329), .ZN(new_n330));
  INV_X1    g144(.A(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n326), .A2(KEYINPUT7), .ZN(new_n332));
  INV_X1    g146(.A(new_n324), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n249), .A2(new_n323), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n333), .B1(KEYINPUT86), .B2(new_n334), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n334), .A2(KEYINPUT86), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n332), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT87), .ZN(new_n338));
  INV_X1    g152(.A(new_n332), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n325), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n333), .A2(new_n334), .A3(new_n339), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT87), .ZN(new_n342));
  NAND4_X1  g156(.A1(new_n337), .A2(new_n340), .A3(new_n321), .A4(new_n342), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n310), .A2(new_n313), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n199), .A2(new_n210), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(new_n314), .ZN(new_n347));
  XNOR2_X1  g161(.A(new_n318), .B(KEYINPUT8), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n286), .B1(new_n343), .B2(new_n350), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n296), .B1(new_n331), .B2(new_n351), .ZN(new_n352));
  AND2_X1   g166(.A1(new_n340), .A2(new_n342), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n353), .A2(new_n349), .A3(new_n321), .A4(new_n337), .ZN(new_n354));
  NAND4_X1  g168(.A1(new_n330), .A2(new_n354), .A3(new_n286), .A4(new_n295), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n294), .B1(new_n352), .B2(new_n355), .ZN(new_n356));
  XNOR2_X1  g170(.A(KEYINPUT9), .B(G234), .ZN(new_n357));
  OAI21_X1  g171(.A(G221), .B1(new_n357), .B2(G902), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n292), .A2(new_n356), .A3(new_n358), .ZN(new_n359));
  NOR2_X1   g173(.A1(G472), .A2(G902), .ZN(new_n360));
  INV_X1    g174(.A(KEYINPUT68), .ZN(new_n361));
  NOR2_X1   g175(.A1(new_n222), .A2(G137), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n224), .A2(G134), .ZN(new_n363));
  OAI21_X1  g177(.A(G131), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  NAND4_X1  g178(.A1(new_n213), .A2(new_n205), .A3(new_n230), .A4(new_n364), .ZN(new_n365));
  AND3_X1   g179(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n366));
  AOI21_X1  g180(.A(KEYINPUT65), .B1(new_n231), .B2(new_n245), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n365), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n307), .A2(new_n308), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n310), .A2(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n368), .A2(new_n370), .ZN(new_n371));
  AND2_X1   g185(.A1(new_n230), .A2(new_n364), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n250), .A2(new_n372), .B1(new_n231), .B2(new_n245), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n373), .A2(KEYINPUT28), .A3(new_n316), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n231), .A2(new_n245), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n316), .A2(new_n365), .A3(new_n375), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT28), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n376), .A2(new_n377), .ZN(new_n378));
  NAND3_X1  g192(.A1(new_n371), .A2(new_n374), .A3(new_n378), .ZN(new_n379));
  NOR2_X1   g193(.A1(G237), .A2(G953), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n380), .A2(G210), .ZN(new_n381));
  XNOR2_X1  g195(.A(new_n381), .B(KEYINPUT27), .ZN(new_n382));
  XOR2_X1   g196(.A(KEYINPUT26), .B(G101), .Z(new_n383));
  XNOR2_X1  g197(.A(new_n382), .B(new_n383), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT31), .ZN(new_n385));
  NAND3_X1  g199(.A1(new_n375), .A2(KEYINPUT30), .A3(new_n365), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n370), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT30), .ZN(new_n388));
  AOI21_X1  g202(.A(new_n387), .B1(new_n388), .B2(new_n368), .ZN(new_n389));
  INV_X1    g203(.A(new_n384), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n390), .A2(new_n376), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n385), .B1(new_n389), .B2(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n316), .B1(new_n373), .B2(KEYINPUT30), .ZN(new_n393));
  INV_X1    g207(.A(new_n365), .ZN(new_n394));
  INV_X1    g208(.A(KEYINPUT65), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n375), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n231), .A2(KEYINPUT65), .A3(new_n245), .ZN(new_n397));
  AOI21_X1  g211(.A(new_n394), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n393), .B1(new_n398), .B2(KEYINPUT30), .ZN(new_n399));
  INV_X1    g213(.A(new_n391), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n399), .A2(KEYINPUT31), .A3(new_n400), .ZN(new_n401));
  AOI221_X4 g215(.A(new_n361), .B1(new_n379), .B2(new_n384), .C1(new_n392), .C2(new_n401), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n392), .A2(new_n401), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n379), .A2(new_n384), .ZN(new_n404));
  AOI21_X1  g218(.A(KEYINPUT68), .B1(new_n403), .B2(new_n404), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n360), .B1(new_n402), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT69), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT32), .ZN(new_n409));
  NOR3_X1   g223(.A1(new_n389), .A2(new_n385), .A3(new_n391), .ZN(new_n410));
  AOI21_X1  g224(.A(KEYINPUT31), .B1(new_n399), .B2(new_n400), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n404), .B1(new_n410), .B2(new_n411), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n361), .ZN(new_n413));
  NAND3_X1  g227(.A1(new_n403), .A2(KEYINPUT68), .A3(new_n404), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n415), .A2(KEYINPUT69), .A3(new_n360), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n408), .A2(new_n409), .A3(new_n416), .ZN(new_n417));
  NAND4_X1  g231(.A1(new_n371), .A2(new_n390), .A3(new_n374), .A4(new_n378), .ZN(new_n418));
  INV_X1    g232(.A(KEYINPUT29), .ZN(new_n419));
  AND2_X1   g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n376), .ZN(new_n421));
  NAND2_X1  g235(.A1(new_n368), .A2(new_n388), .ZN(new_n422));
  AOI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(new_n393), .ZN(new_n423));
  OAI21_X1  g237(.A(KEYINPUT70), .B1(new_n423), .B2(new_n390), .ZN(new_n424));
  INV_X1    g238(.A(KEYINPUT70), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n425), .B(new_n384), .C1(new_n389), .C2(new_n421), .ZN(new_n426));
  AND3_X1   g240(.A1(new_n420), .A2(new_n424), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n378), .A2(KEYINPUT29), .A3(new_n390), .ZN(new_n428));
  INV_X1    g242(.A(KEYINPUT71), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n376), .A2(new_n429), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n375), .A2(new_n365), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n370), .ZN(new_n432));
  NAND4_X1  g246(.A1(new_n316), .A2(KEYINPUT71), .A3(new_n375), .A4(new_n365), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n430), .A2(new_n432), .A3(new_n433), .ZN(new_n434));
  AOI21_X1  g248(.A(new_n428), .B1(KEYINPUT28), .B2(new_n434), .ZN(new_n435));
  OAI21_X1  g249(.A(KEYINPUT72), .B1(new_n435), .B2(G902), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n432), .A2(new_n433), .ZN(new_n437));
  AOI21_X1  g251(.A(KEYINPUT71), .B1(new_n373), .B2(new_n316), .ZN(new_n438));
  OAI21_X1  g252(.A(KEYINPUT28), .B1(new_n437), .B2(new_n438), .ZN(new_n439));
  AOI211_X1 g253(.A(new_n419), .B(new_n384), .C1(new_n376), .C2(new_n377), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n439), .A2(new_n440), .ZN(new_n441));
  INV_X1    g255(.A(KEYINPUT72), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n441), .A2(new_n442), .A3(new_n286), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n436), .A2(new_n443), .ZN(new_n444));
  OAI21_X1  g258(.A(G472), .B1(new_n427), .B2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT73), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g261(.A1(new_n420), .A2(new_n424), .A3(new_n426), .ZN(new_n448));
  NAND3_X1  g262(.A1(new_n448), .A2(new_n436), .A3(new_n443), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(KEYINPUT73), .A3(G472), .ZN(new_n450));
  NAND2_X1  g264(.A1(new_n447), .A2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n360), .ZN(new_n452));
  NOR2_X1   g266(.A1(new_n452), .A2(new_n409), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n453), .B1(new_n402), .B2(new_n405), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT74), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n415), .A2(KEYINPUT74), .A3(new_n453), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n417), .A2(new_n451), .A3(new_n456), .A4(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(G217), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n459), .B1(G234), .B2(new_n286), .ZN(new_n460));
  XNOR2_X1  g274(.A(G125), .B(G140), .ZN(new_n461));
  NAND2_X1  g275(.A1(new_n461), .A2(KEYINPUT16), .ZN(new_n462));
  INV_X1    g276(.A(G140), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n463), .A2(G125), .ZN(new_n464));
  OR2_X1    g278(.A1(new_n464), .A2(KEYINPUT16), .ZN(new_n465));
  NAND3_X1  g279(.A1(new_n462), .A2(G146), .A3(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n466), .A2(KEYINPUT77), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n468));
  NAND4_X1  g282(.A1(new_n462), .A2(new_n468), .A3(new_n465), .A4(G146), .ZN(new_n469));
  AND2_X1   g283(.A1(new_n462), .A2(new_n465), .ZN(new_n470));
  OAI211_X1 g284(.A(new_n467), .B(new_n469), .C1(G146), .C2(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(KEYINPUT24), .B(G110), .ZN(new_n472));
  XNOR2_X1  g286(.A(new_n472), .B(KEYINPUT75), .ZN(new_n473));
  XNOR2_X1  g287(.A(G119), .B(G128), .ZN(new_n474));
  OAI21_X1  g288(.A(KEYINPUT23), .B1(new_n204), .B2(G119), .ZN(new_n475));
  AOI21_X1  g289(.A(KEYINPUT76), .B1(new_n204), .B2(G119), .ZN(new_n476));
  XNOR2_X1  g290(.A(new_n475), .B(new_n476), .ZN(new_n477));
  AOI22_X1  g291(.A1(new_n473), .A2(new_n474), .B1(new_n477), .B2(G110), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n471), .A2(new_n478), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n461), .A2(new_n200), .ZN(new_n480));
  NOR2_X1   g294(.A1(new_n473), .A2(new_n474), .ZN(new_n481));
  NOR2_X1   g295(.A1(new_n477), .A2(G110), .ZN(new_n482));
  OAI211_X1 g296(.A(new_n466), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g297(.A(KEYINPUT22), .B(G137), .ZN(new_n484));
  AND3_X1   g298(.A1(new_n256), .A2(G221), .A3(G234), .ZN(new_n485));
  XOR2_X1   g299(.A(new_n484), .B(new_n485), .Z(new_n486));
  AND3_X1   g300(.A1(new_n479), .A2(new_n483), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n486), .B1(new_n479), .B2(new_n483), .ZN(new_n488));
  NOR2_X1   g302(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(KEYINPUT25), .B1(new_n489), .B2(new_n286), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT25), .ZN(new_n491));
  NOR4_X1   g305(.A1(new_n487), .A2(new_n488), .A3(new_n491), .A4(G902), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n460), .B1(new_n490), .B2(new_n492), .ZN(new_n493));
  NOR2_X1   g307(.A1(new_n460), .A2(G902), .ZN(new_n494));
  XNOR2_X1  g308(.A(new_n494), .B(KEYINPUT78), .ZN(new_n495));
  NAND2_X1  g309(.A1(new_n489), .A2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n493), .A2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n497), .ZN(new_n498));
  NOR3_X1   g312(.A1(new_n357), .A2(new_n459), .A3(G953), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n204), .A2(G143), .ZN(new_n500));
  INV_X1    g314(.A(KEYINPUT13), .ZN(new_n501));
  AOI21_X1  g315(.A(new_n222), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(G128), .B(G143), .ZN(new_n503));
  XOR2_X1   g317(.A(new_n502), .B(new_n503), .Z(new_n504));
  XNOR2_X1  g318(.A(G116), .B(G122), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n505), .B(new_n188), .ZN(new_n506));
  NAND2_X1  g320(.A1(new_n506), .A2(KEYINPUT94), .ZN(new_n507));
  INV_X1    g321(.A(new_n505), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(G107), .ZN(new_n509));
  INV_X1    g323(.A(KEYINPUT94), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n505), .A2(new_n188), .ZN(new_n511));
  NAND3_X1  g325(.A1(new_n509), .A2(new_n510), .A3(new_n511), .ZN(new_n512));
  AOI21_X1  g326(.A(new_n504), .B1(new_n507), .B2(new_n512), .ZN(new_n513));
  XNOR2_X1  g327(.A(new_n503), .B(new_n222), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n299), .A2(KEYINPUT14), .A3(G122), .ZN(new_n515));
  OAI211_X1 g329(.A(G107), .B(new_n515), .C1(new_n508), .C2(KEYINPUT14), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT95), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g332(.A1(new_n505), .A2(KEYINPUT95), .A3(new_n188), .ZN(new_n519));
  NAND4_X1  g333(.A1(new_n514), .A2(new_n516), .A3(new_n518), .A4(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n499), .B1(new_n513), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n507), .A2(new_n512), .ZN(new_n523));
  INV_X1    g337(.A(new_n504), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(new_n499), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n525), .A2(new_n526), .A3(new_n520), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n522), .A2(new_n527), .A3(KEYINPUT96), .A4(new_n286), .ZN(new_n528));
  INV_X1    g342(.A(G478), .ZN(new_n529));
  NOR2_X1   g343(.A1(new_n529), .A2(KEYINPUT15), .ZN(new_n530));
  AND2_X1   g344(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n528), .A2(new_n530), .ZN(new_n532));
  OR2_X1    g346(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(G234), .A2(G237), .ZN(new_n534));
  NAND3_X1  g348(.A1(new_n534), .A2(G902), .A3(G953), .ZN(new_n535));
  XOR2_X1   g349(.A(new_n535), .B(KEYINPUT97), .Z(new_n536));
  XNOR2_X1  g350(.A(KEYINPUT21), .B(G898), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AND3_X1   g352(.A1(new_n534), .A2(G952), .A3(new_n256), .ZN(new_n539));
  INV_X1    g353(.A(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g355(.A(new_n541), .ZN(new_n542));
  NOR2_X1   g356(.A1(new_n533), .A2(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT20), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n380), .A2(G214), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n546), .A2(new_n202), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n380), .A2(G143), .A3(G214), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(KEYINPUT18), .A2(G131), .ZN(new_n550));
  XNOR2_X1  g364(.A(new_n549), .B(new_n550), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n323), .A2(G140), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n463), .A2(G125), .ZN(new_n553));
  OAI21_X1  g367(.A(KEYINPUT88), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n323), .A2(G140), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT88), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n464), .A2(new_n555), .A3(new_n556), .ZN(new_n557));
  NAND3_X1  g371(.A1(new_n554), .A2(G146), .A3(new_n557), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n558), .A2(new_n480), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n551), .A2(new_n559), .ZN(new_n560));
  XNOR2_X1  g374(.A(G113), .B(G122), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n561), .B(G104), .ZN(new_n562));
  XNOR2_X1  g376(.A(new_n562), .B(KEYINPUT92), .ZN(new_n563));
  AOI21_X1  g377(.A(new_n229), .B1(new_n547), .B2(new_n548), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT17), .ZN(new_n565));
  XNOR2_X1  g379(.A(new_n549), .B(G131), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n565), .B1(new_n566), .B2(KEYINPUT17), .ZN(new_n567));
  OAI211_X1 g381(.A(new_n560), .B(new_n563), .C1(new_n567), .C2(new_n471), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n562), .ZN(new_n570));
  INV_X1    g384(.A(KEYINPUT90), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT19), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n571), .B1(new_n461), .B2(new_n572), .ZN(new_n573));
  AND4_X1   g387(.A1(new_n571), .A2(new_n464), .A3(new_n555), .A4(new_n572), .ZN(new_n574));
  NOR2_X1   g388(.A1(new_n573), .A2(new_n574), .ZN(new_n575));
  NAND3_X1  g389(.A1(new_n554), .A2(KEYINPUT19), .A3(new_n557), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT89), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g392(.A1(new_n554), .A2(KEYINPUT89), .A3(KEYINPUT19), .A4(new_n557), .ZN(new_n579));
  AOI211_X1 g393(.A(G146), .B(new_n575), .C1(new_n578), .C2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n549), .A2(G131), .ZN(new_n581));
  OAI21_X1  g395(.A(new_n466), .B1(new_n581), .B2(new_n564), .ZN(new_n582));
  OAI21_X1  g396(.A(new_n560), .B1(new_n580), .B2(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n570), .B1(new_n583), .B2(KEYINPUT91), .ZN(new_n584));
  INV_X1    g398(.A(KEYINPUT91), .ZN(new_n585));
  OAI211_X1 g399(.A(new_n585), .B(new_n560), .C1(new_n580), .C2(new_n582), .ZN(new_n586));
  AOI21_X1  g400(.A(new_n569), .B1(new_n584), .B2(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(G475), .A2(G902), .ZN(new_n588));
  INV_X1    g402(.A(new_n588), .ZN(new_n589));
  OAI211_X1 g403(.A(KEYINPUT93), .B(new_n545), .C1(new_n587), .C2(new_n589), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n560), .B1(new_n567), .B2(new_n471), .ZN(new_n591));
  AND2_X1   g405(.A1(new_n591), .A2(new_n562), .ZN(new_n592));
  OAI21_X1  g406(.A(new_n286), .B1(new_n592), .B2(new_n569), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n593), .A2(G475), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n582), .B1(new_n595), .B2(new_n200), .ZN(new_n596));
  INV_X1    g410(.A(new_n560), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT91), .B1(new_n596), .B2(new_n597), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n598), .A2(new_n562), .A3(new_n586), .ZN(new_n599));
  AOI21_X1  g413(.A(new_n589), .B1(new_n599), .B2(new_n568), .ZN(new_n600));
  INV_X1    g414(.A(KEYINPUT93), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT20), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  AOI211_X1 g416(.A(KEYINPUT93), .B(new_n589), .C1(new_n599), .C2(new_n568), .ZN(new_n603));
  OAI211_X1 g417(.A(new_n590), .B(new_n594), .C1(new_n602), .C2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(KEYINPUT98), .B1(new_n544), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n599), .A2(new_n568), .ZN(new_n606));
  AOI21_X1  g420(.A(new_n601), .B1(new_n606), .B2(new_n588), .ZN(new_n607));
  AOI22_X1  g421(.A1(new_n607), .A2(new_n545), .B1(G475), .B2(new_n593), .ZN(new_n608));
  OAI21_X1  g422(.A(KEYINPUT93), .B1(new_n587), .B2(new_n589), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n600), .A2(new_n601), .ZN(new_n610));
  NAND3_X1  g424(.A1(new_n609), .A2(new_n610), .A3(KEYINPUT20), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT98), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n543), .A2(new_n608), .A3(new_n611), .A4(new_n612), .ZN(new_n613));
  NAND2_X1  g427(.A1(new_n605), .A2(new_n613), .ZN(new_n614));
  NAND4_X1  g428(.A1(new_n359), .A2(new_n458), .A3(new_n498), .A4(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(new_n615), .B(G101), .ZN(G3));
  OAI21_X1  g430(.A(new_n286), .B1(new_n402), .B2(new_n405), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n617), .A2(G472), .ZN(new_n618));
  AND3_X1   g432(.A1(new_n408), .A2(new_n618), .A3(new_n416), .ZN(new_n619));
  INV_X1    g433(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n292), .A2(new_n358), .ZN(new_n621));
  NOR3_X1   g435(.A1(new_n620), .A2(new_n621), .A3(new_n497), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n525), .A2(new_n520), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n623), .A2(KEYINPUT99), .A3(new_n526), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n624), .A2(KEYINPUT33), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n526), .B1(new_n623), .B2(KEYINPUT99), .ZN(new_n626));
  OAI21_X1  g440(.A(KEYINPUT100), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n626), .ZN(new_n628));
  INV_X1    g442(.A(KEYINPUT100), .ZN(new_n629));
  NAND4_X1  g443(.A1(new_n628), .A2(new_n629), .A3(KEYINPUT33), .A4(new_n624), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n522), .A2(new_n527), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n631), .A2(KEYINPUT33), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n529), .A2(G902), .ZN(new_n633));
  NAND4_X1  g447(.A1(new_n627), .A2(new_n630), .A3(new_n632), .A4(new_n633), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n529), .B1(new_n631), .B2(G902), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n604), .A2(new_n636), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n352), .A2(new_n355), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n638), .A2(new_n293), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n637), .A2(new_n542), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n622), .A2(new_n640), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n641), .B(new_n195), .ZN(new_n642));
  XNOR2_X1  g456(.A(KEYINPUT101), .B(KEYINPUT34), .ZN(new_n643));
  XNOR2_X1  g457(.A(new_n642), .B(new_n643), .ZN(G6));
  NAND3_X1  g458(.A1(new_n608), .A2(new_n611), .A3(new_n533), .ZN(new_n645));
  XOR2_X1   g459(.A(new_n541), .B(KEYINPUT102), .Z(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NOR3_X1   g461(.A1(new_n645), .A2(new_n639), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n622), .A2(new_n648), .ZN(new_n649));
  XNOR2_X1  g463(.A(new_n649), .B(new_n188), .ZN(new_n650));
  XOR2_X1   g464(.A(KEYINPUT103), .B(KEYINPUT35), .Z(new_n651));
  XNOR2_X1  g465(.A(new_n650), .B(new_n651), .ZN(G9));
  AOI21_X1  g466(.A(KEYINPUT69), .B1(new_n415), .B2(new_n360), .ZN(new_n653));
  AOI211_X1 g467(.A(new_n407), .B(new_n452), .C1(new_n413), .C2(new_n414), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  NAND2_X1  g469(.A1(new_n479), .A2(new_n483), .ZN(new_n656));
  INV_X1    g470(.A(new_n486), .ZN(new_n657));
  NOR2_X1   g471(.A1(new_n657), .A2(KEYINPUT36), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n656), .B(new_n658), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n495), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n493), .A2(new_n660), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n655), .A2(KEYINPUT104), .A3(new_n618), .A4(new_n661), .ZN(new_n662));
  NAND4_X1  g476(.A1(new_n408), .A2(new_n618), .A3(new_n416), .A4(new_n661), .ZN(new_n663));
  INV_X1    g477(.A(KEYINPUT104), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n359), .A2(new_n662), .A3(new_n665), .A4(new_n614), .ZN(new_n666));
  XNOR2_X1  g480(.A(KEYINPUT37), .B(G110), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT105), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n666), .B(new_n668), .ZN(G12));
  INV_X1    g483(.A(G900), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n536), .A2(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n671), .A2(new_n540), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n645), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n359), .A2(new_n458), .A3(new_n661), .A4(new_n674), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n675), .B(G128), .ZN(G30));
  XNOR2_X1  g490(.A(new_n638), .B(KEYINPUT38), .ZN(new_n677));
  INV_X1    g491(.A(new_n661), .ZN(new_n678));
  AND2_X1   g492(.A1(new_n533), .A2(new_n293), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n677), .A2(new_n604), .A3(new_n678), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n672), .B(KEYINPUT39), .ZN(new_n681));
  AND3_X1   g495(.A1(new_n292), .A2(new_n358), .A3(new_n681), .ZN(new_n682));
  INV_X1    g496(.A(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n680), .B1(new_n683), .B2(KEYINPUT40), .ZN(new_n684));
  INV_X1    g498(.A(KEYINPUT108), .ZN(new_n685));
  NOR3_X1   g499(.A1(new_n653), .A2(new_n654), .A3(KEYINPUT32), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n389), .A2(new_n391), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n434), .A2(new_n384), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT106), .ZN(new_n689));
  NAND2_X1  g503(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND3_X1  g504(.A1(new_n434), .A2(KEYINPUT106), .A3(new_n384), .ZN(new_n691));
  AOI21_X1  g505(.A(new_n687), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  INV_X1    g506(.A(KEYINPUT107), .ZN(new_n693));
  AND2_X1   g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n286), .B1(new_n692), .B2(new_n693), .ZN(new_n695));
  OAI21_X1  g509(.A(G472), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n456), .A2(new_n696), .A3(new_n457), .ZN(new_n697));
  OAI21_X1  g511(.A(new_n685), .B1(new_n686), .B2(new_n697), .ZN(new_n698));
  AND3_X1   g512(.A1(new_n456), .A2(new_n457), .A3(new_n696), .ZN(new_n699));
  NAND3_X1  g513(.A1(new_n699), .A2(KEYINPUT108), .A3(new_n417), .ZN(new_n700));
  NAND2_X1  g514(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n684), .B(new_n701), .C1(KEYINPUT40), .C2(new_n683), .ZN(new_n702));
  XNOR2_X1  g516(.A(new_n702), .B(G143), .ZN(G45));
  NAND3_X1  g517(.A1(new_n604), .A2(new_n636), .A3(new_n672), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n292), .A3(new_n356), .A4(new_n358), .ZN(new_n706));
  INV_X1    g520(.A(new_n706), .ZN(new_n707));
  NAND3_X1  g521(.A1(new_n707), .A2(new_n458), .A3(new_n661), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  OAI21_X1  g523(.A(new_n255), .B1(new_n276), .B2(new_n277), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n289), .B1(new_n710), .B2(new_n280), .ZN(new_n711));
  OAI21_X1  g525(.A(G469), .B1(new_n711), .B2(G902), .ZN(new_n712));
  AND3_X1   g526(.A1(new_n712), .A2(new_n290), .A3(new_n358), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n458), .A2(new_n498), .A3(new_n640), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT41), .B(G113), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n714), .B(new_n715), .ZN(G15));
  NAND4_X1  g530(.A1(new_n458), .A2(new_n498), .A3(new_n648), .A4(new_n713), .ZN(new_n717));
  XNOR2_X1  g531(.A(new_n717), .B(G116), .ZN(G18));
  NAND3_X1  g532(.A1(new_n712), .A2(new_n290), .A3(new_n358), .ZN(new_n719));
  NOR2_X1   g533(.A1(new_n719), .A2(new_n639), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n458), .A2(new_n614), .A3(new_n661), .A4(new_n720), .ZN(new_n721));
  XNOR2_X1  g535(.A(new_n721), .B(G119), .ZN(G21));
  NAND2_X1  g536(.A1(new_n439), .A2(new_n378), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(new_n384), .ZN(new_n724));
  AOI21_X1  g538(.A(new_n452), .B1(new_n403), .B2(new_n724), .ZN(new_n725));
  XOR2_X1   g539(.A(KEYINPUT109), .B(G472), .Z(new_n726));
  AOI211_X1 g540(.A(new_n725), .B(new_n497), .C1(new_n617), .C2(new_n726), .ZN(new_n727));
  AND4_X1   g541(.A1(new_n604), .A2(new_n356), .A3(new_n533), .A4(new_n646), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n713), .A2(new_n727), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g543(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n730));
  NAND4_X1  g544(.A1(new_n604), .A2(new_n356), .A3(new_n533), .A4(new_n646), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n719), .A2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n732), .A2(new_n733), .A3(new_n727), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n730), .A2(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G122), .ZN(G24));
  AOI22_X1  g550(.A1(new_n608), .A2(new_n611), .B1(new_n635), .B2(new_n634), .ZN(new_n737));
  AOI21_X1  g551(.A(KEYINPUT111), .B1(new_n737), .B2(new_n672), .ZN(new_n738));
  AND4_X1   g552(.A1(KEYINPUT111), .A2(new_n604), .A3(new_n636), .A4(new_n672), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  AOI211_X1 g554(.A(new_n725), .B(new_n678), .C1(new_n617), .C2(new_n726), .ZN(new_n741));
  NAND3_X1  g555(.A1(new_n740), .A2(new_n720), .A3(new_n741), .ZN(new_n742));
  XNOR2_X1  g556(.A(new_n742), .B(G125), .ZN(G27));
  NOR2_X1   g557(.A1(new_n638), .A2(new_n294), .ZN(new_n744));
  NAND2_X1  g558(.A1(new_n744), .A2(new_n358), .ZN(new_n745));
  NOR3_X1   g559(.A1(new_n711), .A2(G469), .A3(G902), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n291), .B(KEYINPUT112), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n278), .A2(new_n281), .ZN(new_n748));
  OAI21_X1  g562(.A(new_n747), .B1(new_n748), .B2(new_n285), .ZN(new_n749));
  OAI21_X1  g563(.A(KEYINPUT113), .B1(new_n746), .B2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(new_n747), .ZN(new_n751));
  NOR2_X1   g565(.A1(new_n267), .A2(new_n273), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n751), .B1(new_n752), .B2(G469), .ZN(new_n753));
  INV_X1    g567(.A(KEYINPUT113), .ZN(new_n754));
  NAND3_X1  g568(.A1(new_n290), .A2(new_n753), .A3(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n745), .B1(new_n750), .B2(new_n755), .ZN(new_n756));
  NAND4_X1  g570(.A1(new_n740), .A2(new_n756), .A3(new_n458), .A4(new_n498), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT42), .ZN(new_n758));
  INV_X1    g572(.A(G472), .ZN(new_n759));
  AOI21_X1  g573(.A(new_n442), .B1(new_n441), .B2(new_n286), .ZN(new_n760));
  AOI211_X1 g574(.A(KEYINPUT72), .B(G902), .C1(new_n439), .C2(new_n440), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n760), .A2(new_n761), .ZN(new_n762));
  AOI211_X1 g576(.A(new_n446), .B(new_n759), .C1(new_n762), .C2(new_n448), .ZN(new_n763));
  AOI21_X1  g577(.A(KEYINPUT73), .B1(new_n449), .B2(G472), .ZN(new_n764));
  NOR2_X1   g578(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  AOI21_X1  g579(.A(new_n452), .B1(new_n413), .B2(new_n414), .ZN(new_n766));
  OAI21_X1  g580(.A(new_n454), .B1(new_n766), .B2(KEYINPUT32), .ZN(new_n767));
  OAI211_X1 g581(.A(KEYINPUT42), .B(new_n498), .C1(new_n765), .C2(new_n767), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n737), .A2(KEYINPUT111), .A3(new_n672), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT111), .ZN(new_n770));
  NAND2_X1  g584(.A1(new_n704), .A2(new_n770), .ZN(new_n771));
  NAND2_X1  g585(.A1(new_n769), .A2(new_n771), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n768), .A2(new_n772), .ZN(new_n773));
  AOI22_X1  g587(.A1(new_n757), .A2(new_n758), .B1(new_n773), .B2(new_n756), .ZN(new_n774));
  XOR2_X1   g588(.A(KEYINPUT114), .B(G131), .Z(new_n775));
  XNOR2_X1  g589(.A(new_n774), .B(new_n775), .ZN(G33));
  NAND4_X1  g590(.A1(new_n756), .A2(new_n458), .A3(new_n498), .A4(new_n674), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(G134), .ZN(G36));
  INV_X1    g592(.A(new_n744), .ZN(new_n779));
  AOI21_X1  g593(.A(new_n604), .B1(new_n635), .B2(new_n634), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT43), .ZN(new_n781));
  NAND3_X1  g595(.A1(new_n781), .A2(new_n620), .A3(new_n661), .ZN(new_n782));
  INV_X1    g596(.A(KEYINPUT44), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n784), .B1(new_n783), .B2(new_n782), .ZN(new_n785));
  INV_X1    g599(.A(new_n358), .ZN(new_n786));
  INV_X1    g600(.A(KEYINPUT45), .ZN(new_n787));
  OAI21_X1  g601(.A(G469), .B1(new_n748), .B2(new_n787), .ZN(new_n788));
  NAND2_X1  g602(.A1(new_n274), .A2(new_n283), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n788), .B1(new_n789), .B2(new_n787), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(new_n751), .ZN(new_n791));
  INV_X1    g605(.A(KEYINPUT46), .ZN(new_n792));
  AOI21_X1  g606(.A(new_n746), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OR3_X1    g607(.A1(new_n790), .A2(new_n792), .A3(new_n751), .ZN(new_n794));
  AOI21_X1  g608(.A(new_n786), .B1(new_n793), .B2(new_n794), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n681), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n785), .A2(new_n796), .ZN(new_n797));
  XNOR2_X1  g611(.A(KEYINPUT115), .B(G137), .ZN(new_n798));
  XNOR2_X1  g612(.A(new_n797), .B(new_n798), .ZN(G39));
  INV_X1    g613(.A(KEYINPUT47), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n793), .A2(new_n794), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n800), .B1(new_n801), .B2(new_n786), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n795), .A2(KEYINPUT47), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NOR4_X1   g618(.A1(new_n458), .A2(new_n498), .A3(new_n704), .A4(new_n779), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n804), .A2(new_n805), .ZN(new_n806));
  XNOR2_X1  g620(.A(new_n806), .B(G140), .ZN(G42));
  AND2_X1   g621(.A1(new_n781), .A2(new_n539), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n765), .A2(new_n767), .ZN(new_n809));
  NOR2_X1   g623(.A1(new_n809), .A2(new_n497), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n713), .A2(new_n744), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n808), .A2(new_n810), .A3(new_n812), .ZN(new_n813));
  XNOR2_X1  g627(.A(new_n813), .B(KEYINPUT48), .ZN(new_n814));
  INV_X1    g628(.A(new_n701), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n811), .A2(new_n497), .A3(new_n540), .ZN(new_n816));
  NAND3_X1  g630(.A1(new_n815), .A2(new_n737), .A3(new_n816), .ZN(new_n817));
  INV_X1    g631(.A(G952), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n781), .A2(new_n539), .A3(new_n727), .ZN(new_n819));
  INV_X1    g633(.A(new_n819), .ZN(new_n820));
  AOI211_X1 g634(.A(new_n818), .B(G953), .C1(new_n820), .C2(new_n720), .ZN(new_n821));
  NAND3_X1  g635(.A1(new_n814), .A2(new_n817), .A3(new_n821), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n712), .A2(new_n290), .A3(new_n786), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n802), .A2(new_n803), .A3(new_n823), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n824), .A2(new_n744), .A3(new_n820), .ZN(new_n825));
  NAND3_X1  g639(.A1(new_n808), .A2(new_n741), .A3(new_n812), .ZN(new_n826));
  NOR2_X1   g640(.A1(new_n604), .A2(new_n636), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n815), .A2(new_n816), .A3(new_n827), .ZN(new_n828));
  INV_X1    g642(.A(KEYINPUT50), .ZN(new_n829));
  INV_X1    g643(.A(new_n677), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n830), .A2(new_n713), .A3(new_n294), .ZN(new_n831));
  OR2_X1    g645(.A1(new_n819), .A2(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n829), .B1(new_n832), .B2(KEYINPUT118), .ZN(new_n833));
  OAI211_X1 g647(.A(KEYINPUT118), .B(new_n829), .C1(new_n819), .C2(new_n831), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI211_X1 g649(.A(new_n826), .B(new_n828), .C1(new_n833), .C2(new_n835), .ZN(new_n836));
  OAI21_X1  g650(.A(KEYINPUT51), .B1(new_n825), .B2(new_n836), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n826), .A2(new_n828), .ZN(new_n838));
  INV_X1    g652(.A(new_n833), .ZN(new_n839));
  AOI21_X1  g653(.A(new_n838), .B1(new_n839), .B2(new_n834), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n824), .A2(new_n744), .A3(new_n820), .ZN(new_n842));
  NAND3_X1  g656(.A1(new_n840), .A2(new_n841), .A3(new_n842), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n822), .B1(new_n837), .B2(new_n843), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n678), .A2(new_n604), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n356), .A2(new_n533), .A3(new_n358), .A4(new_n672), .ZN(new_n846));
  AOI211_X1 g660(.A(new_n845), .B(new_n846), .C1(new_n750), .C2(new_n755), .ZN(new_n847));
  NOR3_X1   g661(.A1(new_n686), .A2(new_n697), .A3(new_n685), .ZN(new_n848));
  AOI21_X1  g662(.A(KEYINPUT108), .B1(new_n699), .B2(new_n417), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n847), .B1(new_n848), .B2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(new_n708), .A3(new_n675), .A4(new_n742), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n852));
  OAI211_X1 g666(.A(new_n456), .B(new_n457), .C1(new_n763), .C2(new_n764), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AOI21_X1  g668(.A(new_n678), .B1(new_n854), .B2(new_n417), .ZN(new_n855));
  AOI22_X1  g669(.A1(new_n701), .A2(new_n847), .B1(new_n855), .B2(new_n707), .ZN(new_n856));
  INV_X1    g670(.A(new_n674), .ZN(new_n857));
  NOR3_X1   g671(.A1(new_n621), .A2(new_n857), .A3(new_n639), .ZN(new_n858));
  AND2_X1   g672(.A1(new_n720), .A2(new_n741), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n855), .A2(new_n858), .B1(new_n859), .B2(new_n740), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT52), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n856), .A2(new_n860), .A3(new_n861), .ZN(new_n862));
  AND2_X1   g676(.A1(new_n852), .A2(new_n862), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n735), .A2(new_n666), .A3(new_n714), .A4(new_n717), .ZN(new_n864));
  AOI211_X1 g678(.A(new_n647), .B(new_n639), .C1(new_n637), .C2(new_n645), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n292), .A2(new_n358), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n865), .A2(new_n866), .A3(new_n498), .A4(new_n619), .ZN(new_n867));
  NAND3_X1  g681(.A1(new_n615), .A2(new_n867), .A3(new_n721), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n531), .A2(new_n532), .A3(new_n673), .ZN(new_n869));
  NAND4_X1  g683(.A1(new_n352), .A2(new_n869), .A3(new_n293), .A4(new_n355), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n604), .A2(new_n870), .ZN(new_n871));
  INV_X1    g685(.A(KEYINPUT116), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n871), .A2(new_n872), .ZN(new_n873));
  OAI21_X1  g687(.A(KEYINPUT116), .B1(new_n604), .B2(new_n870), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n873), .A2(new_n874), .ZN(new_n875));
  NAND4_X1  g689(.A1(new_n458), .A2(new_n866), .A3(new_n875), .A4(new_n661), .ZN(new_n876));
  NAND3_X1  g690(.A1(new_n740), .A2(new_n756), .A3(new_n741), .ZN(new_n877));
  NAND3_X1  g691(.A1(new_n777), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NOR4_X1   g692(.A1(new_n864), .A2(new_n774), .A3(new_n868), .A4(new_n878), .ZN(new_n879));
  NAND3_X1  g693(.A1(new_n863), .A2(KEYINPUT53), .A3(new_n879), .ZN(new_n880));
  INV_X1    g694(.A(KEYINPUT53), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n675), .A2(new_n742), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n750), .A2(new_n755), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n846), .A2(new_n845), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n883), .A2(new_n884), .ZN(new_n885));
  AOI21_X1  g699(.A(new_n885), .B1(new_n698), .B2(new_n700), .ZN(new_n886));
  NAND2_X1  g700(.A1(new_n458), .A2(new_n661), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n887), .A2(new_n706), .ZN(new_n888));
  NOR3_X1   g702(.A1(new_n882), .A2(new_n886), .A3(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(KEYINPUT117), .B(KEYINPUT52), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n862), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NOR2_X1   g705(.A1(new_n729), .A2(KEYINPUT110), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n733), .B1(new_n732), .B2(new_n727), .ZN(new_n893));
  OAI21_X1  g707(.A(new_n717), .B1(new_n892), .B2(new_n893), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n666), .A2(new_n714), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n757), .A2(new_n758), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n773), .A2(new_n756), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n897), .A2(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(new_n868), .ZN(new_n900));
  INV_X1    g714(.A(new_n878), .ZN(new_n901));
  NAND4_X1  g715(.A1(new_n896), .A2(new_n899), .A3(new_n900), .A4(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n881), .B1(new_n891), .B2(new_n902), .ZN(new_n903));
  NAND2_X1  g717(.A1(new_n880), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n904), .A2(KEYINPUT54), .ZN(new_n905));
  NOR2_X1   g719(.A1(new_n851), .A2(KEYINPUT52), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n890), .B1(new_n856), .B2(new_n860), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n908), .A2(new_n879), .A3(KEYINPUT53), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n852), .A2(new_n862), .ZN(new_n910));
  OAI21_X1  g724(.A(new_n881), .B1(new_n910), .B2(new_n902), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n909), .A2(new_n911), .ZN(new_n912));
  OR2_X1    g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n844), .A2(new_n905), .A3(new_n913), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n914), .A2(KEYINPUT119), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT119), .ZN(new_n916));
  NAND4_X1  g730(.A1(new_n844), .A2(new_n916), .A3(new_n913), .A4(new_n905), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n818), .A2(new_n256), .ZN(new_n918));
  NAND3_X1  g732(.A1(new_n915), .A2(new_n917), .A3(new_n918), .ZN(new_n919));
  NOR3_X1   g733(.A1(new_n497), .A2(new_n294), .A3(new_n786), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n830), .A2(new_n780), .A3(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n712), .A2(new_n290), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n921), .B1(KEYINPUT49), .B2(new_n922), .ZN(new_n923));
  OAI211_X1 g737(.A(new_n815), .B(new_n923), .C1(KEYINPUT49), .C2(new_n922), .ZN(new_n924));
  NAND2_X1  g738(.A1(new_n919), .A2(new_n924), .ZN(G75));
  NOR2_X1   g739(.A1(new_n256), .A2(G952), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n286), .B1(new_n909), .B2(new_n911), .ZN(new_n928));
  AOI21_X1  g742(.A(KEYINPUT56), .B1(new_n928), .B2(G210), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n322), .A2(new_n329), .ZN(new_n930));
  XNOR2_X1  g744(.A(new_n930), .B(new_n327), .ZN(new_n931));
  XNOR2_X1  g745(.A(new_n931), .B(KEYINPUT55), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n927), .B1(new_n929), .B2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n929), .A2(new_n932), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT120), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND3_X1  g750(.A1(new_n929), .A2(KEYINPUT120), .A3(new_n932), .ZN(new_n937));
  AOI21_X1  g751(.A(new_n933), .B1(new_n936), .B2(new_n937), .ZN(G51));
  XNOR2_X1  g752(.A(new_n912), .B(KEYINPUT54), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n747), .B(KEYINPUT121), .ZN(new_n940));
  XOR2_X1   g754(.A(new_n940), .B(KEYINPUT57), .Z(new_n941));
  NAND2_X1  g755(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n942), .B1(new_n288), .B2(new_n289), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n928), .A2(new_n790), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n926), .B1(new_n943), .B2(new_n944), .ZN(G54));
  NAND3_X1  g759(.A1(new_n928), .A2(KEYINPUT58), .A3(G475), .ZN(new_n946));
  AND2_X1   g760(.A1(new_n946), .A2(new_n587), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n946), .A2(new_n587), .ZN(new_n948));
  NOR3_X1   g762(.A1(new_n947), .A2(new_n948), .A3(new_n926), .ZN(G60));
  AND3_X1   g763(.A1(new_n627), .A2(new_n630), .A3(new_n632), .ZN(new_n950));
  NAND2_X1  g764(.A1(G478), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT59), .ZN(new_n952));
  AND3_X1   g766(.A1(new_n939), .A2(new_n950), .A3(new_n952), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n913), .A2(new_n905), .ZN(new_n954));
  AOI21_X1  g768(.A(new_n950), .B1(new_n954), .B2(new_n952), .ZN(new_n955));
  NOR3_X1   g769(.A1(new_n953), .A2(new_n955), .A3(new_n926), .ZN(G63));
  NAND2_X1  g770(.A1(G217), .A2(G902), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT60), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n912), .A2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n489), .ZN(new_n961));
  NAND3_X1  g775(.A1(new_n960), .A2(KEYINPUT122), .A3(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(KEYINPUT122), .ZN(new_n963));
  AOI21_X1  g777(.A(new_n958), .B1(new_n909), .B2(new_n911), .ZN(new_n964));
  OAI21_X1  g778(.A(new_n963), .B1(new_n964), .B2(new_n489), .ZN(new_n965));
  AOI21_X1  g779(.A(new_n926), .B1(new_n964), .B2(new_n659), .ZN(new_n966));
  NAND4_X1  g780(.A1(new_n962), .A2(new_n965), .A3(new_n966), .A4(KEYINPUT61), .ZN(new_n967));
  INV_X1    g781(.A(KEYINPUT61), .ZN(new_n968));
  AOI21_X1  g782(.A(KEYINPUT53), .B1(new_n863), .B2(new_n879), .ZN(new_n969));
  NOR3_X1   g783(.A1(new_n891), .A2(new_n902), .A3(new_n881), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n659), .B(new_n959), .C1(new_n969), .C2(new_n970), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n927), .ZN(new_n972));
  NOR2_X1   g786(.A1(new_n964), .A2(new_n489), .ZN(new_n973));
  OAI21_X1  g787(.A(new_n968), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n967), .A2(new_n974), .ZN(new_n975));
  INV_X1    g789(.A(KEYINPUT123), .ZN(new_n976));
  NAND2_X1  g790(.A1(new_n975), .A2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n967), .A2(new_n974), .A3(KEYINPUT123), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n977), .A2(new_n978), .ZN(G66));
  INV_X1    g793(.A(G224), .ZN(new_n980));
  OAI21_X1  g794(.A(G953), .B1(new_n537), .B2(new_n980), .ZN(new_n981));
  NOR2_X1   g795(.A1(new_n864), .A2(new_n868), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n981), .B1(new_n982), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n930), .B1(G898), .B2(new_n256), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n983), .B(new_n984), .ZN(G69));
  NAND2_X1  g799(.A1(new_n422), .A2(new_n386), .ZN(new_n986));
  XNOR2_X1  g800(.A(new_n595), .B(KEYINPUT124), .ZN(new_n987));
  XNOR2_X1  g801(.A(new_n986), .B(new_n987), .ZN(new_n988));
  NAND2_X1  g802(.A1(G900), .A2(G953), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT127), .ZN(new_n990));
  NOR2_X1   g804(.A1(new_n882), .A2(new_n888), .ZN(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n990), .B1(new_n797), .B2(new_n992), .ZN(new_n993));
  OAI211_X1 g807(.A(KEYINPUT127), .B(new_n991), .C1(new_n785), .C2(new_n796), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND3_X1  g809(.A1(new_n604), .A2(new_n356), .A3(new_n533), .ZN(new_n996));
  NOR4_X1   g810(.A1(new_n796), .A2(new_n497), .A3(new_n996), .A4(new_n809), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n899), .A2(new_n777), .ZN(new_n998));
  NOR2_X1   g812(.A1(new_n997), .A2(new_n998), .ZN(new_n999));
  NAND3_X1  g813(.A1(new_n995), .A2(new_n999), .A3(new_n806), .ZN(new_n1000));
  OAI211_X1 g814(.A(new_n988), .B(new_n989), .C1(new_n1000), .C2(G953), .ZN(new_n1001));
  AOI21_X1  g815(.A(new_n779), .B1(new_n637), .B2(new_n645), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n682), .A2(new_n458), .A3(new_n498), .A4(new_n1002), .ZN(new_n1003));
  XOR2_X1   g817(.A(new_n1003), .B(KEYINPUT125), .Z(new_n1004));
  OAI21_X1  g818(.A(new_n1004), .B1(new_n785), .B2(new_n796), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1005), .B1(new_n804), .B2(new_n805), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n702), .A2(new_n991), .ZN(new_n1007));
  INV_X1    g821(.A(KEYINPUT62), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1007), .B(new_n1008), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1006), .A2(new_n1009), .ZN(new_n1010));
  INV_X1    g824(.A(KEYINPUT126), .ZN(new_n1011));
  NAND2_X1  g825(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND3_X1  g826(.A1(new_n1006), .A2(new_n1009), .A3(KEYINPUT126), .ZN(new_n1013));
  AOI21_X1  g827(.A(G953), .B1(new_n1012), .B2(new_n1013), .ZN(new_n1014));
  OAI21_X1  g828(.A(new_n1001), .B1(new_n1014), .B2(new_n988), .ZN(new_n1015));
  AOI21_X1  g829(.A(new_n256), .B1(G227), .B2(G900), .ZN(new_n1016));
  NAND2_X1  g830(.A1(new_n1015), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g831(.A(new_n1016), .ZN(new_n1018));
  OAI211_X1 g832(.A(new_n1001), .B(new_n1018), .C1(new_n1014), .C2(new_n988), .ZN(new_n1019));
  NAND2_X1  g833(.A1(new_n1017), .A2(new_n1019), .ZN(G72));
  NAND2_X1  g834(.A1(G472), .A2(G902), .ZN(new_n1021));
  XOR2_X1   g835(.A(new_n1021), .B(KEYINPUT63), .Z(new_n1022));
  INV_X1    g836(.A(new_n982), .ZN(new_n1023));
  OAI21_X1  g837(.A(new_n1022), .B1(new_n1000), .B2(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n1024), .A2(new_n384), .A3(new_n423), .ZN(new_n1025));
  NAND2_X1  g839(.A1(new_n424), .A2(new_n426), .ZN(new_n1026));
  OAI211_X1 g840(.A(new_n904), .B(new_n1022), .C1(new_n687), .C2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1025), .A2(new_n927), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g842(.A1(new_n1012), .A2(new_n982), .A3(new_n1013), .ZN(new_n1029));
  AOI211_X1 g843(.A(new_n384), .B(new_n423), .C1(new_n1029), .C2(new_n1022), .ZN(new_n1030));
  NOR2_X1   g844(.A1(new_n1028), .A2(new_n1030), .ZN(G57));
endmodule


