//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 1 0 1 0 1 1 0 1 1 0 0 0 0 1 1 0 0 0 1 1 0 1 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 1 1 0 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:17 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n674, new_n675,
    new_n676, new_n677, new_n678, new_n679, new_n680, new_n681, new_n682,
    new_n683, new_n684, new_n685, new_n686, new_n687, new_n688, new_n689,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n695, new_n696,
    new_n697, new_n698, new_n699, new_n700, new_n701, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n718,
    new_n719, new_n720, new_n721, new_n722, new_n723, new_n724, new_n725,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n735, new_n736, new_n737, new_n738, new_n739, new_n740,
    new_n741, new_n742, new_n743, new_n744, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1049, new_n1050, new_n1051,
    new_n1052, new_n1053, new_n1054, new_n1055, new_n1056, new_n1057,
    new_n1058, new_n1059, new_n1060, new_n1061, new_n1062, new_n1063,
    new_n1064, new_n1065, new_n1066, new_n1067, new_n1068, new_n1069,
    new_n1070, new_n1071, new_n1072, new_n1073, new_n1074, new_n1075,
    new_n1076, new_n1077, new_n1078, new_n1079, new_n1080, new_n1081,
    new_n1082, new_n1083, new_n1084, new_n1085, new_n1086, new_n1087,
    new_n1088, new_n1089, new_n1090, new_n1091, new_n1093, new_n1094,
    new_n1095, new_n1096, new_n1097, new_n1098, new_n1099, new_n1100,
    new_n1101, new_n1102, new_n1103, new_n1104, new_n1105, new_n1106,
    new_n1107, new_n1108, new_n1109, new_n1110, new_n1111, new_n1112,
    new_n1113, new_n1114, new_n1115, new_n1116, new_n1117, new_n1118,
    new_n1119, new_n1120, new_n1121, new_n1122, new_n1123, new_n1124,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1147, new_n1148, new_n1149,
    new_n1150, new_n1151, new_n1152, new_n1153, new_n1154, new_n1155,
    new_n1156, new_n1157, new_n1158, new_n1159, new_n1160, new_n1161,
    new_n1162, new_n1163, new_n1164, new_n1165, new_n1166, new_n1167,
    new_n1168, new_n1169, new_n1170, new_n1171, new_n1172, new_n1173,
    new_n1174, new_n1175, new_n1176, new_n1177, new_n1178, new_n1179,
    new_n1180, new_n1181, new_n1182, new_n1183, new_n1184, new_n1185,
    new_n1186, new_n1187, new_n1188, new_n1189, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1217, new_n1218, new_n1219, new_n1220, new_n1221, new_n1222,
    new_n1223, new_n1224, new_n1225, new_n1226, new_n1227, new_n1228,
    new_n1229, new_n1230, new_n1231, new_n1232, new_n1233, new_n1234,
    new_n1235, new_n1236, new_n1237, new_n1238, new_n1239, new_n1240,
    new_n1241, new_n1242, new_n1243, new_n1244, new_n1245, new_n1246,
    new_n1247, new_n1248, new_n1249, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1255, new_n1256, new_n1257, new_n1258, new_n1259,
    new_n1260, new_n1261, new_n1262, new_n1263, new_n1264, new_n1265,
    new_n1266, new_n1267, new_n1268, new_n1269, new_n1270, new_n1271,
    new_n1272, new_n1273, new_n1274, new_n1275, new_n1276, new_n1278,
    new_n1279, new_n1280, new_n1281, new_n1282, new_n1283, new_n1284,
    new_n1285, new_n1286, new_n1287, new_n1288, new_n1290, new_n1291,
    new_n1292, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1311, new_n1312, new_n1313, new_n1314, new_n1315, new_n1316,
    new_n1317, new_n1318, new_n1319, new_n1320, new_n1321, new_n1322,
    new_n1323, new_n1324, new_n1325, new_n1326, new_n1327, new_n1328,
    new_n1329, new_n1330, new_n1331, new_n1332, new_n1333, new_n1334,
    new_n1335, new_n1336, new_n1337, new_n1338, new_n1339, new_n1340,
    new_n1341, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1352, new_n1353,
    new_n1354, new_n1355, new_n1356;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0002(.A(G1), .ZN(new_n203));
  INV_X1    g0003(.A(G20), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  INV_X1    g0005(.A(new_n205), .ZN(new_n206));
  XOR2_X1   g0006(.A(KEYINPUT66), .B(G77), .Z(new_n207));
  INV_X1    g0007(.A(G244), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  AOI22_X1  g0009(.A1(G107), .A2(G264), .B1(G116), .B2(G270), .ZN(new_n210));
  AOI22_X1  g0010(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n212));
  NAND2_X1  g0012(.A1(G58), .A2(G232), .ZN(new_n213));
  NAND4_X1  g0013(.A1(new_n210), .A2(new_n211), .A3(new_n212), .A4(new_n213), .ZN(new_n214));
  OAI21_X1  g0014(.A(new_n206), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  XNOR2_X1  g0015(.A(new_n215), .B(KEYINPUT1), .ZN(new_n216));
  OR3_X1    g0016(.A1(new_n206), .A2(KEYINPUT64), .A3(G13), .ZN(new_n217));
  OAI21_X1  g0017(.A(KEYINPUT64), .B1(new_n206), .B2(G13), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI211_X1 g0019(.A(new_n219), .B(G250), .C1(G257), .C2(G264), .ZN(new_n220));
  XOR2_X1   g0020(.A(new_n220), .B(KEYINPUT0), .Z(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n204), .ZN(new_n223));
  NOR2_X1   g0023(.A1(G58), .A2(G68), .ZN(new_n224));
  INV_X1    g0024(.A(KEYINPUT65), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(KEYINPUT65), .B1(G58), .B2(G68), .ZN(new_n227));
  NAND3_X1  g0027(.A1(new_n226), .A2(G50), .A3(new_n227), .ZN(new_n228));
  INV_X1    g0028(.A(new_n228), .ZN(new_n229));
  AOI211_X1 g0029(.A(new_n216), .B(new_n221), .C1(new_n223), .C2(new_n229), .ZN(G361));
  XOR2_X1   g0030(.A(G250), .B(G257), .Z(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XNOR2_X1  g0033(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n235), .B(KEYINPUT69), .ZN(new_n236));
  XNOR2_X1  g0036(.A(G238), .B(G244), .ZN(new_n237));
  INV_X1    g0037(.A(G232), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(KEYINPUT2), .B(G226), .Z(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  INV_X1    g0041(.A(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n236), .B(new_n242), .ZN(G358));
  XNOR2_X1  g0043(.A(G68), .B(G77), .ZN(new_n244));
  INV_X1    g0044(.A(G58), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  XNOR2_X1  g0046(.A(KEYINPUT70), .B(G50), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n246), .B(new_n247), .ZN(new_n248));
  XOR2_X1   g0048(.A(G87), .B(G97), .Z(new_n249));
  XNOR2_X1  g0049(.A(G107), .B(G116), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n248), .B(new_n251), .ZN(G351));
  NAND3_X1  g0052(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n253));
  NAND2_X1  g0053(.A1(new_n253), .A2(new_n222), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n254), .A2(KEYINPUT71), .ZN(new_n255));
  INV_X1    g0055(.A(KEYINPUT71), .ZN(new_n256));
  NAND3_X1  g0056(.A1(new_n253), .A2(new_n256), .A3(new_n222), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G13), .ZN(new_n259));
  NOR3_X1   g0059(.A1(new_n259), .A2(new_n204), .A3(G1), .ZN(new_n260));
  NOR2_X1   g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  OAI211_X1 g0061(.A(new_n261), .B(G50), .C1(G1), .C2(new_n204), .ZN(new_n262));
  XNOR2_X1  g0062(.A(KEYINPUT8), .B(G58), .ZN(new_n263));
  INV_X1    g0063(.A(G33), .ZN(new_n264));
  NOR2_X1   g0064(.A1(new_n264), .A2(G20), .ZN(new_n265));
  INV_X1    g0065(.A(new_n265), .ZN(new_n266));
  INV_X1    g0066(.A(G150), .ZN(new_n267));
  NOR2_X1   g0067(.A1(G20), .A2(G33), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  OAI22_X1  g0069(.A1(new_n263), .A2(new_n266), .B1(new_n267), .B2(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(G50), .ZN(new_n271));
  AOI21_X1  g0071(.A(new_n204), .B1(new_n224), .B2(new_n271), .ZN(new_n272));
  OAI21_X1  g0072(.A(new_n258), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  INV_X1    g0073(.A(new_n260), .ZN(new_n274));
  OAI211_X1 g0074(.A(new_n262), .B(new_n273), .C1(G50), .C2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  AOI21_X1  g0076(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n277));
  INV_X1    g0077(.A(G274), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n203), .B1(G41), .B2(G45), .ZN(new_n279));
  NOR3_X1   g0079(.A1(new_n277), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(new_n279), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n277), .A2(new_n281), .ZN(new_n282));
  AOI21_X1  g0082(.A(new_n280), .B1(G226), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g0083(.A(KEYINPUT3), .B(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G222), .A2(G1698), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n286), .A2(G223), .ZN(new_n287));
  OAI21_X1  g0087(.A(new_n284), .B1(new_n285), .B2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(new_n207), .ZN(new_n289));
  OAI211_X1 g0089(.A(new_n288), .B(new_n277), .C1(new_n289), .C2(new_n284), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n283), .A2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(G190), .ZN(new_n292));
  NOR2_X1   g0092(.A1(new_n291), .A2(new_n292), .ZN(new_n293));
  AOI21_X1  g0093(.A(new_n293), .B1(G200), .B2(new_n291), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n276), .A2(new_n294), .ZN(new_n295));
  XNOR2_X1  g0095(.A(new_n295), .B(KEYINPUT10), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT72), .ZN(new_n297));
  AOI21_X1  g0097(.A(new_n263), .B1(new_n297), .B2(new_n269), .ZN(new_n298));
  OAI21_X1  g0098(.A(new_n298), .B1(new_n297), .B2(new_n269), .ZN(new_n299));
  XNOR2_X1  g0099(.A(KEYINPUT15), .B(G87), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(new_n265), .ZN(new_n302));
  OAI21_X1  g0102(.A(new_n299), .B1(KEYINPUT73), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(KEYINPUT73), .ZN(new_n304));
  OAI21_X1  g0104(.A(new_n304), .B1(new_n204), .B2(new_n207), .ZN(new_n305));
  OAI21_X1  g0105(.A(new_n254), .B1(new_n303), .B2(new_n305), .ZN(new_n306));
  NOR2_X1   g0106(.A1(new_n260), .A2(new_n254), .ZN(new_n307));
  INV_X1    g0107(.A(G77), .ZN(new_n308));
  AOI21_X1  g0108(.A(new_n308), .B1(new_n203), .B2(G20), .ZN(new_n309));
  AOI22_X1  g0109(.A1(new_n307), .A2(new_n309), .B1(new_n207), .B2(new_n260), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n306), .A2(new_n310), .ZN(new_n311));
  NAND2_X1  g0111(.A1(new_n311), .A2(KEYINPUT74), .ZN(new_n312));
  INV_X1    g0112(.A(KEYINPUT74), .ZN(new_n313));
  NAND3_X1  g0113(.A1(new_n306), .A2(new_n313), .A3(new_n310), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n312), .A2(new_n314), .ZN(new_n315));
  NAND3_X1  g0115(.A1(new_n284), .A2(G238), .A3(G1698), .ZN(new_n316));
  NAND3_X1  g0116(.A1(new_n284), .A2(G232), .A3(new_n286), .ZN(new_n317));
  INV_X1    g0117(.A(G107), .ZN(new_n318));
  OAI211_X1 g0118(.A(new_n316), .B(new_n317), .C1(new_n318), .C2(new_n284), .ZN(new_n319));
  NAND2_X1  g0119(.A1(new_n319), .A2(new_n277), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n280), .B1(G244), .B2(new_n282), .ZN(new_n321));
  NAND2_X1  g0121(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NOR2_X1   g0122(.A1(new_n322), .A2(G179), .ZN(new_n323));
  INV_X1    g0123(.A(G169), .ZN(new_n324));
  AOI21_X1  g0124(.A(new_n323), .B1(new_n324), .B2(new_n322), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n315), .A2(new_n325), .ZN(new_n326));
  NAND3_X1  g0126(.A1(new_n320), .A2(G190), .A3(new_n321), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n322), .A2(G200), .ZN(new_n328));
  NAND4_X1  g0128(.A1(new_n312), .A2(new_n314), .A3(new_n327), .A4(new_n328), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n291), .A2(new_n324), .ZN(new_n330));
  INV_X1    g0130(.A(G179), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n283), .A2(new_n331), .A3(new_n290), .ZN(new_n332));
  NAND3_X1  g0132(.A1(new_n275), .A2(new_n330), .A3(new_n332), .ZN(new_n333));
  AND4_X1   g0133(.A1(new_n296), .A2(new_n326), .A3(new_n329), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n282), .A2(G238), .ZN(new_n335));
  NOR2_X1   g0135(.A1(new_n277), .A2(new_n278), .ZN(new_n336));
  INV_X1    g0136(.A(new_n336), .ZN(new_n337));
  OAI21_X1  g0137(.A(new_n335), .B1(new_n279), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(new_n277), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n238), .A2(G1698), .ZN(new_n340));
  OAI211_X1 g0140(.A(new_n284), .B(new_n340), .C1(G226), .C2(G1698), .ZN(new_n341));
  NAND2_X1  g0141(.A1(G33), .A2(G97), .ZN(new_n342));
  AOI21_X1  g0142(.A(new_n339), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g0143(.A(KEYINPUT13), .B1(new_n338), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(new_n343), .ZN(new_n345));
  AOI21_X1  g0145(.A(new_n280), .B1(G238), .B2(new_n282), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT13), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n345), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  NAND2_X1  g0148(.A1(new_n344), .A2(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(G200), .ZN(new_n351));
  NOR2_X1   g0151(.A1(new_n350), .A2(new_n351), .ZN(new_n352));
  OAI22_X1  g0152(.A1(new_n266), .A2(new_n308), .B1(new_n204), .B2(G68), .ZN(new_n353));
  OAI22_X1  g0153(.A1(new_n353), .A2(KEYINPUT75), .B1(new_n271), .B2(new_n269), .ZN(new_n354));
  AND2_X1   g0154(.A1(new_n353), .A2(KEYINPUT75), .ZN(new_n355));
  OAI21_X1  g0155(.A(new_n258), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT11), .ZN(new_n357));
  OR2_X1    g0157(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n356), .A2(new_n357), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT76), .ZN(new_n360));
  OAI22_X1  g0160(.A1(new_n274), .A2(G68), .B1(new_n360), .B2(KEYINPUT12), .ZN(new_n361));
  INV_X1    g0161(.A(KEYINPUT12), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(KEYINPUT76), .B2(new_n362), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n360), .B(KEYINPUT12), .C1(new_n274), .C2(G68), .ZN(new_n364));
  INV_X1    g0164(.A(G68), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n365), .B1(new_n203), .B2(G20), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n363), .A2(new_n364), .B1(new_n307), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g0167(.A1(new_n358), .A2(new_n359), .A3(new_n367), .ZN(new_n368));
  NOR2_X1   g0168(.A1(new_n349), .A2(new_n292), .ZN(new_n369));
  NOR3_X1   g0169(.A1(new_n352), .A2(new_n368), .A3(new_n369), .ZN(new_n370));
  INV_X1    g0170(.A(new_n370), .ZN(new_n371));
  NOR3_X1   g0171(.A1(new_n338), .A2(KEYINPUT13), .A3(new_n343), .ZN(new_n372));
  AOI21_X1  g0172(.A(new_n347), .B1(new_n345), .B2(new_n346), .ZN(new_n373));
  OAI21_X1  g0173(.A(G169), .B1(new_n372), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT14), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n350), .A2(G179), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT14), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n349), .A2(new_n377), .A3(G169), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n375), .A2(new_n376), .A3(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT77), .ZN(new_n381));
  NAND4_X1  g0181(.A1(new_n375), .A2(new_n376), .A3(new_n381), .A4(new_n378), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(new_n368), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n334), .A2(new_n371), .A3(new_n384), .ZN(new_n385));
  NOR2_X1   g0185(.A1(new_n245), .A2(new_n365), .ZN(new_n386));
  OAI21_X1  g0186(.A(G20), .B1(new_n386), .B2(new_n224), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n268), .A2(G159), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  INV_X1    g0189(.A(KEYINPUT7), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n390), .B1(new_n284), .B2(G20), .ZN(new_n391));
  NAND2_X1  g0191(.A1(new_n264), .A2(KEYINPUT3), .ZN(new_n392));
  INV_X1    g0192(.A(KEYINPUT3), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n393), .A2(G33), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n392), .A2(new_n394), .ZN(new_n395));
  NAND3_X1  g0195(.A1(new_n395), .A2(KEYINPUT7), .A3(new_n204), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n391), .A2(new_n396), .ZN(new_n397));
  AOI21_X1  g0197(.A(new_n389), .B1(new_n397), .B2(G68), .ZN(new_n398));
  OAI21_X1  g0198(.A(new_n254), .B1(new_n398), .B2(KEYINPUT16), .ZN(new_n399));
  INV_X1    g0199(.A(KEYINPUT79), .ZN(new_n400));
  INV_X1    g0200(.A(KEYINPUT16), .ZN(new_n401));
  NOR2_X1   g0201(.A1(new_n389), .A2(new_n401), .ZN(new_n402));
  AND3_X1   g0202(.A1(new_n264), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n403));
  INV_X1    g0203(.A(KEYINPUT78), .ZN(new_n404));
  AOI21_X1  g0204(.A(new_n403), .B1(new_n284), .B2(new_n404), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n390), .B1(new_n405), .B2(new_n204), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n392), .A2(new_n394), .A3(new_n404), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n264), .A2(KEYINPUT78), .A3(KEYINPUT3), .ZN(new_n408));
  NAND4_X1  g0208(.A1(new_n407), .A2(new_n390), .A3(new_n204), .A4(new_n408), .ZN(new_n409));
  NAND2_X1  g0209(.A1(new_n409), .A2(G68), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n400), .B(new_n402), .C1(new_n406), .C2(new_n410), .ZN(new_n411));
  OAI21_X1  g0211(.A(new_n402), .B1(new_n406), .B2(new_n410), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n412), .A2(KEYINPUT79), .ZN(new_n413));
  AOI21_X1  g0213(.A(new_n399), .B1(new_n411), .B2(new_n413), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n263), .B1(new_n203), .B2(G20), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n261), .A2(new_n415), .B1(new_n263), .B2(new_n260), .ZN(new_n416));
  INV_X1    g0216(.A(new_n416), .ZN(new_n417));
  OAI21_X1  g0217(.A(KEYINPUT80), .B1(new_n414), .B2(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(new_n254), .ZN(new_n419));
  AOI21_X1  g0219(.A(KEYINPUT7), .B1(new_n395), .B2(new_n204), .ZN(new_n420));
  AOI211_X1 g0220(.A(new_n390), .B(G20), .C1(new_n392), .C2(new_n394), .ZN(new_n421));
  OAI21_X1  g0221(.A(G68), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n389), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  AOI21_X1  g0224(.A(new_n419), .B1(new_n424), .B2(new_n401), .ZN(new_n425));
  INV_X1    g0225(.A(new_n411), .ZN(new_n426));
  NAND3_X1  g0226(.A1(new_n407), .A2(new_n204), .A3(new_n408), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n427), .A2(KEYINPUT7), .ZN(new_n428));
  NAND3_X1  g0228(.A1(new_n428), .A2(G68), .A3(new_n409), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n400), .B1(new_n429), .B2(new_n402), .ZN(new_n430));
  OAI21_X1  g0230(.A(new_n425), .B1(new_n426), .B2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  NAND3_X1  g0232(.A1(new_n431), .A2(new_n432), .A3(new_n416), .ZN(new_n433));
  OR2_X1    g0233(.A1(G223), .A2(G1698), .ZN(new_n434));
  OAI21_X1  g0234(.A(new_n434), .B1(G226), .B2(new_n286), .ZN(new_n435));
  AOI21_X1  g0235(.A(new_n435), .B1(new_n408), .B2(new_n407), .ZN(new_n436));
  INV_X1    g0236(.A(G87), .ZN(new_n437));
  NOR2_X1   g0237(.A1(new_n264), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n277), .B1(new_n436), .B2(new_n438), .ZN(new_n439));
  AOI21_X1  g0239(.A(new_n280), .B1(G232), .B2(new_n282), .ZN(new_n440));
  AND3_X1   g0240(.A1(new_n439), .A2(new_n440), .A3(G179), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n324), .B1(new_n439), .B2(new_n440), .ZN(new_n442));
  NOR2_X1   g0242(.A1(new_n441), .A2(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(new_n443), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n418), .A2(new_n433), .A3(new_n444), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n445), .A2(KEYINPUT18), .ZN(new_n446));
  AOI21_X1  g0246(.A(new_n351), .B1(new_n439), .B2(new_n440), .ZN(new_n447));
  AND2_X1   g0247(.A1(new_n439), .A2(new_n440), .ZN(new_n448));
  AND2_X1   g0248(.A1(KEYINPUT81), .A2(G190), .ZN(new_n449));
  NOR2_X1   g0249(.A1(KEYINPUT81), .A2(G190), .ZN(new_n450));
  NOR2_X1   g0250(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  INV_X1    g0251(.A(new_n451), .ZN(new_n452));
  AOI21_X1  g0252(.A(new_n447), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  NAND3_X1  g0253(.A1(new_n431), .A2(new_n453), .A3(new_n416), .ZN(new_n454));
  XNOR2_X1  g0254(.A(new_n454), .B(KEYINPUT17), .ZN(new_n455));
  INV_X1    g0255(.A(KEYINPUT18), .ZN(new_n456));
  NAND4_X1  g0256(.A1(new_n418), .A2(new_n456), .A3(new_n433), .A4(new_n444), .ZN(new_n457));
  NAND3_X1  g0257(.A1(new_n446), .A2(new_n455), .A3(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n385), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g0260(.A1(G33), .A2(G283), .ZN(new_n461));
  INV_X1    g0261(.A(G97), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n461), .B(new_n204), .C1(G33), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n204), .A2(G116), .ZN(new_n464));
  INV_X1    g0264(.A(new_n464), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n465), .A3(new_n254), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT20), .ZN(new_n467));
  OAI21_X1  g0267(.A(KEYINPUT86), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n464), .B1(new_n222), .B2(new_n253), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT86), .ZN(new_n470));
  NAND4_X1  g0270(.A1(new_n469), .A2(new_n470), .A3(new_n463), .A4(KEYINPUT20), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NAND3_X1  g0272(.A1(new_n468), .A2(new_n471), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n203), .A2(G33), .ZN(new_n474));
  INV_X1    g0274(.A(new_n474), .ZN(new_n475));
  INV_X1    g0275(.A(G116), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n259), .A2(G1), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n307), .A2(new_n477), .B1(new_n478), .B2(new_n464), .ZN(new_n479));
  NAND2_X1  g0279(.A1(new_n473), .A2(new_n479), .ZN(new_n480));
  INV_X1    g0280(.A(G41), .ZN(new_n481));
  OAI211_X1 g0281(.A(new_n203), .B(G45), .C1(new_n481), .C2(KEYINPUT5), .ZN(new_n482));
  INV_X1    g0282(.A(KEYINPUT83), .ZN(new_n483));
  AOI22_X1  g0283(.A1(new_n482), .A2(new_n483), .B1(KEYINPUT5), .B2(new_n481), .ZN(new_n484));
  INV_X1    g0284(.A(G45), .ZN(new_n485));
  NOR2_X1   g0285(.A1(new_n485), .A2(G1), .ZN(new_n486));
  OAI211_X1 g0286(.A(new_n486), .B(KEYINPUT83), .C1(KEYINPUT5), .C2(new_n481), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n484), .A2(new_n487), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n488), .A2(G270), .A3(new_n339), .ZN(new_n489));
  INV_X1    g0289(.A(G264), .ZN(new_n490));
  NAND2_X1  g0290(.A1(new_n490), .A2(G1698), .ZN(new_n491));
  OAI21_X1  g0291(.A(new_n491), .B1(G257), .B2(G1698), .ZN(new_n492));
  AOI21_X1  g0292(.A(new_n492), .B1(new_n408), .B2(new_n407), .ZN(new_n493));
  INV_X1    g0293(.A(G303), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n284), .A2(new_n494), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n277), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND3_X1  g0296(.A1(new_n484), .A2(new_n336), .A3(new_n487), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n489), .A2(new_n496), .A3(new_n497), .ZN(new_n498));
  NAND4_X1  g0298(.A1(new_n480), .A2(new_n498), .A3(KEYINPUT21), .A4(G169), .ZN(new_n499));
  AND2_X1   g0299(.A1(new_n484), .A2(new_n487), .ZN(new_n500));
  AOI21_X1  g0300(.A(new_n277), .B1(new_n484), .B2(new_n487), .ZN(new_n501));
  AOI22_X1  g0301(.A1(new_n336), .A2(new_n500), .B1(new_n501), .B2(G270), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n480), .A2(new_n502), .A3(G179), .A4(new_n496), .ZN(new_n503));
  AND2_X1   g0303(.A1(new_n499), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n480), .A2(new_n498), .A3(G169), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT21), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n498), .A2(G200), .ZN(new_n508));
  INV_X1    g0308(.A(new_n480), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n508), .B(new_n509), .C1(new_n451), .C2(new_n498), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n504), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n511), .A2(KEYINPUT87), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT87), .ZN(new_n513));
  NAND4_X1  g0313(.A1(new_n504), .A2(new_n513), .A3(new_n507), .A4(new_n510), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(G33), .A2(G116), .ZN(new_n516));
  INV_X1    g0316(.A(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n208), .B1(new_n407), .B2(new_n408), .ZN(new_n518));
  AOI21_X1  g0318(.A(new_n517), .B1(new_n518), .B2(G1698), .ZN(new_n519));
  NAND2_X1  g0319(.A1(new_n407), .A2(new_n408), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n520), .A2(G238), .A3(new_n286), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n339), .B1(new_n519), .B2(new_n521), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n486), .A2(new_n278), .ZN(new_n523));
  INV_X1    g0323(.A(G250), .ZN(new_n524));
  OAI21_X1  g0324(.A(new_n524), .B1(new_n485), .B2(G1), .ZN(new_n525));
  NAND3_X1  g0325(.A1(new_n339), .A2(new_n523), .A3(new_n525), .ZN(new_n526));
  INV_X1    g0326(.A(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(G200), .B1(new_n522), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n520), .A2(G244), .A3(G1698), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n521), .A2(new_n529), .A3(new_n516), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(new_n277), .ZN(new_n531));
  NAND3_X1  g0331(.A1(new_n531), .A2(G190), .A3(new_n526), .ZN(new_n532));
  AOI21_X1  g0332(.A(KEYINPUT19), .B1(new_n265), .B2(G97), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n437), .A2(new_n462), .A3(new_n318), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n534), .A2(KEYINPUT85), .ZN(new_n535));
  INV_X1    g0335(.A(KEYINPUT85), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n536), .A2(new_n437), .A3(new_n462), .A4(new_n318), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n535), .A2(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT19), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n539), .B1(new_n342), .B2(new_n204), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n533), .B1(new_n538), .B2(new_n540), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n520), .A2(new_n204), .A3(G68), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n419), .B1(new_n541), .B2(new_n542), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n301), .A2(new_n274), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n274), .A2(new_n255), .A3(new_n257), .A4(new_n474), .ZN(new_n545));
  NOR2_X1   g0345(.A1(new_n545), .A2(new_n437), .ZN(new_n546));
  NOR3_X1   g0346(.A1(new_n543), .A2(new_n544), .A3(new_n546), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n528), .A2(new_n532), .A3(new_n547), .ZN(new_n548));
  INV_X1    g0348(.A(new_n548), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n545), .A2(new_n300), .ZN(new_n550));
  NOR3_X1   g0350(.A1(new_n543), .A2(new_n544), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g0351(.A(G169), .B1(new_n522), .B2(new_n527), .ZN(new_n552));
  NAND3_X1  g0352(.A1(new_n531), .A2(G179), .A3(new_n526), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  INV_X1    g0354(.A(KEYINPUT84), .ZN(new_n555));
  AOI21_X1  g0355(.A(new_n551), .B1(new_n554), .B2(new_n555), .ZN(new_n556));
  NAND3_X1  g0356(.A1(new_n552), .A2(new_n553), .A3(KEYINPUT84), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n549), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n260), .A2(new_n318), .ZN(new_n559));
  INV_X1    g0359(.A(KEYINPUT25), .ZN(new_n560));
  XNOR2_X1  g0360(.A(new_n559), .B(new_n560), .ZN(new_n561));
  OAI21_X1  g0361(.A(new_n561), .B1(new_n318), .B2(new_n545), .ZN(new_n562));
  NAND2_X1  g0362(.A1(KEYINPUT22), .A2(G87), .ZN(new_n563));
  AOI211_X1 g0363(.A(G20), .B(new_n563), .C1(new_n407), .C2(new_n408), .ZN(new_n564));
  NOR2_X1   g0364(.A1(new_n437), .A2(G20), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n565), .A2(new_n392), .A3(new_n394), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT22), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g0368(.A(KEYINPUT23), .ZN(new_n569));
  OAI21_X1  g0369(.A(new_n569), .B1(new_n204), .B2(G107), .ZN(new_n570));
  NAND3_X1  g0370(.A1(new_n318), .A2(KEYINPUT23), .A3(G20), .ZN(new_n571));
  AOI22_X1  g0371(.A1(new_n570), .A2(new_n571), .B1(new_n517), .B2(new_n204), .ZN(new_n572));
  NAND2_X1  g0372(.A1(new_n568), .A2(new_n572), .ZN(new_n573));
  OAI21_X1  g0373(.A(KEYINPUT24), .B1(new_n564), .B2(new_n573), .ZN(new_n574));
  AOI21_X1  g0374(.A(KEYINPUT22), .B1(new_n284), .B2(new_n565), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n570), .A2(new_n571), .ZN(new_n576));
  NAND2_X1  g0376(.A1(new_n517), .A2(new_n204), .ZN(new_n577));
  NAND2_X1  g0377(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n575), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n563), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n520), .A2(new_n204), .A3(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT24), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n579), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n574), .A2(new_n583), .ZN(new_n584));
  AOI21_X1  g0384(.A(new_n562), .B1(new_n584), .B2(new_n254), .ZN(new_n585));
  INV_X1    g0385(.A(G257), .ZN(new_n586));
  NOR2_X1   g0386(.A1(new_n586), .A2(new_n286), .ZN(new_n587));
  INV_X1    g0387(.A(new_n587), .ZN(new_n588));
  INV_X1    g0388(.A(G294), .ZN(new_n589));
  OAI22_X1  g0389(.A1(new_n405), .A2(new_n588), .B1(new_n264), .B2(new_n589), .ZN(new_n590));
  AOI211_X1 g0390(.A(new_n524), .B(G1698), .C1(new_n407), .C2(new_n408), .ZN(new_n591));
  OAI21_X1  g0391(.A(new_n277), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  AOI211_X1 g0392(.A(new_n490), .B(new_n277), .C1(new_n484), .C2(new_n487), .ZN(new_n593));
  INV_X1    g0393(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n592), .A2(new_n594), .A3(new_n497), .ZN(new_n595));
  NAND2_X1  g0395(.A1(new_n595), .A2(G169), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n264), .A2(new_n589), .ZN(new_n597));
  AOI21_X1  g0397(.A(new_n597), .B1(new_n520), .B2(new_n587), .ZN(new_n598));
  NAND3_X1  g0398(.A1(new_n520), .A2(G250), .A3(new_n286), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n593), .B1(new_n600), .B2(new_n277), .ZN(new_n601));
  NAND3_X1  g0401(.A1(new_n601), .A2(G179), .A3(new_n497), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n596), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n585), .B1(new_n603), .B2(KEYINPUT88), .ZN(new_n604));
  AOI21_X1  g0404(.A(new_n324), .B1(new_n601), .B2(new_n497), .ZN(new_n605));
  AOI21_X1  g0405(.A(new_n339), .B1(new_n598), .B2(new_n599), .ZN(new_n606));
  INV_X1    g0406(.A(new_n497), .ZN(new_n607));
  NOR4_X1   g0407(.A1(new_n606), .A2(new_n593), .A3(new_n607), .A4(new_n331), .ZN(new_n608));
  OR3_X1    g0408(.A1(new_n605), .A2(new_n608), .A3(KEYINPUT88), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n604), .A2(new_n609), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n595), .A2(G200), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n601), .A2(G190), .A3(new_n497), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n611), .A2(new_n585), .A3(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n269), .A2(new_n308), .ZN(new_n614));
  INV_X1    g0414(.A(KEYINPUT82), .ZN(new_n615));
  NOR2_X1   g0415(.A1(new_n615), .A2(KEYINPUT6), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT6), .ZN(new_n617));
  NOR2_X1   g0417(.A1(new_n617), .A2(KEYINPUT82), .ZN(new_n618));
  NOR2_X1   g0418(.A1(G97), .A2(G107), .ZN(new_n619));
  AND2_X1   g0419(.A1(G97), .A2(G107), .ZN(new_n620));
  OAI22_X1  g0420(.A1(new_n616), .A2(new_n618), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n617), .A2(KEYINPUT82), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n615), .A2(KEYINPUT6), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n622), .A2(new_n623), .A3(G97), .A4(new_n318), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n621), .A2(new_n624), .ZN(new_n625));
  AOI21_X1  g0425(.A(new_n614), .B1(new_n625), .B2(G20), .ZN(new_n626));
  OAI21_X1  g0426(.A(G107), .B1(new_n420), .B2(new_n421), .ZN(new_n627));
  AOI21_X1  g0427(.A(new_n419), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  NOR2_X1   g0428(.A1(new_n545), .A2(new_n462), .ZN(new_n629));
  NOR2_X1   g0429(.A1(new_n274), .A2(G97), .ZN(new_n630));
  NOR3_X1   g0430(.A1(new_n628), .A2(new_n629), .A3(new_n630), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n520), .A2(G244), .A3(new_n286), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT4), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  NAND4_X1  g0434(.A1(new_n284), .A2(KEYINPUT4), .A3(G244), .A4(new_n286), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n284), .A2(G250), .A3(G1698), .ZN(new_n636));
  NAND3_X1  g0436(.A1(new_n635), .A2(new_n461), .A3(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n637), .ZN(new_n638));
  AOI21_X1  g0438(.A(new_n339), .B1(new_n634), .B2(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n501), .A2(G257), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n640), .A2(new_n497), .ZN(new_n641));
  OAI21_X1  g0441(.A(G200), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  AOI22_X1  g0442(.A1(new_n336), .A2(new_n500), .B1(new_n501), .B2(G257), .ZN(new_n643));
  AOI21_X1  g0443(.A(KEYINPUT4), .B1(new_n518), .B2(new_n286), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n277), .B1(new_n644), .B2(new_n637), .ZN(new_n645));
  NAND3_X1  g0445(.A1(new_n643), .A2(new_n645), .A3(G190), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n631), .A2(new_n642), .A3(new_n646), .ZN(new_n647));
  OAI21_X1  g0447(.A(new_n324), .B1(new_n639), .B2(new_n641), .ZN(new_n648));
  INV_X1    g0448(.A(new_n629), .ZN(new_n649));
  INV_X1    g0449(.A(new_n630), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n318), .B1(new_n391), .B2(new_n396), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n204), .B1(new_n621), .B2(new_n624), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(new_n652), .A3(new_n614), .ZN(new_n653));
  OAI211_X1 g0453(.A(new_n649), .B(new_n650), .C1(new_n653), .C2(new_n419), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n643), .A2(new_n645), .A3(new_n331), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n648), .A2(new_n654), .A3(new_n655), .ZN(new_n656));
  AND3_X1   g0456(.A1(new_n613), .A2(new_n647), .A3(new_n656), .ZN(new_n657));
  NAND4_X1  g0457(.A1(new_n515), .A2(new_n558), .A3(new_n610), .A4(new_n657), .ZN(new_n658));
  NOR2_X1   g0458(.A1(new_n460), .A2(new_n658), .ZN(G372));
  AOI21_X1  g0459(.A(new_n324), .B1(new_n531), .B2(new_n526), .ZN(new_n660));
  AOI211_X1 g0460(.A(new_n331), .B(new_n527), .C1(new_n530), .C2(new_n277), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n555), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g0462(.A(new_n551), .ZN(new_n663));
  NAND3_X1  g0463(.A1(new_n662), .A2(new_n557), .A3(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(new_n656), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(new_n548), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n666), .A2(KEYINPUT26), .ZN(new_n667));
  NOR3_X1   g0467(.A1(new_n564), .A2(new_n573), .A3(KEYINPUT24), .ZN(new_n668));
  AOI21_X1  g0468(.A(new_n582), .B1(new_n579), .B2(new_n581), .ZN(new_n669));
  OAI21_X1  g0469(.A(new_n254), .B1(new_n668), .B2(new_n669), .ZN(new_n670));
  INV_X1    g0470(.A(new_n562), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g0472(.A(new_n672), .B1(new_n605), .B2(new_n608), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n673), .A2(new_n504), .A3(new_n507), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n554), .A2(new_n663), .ZN(new_n675));
  INV_X1    g0475(.A(KEYINPUT89), .ZN(new_n676));
  AOI21_X1  g0476(.A(new_n351), .B1(new_n531), .B2(new_n526), .ZN(new_n677));
  INV_X1    g0477(.A(new_n544), .ZN(new_n678));
  INV_X1    g0478(.A(new_n546), .ZN(new_n679));
  AND2_X1   g0479(.A1(new_n541), .A2(new_n542), .ZN(new_n680));
  OAI211_X1 g0480(.A(new_n678), .B(new_n679), .C1(new_n680), .C2(new_n419), .ZN(new_n681));
  OAI21_X1  g0481(.A(new_n676), .B1(new_n677), .B2(new_n681), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n528), .A2(KEYINPUT89), .A3(new_n547), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n682), .A2(new_n532), .A3(new_n683), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n657), .A2(new_n674), .A3(new_n675), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT26), .ZN(new_n686));
  NAND4_X1  g0486(.A1(new_n684), .A2(new_n686), .A3(new_n665), .A4(new_n675), .ZN(new_n687));
  NAND4_X1  g0487(.A1(new_n667), .A2(new_n685), .A3(new_n675), .A4(new_n687), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n459), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n333), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT90), .ZN(new_n691));
  OR2_X1    g0491(.A1(new_n296), .A2(new_n691), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n296), .A2(new_n691), .ZN(new_n693));
  AND2_X1   g0493(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n443), .B1(new_n431), .B2(new_n416), .ZN(new_n695));
  XNOR2_X1  g0495(.A(new_n695), .B(KEYINPUT18), .ZN(new_n696));
  NOR2_X1   g0496(.A1(new_n370), .A2(new_n326), .ZN(new_n697));
  AOI21_X1  g0497(.A(new_n697), .B1(new_n383), .B2(new_n368), .ZN(new_n698));
  INV_X1    g0498(.A(new_n455), .ZN(new_n699));
  OAI21_X1  g0499(.A(new_n696), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n690), .B1(new_n694), .B2(new_n700), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n689), .A2(new_n701), .ZN(G369));
  NAND2_X1  g0502(.A1(new_n478), .A2(new_n204), .ZN(new_n703));
  OR2_X1    g0503(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n703), .A2(KEYINPUT27), .ZN(new_n705));
  NAND3_X1  g0505(.A1(new_n704), .A2(G213), .A3(new_n705), .ZN(new_n706));
  INV_X1    g0506(.A(G343), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n509), .A2(new_n709), .ZN(new_n710));
  AOI21_X1  g0510(.A(new_n710), .B1(new_n512), .B2(new_n514), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n504), .A2(new_n507), .ZN(new_n712));
  AND2_X1   g0512(.A1(new_n712), .A2(new_n710), .ZN(new_n713));
  OAI21_X1  g0513(.A(G330), .B1(new_n711), .B2(new_n713), .ZN(new_n714));
  NOR2_X1   g0514(.A1(new_n610), .A2(new_n709), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n672), .A2(new_n708), .ZN(new_n716));
  NAND2_X1  g0516(.A1(new_n613), .A2(new_n716), .ZN(new_n717));
  AOI21_X1  g0517(.A(new_n717), .B1(new_n609), .B2(new_n604), .ZN(new_n718));
  NOR2_X1   g0518(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(new_n712), .A3(new_n709), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n603), .A2(new_n672), .A3(new_n709), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n722), .A2(new_n723), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n721), .A2(new_n725), .ZN(G399));
  INV_X1    g0526(.A(new_n219), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n727), .A2(G41), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n538), .A2(G116), .ZN(new_n730));
  NAND3_X1  g0530(.A1(new_n729), .A2(G1), .A3(new_n730), .ZN(new_n731));
  OAI21_X1  g0531(.A(new_n731), .B1(new_n228), .B2(new_n729), .ZN(new_n732));
  XNOR2_X1  g0532(.A(new_n732), .B(KEYINPUT91), .ZN(new_n733));
  XNOR2_X1  g0533(.A(new_n733), .B(KEYINPUT28), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n688), .A2(new_n709), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n735), .A2(KEYINPUT29), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n639), .A2(new_n641), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n498), .A2(new_n331), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n522), .A2(new_n527), .ZN(new_n740));
  NAND4_X1  g0540(.A1(new_n738), .A2(new_n739), .A3(new_n740), .A4(new_n601), .ZN(new_n741));
  INV_X1    g0541(.A(KEYINPUT30), .ZN(new_n742));
  XNOR2_X1  g0542(.A(new_n741), .B(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n595), .B1(new_n639), .B2(new_n641), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n498), .A2(new_n331), .ZN(new_n745));
  OR3_X1    g0545(.A1(new_n740), .A2(new_n745), .A3(KEYINPUT92), .ZN(new_n746));
  OAI21_X1  g0546(.A(KEYINPUT92), .B1(new_n740), .B2(new_n745), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n744), .B1(new_n746), .B2(new_n747), .ZN(new_n748));
  OAI21_X1  g0548(.A(new_n708), .B1(new_n743), .B2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(KEYINPUT31), .ZN(new_n750));
  NAND2_X1  g0550(.A1(new_n749), .A2(new_n750), .ZN(new_n751));
  OAI211_X1 g0551(.A(KEYINPUT31), .B(new_n708), .C1(new_n743), .C2(new_n748), .ZN(new_n752));
  OAI211_X1 g0552(.A(new_n751), .B(new_n752), .C1(new_n658), .C2(new_n708), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G330), .ZN(new_n754));
  AOI21_X1  g0554(.A(KEYINPUT26), .B1(new_n558), .B2(new_n665), .ZN(new_n755));
  AND4_X1   g0555(.A1(KEYINPUT26), .A2(new_n684), .A3(new_n665), .A4(new_n675), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n657), .A2(new_n675), .A3(new_n684), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n712), .B1(new_n604), .B2(new_n609), .ZN(new_n759));
  OAI21_X1  g0559(.A(new_n675), .B1(new_n758), .B2(new_n759), .ZN(new_n760));
  OAI21_X1  g0560(.A(new_n709), .B1(new_n757), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT29), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n737), .A2(new_n754), .A3(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n734), .B1(new_n764), .B2(G1), .ZN(G364));
  NOR2_X1   g0565(.A1(new_n259), .A2(G20), .ZN(new_n766));
  AOI21_X1  g0566(.A(new_n203), .B1(new_n766), .B2(G45), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NOR2_X1   g0568(.A1(new_n728), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR2_X1   g0570(.A1(new_n711), .A2(new_n713), .ZN(new_n771));
  NOR2_X1   g0571(.A1(G13), .A2(G33), .ZN(new_n772));
  INV_X1    g0572(.A(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n773), .A2(G20), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n771), .A2(new_n774), .ZN(new_n775));
  NOR2_X1   g0575(.A1(G179), .A2(G200), .ZN(new_n776));
  INV_X1    g0576(.A(new_n776), .ZN(new_n777));
  NOR3_X1   g0577(.A1(new_n777), .A2(new_n204), .A3(G190), .ZN(new_n778));
  INV_X1    g0578(.A(new_n778), .ZN(new_n779));
  XOR2_X1   g0579(.A(KEYINPUT95), .B(G159), .Z(new_n780));
  NOR2_X1   g0580(.A1(new_n779), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(KEYINPUT32), .ZN(new_n782));
  NOR2_X1   g0582(.A1(new_n204), .A2(new_n331), .ZN(new_n783));
  NAND2_X1  g0583(.A1(new_n783), .A2(new_n351), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n784), .A2(new_n451), .ZN(new_n785));
  INV_X1    g0585(.A(new_n785), .ZN(new_n786));
  OAI22_X1  g0586(.A1(new_n781), .A2(new_n782), .B1(new_n245), .B2(new_n786), .ZN(new_n787));
  AOI211_X1 g0587(.A(new_n395), .B(new_n787), .C1(new_n782), .C2(new_n781), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n783), .A2(G200), .ZN(new_n789));
  NOR2_X1   g0589(.A1(new_n789), .A2(new_n451), .ZN(new_n790));
  NOR2_X1   g0590(.A1(new_n784), .A2(G190), .ZN(new_n791));
  AOI22_X1  g0591(.A1(G50), .A2(new_n790), .B1(new_n791), .B2(new_n289), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n789), .A2(G190), .ZN(new_n793));
  INV_X1    g0593(.A(new_n793), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n788), .B(new_n792), .C1(new_n365), .C2(new_n794), .ZN(new_n795));
  NOR4_X1   g0595(.A1(new_n204), .A2(new_n292), .A3(new_n351), .A4(G179), .ZN(new_n796));
  INV_X1    g0596(.A(new_n796), .ZN(new_n797));
  OR2_X1    g0597(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n798));
  NAND2_X1  g0598(.A1(new_n797), .A2(KEYINPUT96), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n798), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(new_n801));
  NAND2_X1  g0601(.A1(new_n801), .A2(G87), .ZN(new_n802));
  NOR4_X1   g0602(.A1(new_n204), .A2(new_n351), .A3(G179), .A4(G190), .ZN(new_n803));
  XOR2_X1   g0603(.A(new_n803), .B(KEYINPUT97), .Z(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(G107), .ZN(new_n805));
  OAI21_X1  g0605(.A(G20), .B1(new_n777), .B2(new_n292), .ZN(new_n806));
  INV_X1    g0606(.A(KEYINPUT98), .ZN(new_n807));
  OR2_X1    g0607(.A1(new_n806), .A2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n806), .A2(new_n807), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(new_n810), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n811), .A2(G97), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n802), .A2(new_n805), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n791), .ZN(new_n814));
  INV_X1    g0614(.A(G311), .ZN(new_n815));
  NOR2_X1   g0615(.A1(new_n814), .A2(new_n815), .ZN(new_n816));
  AOI211_X1 g0616(.A(new_n284), .B(new_n816), .C1(G329), .C2(new_n778), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT33), .B(G317), .ZN(new_n818));
  XNOR2_X1  g0618(.A(KEYINPUT99), .B(G326), .ZN(new_n819));
  AOI22_X1  g0619(.A1(new_n793), .A2(new_n818), .B1(new_n790), .B2(new_n819), .ZN(new_n820));
  INV_X1    g0620(.A(G322), .ZN(new_n821));
  OAI211_X1 g0621(.A(new_n817), .B(new_n820), .C1(new_n821), .C2(new_n786), .ZN(new_n822));
  AOI22_X1  g0622(.A1(new_n801), .A2(G303), .B1(G283), .B2(new_n804), .ZN(new_n823));
  OAI21_X1  g0623(.A(new_n823), .B1(new_n589), .B2(new_n810), .ZN(new_n824));
  OAI22_X1  g0624(.A1(new_n795), .A2(new_n813), .B1(new_n822), .B2(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n324), .A2(KEYINPUT93), .ZN(new_n826));
  INV_X1    g0626(.A(new_n826), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n204), .B1(KEYINPUT93), .B2(new_n324), .ZN(new_n828));
  AOI21_X1  g0628(.A(new_n222), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n774), .ZN(new_n830));
  XNOR2_X1  g0630(.A(new_n830), .B(KEYINPUT94), .ZN(new_n831));
  INV_X1    g0631(.A(new_n831), .ZN(new_n832));
  NAND3_X1  g0632(.A1(new_n219), .A2(G355), .A3(new_n284), .ZN(new_n833));
  NOR2_X1   g0633(.A1(new_n727), .A2(new_n520), .ZN(new_n834));
  OAI21_X1  g0634(.A(new_n834), .B1(G45), .B2(new_n228), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n248), .A2(new_n485), .ZN(new_n836));
  OAI221_X1 g0636(.A(new_n833), .B1(G116), .B2(new_n219), .C1(new_n835), .C2(new_n836), .ZN(new_n837));
  AOI22_X1  g0637(.A1(new_n825), .A2(new_n829), .B1(new_n832), .B2(new_n837), .ZN(new_n838));
  AOI21_X1  g0638(.A(new_n770), .B1(new_n775), .B2(new_n838), .ZN(new_n839));
  OR3_X1    g0639(.A1(new_n711), .A2(G330), .A3(new_n713), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n769), .B1(new_n840), .B2(new_n714), .ZN(new_n841));
  NOR2_X1   g0641(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT100), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(G396));
  NOR2_X1   g0644(.A1(new_n326), .A2(new_n708), .ZN(new_n845));
  INV_X1    g0645(.A(new_n315), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n329), .B1(new_n846), .B2(new_n709), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n845), .B1(new_n326), .B2(new_n847), .ZN(new_n848));
  NAND3_X1  g0648(.A1(new_n688), .A2(new_n709), .A3(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n849), .A2(KEYINPUT102), .ZN(new_n850));
  INV_X1    g0650(.A(new_n848), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n735), .A2(new_n851), .ZN(new_n852));
  XNOR2_X1  g0652(.A(new_n850), .B(new_n852), .ZN(new_n853));
  AOI21_X1  g0653(.A(new_n769), .B1(new_n853), .B2(new_n754), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n853), .A2(new_n754), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT103), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  NOR3_X1   g0657(.A1(new_n853), .A2(KEYINPUT103), .A3(new_n754), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n854), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  NOR2_X1   g0659(.A1(new_n829), .A2(new_n772), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n770), .B1(new_n308), .B2(new_n860), .ZN(new_n861));
  INV_X1    g0661(.A(new_n829), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n804), .A2(G87), .ZN(new_n863));
  OAI211_X1 g0663(.A(new_n812), .B(new_n863), .C1(new_n318), .C2(new_n800), .ZN(new_n864));
  OAI221_X1 g0664(.A(new_n395), .B1(new_n779), .B2(new_n815), .C1(new_n814), .C2(new_n476), .ZN(new_n865));
  AOI22_X1  g0665(.A1(G303), .A2(new_n790), .B1(new_n793), .B2(G283), .ZN(new_n866));
  OAI21_X1  g0666(.A(new_n866), .B1(new_n589), .B2(new_n786), .ZN(new_n867));
  NOR3_X1   g0667(.A1(new_n864), .A2(new_n865), .A3(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n804), .A2(G68), .ZN(new_n869));
  OAI21_X1  g0669(.A(new_n869), .B1(new_n800), .B2(new_n271), .ZN(new_n870));
  XOR2_X1   g0670(.A(new_n870), .B(KEYINPUT101), .Z(new_n871));
  AOI22_X1  g0671(.A1(G143), .A2(new_n785), .B1(new_n793), .B2(G150), .ZN(new_n872));
  INV_X1    g0672(.A(G137), .ZN(new_n873));
  INV_X1    g0673(.A(new_n790), .ZN(new_n874));
  OAI221_X1 g0674(.A(new_n872), .B1(new_n873), .B2(new_n874), .C1(new_n814), .C2(new_n780), .ZN(new_n875));
  INV_X1    g0675(.A(KEYINPUT34), .ZN(new_n876));
  AND2_X1   g0676(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n875), .A2(new_n876), .ZN(new_n878));
  AOI21_X1  g0678(.A(new_n405), .B1(G132), .B2(new_n778), .ZN(new_n879));
  OAI21_X1  g0679(.A(new_n879), .B1(new_n810), .B2(new_n245), .ZN(new_n880));
  NOR3_X1   g0680(.A1(new_n877), .A2(new_n878), .A3(new_n880), .ZN(new_n881));
  AOI21_X1  g0681(.A(new_n868), .B1(new_n871), .B2(new_n881), .ZN(new_n882));
  OAI221_X1 g0682(.A(new_n861), .B1(new_n862), .B2(new_n882), .C1(new_n848), .C2(new_n773), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n859), .A2(new_n883), .ZN(G384));
  OR2_X1    g0684(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n625), .A2(KEYINPUT35), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n885), .A2(G116), .A3(new_n223), .A4(new_n886), .ZN(new_n887));
  XOR2_X1   g0687(.A(new_n887), .B(KEYINPUT36), .Z(new_n888));
  OR3_X1    g0688(.A1(new_n228), .A2(new_n207), .A3(new_n386), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n271), .A2(G68), .ZN(new_n890));
  AOI211_X1 g0690(.A(new_n203), .B(G13), .C1(new_n889), .C2(new_n890), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n888), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n737), .A2(new_n762), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n893), .A2(new_n459), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n701), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n895), .B(KEYINPUT106), .ZN(new_n896));
  INV_X1    g0696(.A(new_n706), .ZN(new_n897));
  OR2_X1    g0697(.A1(new_n696), .A2(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(new_n845), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n849), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n368), .A2(new_n708), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n384), .A2(new_n371), .A3(new_n901), .ZN(new_n902));
  OAI211_X1 g0702(.A(new_n368), .B(new_n708), .C1(new_n383), .C2(new_n370), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n900), .A2(new_n904), .ZN(new_n905));
  INV_X1    g0705(.A(KEYINPUT38), .ZN(new_n906));
  INV_X1    g0706(.A(new_n454), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n907), .A2(KEYINPUT37), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n418), .A2(new_n433), .A3(new_n897), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n908), .A2(new_n445), .A3(new_n909), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n413), .A2(new_n411), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n429), .A2(new_n423), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n912), .A2(new_n401), .B1(new_n255), .B2(new_n257), .ZN(new_n913));
  AOI21_X1  g0713(.A(new_n417), .B1(new_n911), .B2(new_n913), .ZN(new_n914));
  OAI21_X1  g0714(.A(new_n454), .B1(new_n914), .B2(new_n443), .ZN(new_n915));
  NOR2_X1   g0715(.A1(new_n914), .A2(new_n706), .ZN(new_n916));
  OAI21_X1  g0716(.A(KEYINPUT37), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  AOI221_X4 g0717(.A(new_n906), .B1(new_n910), .B2(new_n917), .C1(new_n458), .C2(new_n916), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n458), .A2(new_n916), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n910), .A2(new_n917), .ZN(new_n920));
  AOI21_X1  g0720(.A(KEYINPUT38), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NOR2_X1   g0721(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n898), .B1(new_n905), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g0723(.A(KEYINPUT39), .B1(new_n918), .B2(new_n921), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n924), .A2(KEYINPUT104), .ZN(new_n925));
  INV_X1    g0725(.A(KEYINPUT105), .ZN(new_n926));
  AND3_X1   g0726(.A1(new_n908), .A2(new_n445), .A3(new_n909), .ZN(new_n927));
  INV_X1    g0727(.A(KEYINPUT37), .ZN(new_n928));
  NOR2_X1   g0728(.A1(new_n907), .A2(new_n695), .ZN(new_n929));
  AOI21_X1  g0729(.A(new_n928), .B1(new_n929), .B2(new_n909), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n926), .B1(new_n927), .B2(new_n930), .ZN(new_n931));
  AND3_X1   g0731(.A1(new_n418), .A2(new_n433), .A3(new_n897), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n444), .B1(new_n414), .B2(new_n417), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n933), .A2(new_n454), .ZN(new_n934));
  OAI21_X1  g0734(.A(KEYINPUT37), .B1(new_n932), .B2(new_n934), .ZN(new_n935));
  NAND3_X1  g0735(.A1(new_n935), .A2(KEYINPUT105), .A3(new_n910), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n909), .B1(new_n696), .B2(new_n455), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND3_X1  g0738(.A1(new_n931), .A2(new_n936), .A3(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n939), .A2(new_n906), .ZN(new_n940));
  INV_X1    g0740(.A(new_n918), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT39), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n940), .A2(new_n941), .A3(new_n942), .ZN(new_n943));
  INV_X1    g0743(.A(KEYINPUT104), .ZN(new_n944));
  OAI211_X1 g0744(.A(new_n944), .B(KEYINPUT39), .C1(new_n918), .C2(new_n921), .ZN(new_n945));
  NAND3_X1  g0745(.A1(new_n925), .A2(new_n943), .A3(new_n945), .ZN(new_n946));
  NOR2_X1   g0746(.A1(new_n384), .A2(new_n708), .ZN(new_n947));
  AOI21_X1  g0747(.A(new_n923), .B1(new_n946), .B2(new_n947), .ZN(new_n948));
  INV_X1    g0748(.A(new_n948), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n896), .B(new_n949), .ZN(new_n950));
  INV_X1    g0750(.A(KEYINPUT107), .ZN(new_n951));
  NAND2_X1  g0751(.A1(new_n935), .A2(new_n910), .ZN(new_n952));
  AOI21_X1  g0752(.A(new_n937), .B1(new_n952), .B2(new_n926), .ZN(new_n953));
  AOI21_X1  g0753(.A(KEYINPUT38), .B1(new_n953), .B2(new_n936), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n951), .B1(new_n954), .B2(new_n918), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n904), .A2(new_n753), .A3(new_n848), .ZN(new_n956));
  INV_X1    g0756(.A(KEYINPUT40), .ZN(new_n957));
  NOR2_X1   g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n940), .A2(new_n941), .A3(KEYINPUT107), .ZN(new_n959));
  NAND3_X1  g0759(.A1(new_n955), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n957), .B1(new_n922), .B2(new_n956), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n459), .A2(new_n753), .ZN(new_n963));
  OAI21_X1  g0763(.A(G330), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  AOI21_X1  g0764(.A(new_n964), .B1(new_n962), .B2(new_n963), .ZN(new_n965));
  NAND2_X1  g0765(.A1(new_n950), .A2(new_n965), .ZN(new_n966));
  NOR2_X1   g0766(.A1(new_n950), .A2(new_n965), .ZN(new_n967));
  INV_X1    g0767(.A(KEYINPUT108), .ZN(new_n968));
  OAI221_X1 g0768(.A(new_n966), .B1(new_n203), .B2(new_n766), .C1(new_n967), .C2(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(new_n967), .ZN(new_n970));
  NOR2_X1   g0770(.A1(new_n970), .A2(KEYINPUT108), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n892), .B1(new_n969), .B2(new_n971), .ZN(G367));
  OAI21_X1  g0772(.A(new_n284), .B1(new_n779), .B2(new_n873), .ZN(new_n973));
  INV_X1    g0773(.A(new_n803), .ZN(new_n974));
  OAI22_X1  g0774(.A1(new_n786), .A2(new_n267), .B1(new_n207), .B2(new_n974), .ZN(new_n975));
  AOI211_X1 g0775(.A(new_n973), .B(new_n975), .C1(G143), .C2(new_n790), .ZN(new_n976));
  INV_X1    g0776(.A(new_n780), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n793), .A2(new_n977), .B1(new_n791), .B2(G50), .ZN(new_n978));
  XNOR2_X1  g0778(.A(new_n978), .B(KEYINPUT112), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n801), .A2(G58), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n811), .A2(G68), .ZN(new_n981));
  NAND4_X1  g0781(.A1(new_n976), .A2(new_n979), .A3(new_n980), .A4(new_n981), .ZN(new_n982));
  AOI22_X1  g0782(.A1(G303), .A2(new_n785), .B1(new_n790), .B2(G311), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT111), .Z(new_n984));
  INV_X1    g0784(.A(KEYINPUT46), .ZN(new_n985));
  OAI21_X1  g0785(.A(new_n985), .B1(new_n800), .B2(new_n476), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n801), .A2(KEYINPUT46), .A3(G116), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n984), .A2(new_n986), .A3(new_n987), .ZN(new_n988));
  INV_X1    g0788(.A(G283), .ZN(new_n989));
  OAI22_X1  g0789(.A1(new_n794), .A2(new_n589), .B1(new_n814), .B2(new_n989), .ZN(new_n990));
  AOI21_X1  g0790(.A(new_n990), .B1(G97), .B2(new_n803), .ZN(new_n991));
  AOI21_X1  g0791(.A(new_n520), .B1(G317), .B2(new_n778), .ZN(new_n992));
  OAI211_X1 g0792(.A(new_n991), .B(new_n992), .C1(new_n318), .C2(new_n810), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n982), .B1(new_n988), .B2(new_n993), .ZN(new_n994));
  XOR2_X1   g0794(.A(new_n994), .B(KEYINPUT47), .Z(new_n995));
  NOR2_X1   g0795(.A1(new_n995), .A2(new_n862), .ZN(new_n996));
  NAND2_X1  g0796(.A1(new_n235), .A2(new_n834), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n831), .B1(new_n727), .B2(new_n301), .ZN(new_n998));
  AOI211_X1 g0798(.A(new_n770), .B(new_n996), .C1(new_n997), .C2(new_n998), .ZN(new_n999));
  INV_X1    g0799(.A(new_n774), .ZN(new_n1000));
  NAND2_X1  g0800(.A1(new_n681), .A2(new_n708), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n684), .A2(new_n675), .A3(new_n1001), .ZN(new_n1002));
  OAI21_X1  g0802(.A(new_n1002), .B1(new_n675), .B2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g0803(.A(new_n999), .B1(new_n1000), .B2(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(new_n1004), .ZN(new_n1005));
  OAI211_X1 g0805(.A(new_n647), .B(new_n656), .C1(new_n631), .C2(new_n709), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n665), .A2(new_n708), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n725), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT45), .ZN(new_n1010));
  XNOR2_X1  g0810(.A(new_n1009), .B(new_n1010), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n1008), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n724), .A2(new_n1012), .ZN(new_n1013));
  XOR2_X1   g0813(.A(new_n1013), .B(KEYINPUT44), .Z(new_n1014));
  NAND2_X1  g0814(.A1(new_n1011), .A2(new_n1014), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1015), .A2(new_n720), .ZN(new_n1016));
  NAND3_X1  g0816(.A1(new_n1011), .A2(new_n1014), .A3(new_n721), .ZN(new_n1017));
  NAND2_X1  g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  INV_X1    g0818(.A(new_n712), .ZN(new_n1019));
  OAI21_X1  g0819(.A(new_n719), .B1(new_n1019), .B2(new_n708), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n722), .ZN(new_n1021));
  XNOR2_X1  g0821(.A(new_n1021), .B(new_n714), .ZN(new_n1022));
  OAI21_X1  g0822(.A(new_n764), .B1(new_n1018), .B2(new_n1022), .ZN(new_n1023));
  XOR2_X1   g0823(.A(new_n728), .B(KEYINPUT41), .Z(new_n1024));
  INV_X1    g0824(.A(new_n1024), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n768), .B1(new_n1023), .B2(new_n1025), .ZN(new_n1026));
  INV_X1    g0826(.A(new_n1026), .ZN(new_n1027));
  NOR2_X1   g0827(.A1(new_n722), .A2(new_n1012), .ZN(new_n1028));
  XNOR2_X1  g0828(.A(new_n1028), .B(KEYINPUT42), .ZN(new_n1029));
  XNOR2_X1  g0829(.A(new_n1008), .B(KEYINPUT109), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n656), .B1(new_n1030), .B2(new_n610), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n709), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  INV_X1    g0833(.A(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n1034), .A2(new_n1035), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT110), .ZN(new_n1037));
  NAND2_X1  g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g0838(.A1(new_n1034), .A2(KEYINPUT110), .A3(new_n1035), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  NOR2_X1   g0840(.A1(new_n721), .A2(new_n1030), .ZN(new_n1041));
  AND2_X1   g0841(.A1(new_n1003), .A2(KEYINPUT43), .ZN(new_n1042));
  OR3_X1    g0842(.A1(new_n1034), .A2(new_n1035), .A3(new_n1042), .ZN(new_n1043));
  AND3_X1   g0843(.A1(new_n1040), .A2(new_n1041), .A3(new_n1043), .ZN(new_n1044));
  AOI21_X1  g0844(.A(new_n1041), .B1(new_n1040), .B2(new_n1043), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n1044), .A2(new_n1045), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n1005), .B1(new_n1027), .B2(new_n1046), .ZN(new_n1047));
  INV_X1    g0847(.A(new_n1047), .ZN(G387));
  NOR2_X1   g0848(.A1(new_n1022), .A2(new_n763), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n1022), .A2(new_n763), .ZN(new_n1051));
  NAND3_X1  g0851(.A1(new_n1050), .A2(new_n728), .A3(new_n1051), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n730), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1053), .A2(new_n219), .A3(new_n284), .ZN(new_n1054));
  OAI21_X1  g0854(.A(new_n1054), .B1(G107), .B2(new_n219), .ZN(new_n1055));
  INV_X1    g0855(.A(new_n834), .ZN(new_n1056));
  AOI211_X1 g0856(.A(G45), .B(new_n1053), .C1(G68), .C2(G77), .ZN(new_n1057));
  NOR2_X1   g0857(.A1(new_n263), .A2(G50), .ZN(new_n1058));
  XNOR2_X1  g0858(.A(new_n1058), .B(KEYINPUT50), .ZN(new_n1059));
  AOI21_X1  g0859(.A(new_n1056), .B1(new_n1057), .B2(new_n1059), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT113), .ZN(new_n1061));
  OR2_X1    g0861(.A1(new_n1060), .A2(new_n1061), .ZN(new_n1062));
  AOI22_X1  g0862(.A1(new_n1060), .A2(new_n1061), .B1(G45), .B2(new_n242), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n1055), .B1(new_n1062), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n769), .B1(new_n1064), .B2(new_n831), .ZN(new_n1065));
  AOI22_X1  g0865(.A1(G317), .A2(new_n785), .B1(new_n791), .B2(G303), .ZN(new_n1066));
  OAI221_X1 g0866(.A(new_n1066), .B1(new_n815), .B2(new_n794), .C1(new_n821), .C2(new_n874), .ZN(new_n1067));
  INV_X1    g0867(.A(KEYINPUT48), .ZN(new_n1068));
  OR2_X1    g0868(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1070));
  AOI22_X1  g0870(.A1(new_n801), .A2(G294), .B1(new_n811), .B2(G283), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n1069), .A2(new_n1070), .A3(new_n1071), .ZN(new_n1072));
  INV_X1    g0872(.A(KEYINPUT49), .ZN(new_n1073));
  OR2_X1    g0873(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1075));
  NOR2_X1   g0875(.A1(new_n974), .A2(new_n476), .ZN(new_n1076));
  AOI211_X1 g0876(.A(new_n520), .B(new_n1076), .C1(new_n778), .C2(new_n819), .ZN(new_n1077));
  NAND3_X1  g0877(.A1(new_n1074), .A2(new_n1075), .A3(new_n1077), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(G50), .A2(new_n785), .B1(new_n791), .B2(G68), .ZN(new_n1079));
  INV_X1    g0879(.A(G159), .ZN(new_n1080));
  OAI221_X1 g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n874), .C1(new_n263), .C2(new_n794), .ZN(new_n1081));
  AOI211_X1 g0881(.A(new_n405), .B(new_n1081), .C1(G150), .C2(new_n778), .ZN(new_n1082));
  NAND2_X1  g0882(.A1(new_n804), .A2(G97), .ZN(new_n1083));
  NAND2_X1  g0883(.A1(new_n811), .A2(new_n301), .ZN(new_n1084));
  NOR2_X1   g0884(.A1(new_n800), .A2(new_n207), .ZN(new_n1085));
  INV_X1    g0885(.A(new_n1085), .ZN(new_n1086));
  NAND4_X1  g0886(.A1(new_n1082), .A2(new_n1083), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n862), .B1(new_n1078), .B2(new_n1087), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1065), .B(new_n1088), .C1(new_n719), .C2(new_n774), .ZN(new_n1089));
  INV_X1    g0889(.A(new_n1022), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n768), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1052), .A2(new_n1091), .ZN(G393));
  INV_X1    g0892(.A(new_n1018), .ZN(new_n1093));
  NOR2_X1   g0893(.A1(new_n1093), .A2(new_n1049), .ZN(new_n1094));
  INV_X1    g0894(.A(KEYINPUT115), .ZN(new_n1095));
  OAI21_X1  g0895(.A(new_n728), .B1(new_n1018), .B2(new_n1050), .ZN(new_n1096));
  OR3_X1    g0896(.A1(new_n1094), .A2(new_n1095), .A3(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1095), .B1(new_n1094), .B2(new_n1096), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1093), .A2(new_n768), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1030), .A2(new_n774), .ZN(new_n1101));
  OAI22_X1  g0901(.A1(new_n1056), .A2(new_n251), .B1(new_n462), .B2(new_n219), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n769), .B1(new_n1102), .B2(new_n831), .ZN(new_n1103));
  XNOR2_X1  g0903(.A(new_n1103), .B(KEYINPUT114), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(G150), .A2(new_n790), .B1(new_n785), .B2(G159), .ZN(new_n1105));
  AOI22_X1  g0905(.A1(new_n801), .A2(G68), .B1(KEYINPUT51), .B2(new_n1105), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n405), .B1(G143), .B2(new_n778), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n263), .ZN(new_n1108));
  AOI22_X1  g0908(.A1(G50), .A2(new_n793), .B1(new_n791), .B2(new_n1108), .ZN(new_n1109));
  AND3_X1   g0909(.A1(new_n863), .A2(new_n1107), .A3(new_n1109), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n811), .A2(G77), .ZN(new_n1111));
  OR2_X1    g0911(.A1(new_n1105), .A2(KEYINPUT51), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1106), .A2(new_n1110), .A3(new_n1111), .A4(new_n1112), .ZN(new_n1113));
  AOI22_X1  g0913(.A1(G311), .A2(new_n785), .B1(new_n790), .B2(G317), .ZN(new_n1114));
  NOR2_X1   g0914(.A1(new_n1114), .A2(KEYINPUT52), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n801), .B2(G283), .ZN(new_n1116));
  OAI221_X1 g0916(.A(new_n395), .B1(new_n779), .B2(new_n821), .C1(new_n814), .C2(new_n589), .ZN(new_n1117));
  AOI21_X1  g0917(.A(new_n1117), .B1(G303), .B2(new_n793), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n811), .A2(G116), .B1(KEYINPUT52), .B2(new_n1114), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n805), .A4(new_n1119), .ZN(new_n1120));
  AND2_X1   g0920(.A1(new_n1113), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g0921(.A(new_n1101), .B(new_n1104), .C1(new_n862), .C2(new_n1121), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1100), .A2(new_n1122), .ZN(new_n1123));
  INV_X1    g0923(.A(new_n1123), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n1099), .A2(new_n1124), .ZN(G390));
  NAND4_X1  g0925(.A1(new_n904), .A2(new_n753), .A3(G330), .A4(new_n848), .ZN(new_n1126));
  XNOR2_X1  g0926(.A(new_n1126), .B(KEYINPUT117), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n753), .A2(G330), .A3(new_n848), .ZN(new_n1128));
  INV_X1    g0928(.A(new_n904), .ZN(new_n1129));
  NAND2_X1  g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  NAND2_X1  g0930(.A1(new_n847), .A2(new_n326), .ZN(new_n1131));
  OAI211_X1 g0931(.A(new_n709), .B(new_n1131), .C1(new_n757), .C2(new_n760), .ZN(new_n1132));
  NAND4_X1  g0932(.A1(new_n1127), .A2(new_n899), .A3(new_n1130), .A4(new_n1132), .ZN(new_n1133));
  NAND2_X1  g0933(.A1(new_n1130), .A2(new_n1126), .ZN(new_n1134));
  NAND2_X1  g0934(.A1(new_n1134), .A2(new_n900), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n894), .B(new_n701), .C1(new_n460), .C2(new_n754), .ZN(new_n1137));
  INV_X1    g0937(.A(new_n1137), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n1136), .A2(new_n1138), .ZN(new_n1139));
  NAND2_X1  g0939(.A1(new_n1132), .A2(new_n899), .ZN(new_n1140));
  AOI21_X1  g0940(.A(new_n947), .B1(new_n1140), .B2(new_n904), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n955), .A2(new_n1141), .A3(new_n959), .ZN(new_n1142));
  INV_X1    g0942(.A(KEYINPUT116), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1142), .A2(new_n1143), .ZN(new_n1144));
  NAND4_X1  g0944(.A1(new_n955), .A2(new_n1141), .A3(new_n959), .A4(KEYINPUT116), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1144), .A2(new_n1145), .ZN(new_n1146));
  INV_X1    g0946(.A(new_n947), .ZN(new_n1147));
  NAND2_X1  g0947(.A1(new_n905), .A2(new_n1147), .ZN(new_n1148));
  NAND4_X1  g0948(.A1(new_n925), .A2(new_n1148), .A3(new_n943), .A4(new_n945), .ZN(new_n1149));
  AOI21_X1  g0949(.A(new_n1126), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1149), .A2(new_n1127), .ZN(new_n1151));
  AOI21_X1  g0951(.A(new_n1151), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1139), .B1(new_n1150), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1137), .B1(new_n1133), .B2(new_n1135), .ZN(new_n1154));
  AND2_X1   g0954(.A1(new_n1149), .A2(new_n1127), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1146), .A2(new_n1155), .ZN(new_n1156));
  AND4_X1   g0956(.A1(new_n925), .A2(new_n1148), .A3(new_n943), .A4(new_n945), .ZN(new_n1157));
  AOI21_X1  g0957(.A(new_n1157), .B1(new_n1144), .B2(new_n1145), .ZN(new_n1158));
  OAI211_X1 g0958(.A(new_n1154), .B(new_n1156), .C1(new_n1126), .C2(new_n1158), .ZN(new_n1159));
  AND3_X1   g0959(.A1(new_n1153), .A2(new_n728), .A3(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(new_n1160), .ZN(new_n1161));
  OR2_X1    g0961(.A1(new_n946), .A2(new_n773), .ZN(new_n1162));
  INV_X1    g0962(.A(new_n860), .ZN(new_n1163));
  OAI21_X1  g0963(.A(new_n769), .B1(new_n1108), .B2(new_n1163), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n801), .A2(G150), .ZN(new_n1165));
  XNOR2_X1  g0965(.A(new_n1165), .B(KEYINPUT53), .ZN(new_n1166));
  AND2_X1   g0966(.A1(new_n778), .A2(G125), .ZN(new_n1167));
  AOI211_X1 g0967(.A(new_n395), .B(new_n1167), .C1(G128), .C2(new_n790), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n811), .A2(G159), .ZN(new_n1169));
  AOI22_X1  g0969(.A1(G132), .A2(new_n785), .B1(new_n793), .B2(G137), .ZN(new_n1170));
  XOR2_X1   g0970(.A(KEYINPUT54), .B(G143), .Z(new_n1171));
  AOI22_X1  g0971(.A1(new_n791), .A2(new_n1171), .B1(G50), .B2(new_n803), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .A4(new_n1172), .ZN(new_n1173));
  AOI22_X1  g0973(.A1(G283), .A2(new_n790), .B1(new_n793), .B2(G107), .ZN(new_n1174));
  OAI21_X1  g0974(.A(new_n1174), .B1(new_n462), .B2(new_n814), .ZN(new_n1175));
  XOR2_X1   g0975(.A(new_n1175), .B(KEYINPUT118), .Z(new_n1176));
  OAI21_X1  g0976(.A(new_n395), .B1(new_n779), .B2(new_n589), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1177), .B1(new_n785), .B2(G116), .ZN(new_n1178));
  NAND4_X1  g0978(.A1(new_n802), .A2(new_n869), .A3(new_n1111), .A4(new_n1178), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n1166), .A2(new_n1173), .B1(new_n1176), .B2(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1164), .B1(new_n1180), .B2(new_n829), .ZN(new_n1181));
  AND2_X1   g0981(.A1(new_n1162), .A2(new_n1181), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1146), .A2(new_n1149), .ZN(new_n1183));
  INV_X1    g0983(.A(new_n1126), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1183), .A2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n767), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1186));
  AOI211_X1 g0986(.A(KEYINPUT119), .B(new_n1182), .C1(new_n1185), .C2(new_n1186), .ZN(new_n1187));
  INV_X1    g0987(.A(KEYINPUT119), .ZN(new_n1188));
  OAI211_X1 g0988(.A(new_n1156), .B(new_n768), .C1(new_n1126), .C2(new_n1158), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1182), .ZN(new_n1190));
  AOI21_X1  g0990(.A(new_n1188), .B1(new_n1189), .B2(new_n1190), .ZN(new_n1191));
  NOR3_X1   g0991(.A1(new_n1187), .A2(new_n1191), .A3(KEYINPUT120), .ZN(new_n1192));
  INV_X1    g0992(.A(KEYINPUT120), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1156), .A2(new_n768), .ZN(new_n1194));
  OAI21_X1  g0994(.A(new_n1190), .B1(new_n1194), .B2(new_n1150), .ZN(new_n1195));
  NAND2_X1  g0995(.A1(new_n1195), .A2(KEYINPUT119), .ZN(new_n1196));
  NAND3_X1  g0996(.A1(new_n1189), .A2(new_n1188), .A3(new_n1190), .ZN(new_n1197));
  AOI21_X1  g0997(.A(new_n1193), .B1(new_n1196), .B2(new_n1197), .ZN(new_n1198));
  OAI21_X1  g0998(.A(new_n1161), .B1(new_n1192), .B2(new_n1198), .ZN(G378));
  NAND3_X1  g0999(.A1(new_n692), .A2(new_n693), .A3(new_n333), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n275), .A2(new_n897), .ZN(new_n1201));
  INV_X1    g1001(.A(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1200), .A2(new_n1202), .ZN(new_n1203));
  NAND4_X1  g1003(.A1(new_n692), .A2(new_n693), .A3(new_n333), .A4(new_n1201), .ZN(new_n1204));
  NAND2_X1  g1004(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1205));
  XNOR2_X1  g1005(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n1206), .ZN(new_n1207));
  NAND2_X1  g1007(.A1(new_n1205), .A2(new_n1207), .ZN(new_n1208));
  NAND3_X1  g1008(.A1(new_n1203), .A2(new_n1204), .A3(new_n1206), .ZN(new_n1209));
  NAND2_X1  g1009(.A1(new_n1208), .A2(new_n1209), .ZN(new_n1210));
  NOR2_X1   g1010(.A1(new_n1210), .A2(new_n773), .ZN(new_n1211));
  NOR2_X1   g1011(.A1(new_n974), .A2(new_n245), .ZN(new_n1212));
  AOI21_X1  g1012(.A(new_n1212), .B1(G107), .B2(new_n785), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G116), .A2(new_n790), .B1(new_n791), .B2(new_n301), .ZN(new_n1214));
  NOR2_X1   g1014(.A1(new_n520), .A2(G41), .ZN(new_n1215));
  AOI22_X1  g1015(.A1(new_n793), .A2(G97), .B1(new_n778), .B2(G283), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1213), .A2(new_n1214), .A3(new_n1215), .A4(new_n1216), .ZN(new_n1217));
  AOI211_X1 g1017(.A(new_n1085), .B(new_n1217), .C1(G68), .C2(new_n811), .ZN(new_n1218));
  XOR2_X1   g1018(.A(new_n1218), .B(KEYINPUT58), .Z(new_n1219));
  NAND2_X1  g1019(.A1(new_n801), .A2(new_n1171), .ZN(new_n1220));
  NAND2_X1  g1020(.A1(new_n811), .A2(G150), .ZN(new_n1221));
  AOI22_X1  g1021(.A1(G128), .A2(new_n785), .B1(new_n793), .B2(G132), .ZN(new_n1222));
  AOI22_X1  g1022(.A1(G125), .A2(new_n790), .B1(new_n791), .B2(G137), .ZN(new_n1223));
  NAND4_X1  g1023(.A1(new_n1220), .A2(new_n1221), .A3(new_n1222), .A4(new_n1223), .ZN(new_n1224));
  NOR2_X1   g1024(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(KEYINPUT59), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n977), .A2(new_n803), .ZN(new_n1227));
  AOI211_X1 g1027(.A(G33), .B(G41), .C1(new_n778), .C2(G124), .ZN(new_n1228));
  NAND3_X1  g1028(.A1(new_n1226), .A2(new_n1227), .A3(new_n1228), .ZN(new_n1229));
  OAI21_X1  g1029(.A(new_n271), .B1(G33), .B2(G41), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n1219), .B1(new_n1225), .B2(new_n1229), .C1(new_n1215), .C2(new_n1230), .ZN(new_n1231));
  INV_X1    g1031(.A(KEYINPUT121), .ZN(new_n1232));
  AOI21_X1  g1032(.A(new_n862), .B1(new_n1231), .B2(new_n1232), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1233), .B1(new_n1232), .B2(new_n1231), .ZN(new_n1234));
  OAI211_X1 g1034(.A(new_n1234), .B(new_n769), .C1(G50), .C2(new_n1163), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1211), .A2(new_n1235), .ZN(new_n1236));
  INV_X1    g1036(.A(new_n1210), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n960), .A2(G330), .A3(new_n961), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1237), .A2(new_n1238), .ZN(new_n1239));
  NAND4_X1  g1039(.A1(new_n1210), .A2(new_n960), .A3(G330), .A4(new_n961), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND2_X1  g1041(.A1(new_n1241), .A2(new_n949), .ZN(new_n1242));
  NAND3_X1  g1042(.A1(new_n1239), .A2(new_n948), .A3(new_n1240), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1242), .A2(new_n1243), .ZN(new_n1244));
  AOI21_X1  g1044(.A(new_n1236), .B1(new_n1244), .B2(new_n768), .ZN(new_n1245));
  AOI22_X1  g1045(.A1(new_n1183), .A2(new_n1184), .B1(new_n1146), .B2(new_n1155), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1137), .B1(new_n1246), .B2(new_n1136), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1243), .ZN(new_n1248));
  AOI21_X1  g1048(.A(new_n948), .B1(new_n1239), .B2(new_n1240), .ZN(new_n1249));
  OAI21_X1  g1049(.A(KEYINPUT57), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  OAI21_X1  g1050(.A(new_n728), .B1(new_n1247), .B2(new_n1250), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(new_n1159), .A2(new_n1138), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT57), .B1(new_n1252), .B2(new_n1244), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n1245), .B1(new_n1251), .B2(new_n1253), .ZN(G375));
  NAND3_X1  g1054(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1139), .A2(new_n1025), .A3(new_n1255), .ZN(new_n1256));
  NAND2_X1  g1056(.A1(new_n1136), .A2(new_n768), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n769), .B1(G68), .B2(new_n1163), .ZN(new_n1258));
  XNOR2_X1  g1058(.A(new_n1258), .B(KEYINPUT122), .ZN(new_n1259));
  AOI22_X1  g1059(.A1(new_n801), .A2(G159), .B1(new_n811), .B2(G50), .ZN(new_n1260));
  OAI22_X1  g1060(.A1(new_n873), .A2(new_n786), .B1(new_n814), .B2(new_n267), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1261), .B1(G132), .B2(new_n790), .ZN(new_n1262));
  AOI21_X1  g1062(.A(new_n405), .B1(G128), .B2(new_n778), .ZN(new_n1263));
  AOI21_X1  g1063(.A(new_n1212), .B1(new_n793), .B2(new_n1171), .ZN(new_n1264));
  NAND4_X1  g1064(.A1(new_n1260), .A2(new_n1262), .A3(new_n1263), .A4(new_n1264), .ZN(new_n1265));
  OAI21_X1  g1065(.A(new_n1084), .B1(new_n989), .B2(new_n786), .ZN(new_n1266));
  XOR2_X1   g1066(.A(new_n1266), .B(KEYINPUT123), .Z(new_n1267));
  NAND2_X1  g1067(.A1(new_n801), .A2(G97), .ZN(new_n1268));
  NAND2_X1  g1068(.A1(new_n804), .A2(G77), .ZN(new_n1269));
  OAI21_X1  g1069(.A(new_n395), .B1(new_n779), .B2(new_n494), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1270), .B1(G107), .B2(new_n791), .ZN(new_n1271));
  AOI22_X1  g1071(.A1(G294), .A2(new_n790), .B1(new_n793), .B2(G116), .ZN(new_n1272));
  NAND4_X1  g1072(.A1(new_n1268), .A2(new_n1269), .A3(new_n1271), .A4(new_n1272), .ZN(new_n1273));
  OAI21_X1  g1073(.A(new_n1265), .B1(new_n1267), .B2(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1259), .B1(new_n1274), .B2(new_n829), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n1275), .B1(new_n904), .B2(new_n773), .ZN(new_n1276));
  NAND3_X1  g1076(.A1(new_n1256), .A2(new_n1257), .A3(new_n1276), .ZN(G381));
  INV_X1    g1077(.A(G384), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(G393), .A2(G396), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1047), .A2(new_n1278), .A3(new_n1279), .ZN(new_n1280));
  NOR3_X1   g1080(.A1(new_n1280), .A2(G390), .A3(G381), .ZN(new_n1281));
  INV_X1    g1081(.A(new_n1245), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1253), .ZN(new_n1283));
  INV_X1    g1083(.A(KEYINPUT57), .ZN(new_n1284));
  AOI21_X1  g1084(.A(new_n1284), .B1(new_n1242), .B2(new_n1243), .ZN(new_n1285));
  AOI21_X1  g1085(.A(new_n729), .B1(new_n1285), .B2(new_n1252), .ZN(new_n1286));
  AOI21_X1  g1086(.A(new_n1282), .B1(new_n1283), .B2(new_n1286), .ZN(new_n1287));
  NOR3_X1   g1087(.A1(new_n1160), .A2(new_n1187), .A3(new_n1191), .ZN(new_n1288));
  NAND3_X1  g1088(.A1(new_n1281), .A2(new_n1287), .A3(new_n1288), .ZN(G407));
  NAND2_X1  g1089(.A1(new_n707), .A2(G213), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1290), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1287), .A2(new_n1288), .A3(new_n1291), .ZN(new_n1292));
  NAND3_X1  g1092(.A1(G407), .A2(G213), .A3(new_n1292), .ZN(G409));
  NAND3_X1  g1093(.A1(new_n1252), .A2(new_n1025), .A3(new_n1244), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1294), .A2(new_n1245), .ZN(new_n1295));
  NAND2_X1  g1095(.A1(new_n1288), .A2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT120), .B1(new_n1187), .B2(new_n1191), .ZN(new_n1297));
  NAND3_X1  g1097(.A1(new_n1196), .A2(new_n1193), .A3(new_n1197), .ZN(new_n1298));
  AOI21_X1  g1098(.A(new_n1160), .B1(new_n1297), .B2(new_n1298), .ZN(new_n1299));
  OAI21_X1  g1099(.A(new_n1296), .B1(new_n1299), .B2(G375), .ZN(new_n1300));
  NAND4_X1  g1100(.A1(new_n1133), .A2(KEYINPUT60), .A3(new_n1135), .A4(new_n1137), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1301), .A2(new_n728), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1139), .A2(KEYINPUT60), .ZN(new_n1303));
  AOI21_X1  g1103(.A(new_n1302), .B1(new_n1303), .B2(new_n1255), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(G384), .A2(KEYINPUT124), .ZN(new_n1305));
  NAND2_X1  g1105(.A1(new_n1257), .A2(new_n1276), .ZN(new_n1306));
  OR3_X1    g1106(.A1(new_n1304), .A2(new_n1305), .A3(new_n1306), .ZN(new_n1307));
  INV_X1    g1107(.A(KEYINPUT124), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1278), .A2(new_n1308), .ZN(new_n1309));
  OAI22_X1  g1109(.A1(new_n1306), .A2(new_n1304), .B1(new_n1309), .B2(new_n1305), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1307), .A2(new_n1310), .ZN(new_n1311));
  INV_X1    g1111(.A(new_n1311), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1300), .A2(new_n1290), .A3(new_n1312), .ZN(new_n1313));
  NAND2_X1  g1113(.A1(new_n1313), .A2(KEYINPUT62), .ZN(new_n1314));
  INV_X1    g1114(.A(KEYINPUT61), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1291), .A2(G2897), .ZN(new_n1316));
  AND3_X1   g1116(.A1(new_n1307), .A2(new_n1310), .A3(new_n1316), .ZN(new_n1317));
  AOI21_X1  g1117(.A(new_n1316), .B1(new_n1307), .B2(new_n1310), .ZN(new_n1318));
  NOR2_X1   g1118(.A1(new_n1317), .A2(new_n1318), .ZN(new_n1319));
  AOI22_X1  g1119(.A1(G378), .A2(new_n1287), .B1(new_n1288), .B2(new_n1295), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n1319), .B1(new_n1320), .B2(new_n1291), .ZN(new_n1321));
  INV_X1    g1121(.A(KEYINPUT62), .ZN(new_n1322));
  NAND4_X1  g1122(.A1(new_n1300), .A2(new_n1322), .A3(new_n1290), .A4(new_n1312), .ZN(new_n1323));
  NAND4_X1  g1123(.A1(new_n1314), .A2(new_n1315), .A3(new_n1321), .A4(new_n1323), .ZN(new_n1324));
  AOI21_X1  g1124(.A(new_n843), .B1(new_n1052), .B2(new_n1091), .ZN(new_n1325));
  OAI21_X1  g1125(.A(KEYINPUT125), .B1(new_n1279), .B2(new_n1325), .ZN(new_n1326));
  INV_X1    g1126(.A(new_n1326), .ZN(new_n1327));
  NAND3_X1  g1127(.A1(G387), .A2(new_n1099), .A3(new_n1124), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(G390), .A2(new_n1047), .ZN(new_n1329));
  AOI21_X1  g1129(.A(new_n1327), .B1(new_n1328), .B2(new_n1329), .ZN(new_n1330));
  INV_X1    g1130(.A(new_n1330), .ZN(new_n1331));
  NOR3_X1   g1131(.A1(new_n1279), .A2(KEYINPUT125), .A3(new_n1325), .ZN(new_n1332));
  OR2_X1    g1132(.A1(new_n1327), .A2(new_n1332), .ZN(new_n1333));
  NAND3_X1  g1133(.A1(new_n1328), .A2(new_n1329), .A3(new_n1333), .ZN(new_n1334));
  AND3_X1   g1134(.A1(new_n1331), .A2(KEYINPUT127), .A3(new_n1334), .ZN(new_n1335));
  AOI21_X1  g1135(.A(KEYINPUT127), .B1(new_n1331), .B2(new_n1334), .ZN(new_n1336));
  NOR2_X1   g1136(.A1(new_n1335), .A2(new_n1336), .ZN(new_n1337));
  NAND2_X1  g1137(.A1(new_n1324), .A2(new_n1337), .ZN(new_n1338));
  AND3_X1   g1138(.A1(new_n1328), .A2(new_n1329), .A3(new_n1333), .ZN(new_n1339));
  NOR2_X1   g1139(.A1(new_n1339), .A2(new_n1330), .ZN(new_n1340));
  INV_X1    g1140(.A(KEYINPUT63), .ZN(new_n1341));
  AOI21_X1  g1141(.A(new_n1340), .B1(new_n1341), .B2(new_n1313), .ZN(new_n1342));
  NAND2_X1  g1142(.A1(G378), .A2(new_n1287), .ZN(new_n1343));
  AOI21_X1  g1143(.A(new_n1291), .B1(new_n1343), .B2(new_n1296), .ZN(new_n1344));
  INV_X1    g1144(.A(KEYINPUT126), .ZN(new_n1345));
  NAND4_X1  g1145(.A1(new_n1344), .A2(new_n1345), .A3(KEYINPUT63), .A4(new_n1312), .ZN(new_n1346));
  OAI21_X1  g1146(.A(KEYINPUT126), .B1(new_n1313), .B2(new_n1341), .ZN(new_n1347));
  NAND2_X1  g1147(.A1(new_n1300), .A2(new_n1290), .ZN(new_n1348));
  AOI21_X1  g1148(.A(KEYINPUT61), .B1(new_n1348), .B2(new_n1319), .ZN(new_n1349));
  NAND4_X1  g1149(.A1(new_n1342), .A2(new_n1346), .A3(new_n1347), .A4(new_n1349), .ZN(new_n1350));
  NAND2_X1  g1150(.A1(new_n1338), .A2(new_n1350), .ZN(G405));
  NAND2_X1  g1151(.A1(G375), .A2(new_n1288), .ZN(new_n1352));
  NAND2_X1  g1152(.A1(new_n1343), .A2(new_n1352), .ZN(new_n1353));
  NAND2_X1  g1153(.A1(new_n1353), .A2(new_n1312), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1343), .A2(new_n1311), .A3(new_n1352), .ZN(new_n1355));
  NAND2_X1  g1155(.A1(new_n1354), .A2(new_n1355), .ZN(new_n1356));
  XNOR2_X1  g1156(.A(new_n1356), .B(new_n1340), .ZN(G402));
endmodule


