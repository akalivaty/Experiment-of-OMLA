//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 0 1 1 1 1 1 0 0 1 0 0 1 1 0 1 0 1 0 0 1 1 0 0 1 1 1 1 0 1 0 0 1 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:55 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n756, new_n758, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n768, new_n769, new_n770, new_n771,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n792, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1004,
    new_n1005, new_n1006, new_n1007, new_n1008, new_n1009, new_n1011,
    new_n1012, new_n1013, new_n1014, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050;
  INV_X1    g000(.A(KEYINPUT87), .ZN(new_n187));
  INV_X1    g001(.A(KEYINPUT80), .ZN(new_n188));
  INV_X1    g002(.A(G104), .ZN(new_n189));
  OAI21_X1  g003(.A(KEYINPUT3), .B1(new_n189), .B2(G107), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  INV_X1    g005(.A(G107), .ZN(new_n192));
  NAND3_X1  g006(.A1(new_n191), .A2(new_n192), .A3(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n189), .A2(G107), .ZN(new_n194));
  NAND3_X1  g008(.A1(new_n190), .A2(new_n193), .A3(new_n194), .ZN(new_n195));
  AND2_X1   g009(.A1(new_n195), .A2(G101), .ZN(new_n196));
  INV_X1    g010(.A(G101), .ZN(new_n197));
  NAND4_X1  g011(.A1(new_n190), .A2(new_n193), .A3(new_n197), .A4(new_n194), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(KEYINPUT4), .ZN(new_n199));
  OAI21_X1  g013(.A(new_n188), .B1(new_n196), .B2(new_n199), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n195), .A2(G101), .ZN(new_n201));
  NAND4_X1  g015(.A1(new_n201), .A2(KEYINPUT80), .A3(KEYINPUT4), .A4(new_n198), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n200), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT4), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n195), .A2(new_n204), .A3(G101), .ZN(new_n205));
  XOR2_X1   g019(.A(KEYINPUT2), .B(G113), .Z(new_n206));
  XNOR2_X1  g020(.A(G116), .B(G119), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g022(.A(KEYINPUT69), .ZN(new_n209));
  NAND3_X1  g023(.A1(new_n208), .A2(KEYINPUT68), .A3(new_n209), .ZN(new_n210));
  INV_X1    g024(.A(G119), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(G116), .ZN(new_n212));
  INV_X1    g026(.A(G116), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(G119), .ZN(new_n214));
  NAND2_X1  g028(.A1(new_n212), .A2(new_n214), .ZN(new_n215));
  XNOR2_X1  g029(.A(KEYINPUT2), .B(G113), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT68), .B1(new_n215), .B2(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n217), .A2(KEYINPUT69), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n206), .A2(new_n207), .ZN(new_n219));
  AND3_X1   g033(.A1(new_n210), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  AOI21_X1  g034(.A(new_n219), .B1(new_n210), .B2(new_n218), .ZN(new_n221));
  OAI211_X1 g035(.A(new_n203), .B(new_n205), .C1(new_n220), .C2(new_n221), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n189), .A2(G107), .ZN(new_n223));
  NOR2_X1   g037(.A1(new_n192), .A2(G104), .ZN(new_n224));
  OAI21_X1  g038(.A(G101), .B1(new_n223), .B2(new_n224), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n198), .A2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n207), .A2(KEYINPUT5), .ZN(new_n228));
  OAI211_X1 g042(.A(new_n228), .B(G113), .C1(KEYINPUT5), .C2(new_n212), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n227), .A2(new_n229), .A3(new_n208), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n222), .A2(new_n230), .ZN(new_n231));
  INV_X1    g045(.A(KEYINPUT6), .ZN(new_n232));
  XNOR2_X1  g046(.A(G110), .B(G122), .ZN(new_n233));
  XOR2_X1   g047(.A(new_n233), .B(KEYINPUT86), .Z(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n231), .A2(new_n232), .A3(new_n235), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n222), .A2(new_n234), .A3(new_n230), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n237), .A2(KEYINPUT6), .ZN(new_n238));
  AOI21_X1  g052(.A(new_n234), .B1(new_n222), .B2(new_n230), .ZN(new_n239));
  OAI211_X1 g053(.A(new_n187), .B(new_n236), .C1(new_n238), .C2(new_n239), .ZN(new_n240));
  INV_X1    g054(.A(new_n239), .ZN(new_n241));
  NAND4_X1  g055(.A1(new_n241), .A2(KEYINPUT87), .A3(KEYINPUT6), .A4(new_n237), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n240), .A2(new_n242), .ZN(new_n243));
  INV_X1    g057(.A(G146), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(G143), .ZN(new_n245));
  INV_X1    g059(.A(G143), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G146), .ZN(new_n247));
  AND2_X1   g061(.A1(new_n245), .A2(new_n247), .ZN(new_n248));
  AND2_X1   g062(.A1(KEYINPUT0), .A2(G128), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n248), .A2(new_n249), .ZN(new_n250));
  INV_X1    g064(.A(KEYINPUT64), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n247), .A2(new_n251), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n246), .A2(KEYINPUT64), .A3(G146), .ZN(new_n253));
  AOI22_X1  g067(.A1(new_n252), .A2(new_n253), .B1(G143), .B2(new_n244), .ZN(new_n254));
  NOR2_X1   g068(.A1(KEYINPUT0), .A2(G128), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n249), .A2(new_n255), .ZN(new_n256));
  INV_X1    g070(.A(new_n256), .ZN(new_n257));
  OAI21_X1  g071(.A(new_n250), .B1(new_n254), .B2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n258), .A2(G125), .ZN(new_n259));
  XNOR2_X1  g073(.A(new_n259), .B(KEYINPUT88), .ZN(new_n260));
  INV_X1    g074(.A(G224), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n261), .A2(G953), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n245), .A2(new_n247), .A3(G128), .ZN(new_n264));
  XNOR2_X1  g078(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n265));
  NOR2_X1   g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AND2_X1   g080(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n267));
  NOR2_X1   g081(.A1(KEYINPUT65), .A2(KEYINPUT1), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n245), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(KEYINPUT66), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  OAI211_X1 g085(.A(new_n245), .B(KEYINPUT66), .C1(new_n267), .C2(new_n268), .ZN(new_n272));
  NAND3_X1  g086(.A1(new_n271), .A2(G128), .A3(new_n272), .ZN(new_n273));
  INV_X1    g087(.A(new_n253), .ZN(new_n274));
  AOI21_X1  g088(.A(KEYINPUT64), .B1(new_n246), .B2(G146), .ZN(new_n275));
  OAI21_X1  g089(.A(new_n245), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n266), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  OAI211_X1 g092(.A(new_n260), .B(new_n263), .C1(G125), .C2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT88), .ZN(new_n280));
  XNOR2_X1  g094(.A(new_n259), .B(new_n280), .ZN(new_n281));
  NOR2_X1   g095(.A1(new_n278), .A2(G125), .ZN(new_n282));
  OAI21_X1  g096(.A(new_n262), .B1(new_n281), .B2(new_n282), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n279), .A2(new_n283), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n243), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g099(.A(G210), .B1(G237), .B2(G902), .ZN(new_n286));
  INV_X1    g100(.A(G902), .ZN(new_n287));
  INV_X1    g101(.A(KEYINPUT7), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n237), .B1(new_n279), .B2(new_n288), .ZN(new_n289));
  OAI21_X1  g103(.A(new_n288), .B1(new_n281), .B2(new_n282), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n234), .B(KEYINPUT8), .ZN(new_n291));
  INV_X1    g105(.A(new_n230), .ZN(new_n292));
  AOI21_X1  g106(.A(new_n227), .B1(new_n208), .B2(new_n229), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n291), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND3_X1  g108(.A1(new_n283), .A2(new_n290), .A3(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(new_n287), .B1(new_n289), .B2(new_n295), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND3_X1  g111(.A1(new_n285), .A2(new_n286), .A3(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(new_n286), .ZN(new_n299));
  INV_X1    g113(.A(new_n284), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n300), .B1(new_n240), .B2(new_n242), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n299), .B1(new_n301), .B2(new_n296), .ZN(new_n302));
  NAND3_X1  g116(.A1(new_n298), .A2(KEYINPUT89), .A3(new_n302), .ZN(new_n303));
  OAI21_X1  g117(.A(G214), .B1(G237), .B2(G902), .ZN(new_n304));
  XOR2_X1   g118(.A(new_n304), .B(KEYINPUT85), .Z(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  INV_X1    g120(.A(KEYINPUT89), .ZN(new_n307));
  NAND4_X1  g121(.A1(new_n285), .A2(new_n307), .A3(new_n286), .A4(new_n297), .ZN(new_n308));
  NAND3_X1  g122(.A1(new_n303), .A2(new_n306), .A3(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(KEYINPUT90), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n309), .A2(new_n310), .ZN(new_n311));
  NAND4_X1  g125(.A1(new_n303), .A2(KEYINPUT90), .A3(new_n308), .A4(new_n306), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  INV_X1    g127(.A(KEYINPUT79), .ZN(new_n314));
  INV_X1    g128(.A(KEYINPUT16), .ZN(new_n315));
  INV_X1    g129(.A(G140), .ZN(new_n316));
  NAND3_X1  g130(.A1(new_n315), .A2(new_n316), .A3(G125), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(KEYINPUT78), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n320), .A2(G140), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n319), .A2(new_n321), .A3(KEYINPUT16), .ZN(new_n322));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(new_n315), .A3(new_n316), .A4(G125), .ZN(new_n324));
  NAND4_X1  g138(.A1(new_n318), .A2(new_n322), .A3(G146), .A4(new_n324), .ZN(new_n325));
  XNOR2_X1  g139(.A(G125), .B(G140), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n326), .A2(new_n244), .ZN(new_n327));
  INV_X1    g141(.A(G128), .ZN(new_n328));
  NAND2_X1  g142(.A1(new_n328), .A2(G119), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT23), .ZN(new_n330));
  OAI21_X1  g144(.A(new_n329), .B1(KEYINPUT77), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n211), .A2(G128), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT77), .B(KEYINPUT23), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n331), .B(new_n332), .C1(new_n333), .C2(new_n329), .ZN(new_n334));
  NOR2_X1   g148(.A1(new_n334), .A2(G110), .ZN(new_n335));
  AND2_X1   g149(.A1(new_n329), .A2(new_n332), .ZN(new_n336));
  XOR2_X1   g150(.A(KEYINPUT24), .B(G110), .Z(new_n337));
  NOR2_X1   g151(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  OAI211_X1 g152(.A(new_n325), .B(new_n327), .C1(new_n335), .C2(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n318), .A2(new_n322), .A3(new_n324), .ZN(new_n340));
  NAND2_X1  g154(.A1(new_n340), .A2(new_n244), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n325), .ZN(new_n342));
  AOI22_X1  g156(.A1(new_n334), .A2(G110), .B1(new_n336), .B2(new_n337), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n342), .A2(new_n343), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n339), .A2(new_n344), .ZN(new_n345));
  XNOR2_X1  g159(.A(KEYINPUT22), .B(G137), .ZN(new_n346));
  INV_X1    g160(.A(G953), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n347), .A2(G221), .A3(G234), .ZN(new_n348));
  XNOR2_X1  g162(.A(new_n346), .B(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(new_n349), .ZN(new_n350));
  NAND2_X1  g164(.A1(new_n345), .A2(new_n350), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n339), .A2(new_n344), .A3(new_n349), .ZN(new_n352));
  NAND3_X1  g166(.A1(new_n351), .A2(new_n287), .A3(new_n352), .ZN(new_n353));
  INV_X1    g167(.A(KEYINPUT25), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NAND4_X1  g169(.A1(new_n351), .A2(KEYINPUT25), .A3(new_n287), .A4(new_n352), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(G217), .ZN(new_n358));
  AOI21_X1  g172(.A(new_n358), .B1(G234), .B2(new_n287), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n314), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  INV_X1    g174(.A(new_n360), .ZN(new_n361));
  NAND3_X1  g175(.A1(new_n357), .A2(new_n314), .A3(new_n359), .ZN(new_n362));
  INV_X1    g176(.A(new_n351), .ZN(new_n363));
  INV_X1    g177(.A(new_n352), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n363), .A2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(new_n359), .A2(G902), .ZN(new_n366));
  NAND2_X1  g180(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n361), .A2(new_n362), .A3(new_n367), .ZN(new_n368));
  INV_X1    g182(.A(KEYINPUT28), .ZN(new_n369));
  AOI22_X1  g183(.A1(new_n276), .A2(new_n256), .B1(new_n249), .B2(new_n248), .ZN(new_n370));
  INV_X1    g184(.A(KEYINPUT11), .ZN(new_n371));
  INV_X1    g185(.A(G134), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n371), .B1(new_n372), .B2(G137), .ZN(new_n373));
  INV_X1    g187(.A(G137), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT11), .A3(G134), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n372), .A2(G137), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n373), .A2(new_n375), .A3(new_n376), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n377), .A2(G131), .ZN(new_n378));
  INV_X1    g192(.A(G131), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n373), .A2(new_n375), .A3(new_n379), .A4(new_n376), .ZN(new_n380));
  NAND2_X1  g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n370), .A2(new_n381), .ZN(new_n382));
  NOR2_X1   g196(.A1(new_n372), .A2(G137), .ZN(new_n383));
  NOR2_X1   g197(.A1(new_n374), .A2(G134), .ZN(new_n384));
  OAI21_X1  g198(.A(G131), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n380), .A2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(KEYINPUT70), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT70), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n380), .A2(new_n385), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n387), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g204(.A(new_n382), .B1(new_n277), .B2(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n219), .ZN(new_n392));
  AOI21_X1  g206(.A(new_n209), .B1(new_n208), .B2(KEYINPUT68), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT68), .ZN(new_n394));
  AOI211_X1 g208(.A(new_n394), .B(KEYINPUT69), .C1(new_n206), .C2(new_n207), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n392), .B1(new_n393), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n210), .A2(new_n218), .A3(new_n219), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n396), .A2(new_n397), .ZN(new_n398));
  OAI21_X1  g212(.A(new_n369), .B1(new_n391), .B2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT73), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n399), .A2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n328), .B1(new_n269), .B2(new_n270), .ZN(new_n402));
  AOI21_X1  g216(.A(new_n254), .B1(new_n402), .B2(new_n272), .ZN(new_n403));
  OAI211_X1 g217(.A(new_n387), .B(new_n389), .C1(new_n403), .C2(new_n266), .ZN(new_n404));
  NAND4_X1  g218(.A1(new_n404), .A2(new_n397), .A3(new_n396), .A4(new_n382), .ZN(new_n405));
  NAND3_X1  g219(.A1(new_n405), .A2(KEYINPUT73), .A3(new_n369), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n401), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g221(.A1(G237), .A2(G953), .ZN(new_n408));
  NAND2_X1  g222(.A1(new_n408), .A2(G210), .ZN(new_n409));
  XOR2_X1   g223(.A(new_n409), .B(KEYINPUT72), .Z(new_n410));
  XNOR2_X1  g224(.A(KEYINPUT26), .B(G101), .ZN(new_n411));
  XNOR2_X1  g225(.A(KEYINPUT71), .B(KEYINPUT27), .ZN(new_n412));
  XNOR2_X1  g226(.A(new_n411), .B(new_n412), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n410), .B(new_n413), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(KEYINPUT29), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n391), .A2(new_n398), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n416), .A2(new_n405), .A3(KEYINPUT75), .ZN(new_n417));
  INV_X1    g231(.A(KEYINPUT75), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n391), .A2(new_n398), .A3(new_n418), .ZN(new_n419));
  NAND3_X1  g233(.A1(new_n417), .A2(KEYINPUT28), .A3(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n420), .A2(KEYINPUT76), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT76), .ZN(new_n422));
  NAND4_X1  g236(.A1(new_n417), .A2(new_n422), .A3(KEYINPUT28), .A4(new_n419), .ZN(new_n423));
  AOI211_X1 g237(.A(new_n407), .B(new_n415), .C1(new_n421), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g238(.A1(new_n391), .A2(new_n398), .ZN(new_n425));
  OAI211_X1 g239(.A(new_n380), .B(new_n385), .C1(new_n403), .C2(new_n266), .ZN(new_n426));
  AOI22_X1  g240(.A1(new_n426), .A2(new_n382), .B1(new_n396), .B2(new_n397), .ZN(new_n427));
  OAI21_X1  g241(.A(KEYINPUT28), .B1(new_n425), .B2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n428), .A2(new_n401), .A3(new_n406), .A4(new_n414), .ZN(new_n429));
  INV_X1    g243(.A(KEYINPUT29), .ZN(new_n430));
  NAND2_X1  g244(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  OAI21_X1  g245(.A(new_n382), .B1(new_n277), .B2(new_n386), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT30), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n432), .A2(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT67), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n404), .A2(KEYINPUT30), .A3(new_n382), .ZN(new_n437));
  NAND3_X1  g251(.A1(new_n432), .A2(KEYINPUT67), .A3(new_n433), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n436), .A2(new_n398), .A3(new_n437), .A4(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(new_n414), .B1(new_n439), .B2(new_n405), .ZN(new_n440));
  OAI21_X1  g254(.A(new_n287), .B1(new_n431), .B2(new_n440), .ZN(new_n441));
  OAI21_X1  g255(.A(G472), .B1(new_n424), .B2(new_n441), .ZN(new_n442));
  NAND3_X1  g256(.A1(new_n439), .A2(new_n405), .A3(new_n414), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT31), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n428), .A2(new_n401), .A3(new_n406), .ZN(new_n445));
  INV_X1    g259(.A(new_n414), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT31), .ZN(new_n448));
  NAND4_X1  g262(.A1(new_n439), .A2(new_n448), .A3(new_n405), .A4(new_n414), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n444), .A2(new_n447), .A3(new_n449), .ZN(new_n450));
  NOR2_X1   g264(.A1(G472), .A2(G902), .ZN(new_n451));
  NAND3_X1  g265(.A1(new_n450), .A2(KEYINPUT32), .A3(new_n451), .ZN(new_n452));
  AND2_X1   g266(.A1(new_n442), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n450), .A2(new_n451), .ZN(new_n454));
  XOR2_X1   g268(.A(KEYINPUT74), .B(KEYINPUT32), .Z(new_n455));
  NAND2_X1  g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  AOI21_X1  g270(.A(new_n368), .B1(new_n453), .B2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(KEYINPUT9), .B(G234), .ZN(new_n458));
  OAI21_X1  g272(.A(G221), .B1(new_n458), .B2(G902), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n245), .A2(KEYINPUT1), .ZN(new_n461));
  AOI22_X1  g275(.A1(new_n461), .A2(G128), .B1(new_n245), .B2(new_n247), .ZN(new_n462));
  OAI211_X1 g276(.A(new_n198), .B(new_n225), .C1(new_n266), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n267), .A2(new_n268), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n248), .A2(new_n464), .A3(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n226), .A2(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(new_n463), .B1(new_n403), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g281(.A1(new_n467), .A2(KEYINPUT12), .A3(new_n381), .ZN(new_n468));
  INV_X1    g282(.A(KEYINPUT81), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n468), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n467), .A2(new_n381), .ZN(new_n471));
  INV_X1    g285(.A(KEYINPUT12), .ZN(new_n472));
  NAND2_X1  g286(.A1(new_n471), .A2(new_n472), .ZN(new_n473));
  NAND4_X1  g287(.A1(new_n467), .A2(KEYINPUT81), .A3(KEYINPUT12), .A4(new_n381), .ZN(new_n474));
  NAND3_X1  g288(.A1(new_n470), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT84), .ZN(new_n476));
  NAND2_X1  g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n203), .A2(new_n370), .A3(new_n205), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  NOR2_X1   g293(.A1(new_n226), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n278), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(new_n381), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n463), .A2(new_n479), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n478), .A2(new_n481), .A3(new_n482), .A4(new_n483), .ZN(new_n484));
  XNOR2_X1  g298(.A(G110), .B(G140), .ZN(new_n485));
  AND2_X1   g299(.A1(new_n347), .A2(G227), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n485), .B(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(new_n487), .ZN(new_n488));
  AND2_X1   g302(.A1(new_n484), .A2(new_n488), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n470), .A2(new_n473), .A3(KEYINPUT84), .A4(new_n474), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n477), .A2(new_n489), .A3(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n480), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n483), .B1(new_n277), .B2(new_n492), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n370), .A2(new_n205), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n494), .B1(new_n200), .B2(new_n202), .ZN(new_n495));
  OAI21_X1  g309(.A(new_n381), .B1(new_n493), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n484), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n487), .ZN(new_n498));
  AOI211_X1 g312(.A(G469), .B(G902), .C1(new_n491), .C2(new_n498), .ZN(new_n499));
  INV_X1    g313(.A(G469), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n475), .A2(new_n484), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n501), .A2(new_n487), .ZN(new_n502));
  INV_X1    g316(.A(KEYINPUT82), .ZN(new_n503));
  NAND2_X1  g317(.A1(new_n489), .A2(new_n496), .ZN(new_n504));
  NAND3_X1  g318(.A1(new_n502), .A2(new_n503), .A3(new_n504), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n488), .B1(new_n475), .B2(new_n484), .ZN(new_n506));
  AND3_X1   g320(.A1(new_n484), .A2(new_n496), .A3(new_n488), .ZN(new_n507));
  OAI21_X1  g321(.A(KEYINPUT82), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n508), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n500), .B1(new_n509), .B2(new_n287), .ZN(new_n510));
  AOI21_X1  g324(.A(new_n499), .B1(new_n510), .B2(KEYINPUT83), .ZN(new_n511));
  INV_X1    g325(.A(KEYINPUT83), .ZN(new_n512));
  AOI21_X1  g326(.A(G902), .B1(new_n505), .B2(new_n508), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n512), .B1(new_n513), .B2(new_n500), .ZN(new_n514));
  AOI21_X1  g328(.A(new_n460), .B1(new_n511), .B2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT102), .ZN(new_n516));
  NOR3_X1   g330(.A1(new_n458), .A2(new_n358), .A3(G953), .ZN(new_n517));
  INV_X1    g331(.A(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n246), .A2(G128), .ZN(new_n519));
  NAND2_X1  g333(.A1(new_n328), .A2(G143), .ZN(new_n520));
  AND3_X1   g334(.A1(new_n519), .A2(new_n520), .A3(new_n372), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT98), .ZN(new_n522));
  NAND4_X1  g336(.A1(new_n522), .A2(new_n246), .A3(KEYINPUT13), .A4(G128), .ZN(new_n523));
  AND2_X1   g337(.A1(new_n523), .A2(G134), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT13), .ZN(new_n525));
  OAI21_X1  g339(.A(new_n525), .B1(new_n328), .B2(G143), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n246), .A2(KEYINPUT13), .A3(G128), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n526), .A2(new_n527), .A3(KEYINPUT98), .A4(new_n520), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n521), .B1(new_n524), .B2(new_n528), .ZN(new_n529));
  INV_X1    g343(.A(KEYINPUT97), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n213), .A2(G122), .ZN(new_n531));
  INV_X1    g345(.A(G122), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n532), .A2(G116), .ZN(new_n533));
  AND3_X1   g347(.A1(new_n531), .A2(new_n533), .A3(new_n192), .ZN(new_n534));
  AOI21_X1  g348(.A(new_n192), .B1(new_n531), .B2(new_n533), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n530), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n531), .A2(new_n533), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n537), .A2(G107), .ZN(new_n538));
  XNOR2_X1  g352(.A(G116), .B(G122), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(new_n192), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(new_n540), .A3(KEYINPUT97), .ZN(new_n541));
  AND3_X1   g355(.A1(new_n529), .A2(new_n536), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g356(.A(new_n372), .B1(new_n519), .B2(new_n520), .ZN(new_n543));
  OAI21_X1  g357(.A(new_n540), .B1(new_n521), .B2(new_n543), .ZN(new_n544));
  INV_X1    g358(.A(KEYINPUT99), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT14), .ZN(new_n546));
  AND3_X1   g360(.A1(new_n531), .A2(new_n533), .A3(new_n546), .ZN(new_n547));
  OAI21_X1  g361(.A(G107), .B1(new_n531), .B2(new_n546), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n545), .B1(new_n547), .B2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n539), .A2(new_n546), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n532), .A2(G116), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n192), .B1(new_n551), .B2(KEYINPUT14), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n550), .A2(KEYINPUT99), .A3(new_n552), .ZN(new_n553));
  AOI21_X1  g367(.A(new_n544), .B1(new_n549), .B2(new_n553), .ZN(new_n554));
  OAI21_X1  g368(.A(new_n518), .B1(new_n542), .B2(new_n554), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT100), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n529), .A2(new_n536), .A3(new_n541), .ZN(new_n557));
  AND2_X1   g371(.A1(new_n549), .A2(new_n553), .ZN(new_n558));
  OAI211_X1 g372(.A(new_n557), .B(new_n517), .C1(new_n558), .C2(new_n544), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n555), .A2(new_n556), .A3(new_n559), .ZN(new_n560));
  OAI211_X1 g374(.A(KEYINPUT100), .B(new_n518), .C1(new_n542), .C2(new_n554), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n560), .A2(new_n287), .A3(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(KEYINPUT101), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g378(.A1(new_n560), .A2(KEYINPUT101), .A3(new_n287), .A4(new_n561), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(G478), .ZN(new_n567));
  NOR2_X1   g381(.A1(new_n567), .A2(KEYINPUT15), .ZN(new_n568));
  INV_X1    g382(.A(new_n568), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n566), .A2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n565), .A2(new_n568), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n516), .B1(new_n570), .B2(new_n571), .ZN(new_n572));
  AOI21_X1  g386(.A(new_n568), .B1(new_n564), .B2(new_n565), .ZN(new_n573));
  INV_X1    g387(.A(new_n571), .ZN(new_n574));
  NOR3_X1   g388(.A1(new_n573), .A2(KEYINPUT102), .A3(new_n574), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n572), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT96), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n326), .B(new_n244), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT91), .ZN(new_n579));
  OR2_X1    g393(.A1(new_n326), .A2(new_n244), .ZN(new_n580));
  INV_X1    g394(.A(KEYINPUT91), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n580), .A2(new_n581), .A3(new_n327), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n579), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(G237), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n584), .A2(new_n347), .A3(G214), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n246), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n408), .A2(G143), .A3(G214), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g402(.A(KEYINPUT18), .ZN(new_n589));
  OAI21_X1  g403(.A(new_n588), .B1(new_n589), .B2(new_n379), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n586), .A2(KEYINPUT18), .A3(G131), .A4(new_n587), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n583), .A2(new_n592), .ZN(new_n593));
  INV_X1    g407(.A(new_n587), .ZN(new_n594));
  AOI21_X1  g408(.A(G143), .B1(new_n408), .B2(G214), .ZN(new_n595));
  OAI211_X1 g409(.A(KEYINPUT17), .B(G131), .C1(new_n594), .C2(new_n595), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n341), .A2(new_n325), .A3(new_n596), .ZN(new_n597));
  AND2_X1   g411(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT94), .ZN(new_n599));
  NAND4_X1  g413(.A1(new_n341), .A2(new_n599), .A3(new_n325), .A4(new_n596), .ZN(new_n600));
  NAND3_X1  g414(.A1(new_n586), .A2(new_n379), .A3(new_n587), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n601), .A2(KEYINPUT92), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n588), .A2(G131), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT17), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT92), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n586), .A2(new_n605), .A3(new_n379), .A4(new_n587), .ZN(new_n606));
  NAND4_X1  g420(.A1(new_n602), .A2(new_n603), .A3(new_n604), .A4(new_n606), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n600), .A2(new_n607), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n593), .B1(new_n598), .B2(new_n608), .ZN(new_n609));
  XNOR2_X1  g423(.A(G113), .B(G122), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(new_n189), .ZN(new_n611));
  INV_X1    g425(.A(new_n611), .ZN(new_n612));
  NOR2_X1   g426(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  AOI22_X1  g427(.A1(new_n579), .A2(new_n582), .B1(new_n590), .B2(new_n591), .ZN(new_n614));
  AND2_X1   g428(.A1(new_n600), .A2(new_n607), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n597), .A2(KEYINPUT94), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n614), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g431(.A(KEYINPUT95), .B1(new_n617), .B2(new_n611), .ZN(new_n618));
  INV_X1    g432(.A(KEYINPUT95), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n609), .A2(new_n619), .A3(new_n612), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n613), .B1(new_n618), .B2(new_n620), .ZN(new_n621));
  OAI21_X1  g435(.A(new_n577), .B1(new_n621), .B2(G902), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n617), .A2(new_n611), .ZN(new_n623));
  NAND3_X1  g437(.A1(new_n616), .A2(new_n607), .A3(new_n600), .ZN(new_n624));
  AOI211_X1 g438(.A(KEYINPUT95), .B(new_n611), .C1(new_n624), .C2(new_n593), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n619), .B1(new_n609), .B2(new_n612), .ZN(new_n626));
  OAI21_X1  g440(.A(new_n623), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n627), .A2(KEYINPUT96), .A3(new_n287), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n622), .A2(G475), .A3(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n602), .A2(new_n603), .A3(new_n606), .ZN(new_n630));
  AND2_X1   g444(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n631));
  NOR2_X1   g445(.A1(KEYINPUT93), .A2(KEYINPUT19), .ZN(new_n632));
  OAI21_X1  g446(.A(new_n326), .B1(new_n631), .B2(new_n632), .ZN(new_n633));
  OAI21_X1  g447(.A(new_n633), .B1(new_n326), .B2(new_n632), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n325), .B1(new_n634), .B2(G146), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n593), .B1(new_n630), .B2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(new_n612), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n623), .A2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  INV_X1    g453(.A(G475), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n640), .A2(new_n287), .ZN(new_n641));
  OAI21_X1  g455(.A(KEYINPUT20), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(KEYINPUT20), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n638), .A2(new_n643), .A3(new_n640), .A4(new_n287), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n629), .A2(new_n645), .ZN(new_n646));
  AND2_X1   g460(.A1(new_n347), .A2(G952), .ZN(new_n647));
  INV_X1    g461(.A(G234), .ZN(new_n648));
  OAI21_X1  g462(.A(new_n647), .B1(new_n648), .B2(new_n584), .ZN(new_n649));
  INV_X1    g463(.A(new_n649), .ZN(new_n650));
  OAI211_X1 g464(.A(G902), .B(G953), .C1(new_n648), .C2(new_n584), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n651), .B(KEYINPUT103), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT21), .B(G898), .ZN(new_n653));
  AOI21_X1  g467(.A(new_n650), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  NOR3_X1   g468(.A1(new_n576), .A2(new_n646), .A3(new_n654), .ZN(new_n655));
  NAND4_X1  g469(.A1(new_n313), .A2(new_n457), .A3(new_n515), .A4(new_n655), .ZN(new_n656));
  XNOR2_X1  g470(.A(KEYINPUT104), .B(G101), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n656), .B(new_n657), .ZN(G3));
  INV_X1    g472(.A(new_n368), .ZN(new_n659));
  AOI21_X1  g473(.A(new_n503), .B1(new_n502), .B2(new_n504), .ZN(new_n660));
  NOR3_X1   g474(.A1(new_n506), .A2(new_n507), .A3(KEYINPUT82), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n287), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n662), .A2(KEYINPUT83), .A3(G469), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n491), .A2(new_n498), .ZN(new_n664));
  NAND3_X1  g478(.A1(new_n664), .A2(new_n500), .A3(new_n287), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n514), .A2(new_n663), .A3(new_n665), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n450), .A2(new_n287), .ZN(new_n667));
  AOI22_X1  g481(.A1(new_n667), .A2(G472), .B1(new_n451), .B2(new_n450), .ZN(new_n668));
  AND4_X1   g482(.A1(new_n659), .A2(new_n666), .A3(new_n459), .A4(new_n668), .ZN(new_n669));
  AOI21_X1  g483(.A(new_n305), .B1(new_n298), .B2(new_n302), .ZN(new_n670));
  INV_X1    g484(.A(new_n654), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT33), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n560), .A2(new_n672), .A3(new_n561), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n555), .A2(KEYINPUT33), .A3(new_n559), .ZN(new_n674));
  NAND4_X1  g488(.A1(new_n673), .A2(G478), .A3(new_n287), .A4(new_n674), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n562), .A2(new_n567), .ZN(new_n676));
  NAND2_X1  g490(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  INV_X1    g491(.A(new_n677), .ZN(new_n678));
  AOI21_X1  g492(.A(new_n678), .B1(new_n629), .B2(new_n645), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n670), .A2(new_n671), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n669), .A2(new_n681), .ZN(new_n682));
  XOR2_X1   g496(.A(KEYINPUT34), .B(G104), .Z(new_n683));
  XNOR2_X1  g497(.A(new_n682), .B(new_n683), .ZN(G6));
  NAND2_X1  g498(.A1(new_n618), .A2(new_n620), .ZN(new_n685));
  AOI21_X1  g499(.A(G902), .B1(new_n685), .B2(new_n623), .ZN(new_n686));
  AOI21_X1  g500(.A(new_n640), .B1(new_n686), .B2(KEYINPUT96), .ZN(new_n687));
  AOI22_X1  g501(.A1(new_n687), .A2(new_n622), .B1(new_n642), .B2(new_n644), .ZN(new_n688));
  NAND4_X1  g502(.A1(new_n670), .A2(new_n671), .A3(new_n688), .A4(new_n576), .ZN(new_n689));
  INV_X1    g503(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g504(.A1(new_n669), .A2(new_n690), .ZN(new_n691));
  XOR2_X1   g505(.A(KEYINPUT35), .B(G107), .Z(new_n692));
  XNOR2_X1  g506(.A(new_n691), .B(new_n692), .ZN(G9));
  NAND2_X1  g507(.A1(new_n667), .A2(G472), .ZN(new_n694));
  OR2_X1    g508(.A1(new_n345), .A2(KEYINPUT105), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n345), .A2(KEYINPUT105), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n695), .A2(new_n696), .ZN(new_n697));
  NOR2_X1   g511(.A1(new_n350), .A2(KEYINPUT36), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n697), .A2(new_n699), .ZN(new_n700));
  NAND3_X1  g514(.A1(new_n695), .A2(new_n698), .A3(new_n696), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n700), .A2(new_n366), .A3(new_n701), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n361), .A2(new_n362), .A3(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n694), .A2(new_n454), .A3(new_n703), .ZN(new_n704));
  XNOR2_X1  g518(.A(new_n704), .B(KEYINPUT106), .ZN(new_n705));
  NAND4_X1  g519(.A1(new_n705), .A2(new_n313), .A3(new_n515), .A4(new_n655), .ZN(new_n706));
  XOR2_X1   g520(.A(KEYINPUT37), .B(G110), .Z(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT107), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n706), .B(new_n708), .ZN(G12));
  NAND3_X1  g523(.A1(new_n456), .A2(new_n442), .A3(new_n452), .ZN(new_n710));
  AND3_X1   g524(.A1(new_n710), .A2(new_n670), .A3(new_n703), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n570), .A2(new_n516), .A3(new_n571), .ZN(new_n712));
  OAI21_X1  g526(.A(KEYINPUT102), .B1(new_n573), .B2(new_n574), .ZN(new_n713));
  NAND4_X1  g527(.A1(new_n629), .A2(new_n645), .A3(new_n712), .A4(new_n713), .ZN(new_n714));
  XNOR2_X1  g528(.A(KEYINPUT108), .B(G900), .ZN(new_n715));
  AOI21_X1  g529(.A(new_n650), .B1(new_n652), .B2(new_n715), .ZN(new_n716));
  OAI21_X1  g530(.A(KEYINPUT109), .B1(new_n714), .B2(new_n716), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT109), .ZN(new_n718));
  INV_X1    g532(.A(new_n716), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n688), .A2(new_n576), .A3(new_n718), .A4(new_n719), .ZN(new_n720));
  AND2_X1   g534(.A1(new_n717), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n711), .A2(new_n721), .A3(new_n515), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G128), .ZN(G30));
  XOR2_X1   g537(.A(new_n716), .B(KEYINPUT39), .Z(new_n724));
  NAND2_X1  g538(.A1(new_n515), .A2(new_n724), .ZN(new_n725));
  OR2_X1    g539(.A1(new_n725), .A2(KEYINPUT40), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n303), .A2(new_n308), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(KEYINPUT38), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n712), .A2(new_n713), .ZN(new_n729));
  NOR2_X1   g543(.A1(new_n688), .A2(new_n729), .ZN(new_n730));
  AND3_X1   g544(.A1(new_n361), .A2(new_n362), .A3(new_n702), .ZN(new_n731));
  NAND3_X1  g545(.A1(new_n730), .A2(new_n306), .A3(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT110), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NOR2_X1   g548(.A1(new_n728), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n725), .A2(KEYINPUT40), .ZN(new_n736));
  NAND2_X1  g550(.A1(new_n732), .A2(new_n733), .ZN(new_n737));
  AND2_X1   g551(.A1(new_n439), .A2(new_n405), .ZN(new_n738));
  NOR2_X1   g552(.A1(new_n738), .A2(new_n446), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n417), .A2(new_n419), .ZN(new_n740));
  OAI21_X1  g554(.A(new_n287), .B1(new_n740), .B2(new_n414), .ZN(new_n741));
  OAI21_X1  g555(.A(G472), .B1(new_n739), .B2(new_n741), .ZN(new_n742));
  NAND3_X1  g556(.A1(new_n456), .A2(new_n742), .A3(new_n452), .ZN(new_n743));
  AND2_X1   g557(.A1(new_n737), .A2(new_n743), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n726), .A2(new_n735), .A3(new_n736), .A4(new_n744), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(G143), .ZN(G45));
  AOI21_X1  g560(.A(new_n731), .B1(new_n453), .B2(new_n456), .ZN(new_n747));
  AOI211_X1 g561(.A(new_n678), .B(new_n716), .C1(new_n629), .C2(new_n645), .ZN(new_n748));
  NAND4_X1  g562(.A1(new_n747), .A2(new_n515), .A3(new_n670), .A4(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G146), .ZN(G48));
  AOI21_X1  g564(.A(new_n500), .B1(new_n664), .B2(new_n287), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n751), .A2(new_n499), .A3(new_n460), .ZN(new_n752));
  NAND3_X1  g566(.A1(new_n457), .A2(new_n681), .A3(new_n752), .ZN(new_n753));
  XNOR2_X1  g567(.A(KEYINPUT41), .B(G113), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n753), .B(new_n754), .ZN(G15));
  NAND3_X1  g569(.A1(new_n690), .A2(new_n457), .A3(new_n752), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G116), .ZN(G18));
  NAND3_X1  g571(.A1(new_n711), .A2(new_n655), .A3(new_n752), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G119), .ZN(G21));
  NAND4_X1  g573(.A1(new_n730), .A2(new_n671), .A3(new_n670), .A4(new_n752), .ZN(new_n760));
  AOI21_X1  g574(.A(new_n407), .B1(new_n421), .B2(new_n423), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(new_n414), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n444), .A2(new_n449), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n451), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n694), .A2(new_n764), .A3(new_n659), .ZN(new_n765));
  OR2_X1    g579(.A1(new_n760), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G122), .ZN(G24));
  NAND2_X1  g581(.A1(new_n670), .A2(new_n752), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n694), .A2(new_n764), .A3(new_n703), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n679), .A2(new_n719), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n768), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  XNOR2_X1  g585(.A(new_n771), .B(new_n320), .ZN(G27));
  INV_X1    g586(.A(KEYINPUT111), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n502), .A2(new_n504), .ZN(new_n774));
  AOI21_X1  g588(.A(new_n500), .B1(new_n774), .B2(new_n287), .ZN(new_n775));
  OAI21_X1  g589(.A(new_n773), .B1(new_n499), .B2(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n506), .A2(new_n507), .ZN(new_n777));
  OAI21_X1  g591(.A(G469), .B1(new_n777), .B2(G902), .ZN(new_n778));
  NAND3_X1  g592(.A1(new_n665), .A2(KEYINPUT111), .A3(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n776), .A2(new_n779), .ZN(new_n780));
  NOR2_X1   g594(.A1(new_n460), .A2(new_n305), .ZN(new_n781));
  AND3_X1   g595(.A1(new_n727), .A2(new_n780), .A3(new_n781), .ZN(new_n782));
  NOR2_X1   g596(.A1(new_n770), .A2(KEYINPUT42), .ZN(new_n783));
  NAND3_X1  g597(.A1(new_n782), .A2(new_n457), .A3(new_n783), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n727), .A2(new_n748), .A3(new_n780), .A4(new_n781), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n442), .A2(new_n452), .ZN(new_n786));
  AOI21_X1  g600(.A(KEYINPUT32), .B1(new_n450), .B2(new_n451), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n659), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  OAI21_X1  g602(.A(KEYINPUT42), .B1(new_n785), .B2(new_n788), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n784), .A2(new_n789), .ZN(new_n790));
  XNOR2_X1  g604(.A(new_n790), .B(new_n379), .ZN(G33));
  NAND3_X1  g605(.A1(new_n782), .A2(new_n721), .A3(new_n457), .ZN(new_n792));
  XNOR2_X1  g606(.A(new_n792), .B(G134), .ZN(G36));
  NOR2_X1   g607(.A1(new_n660), .A2(new_n661), .ZN(new_n794));
  OAI21_X1  g608(.A(G469), .B1(new_n794), .B2(KEYINPUT45), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(KEYINPUT112), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT112), .ZN(new_n797));
  OAI211_X1 g611(.A(new_n797), .B(G469), .C1(new_n794), .C2(KEYINPUT45), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n777), .A2(KEYINPUT45), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n796), .A2(new_n798), .A3(new_n799), .ZN(new_n800));
  NAND2_X1  g614(.A1(G469), .A2(G902), .ZN(new_n801));
  AOI21_X1  g615(.A(KEYINPUT46), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  NOR2_X1   g616(.A1(new_n802), .A2(new_n499), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n800), .A2(KEYINPUT46), .A3(new_n801), .ZN(new_n804));
  NAND2_X1  g618(.A1(new_n803), .A2(new_n804), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n459), .A3(new_n724), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n305), .B1(new_n303), .B2(new_n308), .ZN(new_n807));
  INV_X1    g621(.A(new_n807), .ZN(new_n808));
  NOR2_X1   g622(.A1(new_n668), .A2(new_n731), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n688), .A2(new_n677), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT43), .ZN(new_n811));
  OR3_X1    g625(.A1(new_n646), .A2(KEYINPUT43), .A3(new_n678), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n809), .A2(new_n811), .A3(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT44), .ZN(new_n814));
  AOI21_X1  g628(.A(new_n808), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  OAI21_X1  g629(.A(new_n815), .B1(new_n814), .B2(new_n813), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n806), .A2(new_n816), .ZN(new_n817));
  XNOR2_X1  g631(.A(new_n817), .B(new_n374), .ZN(G39));
  NOR4_X1   g632(.A1(new_n808), .A2(new_n710), .A3(new_n659), .A4(new_n770), .ZN(new_n819));
  AND3_X1   g633(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n459), .ZN(new_n820));
  AOI21_X1  g634(.A(KEYINPUT47), .B1(new_n805), .B2(new_n459), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n819), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  XNOR2_X1  g636(.A(new_n822), .B(G140), .ZN(G42));
  INV_X1    g637(.A(KEYINPUT51), .ZN(new_n824));
  AND3_X1   g638(.A1(new_n811), .A2(new_n812), .A3(new_n650), .ZN(new_n825));
  INV_X1    g639(.A(new_n765), .ZN(new_n826));
  NAND2_X1  g640(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  NOR2_X1   g641(.A1(new_n827), .A2(new_n808), .ZN(new_n828));
  INV_X1    g642(.A(new_n828), .ZN(new_n829));
  NOR2_X1   g643(.A1(new_n820), .A2(new_n821), .ZN(new_n830));
  NOR2_X1   g644(.A1(new_n751), .A2(new_n499), .ZN(new_n831));
  INV_X1    g645(.A(new_n831), .ZN(new_n832));
  OR2_X1    g646(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n832), .A2(KEYINPUT118), .ZN(new_n834));
  NAND3_X1  g648(.A1(new_n833), .A2(new_n460), .A3(new_n834), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n829), .B1(new_n830), .B2(new_n835), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n836), .A2(KEYINPUT119), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n728), .A2(new_n305), .A3(new_n752), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n827), .ZN(new_n839));
  OR2_X1    g653(.A1(KEYINPUT120), .A2(KEYINPUT50), .ZN(new_n840));
  XNOR2_X1  g654(.A(new_n839), .B(new_n840), .ZN(new_n841));
  AND2_X1   g655(.A1(new_n807), .A2(new_n752), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n743), .A2(new_n368), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n842), .A2(new_n650), .A3(new_n843), .ZN(new_n844));
  NOR3_X1   g658(.A1(new_n844), .A2(new_n646), .A3(new_n677), .ZN(new_n845));
  AND3_X1   g659(.A1(new_n694), .A2(new_n764), .A3(new_n703), .ZN(new_n846));
  AND2_X1   g660(.A1(new_n825), .A2(new_n842), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n845), .B1(new_n846), .B2(new_n847), .ZN(new_n848));
  AND2_X1   g662(.A1(new_n841), .A2(new_n848), .ZN(new_n849));
  OAI21_X1  g663(.A(new_n849), .B1(new_n836), .B2(KEYINPUT119), .ZN(new_n850));
  OAI21_X1  g664(.A(new_n824), .B1(new_n837), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n646), .A2(new_n677), .ZN(new_n852));
  OAI221_X1 g666(.A(new_n647), .B1(new_n827), .B2(new_n768), .C1(new_n852), .C2(new_n844), .ZN(new_n853));
  INV_X1    g667(.A(new_n788), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n854), .ZN(new_n855));
  OR2_X1    g669(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n855), .A2(KEYINPUT48), .ZN(new_n857));
  AOI21_X1  g671(.A(new_n853), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(KEYINPUT121), .ZN(new_n859));
  XNOR2_X1  g673(.A(new_n858), .B(new_n859), .ZN(new_n860));
  AND2_X1   g674(.A1(new_n849), .A2(KEYINPUT51), .ZN(new_n861));
  INV_X1    g675(.A(new_n836), .ZN(new_n862));
  AOI21_X1  g676(.A(new_n860), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n851), .A2(new_n863), .ZN(new_n864));
  INV_X1    g678(.A(new_n781), .ZN(new_n865));
  AOI21_X1  g679(.A(new_n865), .B1(new_n303), .B2(new_n308), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n846), .A3(new_n748), .A4(new_n780), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n866), .A2(new_n710), .A3(new_n659), .A4(new_n780), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n717), .A2(new_n720), .ZN(new_n869));
  OAI21_X1  g683(.A(new_n867), .B1(new_n868), .B2(new_n869), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n570), .A2(new_n571), .ZN(new_n871));
  NOR3_X1   g685(.A1(new_n646), .A2(new_n871), .A3(new_n716), .ZN(new_n872));
  NAND2_X1  g686(.A1(new_n807), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g687(.A1(new_n666), .A2(new_n459), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n710), .A2(new_n703), .ZN(new_n875));
  NOR3_X1   g689(.A1(new_n873), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  NOR2_X1   g690(.A1(new_n870), .A2(new_n876), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n854), .A2(new_n748), .A3(new_n780), .A4(new_n866), .ZN(new_n878));
  NAND3_X1  g692(.A1(new_n727), .A2(new_n780), .A3(new_n781), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n710), .A2(new_n659), .ZN(new_n880));
  NOR2_X1   g694(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  AOI22_X1  g695(.A1(new_n878), .A2(KEYINPUT42), .B1(new_n881), .B2(new_n783), .ZN(new_n882));
  NAND3_X1  g696(.A1(new_n710), .A2(new_n670), .A3(new_n703), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n655), .A2(new_n752), .ZN(new_n884));
  NAND3_X1  g698(.A1(new_n710), .A2(new_n659), .A3(new_n752), .ZN(new_n885));
  OAI22_X1  g699(.A1(new_n883), .A2(new_n884), .B1(new_n885), .B2(new_n689), .ZN(new_n886));
  OAI22_X1  g700(.A1(new_n765), .A2(new_n760), .B1(new_n885), .B2(new_n680), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n877), .A2(new_n882), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g703(.A(KEYINPUT113), .B1(new_n688), .B2(new_n678), .ZN(new_n890));
  INV_X1    g704(.A(KEYINPUT113), .ZN(new_n891));
  NAND2_X1  g705(.A1(new_n679), .A2(new_n891), .ZN(new_n892));
  NAND3_X1  g706(.A1(new_n890), .A2(new_n671), .A3(new_n892), .ZN(new_n893));
  AOI21_X1  g707(.A(new_n893), .B1(new_n311), .B2(new_n312), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n669), .B1(new_n894), .B2(KEYINPUT114), .ZN(new_n895));
  INV_X1    g709(.A(new_n893), .ZN(new_n896));
  AND3_X1   g710(.A1(new_n313), .A2(KEYINPUT114), .A3(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n895), .A2(new_n897), .ZN(new_n898));
  AND3_X1   g712(.A1(new_n688), .A2(new_n671), .A3(new_n871), .ZN(new_n899));
  NAND3_X1  g713(.A1(new_n669), .A2(new_n313), .A3(new_n899), .ZN(new_n900));
  NAND3_X1  g714(.A1(new_n706), .A2(new_n656), .A3(new_n900), .ZN(new_n901));
  NOR3_X1   g715(.A1(new_n889), .A2(new_n898), .A3(new_n901), .ZN(new_n902));
  INV_X1    g716(.A(new_n771), .ZN(new_n903));
  AND3_X1   g717(.A1(new_n670), .A2(new_n646), .A3(new_n576), .ZN(new_n904));
  INV_X1    g718(.A(KEYINPUT115), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n731), .A2(new_n905), .A3(new_n719), .ZN(new_n906));
  OAI21_X1  g720(.A(KEYINPUT115), .B1(new_n703), .B2(new_n716), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n460), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n904), .A2(new_n908), .A3(new_n743), .A4(new_n780), .ZN(new_n909));
  NAND4_X1  g723(.A1(new_n722), .A2(new_n749), .A3(new_n903), .A4(new_n909), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT52), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  AND4_X1   g726(.A1(new_n459), .A2(new_n666), .A3(new_n717), .A4(new_n720), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n771), .B1(new_n913), .B2(new_n711), .ZN(new_n914));
  NAND4_X1  g728(.A1(new_n914), .A2(KEYINPUT52), .A3(new_n749), .A4(new_n909), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n912), .A2(new_n915), .ZN(new_n916));
  NAND3_X1  g730(.A1(new_n902), .A2(KEYINPUT53), .A3(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n910), .A2(KEYINPUT116), .A3(KEYINPUT52), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n910), .A2(KEYINPUT116), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(new_n911), .ZN(new_n920));
  AND3_X1   g734(.A1(new_n902), .A2(new_n918), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g735(.A(new_n917), .B1(new_n921), .B2(KEYINPUT53), .ZN(new_n922));
  NAND2_X1  g736(.A1(new_n922), .A2(KEYINPUT54), .ZN(new_n923));
  NAND4_X1  g737(.A1(new_n758), .A2(new_n766), .A3(new_n756), .A4(new_n753), .ZN(new_n924));
  NAND4_X1  g738(.A1(new_n747), .A2(new_n515), .A3(new_n807), .A4(new_n872), .ZN(new_n925));
  NAND3_X1  g739(.A1(new_n792), .A2(new_n925), .A3(new_n867), .ZN(new_n926));
  NOR3_X1   g740(.A1(new_n924), .A2(new_n926), .A3(new_n790), .ZN(new_n927));
  NAND2_X1  g741(.A1(new_n313), .A2(new_n896), .ZN(new_n928));
  INV_X1    g742(.A(KEYINPUT114), .ZN(new_n929));
  NAND2_X1  g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n894), .A2(KEYINPUT114), .ZN(new_n931));
  NAND3_X1  g745(.A1(new_n930), .A2(new_n669), .A3(new_n931), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n706), .A2(new_n656), .A3(new_n900), .ZN(new_n933));
  NAND4_X1  g747(.A1(new_n916), .A2(new_n927), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT53), .ZN(new_n935));
  NAND2_X1  g749(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  INV_X1    g750(.A(KEYINPUT117), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n937), .ZN(new_n938));
  INV_X1    g752(.A(KEYINPUT54), .ZN(new_n939));
  NAND4_X1  g753(.A1(new_n902), .A2(KEYINPUT53), .A3(new_n918), .A4(new_n920), .ZN(new_n940));
  NOR2_X1   g754(.A1(new_n926), .A2(new_n790), .ZN(new_n941));
  NAND4_X1  g755(.A1(new_n933), .A2(new_n941), .A3(new_n932), .A4(new_n888), .ZN(new_n942));
  AND2_X1   g756(.A1(new_n912), .A2(new_n915), .ZN(new_n943));
  OAI211_X1 g757(.A(KEYINPUT117), .B(new_n935), .C1(new_n942), .C2(new_n943), .ZN(new_n944));
  NAND4_X1  g758(.A1(new_n938), .A2(new_n939), .A3(new_n940), .A4(new_n944), .ZN(new_n945));
  NAND2_X1  g759(.A1(new_n923), .A2(new_n945), .ZN(new_n946));
  OAI22_X1  g760(.A1(new_n864), .A2(new_n946), .B1(G952), .B2(G953), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n831), .B(KEYINPUT49), .Z(new_n948));
  NOR3_X1   g762(.A1(new_n948), .A2(new_n865), .A3(new_n810), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n949), .A2(new_n728), .A3(new_n843), .ZN(new_n950));
  NAND2_X1  g764(.A1(new_n947), .A2(new_n950), .ZN(G75));
  XNOR2_X1  g765(.A(new_n243), .B(new_n284), .ZN(new_n952));
  XNOR2_X1  g766(.A(new_n952), .B(KEYINPUT55), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(KEYINPUT56), .ZN(new_n954));
  NAND2_X1  g768(.A1(new_n940), .A2(new_n944), .ZN(new_n955));
  AOI21_X1  g769(.A(KEYINPUT117), .B1(new_n934), .B2(new_n935), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  NAND2_X1  g771(.A1(G210), .A2(G902), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n954), .B1(new_n957), .B2(new_n958), .ZN(new_n959));
  NOR2_X1   g773(.A1(new_n347), .A2(G952), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n959), .A2(new_n961), .ZN(new_n962));
  OAI21_X1  g776(.A(KEYINPUT122), .B1(new_n957), .B2(new_n958), .ZN(new_n963));
  INV_X1    g777(.A(KEYINPUT56), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT122), .ZN(new_n965));
  INV_X1    g779(.A(new_n958), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n965), .B(new_n966), .C1(new_n955), .C2(new_n956), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n963), .A2(new_n964), .A3(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n962), .B1(new_n968), .B2(new_n953), .ZN(G51));
  OAI21_X1  g783(.A(KEYINPUT54), .B1(new_n955), .B2(new_n956), .ZN(new_n970));
  NAND2_X1  g784(.A1(new_n970), .A2(new_n945), .ZN(new_n971));
  XOR2_X1   g785(.A(new_n801), .B(KEYINPUT57), .Z(new_n972));
  NAND2_X1  g786(.A1(new_n971), .A2(new_n972), .ZN(new_n973));
  NAND2_X1  g787(.A1(new_n973), .A2(new_n664), .ZN(new_n974));
  OR3_X1    g788(.A1(new_n957), .A2(new_n287), .A3(new_n800), .ZN(new_n975));
  AOI21_X1  g789(.A(new_n960), .B1(new_n974), .B2(new_n975), .ZN(G54));
  AND2_X1   g790(.A1(KEYINPUT58), .A2(G475), .ZN(new_n977));
  OAI211_X1 g791(.A(G902), .B(new_n977), .C1(new_n955), .C2(new_n956), .ZN(new_n978));
  AND2_X1   g792(.A1(new_n978), .A2(new_n639), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n638), .A2(new_n977), .ZN(new_n980));
  OAI211_X1 g794(.A(G902), .B(new_n980), .C1(new_n955), .C2(new_n956), .ZN(new_n981));
  NAND2_X1  g795(.A1(new_n981), .A2(new_n961), .ZN(new_n982));
  OAI21_X1  g796(.A(KEYINPUT123), .B1(new_n979), .B2(new_n982), .ZN(new_n983));
  NAND2_X1  g797(.A1(new_n978), .A2(new_n639), .ZN(new_n984));
  INV_X1    g798(.A(KEYINPUT123), .ZN(new_n985));
  NAND4_X1  g799(.A1(new_n984), .A2(new_n985), .A3(new_n961), .A4(new_n981), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n983), .A2(new_n986), .ZN(G60));
  NAND2_X1  g801(.A1(new_n673), .A2(new_n674), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(G478), .A2(G902), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT59), .Z(new_n991));
  INV_X1    g805(.A(new_n991), .ZN(new_n992));
  AOI21_X1  g806(.A(new_n989), .B1(new_n946), .B2(new_n992), .ZN(new_n993));
  NAND2_X1  g807(.A1(new_n989), .A2(new_n992), .ZN(new_n994));
  AOI21_X1  g808(.A(new_n994), .B1(new_n970), .B2(new_n945), .ZN(new_n995));
  NOR3_X1   g809(.A1(new_n993), .A2(new_n960), .A3(new_n995), .ZN(G63));
  NAND2_X1  g810(.A1(G217), .A2(G902), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n997), .B(KEYINPUT60), .ZN(new_n998));
  INV_X1    g812(.A(new_n998), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n700), .A2(new_n701), .ZN(new_n1000));
  XOR2_X1   g814(.A(new_n1000), .B(KEYINPUT124), .Z(new_n1001));
  OAI211_X1 g815(.A(new_n999), .B(new_n1001), .C1(new_n955), .C2(new_n956), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n940), .A2(new_n944), .ZN(new_n1003));
  AOI21_X1  g817(.A(new_n998), .B1(new_n1003), .B2(new_n938), .ZN(new_n1004));
  OAI211_X1 g818(.A(new_n961), .B(new_n1002), .C1(new_n1004), .C2(new_n365), .ZN(new_n1005));
  INV_X1    g819(.A(KEYINPUT61), .ZN(new_n1006));
  NAND2_X1  g820(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  OAI22_X1  g821(.A1(new_n957), .A2(new_n998), .B1(new_n364), .B2(new_n363), .ZN(new_n1008));
  NAND4_X1  g822(.A1(new_n1008), .A2(KEYINPUT61), .A3(new_n961), .A4(new_n1002), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1007), .A2(new_n1009), .ZN(G66));
  OAI21_X1  g824(.A(G953), .B1(new_n653), .B2(new_n261), .ZN(new_n1011));
  NOR3_X1   g825(.A1(new_n898), .A2(new_n901), .A3(new_n924), .ZN(new_n1012));
  OAI21_X1  g826(.A(new_n1011), .B1(new_n1012), .B2(G953), .ZN(new_n1013));
  OAI211_X1 g827(.A(new_n240), .B(new_n242), .C1(G898), .C2(new_n347), .ZN(new_n1014));
  XNOR2_X1  g828(.A(new_n1013), .B(new_n1014), .ZN(G69));
  AOI21_X1  g829(.A(new_n347), .B1(G227), .B2(G900), .ZN(new_n1016));
  XOR2_X1   g830(.A(new_n1016), .B(KEYINPUT126), .Z(new_n1017));
  INV_X1    g831(.A(new_n817), .ZN(new_n1018));
  AND2_X1   g832(.A1(new_n822), .A2(new_n1018), .ZN(new_n1019));
  AND2_X1   g833(.A1(new_n854), .A2(new_n904), .ZN(new_n1020));
  NAND4_X1  g834(.A1(new_n805), .A2(new_n459), .A3(new_n724), .A4(new_n1020), .ZN(new_n1021));
  AND2_X1   g835(.A1(new_n914), .A2(new_n749), .ZN(new_n1022));
  AND4_X1   g836(.A1(new_n882), .A2(new_n1021), .A3(new_n792), .A4(new_n1022), .ZN(new_n1023));
  NAND3_X1  g837(.A1(new_n1019), .A2(new_n347), .A3(new_n1023), .ZN(new_n1024));
  NAND3_X1  g838(.A1(new_n436), .A2(new_n437), .A3(new_n438), .ZN(new_n1025));
  XNOR2_X1  g839(.A(new_n1025), .B(new_n634), .ZN(new_n1026));
  NAND2_X1  g840(.A1(G900), .A2(G953), .ZN(new_n1027));
  NAND3_X1  g841(.A1(new_n1024), .A2(new_n1026), .A3(new_n1027), .ZN(new_n1028));
  AOI21_X1  g842(.A(new_n1017), .B1(new_n1028), .B2(KEYINPUT125), .ZN(new_n1029));
  NAND2_X1  g843(.A1(new_n745), .A2(new_n1022), .ZN(new_n1030));
  AND2_X1   g844(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1031));
  NOR2_X1   g845(.A1(new_n1030), .A2(KEYINPUT62), .ZN(new_n1032));
  AOI22_X1  g846(.A1(new_n890), .A2(new_n892), .B1(new_n688), .B2(new_n871), .ZN(new_n1033));
  NOR4_X1   g847(.A1(new_n725), .A2(new_n1033), .A3(new_n808), .A4(new_n880), .ZN(new_n1034));
  NOR3_X1   g848(.A1(new_n1031), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(G953), .B1(new_n1035), .B2(new_n1019), .ZN(new_n1036));
  OAI21_X1  g850(.A(new_n1028), .B1(new_n1036), .B2(new_n1026), .ZN(new_n1037));
  NAND2_X1  g851(.A1(new_n1029), .A2(new_n1037), .ZN(new_n1038));
  OAI221_X1 g852(.A(new_n1028), .B1(KEYINPUT125), .B2(new_n1017), .C1(new_n1036), .C2(new_n1026), .ZN(new_n1039));
  AND2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  NAND3_X1  g854(.A1(new_n1035), .A2(new_n1019), .A3(new_n1012), .ZN(new_n1041));
  XNOR2_X1  g855(.A(KEYINPUT127), .B(KEYINPUT63), .ZN(new_n1042));
  NAND2_X1  g856(.A1(G472), .A2(G902), .ZN(new_n1043));
  XNOR2_X1  g857(.A(new_n1042), .B(new_n1043), .ZN(new_n1044));
  AOI211_X1 g858(.A(new_n446), .B(new_n738), .C1(new_n1041), .C2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g859(.A(new_n738), .B(new_n414), .ZN(new_n1046));
  AND3_X1   g860(.A1(new_n922), .A2(new_n1044), .A3(new_n1046), .ZN(new_n1047));
  NAND2_X1  g861(.A1(new_n738), .A2(new_n446), .ZN(new_n1048));
  NAND3_X1  g862(.A1(new_n1019), .A2(new_n1012), .A3(new_n1023), .ZN(new_n1049));
  AOI21_X1  g863(.A(new_n1048), .B1(new_n1049), .B2(new_n1044), .ZN(new_n1050));
  NOR4_X1   g864(.A1(new_n1045), .A2(new_n1047), .A3(new_n960), .A4(new_n1050), .ZN(G57));
endmodule


