//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 0 0 0 0 1 1 0 1 0 1 1 1 1 1 0 1 0 1 1 0 1 0 0 0 0 0 0 0 1 1 1 0 1 0 1 0 0 0 1 1 0 0 1 0 1 0 0 1 0 0 0 0 1 1 1 1 1 0 1 1 1 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:18 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n679,
    new_n680, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n732, new_n734,
    new_n735, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n744, new_n745, new_n746, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n758, new_n759, new_n760, new_n761, new_n762, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n785, new_n786, new_n787,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n957, new_n958, new_n959, new_n960, new_n961, new_n962,
    new_n963, new_n965, new_n966, new_n967, new_n968, new_n969, new_n970,
    new_n971, new_n972, new_n973, new_n974, new_n975, new_n976, new_n977,
    new_n978, new_n979, new_n981, new_n982, new_n983, new_n984, new_n985,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n995, new_n996, new_n997, new_n998, new_n999, new_n1000,
    new_n1001, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  XNOR2_X1  g001(.A(KEYINPUT69), .B(G902), .ZN(new_n188));
  INV_X1    g002(.A(G146), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G143), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G143), .ZN(new_n192));
  AOI21_X1  g006(.A(new_n191), .B1(new_n192), .B2(G146), .ZN(new_n193));
  NOR3_X1   g007(.A1(new_n189), .A2(KEYINPUT64), .A3(G143), .ZN(new_n194));
  OAI21_X1  g008(.A(new_n190), .B1(new_n193), .B2(new_n194), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n192), .A2(G146), .ZN(new_n196));
  INV_X1    g010(.A(KEYINPUT1), .ZN(new_n197));
  OAI21_X1  g011(.A(G128), .B1(new_n196), .B2(new_n197), .ZN(new_n198));
  NAND3_X1  g012(.A1(new_n195), .A2(KEYINPUT76), .A3(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(KEYINPUT76), .ZN(new_n200));
  OAI21_X1  g014(.A(KEYINPUT64), .B1(new_n189), .B2(G143), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n192), .A3(G146), .ZN(new_n202));
  AOI21_X1  g016(.A(new_n196), .B1(new_n201), .B2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(G128), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n190), .B2(KEYINPUT1), .ZN(new_n205));
  OAI21_X1  g019(.A(new_n200), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(new_n204), .A2(KEYINPUT1), .ZN(new_n207));
  OAI211_X1 g021(.A(new_n190), .B(new_n207), .C1(new_n193), .C2(new_n194), .ZN(new_n208));
  NAND3_X1  g022(.A1(new_n199), .A2(new_n206), .A3(new_n208), .ZN(new_n209));
  INV_X1    g023(.A(G104), .ZN(new_n210));
  OAI21_X1  g024(.A(KEYINPUT3), .B1(new_n210), .B2(G107), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT3), .ZN(new_n212));
  INV_X1    g026(.A(G107), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n212), .A2(new_n213), .A3(G104), .ZN(new_n214));
  INV_X1    g028(.A(G101), .ZN(new_n215));
  NAND2_X1  g029(.A1(new_n210), .A2(G107), .ZN(new_n216));
  NAND4_X1  g030(.A1(new_n211), .A2(new_n214), .A3(new_n215), .A4(new_n216), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n210), .A2(G107), .ZN(new_n218));
  NOR2_X1   g032(.A1(new_n213), .A2(G104), .ZN(new_n219));
  OAI21_X1  g033(.A(G101), .B1(new_n218), .B2(new_n219), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n217), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g035(.A1(new_n209), .A2(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(KEYINPUT10), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n222), .A2(new_n223), .ZN(new_n224));
  NAND3_X1  g038(.A1(new_n211), .A2(new_n214), .A3(new_n216), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G101), .ZN(new_n226));
  NAND3_X1  g040(.A1(new_n226), .A2(KEYINPUT4), .A3(new_n217), .ZN(new_n227));
  NAND2_X1  g041(.A1(KEYINPUT0), .A2(G128), .ZN(new_n228));
  INV_X1    g042(.A(new_n228), .ZN(new_n229));
  OR2_X1    g043(.A1(KEYINPUT0), .A2(G128), .ZN(new_n230));
  AND2_X1   g044(.A1(new_n230), .A2(new_n228), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n192), .A2(G146), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n190), .A2(new_n232), .ZN(new_n233));
  AOI22_X1  g047(.A1(new_n203), .A2(new_n229), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT4), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n225), .A2(new_n235), .A3(G101), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(new_n234), .A3(new_n236), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n197), .B1(G143), .B2(new_n189), .ZN(new_n238));
  OAI21_X1  g052(.A(new_n233), .B1(new_n238), .B2(new_n204), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n208), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n240), .A2(new_n221), .A3(KEYINPUT10), .ZN(new_n241));
  AND2_X1   g055(.A1(new_n237), .A2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT11), .ZN(new_n243));
  INV_X1    g057(.A(G134), .ZN(new_n244));
  OAI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(G137), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n244), .A2(G137), .ZN(new_n246));
  INV_X1    g060(.A(G137), .ZN(new_n247));
  NAND3_X1  g061(.A1(new_n247), .A2(KEYINPUT11), .A3(G134), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n245), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n249), .A2(G131), .ZN(new_n250));
  INV_X1    g064(.A(G131), .ZN(new_n251));
  NAND4_X1  g065(.A1(new_n245), .A2(new_n248), .A3(new_n251), .A4(new_n246), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n250), .A2(new_n252), .ZN(new_n253));
  INV_X1    g067(.A(new_n253), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n224), .A2(new_n242), .A3(new_n254), .ZN(new_n255));
  XNOR2_X1  g069(.A(G110), .B(G140), .ZN(new_n256));
  INV_X1    g070(.A(G227), .ZN(new_n257));
  NOR2_X1   g071(.A1(new_n257), .A2(G953), .ZN(new_n258));
  XNOR2_X1  g072(.A(new_n256), .B(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n259), .ZN(new_n260));
  NAND2_X1  g074(.A1(new_n255), .A2(new_n260), .ZN(new_n261));
  NOR2_X1   g075(.A1(new_n240), .A2(new_n221), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND2_X1  g077(.A1(new_n222), .A2(new_n263), .ZN(new_n264));
  NAND4_X1  g078(.A1(new_n264), .A2(KEYINPUT77), .A3(KEYINPUT12), .A4(new_n253), .ZN(new_n265));
  INV_X1    g079(.A(KEYINPUT77), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n221), .B2(new_n209), .ZN(new_n267));
  NAND2_X1  g081(.A1(new_n253), .A2(KEYINPUT12), .ZN(new_n268));
  OAI21_X1  g082(.A(new_n266), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  AND2_X1   g083(.A1(new_n265), .A2(new_n269), .ZN(new_n270));
  INV_X1    g084(.A(KEYINPUT12), .ZN(new_n271));
  OAI21_X1  g085(.A(new_n253), .B1(new_n267), .B2(KEYINPUT78), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n222), .A2(new_n263), .A3(KEYINPUT78), .ZN(new_n273));
  OAI21_X1  g087(.A(new_n271), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  AOI21_X1  g088(.A(new_n261), .B1(new_n270), .B2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n224), .A2(new_n242), .A3(KEYINPUT79), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT79), .ZN(new_n277));
  AOI21_X1  g091(.A(KEYINPUT10), .B1(new_n209), .B2(new_n221), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n237), .A2(new_n241), .ZN(new_n279));
  OAI21_X1  g093(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n276), .A2(new_n253), .A3(new_n280), .ZN(new_n281));
  AOI21_X1  g095(.A(new_n260), .B1(new_n281), .B2(new_n255), .ZN(new_n282));
  OAI211_X1 g096(.A(new_n187), .B(new_n188), .C1(new_n275), .C2(new_n282), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT80), .ZN(new_n284));
  NAND2_X1  g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n281), .A2(new_n255), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n286), .A2(new_n259), .ZN(new_n287));
  INV_X1    g101(.A(new_n261), .ZN(new_n288));
  INV_X1    g102(.A(KEYINPUT78), .ZN(new_n289));
  AOI21_X1  g103(.A(new_n254), .B1(new_n264), .B2(new_n289), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n267), .A2(KEYINPUT78), .ZN(new_n291));
  AOI21_X1  g105(.A(KEYINPUT12), .B1(new_n290), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g106(.A1(new_n265), .A2(new_n269), .ZN(new_n293));
  OAI21_X1  g107(.A(new_n288), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n287), .A2(new_n294), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n295), .A2(KEYINPUT80), .A3(new_n187), .A4(new_n188), .ZN(new_n296));
  INV_X1    g110(.A(G902), .ZN(new_n297));
  XOR2_X1   g111(.A(new_n259), .B(KEYINPUT75), .Z(new_n298));
  NAND2_X1  g112(.A1(new_n270), .A2(new_n274), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n298), .B1(new_n299), .B2(new_n255), .ZN(new_n300));
  AND2_X1   g114(.A1(new_n288), .A2(new_n281), .ZN(new_n301));
  OAI21_X1  g115(.A(new_n297), .B1(new_n300), .B2(new_n301), .ZN(new_n302));
  AOI22_X1  g116(.A1(new_n285), .A2(new_n296), .B1(new_n302), .B2(G469), .ZN(new_n303));
  XNOR2_X1  g117(.A(KEYINPUT9), .B(G234), .ZN(new_n304));
  OAI21_X1  g118(.A(G221), .B1(new_n304), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  OAI21_X1  g120(.A(G214), .B1(G237), .B2(G902), .ZN(new_n307));
  INV_X1    g121(.A(new_n307), .ZN(new_n308));
  OAI21_X1  g122(.A(G210), .B1(G237), .B2(G902), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  XOR2_X1   g124(.A(KEYINPUT2), .B(G113), .Z(new_n311));
  XNOR2_X1  g125(.A(G116), .B(G119), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n311), .B(new_n312), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n313), .A2(new_n227), .A3(new_n236), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n311), .A2(new_n312), .ZN(new_n315));
  INV_X1    g129(.A(G119), .ZN(new_n316));
  NAND2_X1  g130(.A1(new_n316), .A2(G116), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NOR2_X1   g132(.A1(new_n316), .A2(G116), .ZN(new_n319));
  INV_X1    g133(.A(KEYINPUT5), .ZN(new_n320));
  NOR3_X1   g134(.A1(new_n318), .A2(new_n319), .A3(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(G113), .B1(new_n317), .B2(KEYINPUT5), .ZN(new_n322));
  OAI211_X1 g136(.A(new_n221), .B(new_n315), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n314), .A2(new_n323), .ZN(new_n324));
  XNOR2_X1  g138(.A(G110), .B(G122), .ZN(new_n325));
  INV_X1    g139(.A(new_n325), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n314), .A2(new_n323), .A3(new_n325), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(KEYINPUT6), .A3(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(KEYINPUT6), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n324), .A2(new_n330), .A3(new_n326), .ZN(new_n331));
  NAND3_X1  g145(.A1(new_n233), .A2(new_n228), .A3(new_n230), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT70), .B(G125), .ZN(new_n333));
  OAI211_X1 g147(.A(new_n332), .B(new_n333), .C1(new_n195), .C2(new_n228), .ZN(new_n334));
  AOI22_X1  g148(.A1(new_n203), .A2(new_n207), .B1(new_n198), .B2(new_n233), .ZN(new_n335));
  OAI21_X1  g149(.A(new_n334), .B1(new_n335), .B2(new_n333), .ZN(new_n336));
  INV_X1    g150(.A(G953), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n337), .A2(G224), .ZN(new_n338));
  XNOR2_X1  g152(.A(new_n336), .B(new_n338), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n329), .A2(new_n331), .A3(new_n339), .ZN(new_n340));
  INV_X1    g154(.A(new_n340), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n338), .A2(KEYINPUT7), .ZN(new_n342));
  OAI211_X1 g156(.A(new_n334), .B(new_n342), .C1(new_n335), .C2(new_n333), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n217), .A2(new_n220), .ZN(new_n344));
  NAND2_X1  g158(.A1(new_n322), .A2(KEYINPUT81), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n312), .A2(KEYINPUT5), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT81), .ZN(new_n347));
  OAI211_X1 g161(.A(new_n347), .B(G113), .C1(new_n317), .C2(KEYINPUT5), .ZN(new_n348));
  NAND3_X1  g162(.A1(new_n345), .A2(new_n346), .A3(new_n348), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n344), .B1(new_n349), .B2(new_n315), .ZN(new_n350));
  XNOR2_X1  g164(.A(new_n325), .B(KEYINPUT8), .ZN(new_n351));
  OAI21_X1  g165(.A(new_n315), .B1(new_n321), .B2(new_n322), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(new_n221), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n343), .B1(new_n350), .B2(new_n353), .ZN(new_n354));
  INV_X1    g168(.A(KEYINPUT82), .ZN(new_n355));
  INV_X1    g169(.A(new_n342), .ZN(new_n356));
  AOI21_X1  g170(.A(new_n355), .B1(new_n336), .B2(new_n356), .ZN(new_n357));
  NOR2_X1   g171(.A1(new_n354), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n336), .A2(new_n355), .A3(new_n356), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n358), .A2(new_n328), .A3(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n297), .ZN(new_n361));
  OAI21_X1  g175(.A(new_n310), .B1(new_n341), .B2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(new_n359), .ZN(new_n363));
  NOR3_X1   g177(.A1(new_n363), .A2(new_n354), .A3(new_n357), .ZN(new_n364));
  AOI21_X1  g178(.A(G902), .B1(new_n364), .B2(new_n328), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n365), .A2(new_n309), .A3(new_n340), .ZN(new_n366));
  AOI21_X1  g180(.A(new_n308), .B1(new_n362), .B2(new_n366), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n337), .A2(G952), .ZN(new_n368));
  INV_X1    g182(.A(G234), .ZN(new_n369));
  INV_X1    g183(.A(G237), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n368), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI211_X1 g186(.A(new_n337), .B(new_n188), .C1(G234), .C2(G237), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT21), .B(G898), .ZN(new_n374));
  AOI21_X1  g188(.A(new_n372), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n376), .ZN(new_n377));
  INV_X1    g191(.A(G475), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT85), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n192), .A2(KEYINPUT84), .ZN(new_n380));
  NOR2_X1   g194(.A1(G237), .A2(G953), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n380), .A2(G214), .A3(new_n381), .ZN(new_n382));
  NAND3_X1  g196(.A1(new_n370), .A2(new_n337), .A3(G214), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  XNOR2_X1  g198(.A(KEYINPUT84), .B(G143), .ZN(new_n385));
  OAI211_X1 g199(.A(new_n379), .B(new_n382), .C1(new_n384), .C2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(KEYINPUT18), .A2(G131), .ZN(new_n387));
  XNOR2_X1  g201(.A(new_n386), .B(new_n387), .ZN(new_n388));
  XNOR2_X1  g202(.A(G125), .B(G140), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(new_n189), .ZN(new_n390));
  NOR2_X1   g204(.A1(G125), .A2(G140), .ZN(new_n391));
  AOI21_X1  g205(.A(new_n391), .B1(new_n333), .B2(G140), .ZN(new_n392));
  INV_X1    g206(.A(new_n392), .ZN(new_n393));
  OAI21_X1  g207(.A(new_n390), .B1(new_n393), .B2(new_n189), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n388), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT84), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(G143), .ZN(new_n397));
  AOI22_X1  g211(.A1(new_n397), .A2(new_n380), .B1(new_n381), .B2(G214), .ZN(new_n398));
  NOR2_X1   g212(.A1(new_n396), .A2(G143), .ZN(new_n399));
  NOR2_X1   g213(.A1(new_n383), .A2(new_n399), .ZN(new_n400));
  OAI21_X1  g214(.A(G131), .B1(new_n398), .B2(new_n400), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT17), .ZN(new_n402));
  OAI211_X1 g216(.A(new_n251), .B(new_n382), .C1(new_n384), .C2(new_n385), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND2_X1  g218(.A1(new_n404), .A2(KEYINPUT90), .ZN(new_n405));
  INV_X1    g219(.A(KEYINPUT90), .ZN(new_n406));
  NAND4_X1  g220(.A1(new_n401), .A2(new_n406), .A3(new_n403), .A4(new_n402), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n405), .A2(new_n407), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT16), .ZN(new_n409));
  INV_X1    g223(.A(G140), .ZN(new_n410));
  NAND3_X1  g224(.A1(new_n333), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  OAI21_X1  g225(.A(new_n411), .B1(new_n392), .B2(new_n409), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n412), .A2(new_n189), .ZN(new_n413));
  OAI211_X1 g227(.A(G146), .B(new_n411), .C1(new_n392), .C2(new_n409), .ZN(new_n414));
  OAI211_X1 g228(.A(KEYINPUT17), .B(G131), .C1(new_n398), .C2(new_n400), .ZN(new_n415));
  NAND3_X1  g229(.A1(new_n413), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n395), .B1(new_n408), .B2(new_n416), .ZN(new_n417));
  XNOR2_X1  g231(.A(G113), .B(G122), .ZN(new_n418));
  XNOR2_X1  g232(.A(new_n418), .B(new_n210), .ZN(new_n419));
  INV_X1    g233(.A(new_n419), .ZN(new_n420));
  NAND2_X1  g234(.A1(new_n417), .A2(new_n420), .ZN(new_n421));
  INV_X1    g235(.A(KEYINPUT89), .ZN(new_n422));
  XNOR2_X1  g236(.A(new_n419), .B(new_n422), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n395), .B(new_n423), .C1(new_n408), .C2(new_n416), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n421), .A2(new_n424), .ZN(new_n425));
  AOI21_X1  g239(.A(new_n378), .B1(new_n425), .B2(new_n297), .ZN(new_n426));
  XOR2_X1   g240(.A(KEYINPUT83), .B(KEYINPUT20), .Z(new_n427));
  INV_X1    g241(.A(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(new_n424), .ZN(new_n429));
  AND2_X1   g243(.A1(KEYINPUT70), .A2(G125), .ZN(new_n430));
  NOR2_X1   g244(.A1(KEYINPUT70), .A2(G125), .ZN(new_n431));
  OAI21_X1  g245(.A(G140), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n391), .ZN(new_n433));
  NAND3_X1  g247(.A1(new_n432), .A2(KEYINPUT19), .A3(new_n433), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n389), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n434), .A2(new_n189), .A3(new_n436), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n437), .A2(KEYINPUT87), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT87), .ZN(new_n439));
  NAND4_X1  g253(.A1(new_n434), .A2(new_n439), .A3(new_n189), .A4(new_n436), .ZN(new_n440));
  NAND4_X1  g254(.A1(new_n438), .A2(KEYINPUT88), .A3(new_n414), .A4(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n401), .A2(new_n403), .ZN(new_n442));
  INV_X1    g256(.A(KEYINPUT86), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g258(.A1(new_n401), .A2(KEYINPUT86), .A3(new_n403), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n441), .A2(new_n444), .A3(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n414), .A2(new_n440), .ZN(new_n447));
  INV_X1    g261(.A(new_n447), .ZN(new_n448));
  AOI21_X1  g262(.A(KEYINPUT88), .B1(new_n448), .B2(new_n438), .ZN(new_n449));
  OAI21_X1  g263(.A(new_n395), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n429), .B1(new_n450), .B2(new_n420), .ZN(new_n451));
  NOR2_X1   g265(.A1(G475), .A2(G902), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  OAI21_X1  g267(.A(new_n428), .B1(new_n451), .B2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT20), .ZN(new_n455));
  INV_X1    g269(.A(KEYINPUT88), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n437), .A2(KEYINPUT87), .ZN(new_n457));
  OAI21_X1  g271(.A(new_n456), .B1(new_n457), .B2(new_n447), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n458), .A2(new_n441), .A3(new_n444), .A4(new_n445), .ZN(new_n459));
  AOI21_X1  g273(.A(new_n419), .B1(new_n459), .B2(new_n395), .ZN(new_n460));
  OAI211_X1 g274(.A(new_n455), .B(new_n452), .C1(new_n460), .C2(new_n429), .ZN(new_n461));
  AOI21_X1  g275(.A(new_n426), .B1(new_n454), .B2(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(KEYINPUT13), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n204), .B2(G143), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n192), .A2(KEYINPUT13), .A3(G128), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n204), .A2(G143), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n464), .A2(new_n465), .A3(new_n466), .ZN(new_n467));
  NAND2_X1  g281(.A1(new_n467), .A2(G134), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n192), .A2(G128), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n469), .A2(new_n466), .A3(new_n244), .ZN(new_n470));
  INV_X1    g284(.A(G122), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n471), .A2(G116), .ZN(new_n472));
  INV_X1    g286(.A(G116), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n473), .A2(G122), .ZN(new_n474));
  AOI21_X1  g288(.A(new_n213), .B1(new_n472), .B2(new_n474), .ZN(new_n475));
  AND3_X1   g289(.A1(new_n472), .A2(new_n474), .A3(new_n213), .ZN(new_n476));
  OAI211_X1 g290(.A(new_n468), .B(new_n470), .C1(new_n475), .C2(new_n476), .ZN(new_n477));
  NOR2_X1   g291(.A1(new_n204), .A2(G143), .ZN(new_n478));
  NOR2_X1   g292(.A1(new_n192), .A2(G128), .ZN(new_n479));
  OAI21_X1  g293(.A(G134), .B1(new_n478), .B2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n480), .A2(new_n470), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n473), .A2(KEYINPUT14), .A3(G122), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n472), .A2(new_n474), .ZN(new_n483));
  OAI211_X1 g297(.A(G107), .B(new_n482), .C1(new_n483), .C2(KEYINPUT14), .ZN(new_n484));
  XNOR2_X1  g298(.A(G116), .B(G122), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(new_n213), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n481), .A2(new_n484), .A3(new_n486), .ZN(new_n487));
  INV_X1    g301(.A(G217), .ZN(new_n488));
  NOR3_X1   g302(.A1(new_n304), .A2(new_n488), .A3(G953), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n477), .A2(new_n487), .A3(new_n489), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  AOI21_X1  g305(.A(new_n489), .B1(new_n477), .B2(new_n487), .ZN(new_n492));
  OAI21_X1  g306(.A(new_n188), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G478), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n494), .A2(KEYINPUT15), .ZN(new_n495));
  XNOR2_X1  g309(.A(new_n493), .B(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n462), .A2(new_n497), .ZN(new_n498));
  NOR4_X1   g312(.A1(new_n303), .A2(new_n306), .A3(new_n377), .A4(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n488), .B1(new_n188), .B2(G234), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  NOR2_X1   g315(.A1(KEYINPUT74), .A2(KEYINPUT25), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n337), .A2(G221), .A3(G234), .ZN(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(KEYINPUT72), .ZN(new_n504));
  XNOR2_X1  g318(.A(KEYINPUT22), .B(G137), .ZN(new_n505));
  XNOR2_X1  g319(.A(new_n504), .B(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  NAND2_X1  g321(.A1(new_n316), .A2(G128), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n204), .A2(G119), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g324(.A(KEYINPUT24), .B(G110), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT71), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n510), .A2(new_n511), .A3(KEYINPUT71), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n204), .A2(KEYINPUT23), .A3(G119), .ZN(new_n516));
  INV_X1    g330(.A(new_n509), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n508), .B(new_n516), .C1(new_n517), .C2(KEYINPUT23), .ZN(new_n518));
  OAI211_X1 g332(.A(new_n514), .B(new_n515), .C1(G110), .C2(new_n518), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n519), .A2(new_n414), .A3(new_n390), .ZN(new_n520));
  INV_X1    g334(.A(new_n520), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n518), .A2(G110), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n510), .B2(new_n511), .ZN(new_n523));
  AOI21_X1  g337(.A(new_n523), .B1(new_n413), .B2(new_n414), .ZN(new_n524));
  OAI21_X1  g338(.A(KEYINPUT73), .B1(new_n521), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n413), .A2(new_n414), .ZN(new_n526));
  INV_X1    g340(.A(new_n523), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT73), .ZN(new_n529));
  NAND3_X1  g343(.A1(new_n528), .A2(new_n529), .A3(new_n520), .ZN(new_n530));
  AOI21_X1  g344(.A(new_n507), .B1(new_n525), .B2(new_n530), .ZN(new_n531));
  NAND2_X1  g345(.A1(new_n528), .A2(new_n520), .ZN(new_n532));
  AOI21_X1  g346(.A(new_n506), .B1(new_n532), .B2(KEYINPUT73), .ZN(new_n533));
  OR2_X1    g347(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n188), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n502), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  NOR4_X1   g350(.A1(new_n531), .A2(new_n533), .A3(new_n535), .A4(new_n502), .ZN(new_n537));
  INV_X1    g351(.A(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n501), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NOR2_X1   g353(.A1(new_n531), .A2(new_n533), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n500), .A2(G902), .ZN(new_n541));
  AND2_X1   g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  OR2_X1    g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n234), .A2(new_n253), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n247), .A2(G134), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n244), .A2(G137), .ZN(new_n546));
  OAI21_X1  g360(.A(G131), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n252), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n240), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n544), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n550), .A2(new_n313), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n551), .A2(KEYINPUT28), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n550), .A2(new_n313), .ZN(new_n553));
  AOI22_X1  g367(.A1(new_n253), .A2(new_n234), .B1(new_n240), .B2(new_n548), .ZN(new_n554));
  INV_X1    g368(.A(new_n313), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n552), .B1(new_n557), .B2(KEYINPUT28), .ZN(new_n558));
  NAND2_X1  g372(.A1(new_n381), .A2(G210), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n559), .B(KEYINPUT27), .ZN(new_n560));
  XNOR2_X1  g374(.A(KEYINPUT26), .B(G101), .ZN(new_n561));
  XNOR2_X1  g375(.A(new_n560), .B(new_n561), .ZN(new_n562));
  AOI21_X1  g376(.A(KEYINPUT29), .B1(new_n558), .B2(new_n562), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT67), .ZN(new_n564));
  INV_X1    g378(.A(new_n562), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n544), .A2(new_n549), .A3(KEYINPUT30), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n566), .A2(new_n313), .ZN(new_n567));
  OAI21_X1  g381(.A(KEYINPUT65), .B1(new_n554), .B2(KEYINPUT30), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT65), .ZN(new_n569));
  INV_X1    g383(.A(KEYINPUT30), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n550), .A2(new_n569), .A3(new_n570), .ZN(new_n571));
  AOI21_X1  g385(.A(new_n567), .B1(new_n568), .B2(new_n571), .ZN(new_n572));
  OAI211_X1 g386(.A(new_n564), .B(new_n565), .C1(new_n572), .C2(new_n551), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n568), .A2(new_n571), .ZN(new_n574));
  AOI21_X1  g388(.A(new_n555), .B1(new_n554), .B2(KEYINPUT30), .ZN(new_n575));
  AOI21_X1  g389(.A(new_n551), .B1(new_n574), .B2(new_n575), .ZN(new_n576));
  OAI21_X1  g390(.A(KEYINPUT67), .B1(new_n576), .B2(new_n562), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n563), .A2(new_n573), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n578), .A2(KEYINPUT68), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT68), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n563), .A2(new_n577), .A3(new_n580), .A4(new_n573), .ZN(new_n581));
  NAND3_X1  g395(.A1(new_n558), .A2(KEYINPUT29), .A3(new_n562), .ZN(new_n582));
  NAND4_X1  g396(.A1(new_n579), .A2(new_n581), .A3(new_n582), .A4(new_n188), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(G472), .ZN(new_n584));
  INV_X1    g398(.A(G472), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(new_n297), .ZN(new_n586));
  INV_X1    g400(.A(KEYINPUT31), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n556), .A2(new_n562), .ZN(new_n588));
  OAI21_X1  g402(.A(new_n587), .B1(new_n572), .B2(new_n588), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n569), .B1(new_n550), .B2(new_n570), .ZN(new_n590));
  AOI211_X1 g404(.A(KEYINPUT65), .B(KEYINPUT30), .C1(new_n544), .C2(new_n549), .ZN(new_n591));
  OAI21_X1  g405(.A(new_n575), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(new_n588), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(KEYINPUT31), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g408(.A1(new_n589), .A2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT28), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n556), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n557), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n597), .B1(new_n598), .B2(new_n596), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(new_n565), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n586), .B1(new_n595), .B2(new_n600), .ZN(new_n601));
  OAI21_X1  g415(.A(KEYINPUT66), .B1(new_n601), .B2(KEYINPUT32), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n601), .A2(KEYINPUT32), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT66), .ZN(new_n604));
  INV_X1    g418(.A(KEYINPUT32), .ZN(new_n605));
  AOI22_X1  g419(.A1(new_n589), .A2(new_n594), .B1(new_n599), .B2(new_n565), .ZN(new_n606));
  OAI211_X1 g420(.A(new_n604), .B(new_n605), .C1(new_n606), .C2(new_n586), .ZN(new_n607));
  AND3_X1   g421(.A1(new_n602), .A2(new_n603), .A3(new_n607), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n543), .B1(new_n584), .B2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n499), .A2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(G101), .ZN(G3));
  AOI21_X1  g425(.A(new_n535), .B1(new_n595), .B2(new_n600), .ZN(new_n612));
  OAI22_X1  g426(.A1(new_n612), .A2(new_n585), .B1(new_n586), .B2(new_n606), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n543), .A2(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n285), .A2(new_n296), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n302), .A2(G469), .ZN(new_n616));
  AOI21_X1  g430(.A(new_n306), .B1(new_n615), .B2(new_n616), .ZN(new_n617));
  AOI21_X1  g431(.A(KEYINPUT92), .B1(new_n493), .B2(new_n494), .ZN(new_n618));
  INV_X1    g432(.A(new_n468), .ZN(new_n619));
  OAI21_X1  g433(.A(new_n470), .B1(new_n476), .B2(new_n475), .ZN(new_n620));
  AND3_X1   g434(.A1(new_n469), .A2(new_n466), .A3(new_n244), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n244), .B1(new_n469), .B2(new_n466), .ZN(new_n622));
  OAI21_X1  g436(.A(new_n486), .B1(new_n621), .B2(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n482), .A2(G107), .ZN(new_n624));
  INV_X1    g438(.A(KEYINPUT14), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n624), .B1(new_n625), .B2(new_n485), .ZN(new_n626));
  OAI22_X1  g440(.A1(new_n619), .A2(new_n620), .B1(new_n623), .B2(new_n626), .ZN(new_n627));
  INV_X1    g441(.A(new_n489), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n629), .A2(new_n490), .ZN(new_n630));
  INV_X1    g444(.A(new_n475), .ZN(new_n631));
  AOI21_X1  g445(.A(new_n621), .B1(new_n631), .B2(new_n486), .ZN(new_n632));
  AOI22_X1  g446(.A1(new_n480), .A2(new_n470), .B1(new_n213), .B2(new_n485), .ZN(new_n633));
  AOI22_X1  g447(.A1(new_n632), .A2(new_n468), .B1(new_n633), .B2(new_n484), .ZN(new_n634));
  OAI21_X1  g448(.A(KEYINPUT91), .B1(new_n634), .B2(new_n489), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n630), .A2(new_n635), .A3(KEYINPUT33), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT33), .ZN(new_n637));
  OAI211_X1 g451(.A(new_n629), .B(new_n490), .C1(KEYINPUT91), .C2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n636), .A2(new_n638), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n535), .A2(new_n494), .ZN(new_n640));
  AOI21_X1  g454(.A(new_n618), .B1(new_n639), .B2(new_n640), .ZN(new_n641));
  INV_X1    g455(.A(new_n640), .ZN(new_n642));
  AOI211_X1 g456(.A(KEYINPUT92), .B(new_n642), .C1(new_n636), .C2(new_n638), .ZN(new_n643));
  OAI21_X1  g457(.A(KEYINPUT93), .B1(new_n641), .B2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(KEYINPUT92), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n639), .A2(new_n645), .A3(new_n640), .ZN(new_n646));
  INV_X1    g460(.A(KEYINPUT93), .ZN(new_n647));
  AOI21_X1  g461(.A(new_n642), .B1(new_n636), .B2(new_n638), .ZN(new_n648));
  OAI211_X1 g462(.A(new_n646), .B(new_n647), .C1(new_n648), .C2(new_n618), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n644), .A2(new_n649), .ZN(new_n650));
  NOR3_X1   g464(.A1(new_n377), .A2(new_n462), .A3(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n614), .A2(new_n617), .A3(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(KEYINPUT34), .B(G104), .Z(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(G6));
  INV_X1    g468(.A(KEYINPUT94), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n426), .B(new_n655), .ZN(new_n656));
  NAND2_X1  g470(.A1(new_n450), .A2(new_n420), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n657), .A2(new_n424), .ZN(new_n658));
  NAND3_X1  g472(.A1(new_n658), .A2(new_n452), .A3(new_n427), .ZN(new_n659));
  NAND2_X1  g473(.A1(new_n659), .A2(new_n454), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  NOR3_X1   g475(.A1(new_n661), .A2(new_n377), .A3(new_n497), .ZN(new_n662));
  NAND3_X1  g476(.A1(new_n614), .A2(new_n617), .A3(new_n662), .ZN(new_n663));
  XOR2_X1   g477(.A(KEYINPUT35), .B(G107), .Z(new_n664));
  XNOR2_X1  g478(.A(new_n663), .B(new_n664), .ZN(G9));
  INV_X1    g479(.A(new_n502), .ZN(new_n666));
  AOI21_X1  g480(.A(new_n666), .B1(new_n540), .B2(new_n188), .ZN(new_n667));
  OAI21_X1  g481(.A(new_n500), .B1(new_n667), .B2(new_n537), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n506), .A2(KEYINPUT36), .ZN(new_n669));
  XNOR2_X1  g483(.A(new_n532), .B(new_n669), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n541), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n668), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR2_X1   g487(.A1(new_n673), .A2(new_n613), .ZN(new_n674));
  INV_X1    g488(.A(KEYINPUT95), .ZN(new_n675));
  NAND2_X1  g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  OAI21_X1  g490(.A(KEYINPUT95), .B1(new_n673), .B2(new_n613), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n499), .A2(new_n676), .A3(new_n677), .ZN(new_n678));
  XOR2_X1   g492(.A(KEYINPUT37), .B(G110), .Z(new_n679));
  XNOR2_X1  g493(.A(new_n679), .B(KEYINPUT96), .ZN(new_n680));
  XNOR2_X1  g494(.A(new_n678), .B(new_n680), .ZN(G12));
  NAND2_X1  g495(.A1(new_n672), .A2(new_n367), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n682), .B1(new_n584), .B2(new_n608), .ZN(new_n683));
  INV_X1    g497(.A(G900), .ZN(new_n684));
  AOI21_X1  g498(.A(new_n372), .B1(new_n373), .B2(new_n684), .ZN(new_n685));
  INV_X1    g499(.A(new_n685), .ZN(new_n686));
  NAND4_X1  g500(.A1(new_n656), .A2(new_n496), .A3(new_n660), .A4(new_n686), .ZN(new_n687));
  NOR3_X1   g501(.A1(new_n303), .A2(new_n687), .A3(new_n306), .ZN(new_n688));
  NAND2_X1  g502(.A1(new_n683), .A2(new_n688), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT97), .B(G128), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G30));
  INV_X1    g505(.A(new_n426), .ZN(new_n692));
  AOI21_X1  g506(.A(new_n427), .B1(new_n658), .B2(new_n452), .ZN(new_n693));
  INV_X1    g507(.A(new_n461), .ZN(new_n694));
  OAI21_X1  g508(.A(new_n692), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  AOI21_X1  g509(.A(new_n565), .B1(new_n592), .B2(new_n556), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n557), .A2(new_n562), .ZN(new_n697));
  OAI21_X1  g511(.A(KEYINPUT98), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  INV_X1    g512(.A(new_n697), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT98), .ZN(new_n700));
  OAI211_X1 g514(.A(new_n699), .B(new_n700), .C1(new_n576), .C2(new_n565), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n698), .A2(new_n297), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(G472), .ZN(new_n703));
  NAND4_X1  g517(.A1(new_n602), .A2(new_n703), .A3(new_n603), .A4(new_n607), .ZN(new_n704));
  INV_X1    g518(.A(KEYINPUT99), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  AOI22_X1  g520(.A1(new_n702), .A2(G472), .B1(new_n601), .B2(KEYINPUT32), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n707), .A2(KEYINPUT99), .A3(new_n602), .A4(new_n607), .ZN(new_n708));
  NAND2_X1  g522(.A1(new_n706), .A2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n362), .A2(new_n366), .ZN(new_n710));
  XNOR2_X1  g524(.A(new_n710), .B(KEYINPUT38), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n672), .A2(new_n308), .A3(new_n497), .ZN(new_n712));
  AND4_X1   g526(.A1(new_n695), .A2(new_n709), .A3(new_n711), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n685), .B(KEYINPUT39), .ZN(new_n714));
  OR3_X1    g528(.A1(new_n303), .A2(new_n306), .A3(new_n714), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n715), .A2(KEYINPUT40), .ZN(new_n717));
  NAND3_X1  g531(.A1(new_n713), .A2(new_n716), .A3(new_n717), .ZN(new_n718));
  XNOR2_X1  g532(.A(new_n718), .B(G143), .ZN(G45));
  NAND4_X1  g533(.A1(new_n695), .A2(new_n644), .A3(new_n649), .A4(new_n686), .ZN(new_n720));
  NOR3_X1   g534(.A1(new_n303), .A2(new_n720), .A3(new_n306), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n683), .A2(new_n721), .ZN(new_n722));
  XNOR2_X1  g536(.A(new_n722), .B(G146), .ZN(G48));
  NAND2_X1  g537(.A1(new_n295), .A2(new_n188), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(G469), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n615), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n726), .A2(new_n306), .ZN(new_n727));
  NAND3_X1  g541(.A1(new_n609), .A2(new_n651), .A3(new_n727), .ZN(new_n728));
  XNOR2_X1  g542(.A(KEYINPUT41), .B(G113), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(KEYINPUT100), .ZN(new_n730));
  XNOR2_X1  g544(.A(new_n728), .B(new_n730), .ZN(G15));
  NAND3_X1  g545(.A1(new_n609), .A2(new_n662), .A3(new_n727), .ZN(new_n732));
  XNOR2_X1  g546(.A(new_n732), .B(G116), .ZN(G18));
  NOR2_X1   g547(.A1(new_n498), .A2(new_n375), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n683), .A2(new_n727), .A3(new_n734), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G119), .ZN(G21));
  NAND2_X1  g550(.A1(new_n599), .A2(KEYINPUT101), .ZN(new_n737));
  INV_X1    g551(.A(KEYINPUT101), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n558), .A2(new_n738), .ZN(new_n739));
  NAND3_X1  g553(.A1(new_n737), .A2(new_n739), .A3(new_n565), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n586), .B1(new_n740), .B2(new_n595), .ZN(new_n741));
  INV_X1    g555(.A(KEYINPUT102), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n742), .B1(new_n612), .B2(new_n585), .ZN(new_n743));
  OAI211_X1 g557(.A(KEYINPUT102), .B(G472), .C1(new_n606), .C2(new_n535), .ZN(new_n744));
  AOI21_X1  g558(.A(new_n741), .B1(new_n743), .B2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n539), .A2(new_n542), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  INV_X1    g561(.A(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT103), .ZN(new_n749));
  NAND4_X1  g563(.A1(new_n695), .A2(new_n749), .A3(new_n367), .A4(new_n496), .ZN(new_n750));
  AND4_X1   g564(.A1(new_n297), .A2(new_n340), .A3(new_n309), .A4(new_n360), .ZN(new_n751));
  AOI21_X1  g565(.A(new_n309), .B1(new_n365), .B2(new_n340), .ZN(new_n752));
  OAI211_X1 g566(.A(new_n307), .B(new_n496), .C1(new_n751), .C2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(KEYINPUT103), .B1(new_n753), .B2(new_n462), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n750), .A2(new_n754), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n748), .A2(new_n727), .A3(new_n376), .A4(new_n755), .ZN(new_n756));
  XNOR2_X1  g570(.A(new_n756), .B(G122), .ZN(G24));
  NOR3_X1   g571(.A1(new_n462), .A2(new_n650), .A3(new_n685), .ZN(new_n758));
  AND3_X1   g572(.A1(new_n745), .A2(new_n672), .A3(new_n758), .ZN(new_n759));
  AND4_X1   g573(.A1(new_n305), .A2(new_n615), .A3(new_n367), .A4(new_n725), .ZN(new_n760));
  NAND2_X1  g574(.A1(new_n759), .A2(new_n760), .ZN(new_n761));
  XNOR2_X1  g575(.A(KEYINPUT104), .B(G125), .ZN(new_n762));
  XNOR2_X1  g576(.A(new_n761), .B(new_n762), .ZN(G27));
  XNOR2_X1  g577(.A(new_n601), .B(new_n605), .ZN(new_n764));
  AOI21_X1  g578(.A(new_n543), .B1(new_n764), .B2(new_n584), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n758), .A2(KEYINPUT42), .ZN(new_n766));
  NAND2_X1  g580(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(G469), .A2(G902), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT105), .Z(new_n769));
  NOR2_X1   g583(.A1(new_n300), .A2(new_n301), .ZN(new_n770));
  AOI21_X1  g584(.A(new_n769), .B1(new_n770), .B2(G469), .ZN(new_n771));
  AOI21_X1  g585(.A(new_n306), .B1(new_n615), .B2(new_n771), .ZN(new_n772));
  NAND3_X1  g586(.A1(new_n362), .A2(new_n307), .A3(new_n366), .ZN(new_n773));
  INV_X1    g587(.A(new_n773), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  OAI21_X1  g589(.A(KEYINPUT107), .B1(new_n767), .B2(new_n775), .ZN(new_n776));
  INV_X1    g590(.A(new_n775), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT107), .ZN(new_n778));
  NAND4_X1  g592(.A1(new_n777), .A2(new_n778), .A3(new_n765), .A4(new_n766), .ZN(new_n779));
  INV_X1    g593(.A(new_n609), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n780), .A2(new_n775), .A3(new_n720), .ZN(new_n781));
  XOR2_X1   g595(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n782));
  OAI211_X1 g596(.A(new_n776), .B(new_n779), .C1(new_n781), .C2(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(G131), .ZN(G33));
  INV_X1    g598(.A(new_n687), .ZN(new_n785));
  NAND3_X1  g599(.A1(new_n777), .A2(new_n609), .A3(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(KEYINPUT108), .ZN(new_n787));
  XNOR2_X1  g601(.A(new_n787), .B(G134), .ZN(G36));
  NAND3_X1  g602(.A1(new_n462), .A2(new_n644), .A3(new_n649), .ZN(new_n789));
  XNOR2_X1  g603(.A(new_n789), .B(KEYINPUT43), .ZN(new_n790));
  OR2_X1    g604(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(KEYINPUT110), .ZN(new_n792));
  AND4_X1   g606(.A1(new_n613), .A2(new_n791), .A3(new_n672), .A4(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n773), .B1(new_n793), .B2(KEYINPUT44), .ZN(new_n794));
  INV_X1    g608(.A(new_n769), .ZN(new_n795));
  OAI21_X1  g609(.A(G469), .B1(new_n770), .B2(KEYINPUT45), .ZN(new_n796));
  INV_X1    g610(.A(KEYINPUT109), .ZN(new_n797));
  AND2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n770), .A2(KEYINPUT45), .ZN(new_n799));
  OAI21_X1  g613(.A(new_n799), .B1(new_n796), .B2(new_n797), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n795), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  INV_X1    g615(.A(KEYINPUT46), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n801), .A2(new_n802), .ZN(new_n803));
  OAI211_X1 g617(.A(KEYINPUT46), .B(new_n795), .C1(new_n798), .C2(new_n800), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n803), .A2(new_n615), .A3(new_n804), .ZN(new_n805));
  NAND2_X1  g619(.A1(new_n805), .A2(new_n305), .ZN(new_n806));
  NOR2_X1   g620(.A1(new_n806), .A2(new_n714), .ZN(new_n807));
  OAI211_X1 g621(.A(new_n794), .B(new_n807), .C1(KEYINPUT44), .C2(new_n793), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(G137), .ZN(G39));
  NAND2_X1  g623(.A1(new_n584), .A2(new_n608), .ZN(new_n810));
  NOR4_X1   g624(.A1(new_n810), .A2(new_n746), .A3(new_n720), .A4(new_n773), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n805), .A2(KEYINPUT47), .A3(new_n305), .ZN(new_n812));
  INV_X1    g626(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g627(.A(KEYINPUT47), .B1(new_n805), .B2(new_n305), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n811), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  XNOR2_X1  g629(.A(new_n815), .B(G140), .ZN(G42));
  XOR2_X1   g630(.A(new_n726), .B(KEYINPUT49), .Z(new_n817));
  NAND3_X1  g631(.A1(new_n746), .A2(new_n305), .A3(new_n307), .ZN(new_n818));
  NOR3_X1   g632(.A1(new_n818), .A2(new_n711), .A3(new_n789), .ZN(new_n819));
  INV_X1    g633(.A(new_n709), .ZN(new_n820));
  NAND3_X1  g634(.A1(new_n817), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  INV_X1    g635(.A(new_n727), .ZN(new_n822));
  NOR2_X1   g636(.A1(new_n822), .A2(new_n773), .ZN(new_n823));
  AND4_X1   g637(.A1(new_n746), .A2(new_n823), .A3(new_n372), .A4(new_n820), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n462), .A2(new_n650), .ZN(new_n825));
  NAND2_X1  g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  OR3_X1    g640(.A1(new_n790), .A2(KEYINPUT116), .A3(new_n371), .ZN(new_n827));
  OAI21_X1  g641(.A(KEYINPUT116), .B1(new_n790), .B2(new_n371), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n747), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n829), .A2(new_n760), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n826), .A2(new_n368), .A3(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n827), .A2(new_n828), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n832), .A2(new_n765), .A3(new_n823), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n833), .A2(KEYINPUT48), .ZN(new_n834));
  NAND2_X1  g648(.A1(new_n833), .A2(KEYINPUT48), .ZN(new_n835));
  AOI21_X1  g649(.A(new_n831), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT118), .ZN(new_n837));
  NOR2_X1   g651(.A1(new_n837), .A2(KEYINPUT50), .ZN(new_n838));
  INV_X1    g652(.A(new_n838), .ZN(new_n839));
  NOR3_X1   g653(.A1(new_n822), .A2(new_n307), .A3(new_n711), .ZN(new_n840));
  AND3_X1   g654(.A1(new_n829), .A2(new_n839), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g655(.A(new_n839), .B1(new_n829), .B2(new_n840), .ZN(new_n842));
  OR2_X1    g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n832), .A2(new_n823), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n745), .A2(new_n672), .ZN(new_n845));
  AND2_X1   g659(.A1(new_n462), .A2(new_n650), .ZN(new_n846));
  AOI22_X1  g660(.A1(new_n844), .A2(new_n845), .B1(new_n824), .B2(new_n846), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n847), .ZN(new_n848));
  NAND2_X1  g662(.A1(new_n829), .A2(new_n774), .ZN(new_n849));
  NOR2_X1   g663(.A1(new_n813), .A2(new_n814), .ZN(new_n850));
  INV_X1    g664(.A(new_n726), .ZN(new_n851));
  NAND2_X1  g665(.A1(new_n851), .A2(new_n306), .ZN(new_n852));
  AOI21_X1  g666(.A(new_n849), .B1(new_n850), .B2(new_n852), .ZN(new_n853));
  OAI21_X1  g667(.A(new_n836), .B1(new_n848), .B2(new_n853), .ZN(new_n854));
  INV_X1    g668(.A(KEYINPUT117), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n855), .B1(new_n813), .B2(new_n814), .ZN(new_n856));
  INV_X1    g670(.A(new_n814), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n857), .A2(KEYINPUT117), .A3(new_n812), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n856), .A2(new_n858), .A3(new_n852), .ZN(new_n859));
  OAI211_X1 g673(.A(new_n843), .B(new_n847), .C1(new_n859), .C2(new_n849), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT51), .ZN(new_n861));
  AOI21_X1  g675(.A(new_n854), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g676(.A(KEYINPUT53), .ZN(new_n863));
  NAND4_X1  g677(.A1(new_n678), .A2(new_n728), .A3(new_n610), .A4(new_n652), .ZN(new_n864));
  XNOR2_X1  g678(.A(new_n496), .B(KEYINPUT111), .ZN(new_n865));
  NOR3_X1   g679(.A1(new_n377), .A2(new_n695), .A3(new_n865), .ZN(new_n866));
  NAND3_X1  g680(.A1(new_n614), .A2(new_n617), .A3(new_n866), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n732), .A2(new_n756), .A3(new_n735), .A4(new_n867), .ZN(new_n868));
  NAND2_X1  g682(.A1(new_n865), .A2(new_n686), .ZN(new_n869));
  NOR3_X1   g683(.A1(new_n673), .A2(new_n661), .A3(new_n869), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n870), .A2(new_n810), .A3(new_n617), .ZN(new_n871));
  NAND2_X1  g685(.A1(new_n759), .A2(new_n772), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n773), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  NOR3_X1   g687(.A1(new_n864), .A2(new_n868), .A3(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n668), .A2(new_n671), .A3(new_n686), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n875), .A2(KEYINPUT112), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT112), .ZN(new_n877));
  NAND4_X1  g691(.A1(new_n668), .A2(new_n877), .A3(new_n671), .A4(new_n686), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n876), .A2(new_n878), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n709), .A2(new_n755), .A3(new_n772), .A4(new_n879), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n880), .A2(new_n689), .A3(new_n722), .A4(new_n761), .ZN(new_n881));
  NAND2_X1  g695(.A1(new_n881), .A2(KEYINPUT52), .ZN(new_n882));
  NAND4_X1  g696(.A1(new_n874), .A2(new_n783), .A3(new_n787), .A4(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT113), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n881), .A2(new_n884), .ZN(new_n885));
  AOI22_X1  g699(.A1(new_n706), .A2(new_n708), .B1(new_n876), .B2(new_n878), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n772), .A2(new_n755), .ZN(new_n887));
  AOI22_X1  g701(.A1(new_n886), .A2(new_n887), .B1(new_n683), .B2(new_n721), .ZN(new_n888));
  AOI22_X1  g702(.A1(new_n683), .A2(new_n688), .B1(new_n759), .B2(new_n760), .ZN(new_n889));
  NAND3_X1  g703(.A1(new_n888), .A2(KEYINPUT113), .A3(new_n889), .ZN(new_n890));
  AOI21_X1  g704(.A(KEYINPUT52), .B1(new_n885), .B2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n863), .B1(new_n883), .B2(new_n891), .ZN(new_n892));
  INV_X1    g706(.A(KEYINPUT114), .ZN(new_n893));
  AND3_X1   g707(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n890), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n893), .B1(new_n894), .B2(new_n891), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n864), .A2(new_n868), .ZN(new_n896));
  INV_X1    g710(.A(new_n873), .ZN(new_n897));
  NAND4_X1  g711(.A1(new_n787), .A2(new_n896), .A3(new_n783), .A4(new_n897), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT52), .ZN(new_n900));
  AND4_X1   g714(.A1(KEYINPUT113), .A2(new_n889), .A3(new_n722), .A4(new_n880), .ZN(new_n901));
  AOI21_X1  g715(.A(KEYINPUT113), .B1(new_n888), .B2(new_n889), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n900), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g717(.A1(new_n885), .A2(KEYINPUT52), .A3(new_n890), .ZN(new_n904));
  NAND3_X1  g718(.A1(new_n903), .A2(KEYINPUT114), .A3(new_n904), .ZN(new_n905));
  NAND3_X1  g719(.A1(new_n895), .A2(new_n899), .A3(new_n905), .ZN(new_n906));
  OAI21_X1  g720(.A(new_n892), .B1(new_n906), .B2(new_n863), .ZN(new_n907));
  NAND2_X1  g721(.A1(new_n907), .A2(KEYINPUT54), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n883), .A2(new_n863), .A3(new_n891), .ZN(new_n909));
  AOI21_X1  g723(.A(new_n909), .B1(new_n906), .B2(new_n863), .ZN(new_n910));
  XNOR2_X1  g724(.A(KEYINPUT115), .B(KEYINPUT54), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  NAND4_X1  g726(.A1(new_n862), .A2(KEYINPUT119), .A3(new_n908), .A4(new_n912), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n913), .B1(G952), .B2(G953), .ZN(new_n914));
  AND2_X1   g728(.A1(new_n908), .A2(new_n912), .ZN(new_n915));
  AOI21_X1  g729(.A(KEYINPUT119), .B1(new_n915), .B2(new_n862), .ZN(new_n916));
  OAI21_X1  g730(.A(new_n821), .B1(new_n914), .B2(new_n916), .ZN(G75));
  NAND2_X1  g731(.A1(new_n906), .A2(new_n863), .ZN(new_n918));
  INV_X1    g732(.A(new_n909), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND3_X1  g734(.A1(new_n920), .A2(new_n535), .A3(new_n310), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n329), .A2(new_n331), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(new_n339), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT55), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n925), .A2(KEYINPUT56), .ZN(new_n926));
  AND3_X1   g740(.A1(new_n921), .A2(new_n924), .A3(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n924), .B1(new_n921), .B2(new_n926), .ZN(new_n928));
  NOR2_X1   g742(.A1(new_n337), .A2(G952), .ZN(new_n929));
  NOR3_X1   g743(.A1(new_n927), .A2(new_n928), .A3(new_n929), .ZN(G51));
  AND2_X1   g744(.A1(new_n910), .A2(new_n911), .ZN(new_n931));
  NOR2_X1   g745(.A1(new_n910), .A2(new_n911), .ZN(new_n932));
  NOR2_X1   g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n769), .B(KEYINPUT57), .Z(new_n934));
  OAI21_X1  g748(.A(new_n295), .B1(new_n933), .B2(new_n934), .ZN(new_n935));
  OR4_X1    g749(.A1(new_n188), .A2(new_n910), .A3(new_n798), .A4(new_n800), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n929), .B1(new_n935), .B2(new_n936), .ZN(G54));
  INV_X1    g751(.A(KEYINPUT58), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n378), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n903), .A2(new_n904), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n898), .B1(new_n940), .B2(new_n893), .ZN(new_n941));
  AOI21_X1  g755(.A(KEYINPUT53), .B1(new_n941), .B2(new_n905), .ZN(new_n942));
  OAI211_X1 g756(.A(new_n535), .B(new_n939), .C1(new_n942), .C2(new_n909), .ZN(new_n943));
  NAND2_X1  g757(.A1(new_n943), .A2(new_n451), .ZN(new_n944));
  NOR3_X1   g758(.A1(new_n451), .A2(new_n938), .A3(new_n378), .ZN(new_n945));
  OAI211_X1 g759(.A(new_n535), .B(new_n945), .C1(new_n942), .C2(new_n909), .ZN(new_n946));
  INV_X1    g760(.A(KEYINPUT121), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g762(.A(new_n929), .ZN(new_n949));
  NAND4_X1  g763(.A1(new_n920), .A2(KEYINPUT121), .A3(new_n535), .A4(new_n945), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n944), .A2(new_n948), .A3(new_n949), .A4(new_n950), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT122), .ZN(new_n952));
  NAND2_X1  g766(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  AOI21_X1  g767(.A(new_n929), .B1(new_n943), .B2(new_n451), .ZN(new_n954));
  NAND4_X1  g768(.A1(new_n954), .A2(KEYINPUT122), .A3(new_n948), .A4(new_n950), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(new_n955), .ZN(G60));
  NAND2_X1  g770(.A1(G478), .A2(G902), .ZN(new_n957));
  XOR2_X1   g771(.A(new_n957), .B(KEYINPUT59), .Z(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n639), .A2(new_n959), .ZN(new_n960));
  OAI21_X1  g774(.A(new_n949), .B1(new_n933), .B2(new_n960), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n908), .A2(new_n912), .ZN(new_n962));
  AOI21_X1  g776(.A(new_n639), .B1(new_n962), .B2(new_n959), .ZN(new_n963));
  NOR2_X1   g777(.A1(new_n961), .A2(new_n963), .ZN(G63));
  NAND2_X1  g778(.A1(G217), .A2(G902), .ZN(new_n965));
  XOR2_X1   g779(.A(new_n965), .B(KEYINPUT123), .Z(new_n966));
  XOR2_X1   g780(.A(new_n966), .B(KEYINPUT60), .Z(new_n967));
  INV_X1    g781(.A(new_n967), .ZN(new_n968));
  AOI21_X1  g782(.A(new_n968), .B1(new_n918), .B2(new_n919), .ZN(new_n969));
  XNOR2_X1  g783(.A(new_n670), .B(KEYINPUT124), .ZN(new_n970));
  AOI21_X1  g784(.A(new_n929), .B1(new_n969), .B2(new_n970), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n534), .B1(new_n910), .B2(new_n968), .ZN(new_n972));
  INV_X1    g786(.A(KEYINPUT125), .ZN(new_n973));
  INV_X1    g787(.A(KEYINPUT61), .ZN(new_n974));
  OAI211_X1 g788(.A(new_n971), .B(new_n972), .C1(new_n973), .C2(new_n974), .ZN(new_n975));
  OAI211_X1 g789(.A(new_n967), .B(new_n970), .C1(new_n942), .C2(new_n909), .ZN(new_n976));
  NAND3_X1  g790(.A1(new_n972), .A2(new_n949), .A3(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n973), .A3(new_n949), .ZN(new_n978));
  NAND3_X1  g792(.A1(new_n977), .A2(KEYINPUT61), .A3(new_n978), .ZN(new_n979));
  AND2_X1   g793(.A1(new_n975), .A2(new_n979), .ZN(G66));
  INV_X1    g794(.A(G224), .ZN(new_n981));
  OAI21_X1  g795(.A(G953), .B1(new_n374), .B2(new_n981), .ZN(new_n982));
  OAI21_X1  g796(.A(new_n982), .B1(new_n896), .B2(G953), .ZN(new_n983));
  OAI21_X1  g797(.A(new_n922), .B1(G898), .B2(new_n337), .ZN(new_n984));
  XNOR2_X1  g798(.A(new_n984), .B(KEYINPUT126), .ZN(new_n985));
  XNOR2_X1  g799(.A(new_n983), .B(new_n985), .ZN(G69));
  AND2_X1   g800(.A1(new_n808), .A2(new_n815), .ZN(new_n987));
  NAND2_X1  g801(.A1(new_n889), .A2(new_n722), .ZN(new_n988));
  INV_X1    g802(.A(new_n988), .ZN(new_n989));
  NAND2_X1  g803(.A1(new_n989), .A2(new_n718), .ZN(new_n990));
  XOR2_X1   g804(.A(new_n990), .B(KEYINPUT62), .Z(new_n991));
  NOR2_X1   g805(.A1(new_n695), .A2(new_n865), .ZN(new_n992));
  OAI21_X1  g806(.A(new_n774), .B1(new_n992), .B2(new_n825), .ZN(new_n993));
  OR3_X1    g807(.A1(new_n780), .A2(new_n715), .A3(new_n993), .ZN(new_n994));
  NAND3_X1  g808(.A1(new_n987), .A2(new_n991), .A3(new_n994), .ZN(new_n995));
  NAND2_X1  g809(.A1(new_n995), .A2(new_n337), .ZN(new_n996));
  NAND2_X1  g810(.A1(new_n574), .A2(new_n566), .ZN(new_n997));
  NAND2_X1  g811(.A1(new_n434), .A2(new_n436), .ZN(new_n998));
  XNOR2_X1  g812(.A(new_n997), .B(new_n998), .ZN(new_n999));
  INV_X1    g813(.A(new_n999), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n996), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g815(.A1(new_n337), .A2(G900), .ZN(new_n1002));
  NAND3_X1  g816(.A1(new_n807), .A2(new_n755), .A3(new_n765), .ZN(new_n1003));
  AND3_X1   g817(.A1(new_n787), .A2(new_n783), .A3(new_n989), .ZN(new_n1004));
  NAND3_X1  g818(.A1(new_n987), .A2(new_n1003), .A3(new_n1004), .ZN(new_n1005));
  AOI21_X1  g819(.A(new_n1002), .B1(new_n1005), .B2(new_n337), .ZN(new_n1006));
  OAI21_X1  g820(.A(new_n1001), .B1(new_n1006), .B2(new_n1000), .ZN(new_n1007));
  OAI21_X1  g821(.A(G953), .B1(new_n257), .B2(new_n684), .ZN(new_n1008));
  XNOR2_X1  g822(.A(new_n1008), .B(KEYINPUT127), .ZN(new_n1009));
  XNOR2_X1  g823(.A(new_n1007), .B(new_n1009), .ZN(G72));
  NAND2_X1  g824(.A1(G472), .A2(G902), .ZN(new_n1011));
  XOR2_X1   g825(.A(new_n1011), .B(KEYINPUT63), .Z(new_n1012));
  INV_X1    g826(.A(new_n896), .ZN(new_n1013));
  OAI21_X1  g827(.A(new_n1012), .B1(new_n995), .B2(new_n1013), .ZN(new_n1014));
  AOI21_X1  g828(.A(new_n929), .B1(new_n1014), .B2(new_n696), .ZN(new_n1015));
  OAI211_X1 g829(.A(new_n577), .B(new_n573), .C1(new_n572), .C2(new_n588), .ZN(new_n1016));
  NAND3_X1  g830(.A1(new_n907), .A2(new_n1012), .A3(new_n1016), .ZN(new_n1017));
  OAI21_X1  g831(.A(new_n1012), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1018));
  NAND3_X1  g832(.A1(new_n1018), .A2(new_n565), .A3(new_n576), .ZN(new_n1019));
  AND3_X1   g833(.A1(new_n1015), .A2(new_n1017), .A3(new_n1019), .ZN(G57));
endmodule


