//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 0 1 1 1 1 1 1 0 1 1 0 0 0 1 1 0 0 1 1 0 0 0 1 0 1 0 1 0 1 0 0 0 0 1 1 1 1 1 1 0 1 0 0 0 0 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:06 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n453, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n524, new_n525,
    new_n526, new_n527, new_n528, new_n529, new_n530, new_n531, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n555, new_n556, new_n557, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n568, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n604, new_n607, new_n608, new_n610, new_n611, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n826, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1184,
    new_n1185, new_n1186;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT64), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XOR2_X1   g011(.A(KEYINPUT65), .B(G96), .Z(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G221), .A2(G220), .A3(G218), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT66), .ZN(new_n451));
  XNOR2_X1  g026(.A(new_n451), .B(KEYINPUT2), .ZN(new_n452));
  NAND4_X1  g027(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n453));
  NOR2_X1   g028(.A1(new_n452), .A2(new_n453), .ZN(G325));
  INV_X1    g029(.A(G325), .ZN(G261));
  NAND2_X1  g030(.A1(new_n452), .A2(G2106), .ZN(new_n456));
  NAND2_X1  g031(.A1(new_n453), .A2(G567), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n456), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  XNOR2_X1  g034(.A(KEYINPUT3), .B(G2104), .ZN(new_n460));
  INV_X1    g035(.A(G2105), .ZN(new_n461));
  NAND3_X1  g036(.A1(new_n460), .A2(G137), .A3(new_n461), .ZN(new_n462));
  INV_X1    g037(.A(G2104), .ZN(new_n463));
  NOR2_X1   g038(.A1(new_n463), .A2(G2105), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(G101), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n462), .A2(new_n465), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n463), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT67), .ZN(new_n471));
  NAND2_X1  g046(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g047(.A1(G113), .A2(G2104), .ZN(new_n473));
  NAND4_X1  g048(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT67), .A4(G125), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n472), .A2(new_n473), .A3(new_n474), .ZN(new_n475));
  AOI21_X1  g050(.A(new_n466), .B1(new_n475), .B2(G2105), .ZN(G160));
  NAND2_X1  g051(.A1(new_n460), .A2(G2105), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(new_n478));
  NAND2_X1  g053(.A1(new_n478), .A2(G124), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n467), .A2(new_n469), .ZN(new_n480));
  NOR2_X1   g055(.A1(new_n480), .A2(G2105), .ZN(new_n481));
  NAND2_X1  g056(.A1(new_n481), .A2(G136), .ZN(new_n482));
  OR2_X1    g057(.A1(G100), .A2(G2105), .ZN(new_n483));
  OAI211_X1 g058(.A(new_n483), .B(G2104), .C1(G112), .C2(new_n461), .ZN(new_n484));
  NAND3_X1  g059(.A1(new_n479), .A2(new_n482), .A3(new_n484), .ZN(new_n485));
  INV_X1    g060(.A(new_n485), .ZN(G162));
  NAND3_X1  g061(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n487));
  NAND2_X1  g062(.A1(G114), .A2(G2104), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n487), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g064(.A1(new_n489), .A2(G2105), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n467), .A2(new_n469), .A3(G138), .A4(new_n461), .ZN(new_n491));
  INV_X1    g066(.A(KEYINPUT4), .ZN(new_n492));
  NAND3_X1  g067(.A1(new_n491), .A2(KEYINPUT68), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n464), .A2(G102), .ZN(new_n494));
  XNOR2_X1  g069(.A(KEYINPUT68), .B(KEYINPUT4), .ZN(new_n495));
  NAND4_X1  g070(.A1(new_n460), .A2(new_n495), .A3(G138), .A4(new_n461), .ZN(new_n496));
  NAND4_X1  g071(.A1(new_n490), .A2(new_n493), .A3(new_n494), .A4(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT70), .ZN(new_n499));
  XNOR2_X1  g074(.A(KEYINPUT69), .B(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT6), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n499), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  INV_X1    g077(.A(KEYINPUT69), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n503), .A2(G651), .ZN(new_n504));
  INV_X1    g079(.A(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n505), .A2(KEYINPUT69), .ZN(new_n506));
  OAI211_X1 g081(.A(KEYINPUT70), .B(KEYINPUT6), .C1(new_n504), .C2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n501), .A2(G651), .ZN(new_n508));
  NAND4_X1  g083(.A1(new_n502), .A2(G543), .A3(new_n507), .A4(new_n508), .ZN(new_n509));
  INV_X1    g084(.A(G50), .ZN(new_n510));
  INV_X1    g085(.A(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  AOI22_X1  g091(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n517));
  INV_X1    g092(.A(new_n500), .ZN(new_n518));
  OAI22_X1  g093(.A1(new_n509), .A2(new_n510), .B1(new_n517), .B2(new_n518), .ZN(new_n519));
  NAND4_X1  g094(.A1(new_n502), .A2(new_n516), .A3(new_n507), .A4(new_n508), .ZN(new_n520));
  XOR2_X1   g095(.A(KEYINPUT71), .B(G88), .Z(new_n521));
  NOR2_X1   g096(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NOR2_X1   g097(.A1(new_n519), .A2(new_n522), .ZN(G166));
  AND3_X1   g098(.A1(new_n502), .A2(new_n508), .A3(new_n507), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G89), .ZN(new_n525));
  INV_X1    g100(.A(G63), .ZN(new_n526));
  OAI21_X1  g101(.A(new_n525), .B1(new_n526), .B2(new_n505), .ZN(new_n527));
  INV_X1    g102(.A(new_n509), .ZN(new_n528));
  AOI22_X1  g103(.A1(new_n527), .A2(new_n516), .B1(G51), .B2(new_n528), .ZN(new_n529));
  NAND3_X1  g104(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n530));
  XNOR2_X1  g105(.A(new_n530), .B(KEYINPUT7), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n529), .A2(new_n531), .ZN(G286));
  INV_X1    g107(.A(G286), .ZN(G168));
  NAND2_X1  g108(.A1(G77), .A2(G543), .ZN(new_n534));
  INV_X1    g109(.A(G64), .ZN(new_n535));
  OAI21_X1  g110(.A(new_n534), .B1(new_n515), .B2(new_n535), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n536), .A2(new_n500), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT72), .ZN(new_n538));
  XNOR2_X1  g113(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g114(.A(G52), .ZN(new_n540));
  INV_X1    g115(.A(G90), .ZN(new_n541));
  OAI22_X1  g116(.A1(new_n540), .A2(new_n509), .B1(new_n520), .B2(new_n541), .ZN(new_n542));
  NOR2_X1   g117(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  INV_X1    g118(.A(KEYINPUT73), .ZN(new_n544));
  XNOR2_X1  g119(.A(new_n543), .B(new_n544), .ZN(G171));
  INV_X1    g120(.A(G81), .ZN(new_n546));
  AOI22_X1  g121(.A1(new_n516), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n547));
  OAI22_X1  g122(.A1(new_n520), .A2(new_n546), .B1(new_n547), .B2(new_n518), .ZN(new_n548));
  XOR2_X1   g123(.A(KEYINPUT74), .B(G43), .Z(new_n549));
  NOR2_X1   g124(.A1(new_n509), .A2(new_n549), .ZN(new_n550));
  NOR2_X1   g125(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n551), .A2(G860), .ZN(G153));
  AND3_X1   g127(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n553), .A2(G36), .ZN(G176));
  NAND2_X1  g129(.A1(G1), .A2(G3), .ZN(new_n555));
  XNOR2_X1  g130(.A(new_n555), .B(KEYINPUT8), .ZN(new_n556));
  NAND2_X1  g131(.A1(new_n553), .A2(new_n556), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n557), .B(KEYINPUT75), .ZN(G188));
  NAND2_X1  g133(.A1(new_n516), .A2(G65), .ZN(new_n559));
  NAND2_X1  g134(.A1(G78), .A2(G543), .ZN(new_n560));
  AOI21_X1  g135(.A(new_n505), .B1(new_n559), .B2(new_n560), .ZN(new_n561));
  INV_X1    g136(.A(G91), .ZN(new_n562));
  NOR2_X1   g137(.A1(new_n520), .A2(new_n562), .ZN(new_n563));
  INV_X1    g138(.A(KEYINPUT9), .ZN(new_n564));
  NAND4_X1  g139(.A1(new_n524), .A2(new_n564), .A3(G53), .A4(G543), .ZN(new_n565));
  INV_X1    g140(.A(G53), .ZN(new_n566));
  OAI21_X1  g141(.A(KEYINPUT9), .B1(new_n509), .B2(new_n566), .ZN(new_n567));
  AOI211_X1 g142(.A(new_n561), .B(new_n563), .C1(new_n565), .C2(new_n567), .ZN(new_n568));
  INV_X1    g143(.A(new_n568), .ZN(G299));
  XNOR2_X1  g144(.A(new_n543), .B(KEYINPUT73), .ZN(G301));
  INV_X1    g145(.A(G166), .ZN(G303));
  OAI21_X1  g146(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n572));
  INV_X1    g147(.A(G87), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n520), .B2(new_n573), .ZN(new_n574));
  INV_X1    g149(.A(G49), .ZN(new_n575));
  NOR2_X1   g150(.A1(new_n509), .A2(new_n575), .ZN(new_n576));
  NOR2_X1   g151(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  INV_X1    g152(.A(new_n577), .ZN(G288));
  INV_X1    g153(.A(G48), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n516), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n580));
  OAI22_X1  g155(.A1(new_n509), .A2(new_n579), .B1(new_n580), .B2(new_n518), .ZN(new_n581));
  INV_X1    g156(.A(G86), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n520), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g158(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  INV_X1    g159(.A(new_n584), .ZN(G305));
  INV_X1    g160(.A(G47), .ZN(new_n586));
  AOI22_X1  g161(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n587));
  OAI22_X1  g162(.A1(new_n509), .A2(new_n586), .B1(new_n587), .B2(new_n518), .ZN(new_n588));
  INV_X1    g163(.A(G85), .ZN(new_n589));
  NOR2_X1   g164(.A1(new_n520), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g165(.A1(new_n588), .A2(new_n590), .ZN(new_n591));
  INV_X1    g166(.A(new_n591), .ZN(G290));
  INV_X1    g167(.A(G92), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n520), .A2(new_n593), .ZN(new_n594));
  XNOR2_X1  g169(.A(new_n594), .B(KEYINPUT10), .ZN(new_n595));
  NAND2_X1  g170(.A1(new_n528), .A2(G54), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n516), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n597));
  OR2_X1    g172(.A1(new_n597), .A2(new_n505), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G284));
  OAI21_X1  g177(.A(new_n601), .B1(G171), .B2(new_n600), .ZN(G321));
  NAND2_X1  g178(.A1(G299), .A2(new_n600), .ZN(new_n604));
  OAI21_X1  g179(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G297));
  OAI21_X1  g180(.A(new_n604), .B1(G168), .B2(new_n600), .ZN(G280));
  AND3_X1   g181(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n607));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n607), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND2_X1  g184(.A1(new_n607), .A2(new_n608), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(G868), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n611), .B1(G868), .B2(new_n551), .ZN(G323));
  XNOR2_X1  g187(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g188(.A1(new_n461), .A2(G111), .ZN(new_n614));
  AOI21_X1  g189(.A(new_n463), .B1(new_n614), .B2(KEYINPUT77), .ZN(new_n615));
  OAI221_X1 g190(.A(new_n615), .B1(KEYINPUT77), .B2(new_n614), .C1(G99), .C2(G2105), .ZN(new_n616));
  AOI22_X1  g191(.A1(new_n478), .A2(G123), .B1(new_n481), .B2(G135), .ZN(new_n617));
  NAND2_X1  g192(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g193(.A(G2096), .ZN(new_n619));
  XNOR2_X1  g194(.A(new_n618), .B(new_n619), .ZN(new_n620));
  NAND2_X1  g195(.A1(new_n460), .A2(new_n464), .ZN(new_n621));
  XOR2_X1   g196(.A(new_n621), .B(KEYINPUT12), .Z(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT76), .B(KEYINPUT13), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(G2100), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n622), .B(new_n624), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n620), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(KEYINPUT15), .B(G2430), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(G2435), .ZN(new_n628));
  XOR2_X1   g203(.A(G2427), .B(G2438), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  NAND2_X1  g205(.A1(new_n630), .A2(KEYINPUT14), .ZN(new_n631));
  XNOR2_X1  g206(.A(G2451), .B(G2454), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT78), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT16), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n631), .B(new_n634), .ZN(new_n635));
  XOR2_X1   g210(.A(G2443), .B(G2446), .Z(new_n636));
  XNOR2_X1  g211(.A(new_n635), .B(new_n636), .ZN(new_n637));
  XOR2_X1   g212(.A(G1341), .B(G1348), .Z(new_n638));
  XNOR2_X1  g213(.A(new_n637), .B(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(G14), .ZN(G401));
  XNOR2_X1  g215(.A(G2067), .B(G2678), .ZN(new_n641));
  XNOR2_X1  g216(.A(G2072), .B(G2078), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(G2084), .B(G2090), .Z(new_n644));
  NOR2_X1   g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT79), .ZN(new_n646));
  INV_X1    g221(.A(new_n641), .ZN(new_n647));
  XOR2_X1   g222(.A(new_n642), .B(KEYINPUT17), .Z(new_n648));
  OAI21_X1  g223(.A(new_n646), .B1(new_n647), .B2(new_n648), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n648), .A2(new_n647), .A3(new_n644), .ZN(new_n650));
  NAND3_X1  g225(.A1(new_n644), .A2(new_n641), .A3(new_n642), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n651), .B(KEYINPUT18), .Z(new_n652));
  NAND3_X1  g227(.A1(new_n649), .A2(new_n650), .A3(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(new_n653), .B(KEYINPUT80), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(new_n619), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(G2100), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(new_n657), .B(KEYINPUT19), .ZN(new_n658));
  XOR2_X1   g233(.A(G1956), .B(G2474), .Z(new_n659));
  XOR2_X1   g234(.A(G1961), .B(G1966), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n659), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n658), .ZN(new_n663));
  NOR2_X1   g238(.A1(new_n659), .A2(new_n660), .ZN(new_n664));
  AOI22_X1  g239(.A1(new_n662), .A2(KEYINPUT20), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g241(.A1(new_n666), .A2(new_n658), .A3(new_n661), .ZN(new_n667));
  OAI211_X1 g242(.A(new_n665), .B(new_n667), .C1(KEYINPUT20), .C2(new_n662), .ZN(new_n668));
  XOR2_X1   g243(.A(G1991), .B(G1996), .Z(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(G1981), .B(G1986), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n670), .B(new_n671), .ZN(new_n672));
  XOR2_X1   g247(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n673));
  XNOR2_X1  g248(.A(new_n672), .B(new_n673), .ZN(G229));
  INV_X1    g249(.A(G29), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n675), .A2(G27), .ZN(new_n676));
  OAI21_X1  g251(.A(new_n676), .B1(G164), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g252(.A1(new_n677), .A2(G2078), .ZN(new_n678));
  NAND2_X1  g253(.A1(G168), .A2(G16), .ZN(new_n679));
  OAI211_X1 g254(.A(new_n679), .B(KEYINPUT90), .C1(G16), .C2(G21), .ZN(new_n680));
  INV_X1    g255(.A(G16), .ZN(new_n681));
  OR3_X1    g256(.A1(G286), .A2(KEYINPUT90), .A3(new_n681), .ZN(new_n682));
  NAND2_X1  g257(.A1(new_n680), .A2(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n683), .A2(KEYINPUT91), .ZN(new_n684));
  INV_X1    g259(.A(KEYINPUT91), .ZN(new_n685));
  NAND3_X1  g260(.A1(new_n680), .A2(new_n685), .A3(new_n682), .ZN(new_n686));
  NAND3_X1  g261(.A1(new_n684), .A2(G1966), .A3(new_n686), .ZN(new_n687));
  XNOR2_X1  g262(.A(new_n687), .B(KEYINPUT92), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n616), .A2(new_n617), .A3(G29), .ZN(new_n689));
  XNOR2_X1  g264(.A(KEYINPUT93), .B(KEYINPUT30), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G28), .ZN(new_n691));
  NOR2_X1   g266(.A1(G29), .A2(G32), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n464), .A2(G105), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n460), .A2(new_n461), .ZN(new_n694));
  INV_X1    g269(.A(G141), .ZN(new_n695));
  INV_X1    g270(.A(G129), .ZN(new_n696));
  OAI221_X1 g271(.A(new_n693), .B1(new_n694), .B2(new_n695), .C1(new_n696), .C2(new_n477), .ZN(new_n697));
  NAND3_X1  g272(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n698), .B(KEYINPUT89), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(new_n700));
  AND2_X1   g275(.A1(new_n700), .A2(KEYINPUT26), .ZN(new_n701));
  NOR2_X1   g276(.A1(new_n700), .A2(KEYINPUT26), .ZN(new_n702));
  NOR3_X1   g277(.A1(new_n697), .A2(new_n701), .A3(new_n702), .ZN(new_n703));
  AOI21_X1  g278(.A(new_n692), .B1(new_n703), .B2(G29), .ZN(new_n704));
  INV_X1    g279(.A(new_n704), .ZN(new_n705));
  XOR2_X1   g280(.A(KEYINPUT27), .B(G1996), .Z(new_n706));
  INV_X1    g281(.A(new_n706), .ZN(new_n707));
  OAI221_X1 g282(.A(new_n689), .B1(G29), .B2(new_n691), .C1(new_n705), .C2(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n675), .A2(G35), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G162), .B2(new_n675), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT95), .B(KEYINPUT29), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n711), .B(KEYINPUT96), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n710), .B(new_n712), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G2090), .ZN(new_n714));
  OR2_X1    g289(.A1(KEYINPUT24), .A2(G34), .ZN(new_n715));
  NAND2_X1  g290(.A1(KEYINPUT24), .A2(G34), .ZN(new_n716));
  NAND3_X1  g291(.A1(new_n715), .A2(new_n675), .A3(new_n716), .ZN(new_n717));
  OAI21_X1  g292(.A(new_n717), .B1(G160), .B2(new_n675), .ZN(new_n718));
  OR2_X1    g293(.A1(new_n718), .A2(G2084), .ZN(new_n719));
  NAND2_X1  g294(.A1(new_n714), .A2(new_n719), .ZN(new_n720));
  AOI211_X1 g295(.A(new_n708), .B(new_n720), .C1(new_n705), .C2(new_n707), .ZN(new_n721));
  NAND2_X1  g296(.A1(new_n681), .A2(G19), .ZN(new_n722));
  OAI21_X1  g297(.A(new_n722), .B1(new_n551), .B2(new_n681), .ZN(new_n723));
  XOR2_X1   g298(.A(new_n723), .B(G1341), .Z(new_n724));
  NAND2_X1  g299(.A1(new_n675), .A2(G26), .ZN(new_n725));
  INV_X1    g300(.A(G128), .ZN(new_n726));
  NOR2_X1   g301(.A1(new_n477), .A2(new_n726), .ZN(new_n727));
  NAND3_X1  g302(.A1(new_n481), .A2(KEYINPUT85), .A3(G140), .ZN(new_n728));
  INV_X1    g303(.A(KEYINPUT85), .ZN(new_n729));
  INV_X1    g304(.A(G140), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n694), .B2(new_n730), .ZN(new_n731));
  AOI21_X1  g306(.A(new_n727), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  OAI21_X1  g307(.A(G2104), .B1(new_n461), .B2(G116), .ZN(new_n733));
  INV_X1    g308(.A(G104), .ZN(new_n734));
  AOI21_X1  g309(.A(new_n733), .B1(new_n734), .B2(new_n461), .ZN(new_n735));
  INV_X1    g310(.A(new_n735), .ZN(new_n736));
  AND2_X1   g311(.A1(new_n732), .A2(new_n736), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n725), .B1(new_n737), .B2(new_n675), .ZN(new_n738));
  MUX2_X1   g313(.A(new_n725), .B(new_n738), .S(KEYINPUT28), .Z(new_n739));
  INV_X1    g314(.A(G2067), .ZN(new_n740));
  XNOR2_X1  g315(.A(new_n739), .B(new_n740), .ZN(new_n741));
  NAND3_X1  g316(.A1(new_n721), .A2(new_n724), .A3(new_n741), .ZN(new_n742));
  AND2_X1   g317(.A1(new_n681), .A2(G20), .ZN(new_n743));
  AOI21_X1  g318(.A(new_n743), .B1(G299), .B2(G16), .ZN(new_n744));
  MUX2_X1   g319(.A(new_n743), .B(new_n744), .S(KEYINPUT23), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT97), .B(G1956), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n745), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g322(.A1(new_n718), .A2(G2084), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n677), .A2(G2078), .ZN(new_n749));
  OAI211_X1 g324(.A(new_n748), .B(new_n749), .C1(new_n713), .C2(G2090), .ZN(new_n750));
  NAND2_X1  g325(.A1(new_n464), .A2(G103), .ZN(new_n751));
  INV_X1    g326(.A(KEYINPUT86), .ZN(new_n752));
  XNOR2_X1  g327(.A(new_n751), .B(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n753), .A2(KEYINPUT25), .ZN(new_n754));
  XNOR2_X1  g329(.A(new_n751), .B(KEYINPUT86), .ZN(new_n755));
  INV_X1    g330(.A(KEYINPUT25), .ZN(new_n756));
  NAND2_X1  g331(.A1(new_n755), .A2(new_n756), .ZN(new_n757));
  NAND3_X1  g332(.A1(new_n481), .A2(KEYINPUT87), .A3(G139), .ZN(new_n758));
  INV_X1    g333(.A(KEYINPUT87), .ZN(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  OAI21_X1  g335(.A(new_n759), .B1(new_n694), .B2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n758), .A2(new_n761), .ZN(new_n762));
  NAND3_X1  g337(.A1(new_n754), .A2(new_n757), .A3(new_n762), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT88), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  NAND4_X1  g340(.A1(new_n754), .A2(new_n757), .A3(new_n762), .A4(KEYINPUT88), .ZN(new_n766));
  NAND2_X1  g341(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n460), .A2(G127), .ZN(new_n768));
  NAND2_X1  g343(.A1(G115), .A2(G2104), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n461), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  INV_X1    g345(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g346(.A1(new_n767), .A2(new_n771), .ZN(new_n772));
  MUX2_X1   g347(.A(G33), .B(new_n772), .S(G29), .Z(new_n773));
  AOI21_X1  g348(.A(new_n750), .B1(new_n773), .B2(G2072), .ZN(new_n774));
  OAI211_X1 g349(.A(new_n747), .B(new_n774), .C1(G2072), .C2(new_n773), .ZN(new_n775));
  XOR2_X1   g350(.A(KEYINPUT31), .B(G11), .Z(new_n776));
  NAND2_X1  g351(.A1(new_n681), .A2(G4), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(new_n607), .B2(new_n681), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G1348), .ZN(new_n779));
  NOR4_X1   g354(.A1(new_n742), .A2(new_n775), .A3(new_n776), .A4(new_n779), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n684), .A2(new_n686), .ZN(new_n781));
  INV_X1    g356(.A(G1966), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  INV_X1    g358(.A(G5), .ZN(new_n784));
  AOI21_X1  g359(.A(KEYINPUT94), .B1(new_n784), .B2(new_n681), .ZN(new_n785));
  AND3_X1   g360(.A1(new_n784), .A2(new_n681), .A3(KEYINPUT94), .ZN(new_n786));
  AOI211_X1 g361(.A(new_n785), .B(new_n786), .C1(G171), .C2(G16), .ZN(new_n787));
  XNOR2_X1  g362(.A(new_n787), .B(G1961), .ZN(new_n788));
  NOR2_X1   g363(.A1(new_n745), .A2(new_n746), .ZN(new_n789));
  NOR2_X1   g364(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n688), .A2(new_n780), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n481), .A2(G131), .ZN(new_n792));
  XOR2_X1   g367(.A(new_n792), .B(KEYINPUT81), .Z(new_n793));
  INV_X1    g368(.A(G95), .ZN(new_n794));
  AND3_X1   g369(.A1(new_n794), .A2(new_n461), .A3(KEYINPUT82), .ZN(new_n795));
  AOI21_X1  g370(.A(KEYINPUT82), .B1(new_n794), .B2(new_n461), .ZN(new_n796));
  OAI221_X1 g371(.A(G2104), .B1(G107), .B2(new_n461), .C1(new_n795), .C2(new_n796), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n478), .A2(G119), .ZN(new_n798));
  NAND3_X1  g373(.A1(new_n793), .A2(new_n797), .A3(new_n798), .ZN(new_n799));
  MUX2_X1   g374(.A(G25), .B(new_n799), .S(G29), .Z(new_n800));
  XNOR2_X1  g375(.A(KEYINPUT35), .B(G1991), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n800), .B(new_n801), .ZN(new_n802));
  NAND2_X1  g377(.A1(new_n681), .A2(G22), .ZN(new_n803));
  OAI21_X1  g378(.A(new_n803), .B1(G166), .B2(new_n681), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n804), .B(G1971), .ZN(new_n805));
  NAND2_X1  g380(.A1(new_n681), .A2(G23), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n806), .B1(new_n577), .B2(new_n681), .ZN(new_n807));
  XOR2_X1   g382(.A(new_n807), .B(KEYINPUT33), .Z(new_n808));
  AOI21_X1  g383(.A(new_n805), .B1(new_n808), .B2(G1976), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n681), .A2(G6), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(new_n584), .B2(new_n681), .ZN(new_n811));
  XOR2_X1   g386(.A(KEYINPUT32), .B(G1981), .Z(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n813), .C1(G1976), .C2(new_n808), .ZN(new_n814));
  AOI21_X1  g389(.A(new_n802), .B1(new_n814), .B2(KEYINPUT34), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n681), .A2(G24), .ZN(new_n816));
  OAI21_X1  g391(.A(new_n816), .B1(new_n591), .B2(new_n681), .ZN(new_n817));
  XOR2_X1   g392(.A(KEYINPUT83), .B(G1986), .Z(new_n818));
  XNOR2_X1  g393(.A(new_n817), .B(new_n818), .ZN(new_n819));
  OAI211_X1 g394(.A(new_n815), .B(new_n819), .C1(KEYINPUT34), .C2(new_n814), .ZN(new_n820));
  OAI21_X1  g395(.A(KEYINPUT36), .B1(new_n820), .B2(KEYINPUT84), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n820), .A2(KEYINPUT84), .ZN(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n820), .A2(KEYINPUT84), .A3(KEYINPUT36), .ZN(new_n824));
  AOI211_X1 g399(.A(new_n678), .B(new_n791), .C1(new_n823), .C2(new_n824), .ZN(G311));
  AOI21_X1  g400(.A(new_n791), .B1(new_n823), .B2(new_n824), .ZN(new_n826));
  OAI21_X1  g401(.A(new_n826), .B1(G2078), .B2(new_n677), .ZN(G150));
  INV_X1    g402(.A(G55), .ZN(new_n828));
  AOI22_X1  g403(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n829));
  OAI22_X1  g404(.A1(new_n509), .A2(new_n828), .B1(new_n829), .B2(new_n518), .ZN(new_n830));
  INV_X1    g405(.A(G93), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n520), .A2(new_n831), .ZN(new_n832));
  OR2_X1    g407(.A1(new_n830), .A2(new_n832), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n833), .A2(G860), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT98), .ZN(new_n835));
  XNOR2_X1  g410(.A(new_n835), .B(KEYINPUT37), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n607), .A2(G559), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n837), .B(KEYINPUT38), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n833), .A2(new_n551), .ZN(new_n839));
  NOR2_X1   g414(.A1(new_n830), .A2(new_n832), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n840), .B1(new_n548), .B2(new_n550), .ZN(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n841), .ZN(new_n842));
  XNOR2_X1  g417(.A(new_n842), .B(KEYINPUT39), .ZN(new_n843));
  XNOR2_X1  g418(.A(new_n838), .B(new_n843), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n836), .B1(new_n844), .B2(G860), .ZN(G145));
  XNOR2_X1  g420(.A(new_n618), .B(G160), .ZN(new_n846));
  INV_X1    g421(.A(new_n703), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n799), .B(new_n485), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  INV_X1    g425(.A(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n772), .A2(new_n737), .ZN(new_n852));
  INV_X1    g427(.A(new_n737), .ZN(new_n853));
  NAND3_X1  g428(.A1(new_n767), .A2(new_n853), .A3(new_n771), .ZN(new_n854));
  NAND3_X1  g429(.A1(new_n852), .A2(G164), .A3(new_n854), .ZN(new_n855));
  AOI211_X1 g430(.A(new_n770), .B(new_n737), .C1(new_n765), .C2(new_n766), .ZN(new_n856));
  AOI21_X1  g431(.A(new_n853), .B1(new_n767), .B2(new_n771), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n497), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(new_n622), .ZN(new_n859));
  NAND3_X1  g434(.A1(new_n855), .A2(new_n858), .A3(new_n859), .ZN(new_n860));
  INV_X1    g435(.A(new_n860), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n859), .B1(new_n855), .B2(new_n858), .ZN(new_n862));
  NAND2_X1  g437(.A1(new_n478), .A2(G130), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n481), .A2(G142), .ZN(new_n864));
  OR2_X1    g439(.A1(G106), .A2(G2105), .ZN(new_n865));
  OAI211_X1 g440(.A(new_n865), .B(G2104), .C1(G118), .C2(new_n461), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n864), .A3(new_n866), .ZN(new_n867));
  NOR3_X1   g442(.A1(new_n861), .A2(new_n862), .A3(new_n867), .ZN(new_n868));
  INV_X1    g443(.A(new_n867), .ZN(new_n869));
  NAND2_X1  g444(.A1(new_n855), .A2(new_n858), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n870), .A2(new_n622), .ZN(new_n871));
  AOI21_X1  g446(.A(new_n869), .B1(new_n871), .B2(new_n860), .ZN(new_n872));
  OAI21_X1  g447(.A(new_n851), .B1(new_n868), .B2(new_n872), .ZN(new_n873));
  INV_X1    g448(.A(G37), .ZN(new_n874));
  OAI21_X1  g449(.A(new_n867), .B1(new_n861), .B2(new_n862), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n871), .A2(new_n869), .A3(new_n860), .ZN(new_n876));
  NAND3_X1  g451(.A1(new_n875), .A2(new_n876), .A3(new_n850), .ZN(new_n877));
  NAND3_X1  g452(.A1(new_n873), .A2(new_n874), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g453(.A1(new_n878), .A2(KEYINPUT99), .ZN(new_n879));
  INV_X1    g454(.A(KEYINPUT99), .ZN(new_n880));
  NAND4_X1  g455(.A1(new_n873), .A2(new_n880), .A3(new_n874), .A4(new_n877), .ZN(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g458(.A1(new_n833), .A2(G868), .ZN(new_n884));
  XNOR2_X1  g459(.A(new_n577), .B(KEYINPUT100), .ZN(new_n885));
  XNOR2_X1  g460(.A(new_n885), .B(G290), .ZN(new_n886));
  XOR2_X1   g461(.A(G166), .B(new_n584), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n887), .A2(KEYINPUT101), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n886), .A2(new_n888), .ZN(new_n889));
  OR2_X1    g464(.A1(new_n887), .A2(KEYINPUT101), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n890), .A2(new_n886), .A3(new_n888), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  XOR2_X1   g467(.A(new_n892), .B(KEYINPUT42), .Z(new_n893));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n894));
  AND2_X1   g469(.A1(new_n839), .A2(new_n841), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n610), .B(new_n895), .ZN(new_n896));
  INV_X1    g471(.A(KEYINPUT41), .ZN(new_n897));
  NAND2_X1  g472(.A1(new_n599), .A2(new_n568), .ZN(new_n898));
  INV_X1    g473(.A(new_n898), .ZN(new_n899));
  NOR2_X1   g474(.A1(new_n599), .A2(new_n568), .ZN(new_n900));
  OAI21_X1  g475(.A(new_n897), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n607), .A2(G299), .ZN(new_n902));
  NAND3_X1  g477(.A1(new_n902), .A2(KEYINPUT41), .A3(new_n898), .ZN(new_n903));
  AOI21_X1  g478(.A(new_n896), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n902), .A2(new_n898), .ZN(new_n905));
  AND2_X1   g480(.A1(new_n896), .A2(new_n905), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n894), .B1(new_n904), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n893), .A2(new_n907), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n904), .A2(new_n906), .A3(new_n894), .ZN(new_n909));
  XNOR2_X1  g484(.A(new_n908), .B(new_n909), .ZN(new_n910));
  AOI21_X1  g485(.A(new_n884), .B1(new_n910), .B2(G868), .ZN(G295));
  AOI21_X1  g486(.A(new_n884), .B1(new_n910), .B2(G868), .ZN(G331));
  INV_X1    g487(.A(KEYINPUT103), .ZN(new_n913));
  NAND2_X1  g488(.A1(new_n901), .A2(new_n903), .ZN(new_n914));
  NAND2_X1  g489(.A1(G171), .A2(new_n895), .ZN(new_n915));
  NAND2_X1  g490(.A1(G301), .A2(new_n842), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n917), .A2(G286), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n914), .A2(new_n918), .A3(new_n919), .ZN(new_n920));
  AND3_X1   g495(.A1(new_n915), .A2(new_n916), .A3(G168), .ZN(new_n921));
  AOI21_X1  g496(.A(G168), .B1(new_n915), .B2(new_n916), .ZN(new_n922));
  OAI21_X1  g497(.A(new_n905), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n913), .B1(new_n920), .B2(new_n923), .ZN(new_n924));
  NOR2_X1   g499(.A1(new_n921), .A2(new_n922), .ZN(new_n925));
  AOI21_X1  g500(.A(KEYINPUT103), .B1(new_n925), .B2(new_n914), .ZN(new_n926));
  NOR3_X1   g501(.A1(new_n924), .A2(new_n926), .A3(new_n892), .ZN(new_n927));
  NOR2_X1   g502(.A1(new_n927), .A2(G37), .ZN(new_n928));
  OAI21_X1  g503(.A(new_n892), .B1(new_n924), .B2(new_n926), .ZN(new_n929));
  AOI21_X1  g504(.A(KEYINPUT43), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  AOI22_X1  g505(.A1(new_n920), .A2(new_n923), .B1(new_n889), .B2(new_n891), .ZN(new_n931));
  INV_X1    g506(.A(KEYINPUT43), .ZN(new_n932));
  NOR4_X1   g507(.A1(new_n927), .A2(new_n931), .A3(new_n932), .A4(G37), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT44), .B1(new_n930), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(KEYINPUT44), .ZN(new_n935));
  AOI21_X1  g510(.A(new_n932), .B1(new_n928), .B2(new_n929), .ZN(new_n936));
  NOR4_X1   g511(.A1(new_n927), .A2(new_n931), .A3(KEYINPUT43), .A4(G37), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n935), .B1(new_n936), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  NAND2_X1  g514(.A1(new_n475), .A2(G2105), .ZN(new_n940));
  INV_X1    g515(.A(new_n466), .ZN(new_n941));
  AND4_X1   g516(.A1(KEYINPUT104), .A2(new_n940), .A3(G40), .A4(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT104), .B1(G160), .B2(G40), .ZN(new_n943));
  NOR2_X1   g518(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  INV_X1    g519(.A(G1384), .ZN(new_n945));
  INV_X1    g520(.A(new_n488), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n946), .B1(new_n460), .B2(G126), .ZN(new_n947));
  OAI211_X1 g522(.A(new_n496), .B(new_n494), .C1(new_n947), .C2(new_n461), .ZN(new_n948));
  INV_X1    g523(.A(new_n493), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n945), .B1(new_n948), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(KEYINPUT45), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n950), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g527(.A1(new_n944), .A2(new_n952), .ZN(new_n953));
  INV_X1    g528(.A(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n954), .A2(G1996), .ZN(new_n955));
  INV_X1    g530(.A(KEYINPUT126), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n956), .A2(KEYINPUT46), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n955), .B(new_n957), .Z(new_n958));
  NAND2_X1  g533(.A1(new_n853), .A2(G2067), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n737), .A2(new_n740), .ZN(new_n960));
  AND2_X1   g535(.A1(new_n959), .A2(new_n960), .ZN(new_n961));
  INV_X1    g536(.A(new_n961), .ZN(new_n962));
  OAI21_X1  g537(.A(new_n953), .B1(new_n962), .B2(new_n847), .ZN(new_n963));
  OAI211_X1 g538(.A(new_n958), .B(new_n963), .C1(new_n956), .C2(KEYINPUT46), .ZN(new_n964));
  XOR2_X1   g539(.A(KEYINPUT127), .B(KEYINPUT47), .Z(new_n965));
  XNOR2_X1  g540(.A(new_n964), .B(new_n965), .ZN(new_n966));
  XNOR2_X1  g541(.A(new_n703), .B(G1996), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n961), .A2(new_n967), .ZN(new_n968));
  NOR2_X1   g543(.A1(new_n799), .A2(new_n801), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(new_n960), .B1(new_n968), .B2(new_n970), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n953), .ZN(new_n972));
  NOR3_X1   g547(.A1(new_n954), .A2(G1986), .A3(G290), .ZN(new_n973));
  XOR2_X1   g548(.A(new_n973), .B(KEYINPUT48), .Z(new_n974));
  AND2_X1   g549(.A1(new_n799), .A2(new_n801), .ZN(new_n975));
  NOR3_X1   g550(.A1(new_n968), .A2(new_n969), .A3(new_n975), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n974), .B1(new_n976), .B2(new_n954), .ZN(new_n977));
  AND3_X1   g552(.A1(new_n966), .A2(new_n972), .A3(new_n977), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT63), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT52), .ZN(new_n980));
  INV_X1    g555(.A(G8), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n940), .A2(G40), .A3(new_n941), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT104), .ZN(new_n983));
  NAND2_X1  g558(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  NAND3_X1  g559(.A1(G160), .A2(KEYINPUT104), .A3(G40), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  INV_X1    g561(.A(new_n950), .ZN(new_n987));
  AOI21_X1  g562(.A(new_n981), .B1(new_n986), .B2(new_n987), .ZN(new_n988));
  NAND2_X1  g563(.A1(new_n577), .A2(G1976), .ZN(new_n989));
  AOI21_X1  g564(.A(new_n980), .B1(new_n988), .B2(new_n989), .ZN(new_n990));
  INV_X1    g565(.A(G1976), .ZN(new_n991));
  AOI21_X1  g566(.A(KEYINPUT52), .B1(G288), .B2(new_n991), .ZN(new_n992));
  NAND3_X1  g567(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(new_n993), .ZN(new_n994));
  XNOR2_X1  g569(.A(KEYINPUT109), .B(G1981), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n584), .A2(new_n995), .ZN(new_n996));
  XNOR2_X1  g571(.A(KEYINPUT110), .B(G86), .ZN(new_n997));
  NOR2_X1   g572(.A1(new_n520), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(G1981), .B1(new_n581), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n996), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1000), .A2(new_n1001), .ZN(new_n1002));
  NAND3_X1  g577(.A1(new_n996), .A2(KEYINPUT49), .A3(new_n999), .ZN(new_n1003));
  NAND3_X1  g578(.A1(new_n1002), .A2(new_n988), .A3(new_n1003), .ZN(new_n1004));
  NAND2_X1  g579(.A1(new_n1004), .A2(KEYINPUT111), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT111), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(new_n1006), .A3(new_n988), .A4(new_n1003), .ZN(new_n1007));
  AOI211_X1 g582(.A(new_n990), .B(new_n994), .C1(new_n1005), .C2(new_n1007), .ZN(new_n1008));
  OAI211_X1 g583(.A(KEYINPUT55), .B(G8), .C1(new_n519), .C2(new_n522), .ZN(new_n1009));
  OR2_X1    g584(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT55), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1011), .B1(G166), .B2(new_n981), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(KEYINPUT107), .ZN(new_n1013));
  NAND3_X1  g588(.A1(new_n1010), .A2(new_n1012), .A3(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(new_n1014), .ZN(new_n1015));
  AND3_X1   g590(.A1(new_n497), .A2(KEYINPUT50), .A3(new_n945), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT50), .B1(new_n497), .B2(new_n945), .ZN(new_n1017));
  OAI22_X1  g592(.A1(new_n942), .A2(new_n943), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  OR2_X1    g593(.A1(new_n1018), .A2(KEYINPUT112), .ZN(new_n1019));
  AOI21_X1  g594(.A(G2090), .B1(new_n1018), .B2(KEYINPUT112), .ZN(new_n1020));
  XOR2_X1   g595(.A(KEYINPUT106), .B(G1971), .Z(new_n1021));
  INV_X1    g596(.A(KEYINPUT105), .ZN(new_n1022));
  AND3_X1   g597(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n1023));
  AOI21_X1  g598(.A(KEYINPUT45), .B1(new_n497), .B2(new_n945), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1022), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  NAND2_X1  g600(.A1(new_n952), .A2(KEYINPUT105), .ZN(new_n1026));
  NAND3_X1  g601(.A1(new_n1025), .A2(new_n986), .A3(new_n1026), .ZN(new_n1027));
  AOI22_X1  g602(.A1(new_n1019), .A2(new_n1020), .B1(new_n1021), .B2(new_n1027), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1015), .B1(new_n1028), .B2(new_n981), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT50), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n950), .A2(new_n1030), .ZN(new_n1031));
  NAND3_X1  g606(.A1(new_n497), .A2(KEYINPUT50), .A3(new_n945), .ZN(new_n1032));
  AOI22_X1  g607(.A1(new_n984), .A2(new_n985), .B1(new_n1031), .B2(new_n1032), .ZN(new_n1033));
  INV_X1    g608(.A(G2090), .ZN(new_n1034));
  AOI22_X1  g609(.A1(new_n1027), .A2(new_n1021), .B1(new_n1033), .B2(new_n1034), .ZN(new_n1035));
  NOR2_X1   g610(.A1(new_n1035), .A2(new_n981), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1014), .ZN(new_n1037));
  INV_X1    g612(.A(KEYINPUT108), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1037), .A2(new_n1038), .ZN(new_n1039));
  AOI21_X1  g614(.A(KEYINPUT108), .B1(new_n1036), .B2(new_n1014), .ZN(new_n1040));
  OAI211_X1 g615(.A(new_n1008), .B(new_n1029), .C1(new_n1039), .C2(new_n1040), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n497), .A2(KEYINPUT45), .A3(new_n945), .ZN(new_n1042));
  NAND2_X1  g617(.A1(new_n952), .A2(new_n1042), .ZN(new_n1043));
  OAI21_X1  g618(.A(new_n782), .B1(new_n944), .B2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1045));
  INV_X1    g620(.A(G2084), .ZN(new_n1046));
  NAND3_X1  g621(.A1(new_n986), .A2(new_n1045), .A3(new_n1046), .ZN(new_n1047));
  AOI21_X1  g622(.A(new_n981), .B1(new_n1044), .B2(new_n1047), .ZN(new_n1048));
  NAND2_X1  g623(.A1(new_n1048), .A2(G168), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n979), .B1(new_n1041), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1005), .A2(new_n1007), .ZN(new_n1051));
  INV_X1    g626(.A(new_n990), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1015), .B1(new_n1035), .B2(new_n981), .ZN(new_n1053));
  NAND4_X1  g628(.A1(new_n1051), .A2(new_n1052), .A3(new_n993), .A4(new_n1053), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT113), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n979), .B1(new_n1054), .B2(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(new_n1037), .B(new_n1038), .ZN(new_n1057));
  INV_X1    g632(.A(new_n1049), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1008), .A2(KEYINPUT113), .A3(new_n1053), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1056), .A2(new_n1057), .A3(new_n1058), .A4(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1050), .A2(new_n1060), .ZN(new_n1061));
  INV_X1    g636(.A(new_n1057), .ZN(new_n1062));
  NAND3_X1  g637(.A1(new_n1051), .A2(new_n991), .A3(new_n577), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(new_n996), .ZN(new_n1064));
  AOI22_X1  g639(.A1(new_n1062), .A2(new_n1008), .B1(new_n1064), .B2(new_n988), .ZN(new_n1065));
  NAND2_X1  g640(.A1(new_n1061), .A2(new_n1065), .ZN(new_n1066));
  OAI211_X1 g641(.A(new_n952), .B(new_n1042), .C1(new_n942), .C2(new_n943), .ZN(new_n1067));
  AOI22_X1  g642(.A1(new_n1033), .A2(new_n1046), .B1(new_n1067), .B2(new_n782), .ZN(new_n1068));
  NOR3_X1   g643(.A1(new_n1068), .A2(new_n981), .A3(G168), .ZN(new_n1069));
  INV_X1    g644(.A(new_n1069), .ZN(new_n1070));
  AOI21_X1  g645(.A(new_n981), .B1(new_n1068), .B2(G168), .ZN(new_n1071));
  AOI21_X1  g646(.A(KEYINPUT51), .B1(new_n1071), .B2(KEYINPUT122), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1044), .A2(new_n1047), .ZN(new_n1073));
  OAI211_X1 g648(.A(KEYINPUT122), .B(G8), .C1(new_n1073), .C2(G286), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  NOR2_X1   g650(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1076));
  OAI21_X1  g651(.A(new_n1070), .B1(new_n1072), .B2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(KEYINPUT123), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT62), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1080));
  NOR2_X1   g655(.A1(G168), .A2(new_n981), .ZN(new_n1081));
  OAI211_X1 g656(.A(KEYINPUT122), .B(KEYINPUT51), .C1(new_n1081), .C2(new_n1048), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1080), .A2(new_n1082), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n1084));
  NAND3_X1  g659(.A1(new_n1083), .A2(new_n1084), .A3(new_n1070), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1078), .A2(new_n1079), .A3(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1084), .B1(new_n1083), .B2(new_n1070), .ZN(new_n1087));
  AOI211_X1 g662(.A(KEYINPUT123), .B(new_n1069), .C1(new_n1080), .C2(new_n1082), .ZN(new_n1088));
  OAI21_X1  g663(.A(KEYINPUT62), .B1(new_n1087), .B2(new_n1088), .ZN(new_n1089));
  NAND2_X1  g664(.A1(new_n1086), .A2(new_n1089), .ZN(new_n1090));
  INV_X1    g665(.A(new_n1067), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT53), .ZN(new_n1092));
  NOR2_X1   g667(.A1(new_n1092), .A2(G2078), .ZN(new_n1093));
  INV_X1    g668(.A(G1961), .ZN(new_n1094));
  AOI22_X1  g669(.A1(new_n1091), .A2(new_n1093), .B1(new_n1094), .B2(new_n1018), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n1092), .B1(new_n1027), .B2(G2078), .ZN(new_n1096));
  AOI21_X1  g671(.A(G301), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1097), .ZN(new_n1098));
  INV_X1    g673(.A(KEYINPUT54), .ZN(new_n1099));
  INV_X1    g674(.A(new_n1043), .ZN(new_n1100));
  NOR3_X1   g675(.A1(new_n982), .A2(new_n1092), .A3(G2078), .ZN(new_n1101));
  AOI22_X1  g676(.A1(new_n1018), .A2(new_n1094), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1102));
  AND3_X1   g677(.A1(new_n1096), .A2(G301), .A3(new_n1102), .ZN(new_n1103));
  OAI21_X1  g678(.A(new_n1099), .B1(new_n1103), .B2(new_n1097), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT124), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  OAI211_X1 g681(.A(KEYINPUT124), .B(new_n1099), .C1(new_n1103), .C2(new_n1097), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1095), .A2(new_n1096), .A3(G301), .ZN(new_n1109));
  AND2_X1   g684(.A1(new_n1096), .A2(new_n1102), .ZN(new_n1110));
  OAI211_X1 g685(.A(KEYINPUT54), .B(new_n1109), .C1(new_n1110), .C2(G301), .ZN(new_n1111));
  OAI211_X1 g686(.A(new_n1108), .B(new_n1111), .C1(new_n1087), .C2(new_n1088), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT118), .ZN(new_n1113));
  OAI211_X1 g688(.A(new_n740), .B(new_n987), .C1(new_n942), .C2(new_n943), .ZN(new_n1114));
  NAND2_X1  g689(.A1(new_n1114), .A2(KEYINPUT117), .ZN(new_n1115));
  INV_X1    g690(.A(G1348), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1018), .A2(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(KEYINPUT117), .ZN(new_n1118));
  NAND4_X1  g693(.A1(new_n986), .A2(new_n1118), .A3(new_n740), .A4(new_n987), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1115), .A2(new_n1117), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n607), .ZN(new_n1121));
  INV_X1    g696(.A(new_n567), .ZN(new_n1122));
  NOR3_X1   g697(.A1(new_n509), .A2(KEYINPUT9), .A3(new_n566), .ZN(new_n1123));
  OAI21_X1  g698(.A(KEYINPUT115), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  INV_X1    g699(.A(KEYINPUT116), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT57), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1124), .A2(new_n1125), .A3(new_n1126), .ZN(new_n1127));
  INV_X1    g702(.A(KEYINPUT115), .ZN(new_n1128));
  AOI21_X1  g703(.A(new_n1128), .B1(new_n565), .B2(new_n567), .ZN(new_n1129));
  OAI21_X1  g704(.A(KEYINPUT116), .B1(new_n1129), .B2(KEYINPUT57), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1127), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1131), .A2(G299), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1127), .A2(new_n1130), .A3(new_n568), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI21_X1  g709(.A(KEYINPUT114), .B1(new_n1033), .B2(G1956), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT114), .ZN(new_n1136));
  INV_X1    g711(.A(G1956), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1018), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1138));
  AND3_X1   g713(.A1(new_n1025), .A2(new_n986), .A3(new_n1026), .ZN(new_n1139));
  XNOR2_X1  g714(.A(KEYINPUT56), .B(G2072), .ZN(new_n1140));
  AOI22_X1  g715(.A1(new_n1135), .A2(new_n1138), .B1(new_n1139), .B2(new_n1140), .ZN(new_n1141));
  AOI21_X1  g716(.A(new_n1121), .B1(new_n1134), .B2(new_n1141), .ZN(new_n1142));
  NOR2_X1   g717(.A1(new_n1141), .A2(new_n1134), .ZN(new_n1143));
  OAI21_X1  g718(.A(new_n1113), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AND3_X1   g719(.A1(new_n1127), .A2(new_n568), .A3(new_n1130), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n568), .B1(new_n1127), .B2(new_n1130), .ZN(new_n1146));
  NOR2_X1   g721(.A1(new_n1145), .A2(new_n1146), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1025), .A2(new_n986), .A3(new_n1026), .A4(new_n1140), .ZN(new_n1148));
  AND3_X1   g723(.A1(new_n1018), .A2(new_n1136), .A3(new_n1137), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1136), .B1(new_n1018), .B2(new_n1137), .ZN(new_n1150));
  OAI21_X1  g725(.A(new_n1148), .B1(new_n1149), .B2(new_n1150), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  NOR2_X1   g727(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1153));
  OAI211_X1 g728(.A(KEYINPUT118), .B(new_n1152), .C1(new_n1153), .C2(new_n1121), .ZN(new_n1154));
  NAND2_X1  g729(.A1(new_n1144), .A2(new_n1154), .ZN(new_n1155));
  XOR2_X1   g730(.A(KEYINPUT120), .B(KEYINPUT61), .Z(new_n1156));
  NAND2_X1  g731(.A1(new_n1141), .A2(new_n1134), .ZN(new_n1157));
  AOI21_X1  g732(.A(new_n1156), .B1(new_n1157), .B2(new_n1152), .ZN(new_n1158));
  AND2_X1   g733(.A1(new_n1115), .A2(new_n1119), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT60), .ZN(new_n1160));
  NAND4_X1  g735(.A1(new_n1159), .A2(new_n1160), .A3(new_n607), .A4(new_n1117), .ZN(new_n1161));
  XOR2_X1   g736(.A(KEYINPUT58), .B(G1341), .Z(new_n1162));
  OAI21_X1  g737(.A(new_n1162), .B1(new_n944), .B2(new_n950), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(new_n1027), .B2(G1996), .ZN(new_n1164));
  OR2_X1    g739(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g740(.A1(KEYINPUT119), .A2(KEYINPUT59), .ZN(new_n1166));
  NAND4_X1  g741(.A1(new_n1164), .A2(new_n551), .A3(new_n1165), .A4(new_n1166), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n1164), .A2(new_n551), .ZN(new_n1168));
  OAI211_X1 g743(.A(new_n1161), .B(new_n1167), .C1(new_n1168), .C2(new_n1165), .ZN(new_n1169));
  NAND3_X1  g744(.A1(new_n1159), .A2(new_n599), .A3(new_n1117), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n1160), .B1(new_n1170), .B2(new_n1121), .ZN(new_n1171));
  NOR3_X1   g746(.A1(new_n1158), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  OR2_X1    g747(.A1(new_n1157), .A2(KEYINPUT121), .ZN(new_n1173));
  NAND2_X1  g748(.A1(new_n1157), .A2(KEYINPUT121), .ZN(new_n1174));
  NAND4_X1  g749(.A1(new_n1173), .A2(KEYINPUT61), .A3(new_n1174), .A4(new_n1152), .ZN(new_n1175));
  AOI21_X1  g750(.A(new_n1155), .B1(new_n1172), .B2(new_n1175), .ZN(new_n1176));
  OAI22_X1  g751(.A1(new_n1090), .A2(new_n1098), .B1(new_n1112), .B2(new_n1176), .ZN(new_n1177));
  XNOR2_X1  g752(.A(new_n1041), .B(KEYINPUT125), .ZN(new_n1178));
  AOI21_X1  g753(.A(new_n1066), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  XNOR2_X1  g754(.A(new_n591), .B(G1986), .ZN(new_n1180));
  AOI21_X1  g755(.A(new_n954), .B1(new_n976), .B2(new_n1180), .ZN(new_n1181));
  OAI21_X1  g756(.A(new_n978), .B1(new_n1179), .B2(new_n1181), .ZN(G329));
  assign    G231 = 1'b0;
  OR2_X1    g757(.A1(G227), .A2(G401), .ZN(new_n1184));
  AOI21_X1  g758(.A(new_n1184), .B1(new_n879), .B2(new_n881), .ZN(new_n1185));
  NOR2_X1   g759(.A1(G229), .A2(new_n458), .ZN(new_n1186));
  OAI211_X1 g760(.A(new_n1185), .B(new_n1186), .C1(new_n936), .C2(new_n937), .ZN(G225));
  INV_X1    g761(.A(G225), .ZN(G308));
endmodule


