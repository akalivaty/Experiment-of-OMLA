

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591;

  INV_X1 U323 ( .A(KEYINPUT90), .ZN(n314) );
  XNOR2_X1 U324 ( .A(KEYINPUT120), .B(KEYINPUT54), .ZN(n291) );
  INV_X1 U325 ( .A(KEYINPUT46), .ZN(n457) );
  INV_X1 U326 ( .A(KEYINPUT98), .ZN(n397) );
  XNOR2_X1 U327 ( .A(KEYINPUT32), .B(KEYINPUT72), .ZN(n439) );
  XNOR2_X1 U328 ( .A(n315), .B(n314), .ZN(n316) );
  XNOR2_X1 U329 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U330 ( .A(n414), .B(n316), .ZN(n319) );
  XNOR2_X1 U331 ( .A(n450), .B(n449), .ZN(n581) );
  XOR2_X1 U332 ( .A(n328), .B(n344), .Z(n526) );
  XNOR2_X1 U333 ( .A(KEYINPUT58), .B(G190GAT), .ZN(n477) );
  XNOR2_X1 U334 ( .A(n453), .B(n452), .ZN(n454) );
  XNOR2_X1 U335 ( .A(n478), .B(n477), .ZN(G1351GAT) );
  XOR2_X1 U336 ( .A(KEYINPUT81), .B(KEYINPUT24), .Z(n293) );
  XNOR2_X1 U337 ( .A(G218GAT), .B(KEYINPUT22), .ZN(n292) );
  XNOR2_X1 U338 ( .A(n293), .B(n292), .ZN(n312) );
  XOR2_X1 U339 ( .A(KEYINPUT82), .B(KEYINPUT23), .Z(n295) );
  NAND2_X1 U340 ( .A1(G228GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U341 ( .A(n295), .B(n294), .ZN(n296) );
  XOR2_X1 U342 ( .A(n296), .B(G204GAT), .Z(n301) );
  XNOR2_X1 U343 ( .A(G155GAT), .B(KEYINPUT3), .ZN(n297) );
  XNOR2_X1 U344 ( .A(n297), .B(KEYINPUT2), .ZN(n356) );
  XOR2_X1 U345 ( .A(G197GAT), .B(KEYINPUT21), .Z(n299) );
  XNOR2_X1 U346 ( .A(G211GAT), .B(KEYINPUT80), .ZN(n298) );
  XNOR2_X1 U347 ( .A(n299), .B(n298), .ZN(n322) );
  XNOR2_X1 U348 ( .A(n356), .B(n322), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(G141GAT), .B(G22GAT), .Z(n424) );
  XOR2_X1 U351 ( .A(n302), .B(n424), .Z(n310) );
  XOR2_X1 U352 ( .A(G162GAT), .B(G50GAT), .Z(n401) );
  INV_X1 U353 ( .A(G78GAT), .ZN(n303) );
  NAND2_X1 U354 ( .A1(KEYINPUT71), .A2(n303), .ZN(n306) );
  INV_X1 U355 ( .A(KEYINPUT71), .ZN(n304) );
  NAND2_X1 U356 ( .A1(n304), .A2(G78GAT), .ZN(n305) );
  NAND2_X1 U357 ( .A1(n306), .A2(n305), .ZN(n308) );
  XNOR2_X1 U358 ( .A(G148GAT), .B(G106GAT), .ZN(n307) );
  XNOR2_X1 U359 ( .A(n308), .B(n307), .ZN(n440) );
  XNOR2_X1 U360 ( .A(n401), .B(n440), .ZN(n309) );
  XNOR2_X1 U361 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U362 ( .A(n312), .B(n311), .Z(n471) );
  XOR2_X1 U363 ( .A(KEYINPUT28), .B(n471), .Z(n518) );
  XNOR2_X1 U364 ( .A(G218GAT), .B(G36GAT), .ZN(n313) );
  XNOR2_X1 U365 ( .A(n313), .B(G190GAT), .ZN(n414) );
  NAND2_X1 U366 ( .A1(G226GAT), .A2(G233GAT), .ZN(n315) );
  XOR2_X1 U367 ( .A(G8GAT), .B(G169GAT), .Z(n431) );
  XNOR2_X1 U368 ( .A(n431), .B(KEYINPUT88), .ZN(n317) );
  XNOR2_X1 U369 ( .A(n317), .B(KEYINPUT89), .ZN(n318) );
  XOR2_X1 U370 ( .A(n319), .B(n318), .Z(n324) );
  XOR2_X1 U371 ( .A(G204GAT), .B(G176GAT), .Z(n321) );
  XNOR2_X1 U372 ( .A(G92GAT), .B(G64GAT), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n321), .B(n320), .ZN(n443) );
  XNOR2_X1 U374 ( .A(n322), .B(n443), .ZN(n323) );
  XNOR2_X1 U375 ( .A(n324), .B(n323), .ZN(n328) );
  XOR2_X1 U376 ( .A(KEYINPUT78), .B(KEYINPUT17), .Z(n326) );
  XNOR2_X1 U377 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n325) );
  XNOR2_X1 U378 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U379 ( .A(G183GAT), .B(n327), .ZN(n344) );
  INV_X1 U380 ( .A(n526), .ZN(n501) );
  XOR2_X1 U381 ( .A(G120GAT), .B(G71GAT), .Z(n437) );
  XOR2_X1 U382 ( .A(KEYINPUT65), .B(G99GAT), .Z(n330) );
  XNOR2_X1 U383 ( .A(G43GAT), .B(G190GAT), .ZN(n329) );
  XNOR2_X1 U384 ( .A(n330), .B(n329), .ZN(n331) );
  XNOR2_X1 U385 ( .A(n437), .B(n331), .ZN(n333) );
  AND2_X1 U386 ( .A1(G227GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n335) );
  INV_X1 U388 ( .A(KEYINPUT79), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n339) );
  XOR2_X1 U390 ( .A(G113GAT), .B(G127GAT), .Z(n337) );
  XNOR2_X1 U391 ( .A(G134GAT), .B(KEYINPUT0), .ZN(n336) );
  XNOR2_X1 U392 ( .A(n337), .B(n336), .ZN(n360) );
  XNOR2_X1 U393 ( .A(n360), .B(KEYINPUT77), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n343) );
  XOR2_X1 U395 ( .A(KEYINPUT20), .B(G169GAT), .Z(n341) );
  XNOR2_X1 U396 ( .A(G15GAT), .B(G176GAT), .ZN(n340) );
  XNOR2_X1 U397 ( .A(n341), .B(n340), .ZN(n342) );
  XNOR2_X1 U398 ( .A(n343), .B(n342), .ZN(n345) );
  XOR2_X1 U399 ( .A(n345), .B(n344), .Z(n350) );
  INV_X1 U400 ( .A(n350), .ZN(n503) );
  NOR2_X1 U401 ( .A1(n501), .A2(n503), .ZN(n347) );
  INV_X1 U402 ( .A(n471), .ZN(n346) );
  NOR2_X1 U403 ( .A1(n347), .A2(n346), .ZN(n348) );
  XNOR2_X1 U404 ( .A(n348), .B(KEYINPUT25), .ZN(n353) );
  XNOR2_X1 U405 ( .A(KEYINPUT91), .B(KEYINPUT27), .ZN(n349) );
  XOR2_X1 U406 ( .A(n526), .B(n349), .Z(n377) );
  NOR2_X1 U407 ( .A1(n350), .A2(n471), .ZN(n351) );
  XNOR2_X1 U408 ( .A(KEYINPUT26), .B(n351), .ZN(n574) );
  NAND2_X1 U409 ( .A1(n377), .A2(n574), .ZN(n352) );
  NAND2_X1 U410 ( .A1(n353), .A2(n352), .ZN(n375) );
  XOR2_X1 U411 ( .A(KEYINPUT5), .B(G57GAT), .Z(n355) );
  XNOR2_X1 U412 ( .A(KEYINPUT1), .B(KEYINPUT6), .ZN(n354) );
  XNOR2_X1 U413 ( .A(n355), .B(n354), .ZN(n374) );
  XOR2_X1 U414 ( .A(G85GAT), .B(G162GAT), .Z(n358) );
  XNOR2_X1 U415 ( .A(G120GAT), .B(n356), .ZN(n357) );
  XNOR2_X1 U416 ( .A(n358), .B(n357), .ZN(n359) );
  XNOR2_X1 U417 ( .A(G29GAT), .B(n359), .ZN(n372) );
  XOR2_X1 U418 ( .A(n360), .B(KEYINPUT4), .Z(n362) );
  NAND2_X1 U419 ( .A1(G225GAT), .A2(G233GAT), .ZN(n361) );
  XNOR2_X1 U420 ( .A(n362), .B(n361), .ZN(n366) );
  XOR2_X1 U421 ( .A(KEYINPUT83), .B(KEYINPUT87), .Z(n364) );
  XNOR2_X1 U422 ( .A(KEYINPUT85), .B(KEYINPUT86), .ZN(n363) );
  XNOR2_X1 U423 ( .A(n364), .B(n363), .ZN(n365) );
  XNOR2_X1 U424 ( .A(n366), .B(n365), .ZN(n370) );
  XOR2_X1 U425 ( .A(KEYINPUT84), .B(G1GAT), .Z(n368) );
  XNOR2_X1 U426 ( .A(G148GAT), .B(G141GAT), .ZN(n367) );
  XNOR2_X1 U427 ( .A(n368), .B(n367), .ZN(n369) );
  XNOR2_X1 U428 ( .A(n370), .B(n369), .ZN(n371) );
  XNOR2_X1 U429 ( .A(n372), .B(n371), .ZN(n373) );
  XOR2_X1 U430 ( .A(n374), .B(n373), .Z(n524) );
  INV_X1 U431 ( .A(n524), .ZN(n572) );
  NAND2_X1 U432 ( .A1(n375), .A2(n572), .ZN(n376) );
  XNOR2_X1 U433 ( .A(n376), .B(KEYINPUT92), .ZN(n379) );
  NAND2_X1 U434 ( .A1(n524), .A2(n377), .ZN(n547) );
  NOR2_X1 U435 ( .A1(n518), .A2(n547), .ZN(n532) );
  NAND2_X1 U436 ( .A1(n532), .A2(n503), .ZN(n378) );
  NAND2_X1 U437 ( .A1(n379), .A2(n378), .ZN(n380) );
  XOR2_X1 U438 ( .A(KEYINPUT93), .B(n380), .Z(n482) );
  XOR2_X1 U439 ( .A(G78GAT), .B(G211GAT), .Z(n382) );
  XNOR2_X1 U440 ( .A(G127GAT), .B(G155GAT), .ZN(n381) );
  XNOR2_X1 U441 ( .A(n382), .B(n381), .ZN(n396) );
  XOR2_X1 U442 ( .A(G1GAT), .B(G15GAT), .Z(n432) );
  XNOR2_X1 U443 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n383) );
  XNOR2_X1 U444 ( .A(n383), .B(KEYINPUT70), .ZN(n444) );
  XOR2_X1 U445 ( .A(n432), .B(n444), .Z(n385) );
  XNOR2_X1 U446 ( .A(G183GAT), .B(G71GAT), .ZN(n384) );
  XNOR2_X1 U447 ( .A(n385), .B(n384), .ZN(n389) );
  XOR2_X1 U448 ( .A(KEYINPUT12), .B(KEYINPUT75), .Z(n387) );
  NAND2_X1 U449 ( .A1(G231GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U450 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U451 ( .A(n389), .B(n388), .Z(n394) );
  XOR2_X1 U452 ( .A(KEYINPUT14), .B(G64GAT), .Z(n391) );
  XNOR2_X1 U453 ( .A(G22GAT), .B(G8GAT), .ZN(n390) );
  XNOR2_X1 U454 ( .A(n391), .B(n390), .ZN(n392) );
  XNOR2_X1 U455 ( .A(n392), .B(KEYINPUT15), .ZN(n393) );
  XNOR2_X1 U456 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U457 ( .A(n396), .B(n395), .Z(n557) );
  NAND2_X1 U458 ( .A1(n482), .A2(n557), .ZN(n398) );
  XNOR2_X1 U459 ( .A(n398), .B(n397), .ZN(n417) );
  XOR2_X1 U460 ( .A(G92GAT), .B(KEYINPUT64), .Z(n400) );
  XNOR2_X1 U461 ( .A(KEYINPUT11), .B(KEYINPUT73), .ZN(n399) );
  XNOR2_X1 U462 ( .A(n400), .B(n399), .ZN(n405) );
  XOR2_X1 U463 ( .A(G106GAT), .B(KEYINPUT67), .Z(n403) );
  XOR2_X1 U464 ( .A(G85GAT), .B(G99GAT), .Z(n448) );
  XNOR2_X1 U465 ( .A(n401), .B(n448), .ZN(n402) );
  XNOR2_X1 U466 ( .A(n403), .B(n402), .ZN(n404) );
  XOR2_X1 U467 ( .A(n405), .B(n404), .Z(n407) );
  NAND2_X1 U468 ( .A1(G232GAT), .A2(G233GAT), .ZN(n406) );
  XNOR2_X1 U469 ( .A(n407), .B(n406), .ZN(n411) );
  XOR2_X1 U470 ( .A(KEYINPUT74), .B(KEYINPUT9), .Z(n409) );
  XNOR2_X1 U471 ( .A(G134GAT), .B(KEYINPUT10), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n409), .B(n408), .ZN(n410) );
  XOR2_X1 U473 ( .A(n411), .B(n410), .Z(n416) );
  XOR2_X1 U474 ( .A(G43GAT), .B(KEYINPUT7), .Z(n413) );
  XNOR2_X1 U475 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n412) );
  XNOR2_X1 U476 ( .A(n413), .B(n412), .ZN(n423) );
  XNOR2_X1 U477 ( .A(n423), .B(n414), .ZN(n415) );
  XOR2_X1 U478 ( .A(n416), .B(n415), .Z(n561) );
  XOR2_X1 U479 ( .A(KEYINPUT36), .B(n561), .Z(n587) );
  NAND2_X1 U480 ( .A1(n417), .A2(n587), .ZN(n418) );
  XNOR2_X1 U481 ( .A(n418), .B(KEYINPUT37), .ZN(n420) );
  XNOR2_X1 U482 ( .A(KEYINPUT99), .B(KEYINPUT100), .ZN(n419) );
  XNOR2_X1 U483 ( .A(n420), .B(n419), .ZN(n496) );
  XOR2_X1 U484 ( .A(G197GAT), .B(G50GAT), .Z(n422) );
  XNOR2_X1 U485 ( .A(G113GAT), .B(G36GAT), .ZN(n421) );
  XNOR2_X1 U486 ( .A(n422), .B(n421), .ZN(n436) );
  XOR2_X1 U487 ( .A(n424), .B(n423), .Z(n426) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n425) );
  XNOR2_X1 U489 ( .A(n426), .B(n425), .ZN(n430) );
  XOR2_X1 U490 ( .A(KEYINPUT69), .B(KEYINPUT30), .Z(n428) );
  XNOR2_X1 U491 ( .A(KEYINPUT29), .B(KEYINPUT68), .ZN(n427) );
  XNOR2_X1 U492 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U493 ( .A(n430), .B(n429), .Z(n434) );
  XNOR2_X1 U494 ( .A(n432), .B(n431), .ZN(n433) );
  XNOR2_X1 U495 ( .A(n434), .B(n433), .ZN(n435) );
  XOR2_X1 U496 ( .A(n436), .B(n435), .Z(n549) );
  XNOR2_X1 U497 ( .A(n437), .B(KEYINPUT33), .ZN(n438) );
  XNOR2_X1 U498 ( .A(n438), .B(KEYINPUT31), .ZN(n442) );
  XOR2_X1 U499 ( .A(n442), .B(n441), .Z(n446) );
  XNOR2_X1 U500 ( .A(n444), .B(n443), .ZN(n445) );
  XNOR2_X1 U501 ( .A(n446), .B(n445), .ZN(n450) );
  NAND2_X1 U502 ( .A1(G230GAT), .A2(G233GAT), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XNOR2_X1 U504 ( .A(n581), .B(KEYINPUT41), .ZN(n456) );
  XNOR2_X1 U505 ( .A(n456), .B(KEYINPUT103), .ZN(n564) );
  NAND2_X1 U506 ( .A1(n549), .A2(n564), .ZN(n511) );
  NOR2_X1 U507 ( .A1(n496), .A2(n511), .ZN(n451) );
  XNOR2_X1 U508 ( .A(KEYINPUT108), .B(n451), .ZN(n530) );
  NAND2_X1 U509 ( .A1(n518), .A2(n530), .ZN(n455) );
  XOR2_X1 U510 ( .A(KEYINPUT112), .B(KEYINPUT44), .Z(n453) );
  XNOR2_X1 U511 ( .A(G106GAT), .B(KEYINPUT111), .ZN(n452) );
  XNOR2_X1 U512 ( .A(n455), .B(n454), .ZN(G1339GAT) );
  XOR2_X1 U513 ( .A(KEYINPUT121), .B(KEYINPUT122), .Z(n474) );
  XOR2_X1 U514 ( .A(KEYINPUT47), .B(KEYINPUT113), .Z(n462) );
  NOR2_X1 U515 ( .A1(n549), .A2(n456), .ZN(n458) );
  XNOR2_X1 U516 ( .A(n458), .B(n457), .ZN(n460) );
  INV_X1 U517 ( .A(n561), .ZN(n542) );
  INV_X1 U518 ( .A(n557), .ZN(n585) );
  NOR2_X1 U519 ( .A1(n542), .A2(n585), .ZN(n459) );
  NAND2_X1 U520 ( .A1(n460), .A2(n459), .ZN(n461) );
  XNOR2_X1 U521 ( .A(n462), .B(n461), .ZN(n468) );
  INV_X1 U522 ( .A(n549), .ZN(n576) );
  INV_X1 U523 ( .A(n581), .ZN(n479) );
  XOR2_X1 U524 ( .A(KEYINPUT66), .B(KEYINPUT45), .Z(n464) );
  NAND2_X1 U525 ( .A1(n585), .A2(n587), .ZN(n463) );
  XNOR2_X1 U526 ( .A(n464), .B(n463), .ZN(n465) );
  NAND2_X1 U527 ( .A1(n479), .A2(n465), .ZN(n466) );
  NOR2_X1 U528 ( .A1(n576), .A2(n466), .ZN(n467) );
  NOR2_X1 U529 ( .A1(n468), .A2(n467), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n469), .B(KEYINPUT48), .ZN(n546) );
  NOR2_X1 U531 ( .A1(n501), .A2(n546), .ZN(n470) );
  XNOR2_X1 U532 ( .A(n470), .B(n291), .ZN(n571) );
  AND2_X1 U533 ( .A1(n572), .A2(n471), .ZN(n472) );
  NAND2_X1 U534 ( .A1(n571), .A2(n472), .ZN(n473) );
  XNOR2_X1 U535 ( .A(n474), .B(n473), .ZN(n475) );
  XOR2_X1 U536 ( .A(KEYINPUT55), .B(n475), .Z(n476) );
  NOR2_X2 U537 ( .A1(n503), .A2(n476), .ZN(n569) );
  NAND2_X1 U538 ( .A1(n569), .A2(n542), .ZN(n478) );
  XOR2_X1 U539 ( .A(KEYINPUT95), .B(KEYINPUT34), .Z(n486) );
  NAND2_X1 U540 ( .A1(n479), .A2(n576), .ZN(n495) );
  XNOR2_X1 U541 ( .A(KEYINPUT76), .B(KEYINPUT16), .ZN(n481) );
  NOR2_X1 U542 ( .A1(n542), .A2(n557), .ZN(n480) );
  XNOR2_X1 U543 ( .A(n481), .B(n480), .ZN(n483) );
  NAND2_X1 U544 ( .A1(n483), .A2(n482), .ZN(n510) );
  NOR2_X1 U545 ( .A1(n495), .A2(n510), .ZN(n484) );
  XNOR2_X1 U546 ( .A(KEYINPUT94), .B(n484), .ZN(n492) );
  NAND2_X1 U547 ( .A1(n524), .A2(n492), .ZN(n485) );
  XNOR2_X1 U548 ( .A(n486), .B(n485), .ZN(n487) );
  XNOR2_X1 U549 ( .A(G1GAT), .B(n487), .ZN(G1324GAT) );
  NAND2_X1 U550 ( .A1(n492), .A2(n526), .ZN(n488) );
  XNOR2_X1 U551 ( .A(n488), .B(KEYINPUT96), .ZN(n489) );
  XNOR2_X1 U552 ( .A(G8GAT), .B(n489), .ZN(G1325GAT) );
  XOR2_X1 U553 ( .A(G15GAT), .B(KEYINPUT35), .Z(n491) );
  INV_X1 U554 ( .A(n503), .ZN(n533) );
  NAND2_X1 U555 ( .A1(n533), .A2(n492), .ZN(n490) );
  XNOR2_X1 U556 ( .A(n491), .B(n490), .ZN(G1326GAT) );
  XOR2_X1 U557 ( .A(G22GAT), .B(KEYINPUT97), .Z(n494) );
  NAND2_X1 U558 ( .A1(n518), .A2(n492), .ZN(n493) );
  XNOR2_X1 U559 ( .A(n494), .B(n493), .ZN(G1327GAT) );
  NOR2_X1 U560 ( .A1(n496), .A2(n495), .ZN(n498) );
  XNOR2_X1 U561 ( .A(KEYINPUT101), .B(KEYINPUT38), .ZN(n497) );
  XNOR2_X1 U562 ( .A(n498), .B(n497), .ZN(n507) );
  NOR2_X1 U563 ( .A1(n507), .A2(n572), .ZN(n500) );
  XNOR2_X1 U564 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n499) );
  XNOR2_X1 U565 ( .A(n500), .B(n499), .ZN(G1328GAT) );
  NOR2_X1 U566 ( .A1(n501), .A2(n507), .ZN(n502) );
  XOR2_X1 U567 ( .A(G36GAT), .B(n502), .Z(G1329GAT) );
  NOR2_X1 U568 ( .A1(n507), .A2(n503), .ZN(n504) );
  XOR2_X1 U569 ( .A(KEYINPUT40), .B(n504), .Z(n505) );
  XNOR2_X1 U570 ( .A(G43GAT), .B(n505), .ZN(G1330GAT) );
  INV_X1 U571 ( .A(n518), .ZN(n506) );
  NOR2_X1 U572 ( .A1(n507), .A2(n506), .ZN(n508) );
  XOR2_X1 U573 ( .A(KEYINPUT102), .B(n508), .Z(n509) );
  XNOR2_X1 U574 ( .A(G50GAT), .B(n509), .ZN(G1331GAT) );
  XNOR2_X1 U575 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n513) );
  NOR2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n519) );
  NAND2_X1 U577 ( .A1(n524), .A2(n519), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n513), .B(n512), .ZN(G1332GAT) );
  XOR2_X1 U579 ( .A(KEYINPUT104), .B(KEYINPUT105), .Z(n515) );
  NAND2_X1 U580 ( .A1(n519), .A2(n526), .ZN(n514) );
  XNOR2_X1 U581 ( .A(n515), .B(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G64GAT), .B(n516), .ZN(G1333GAT) );
  NAND2_X1 U583 ( .A1(n519), .A2(n533), .ZN(n517) );
  XNOR2_X1 U584 ( .A(n517), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U585 ( .A(KEYINPUT106), .B(KEYINPUT43), .Z(n521) );
  NAND2_X1 U586 ( .A1(n519), .A2(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(n521), .B(n520), .ZN(n523) );
  XOR2_X1 U588 ( .A(G78GAT), .B(KEYINPUT107), .Z(n522) );
  XNOR2_X1 U589 ( .A(n523), .B(n522), .ZN(G1335GAT) );
  NAND2_X1 U590 ( .A1(n524), .A2(n530), .ZN(n525) );
  XNOR2_X1 U591 ( .A(G85GAT), .B(n525), .ZN(G1336GAT) );
  XOR2_X1 U592 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n528) );
  NAND2_X1 U593 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U594 ( .A(n528), .B(n527), .ZN(n529) );
  XNOR2_X1 U595 ( .A(G92GAT), .B(n529), .ZN(G1337GAT) );
  NAND2_X1 U596 ( .A1(n530), .A2(n533), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n531), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  NOR2_X1 U599 ( .A1(n546), .A2(n534), .ZN(n543) );
  NAND2_X1 U600 ( .A1(n576), .A2(n543), .ZN(n535) );
  XNOR2_X1 U601 ( .A(n535), .B(KEYINPUT114), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G113GAT), .B(n536), .ZN(G1340GAT) );
  XOR2_X1 U603 ( .A(G120GAT), .B(KEYINPUT49), .Z(n538) );
  NAND2_X1 U604 ( .A1(n543), .A2(n564), .ZN(n537) );
  XNOR2_X1 U605 ( .A(n538), .B(n537), .ZN(G1341GAT) );
  XOR2_X1 U606 ( .A(KEYINPUT50), .B(KEYINPUT115), .Z(n540) );
  NAND2_X1 U607 ( .A1(n543), .A2(n585), .ZN(n539) );
  XNOR2_X1 U608 ( .A(n540), .B(n539), .ZN(n541) );
  XNOR2_X1 U609 ( .A(G127GAT), .B(n541), .ZN(G1342GAT) );
  XOR2_X1 U610 ( .A(G134GAT), .B(KEYINPUT51), .Z(n545) );
  NAND2_X1 U611 ( .A1(n543), .A2(n542), .ZN(n544) );
  XNOR2_X1 U612 ( .A(n545), .B(n544), .ZN(G1343GAT) );
  NOR2_X1 U613 ( .A1(n547), .A2(n546), .ZN(n548) );
  NAND2_X1 U614 ( .A1(n548), .A2(n574), .ZN(n560) );
  NOR2_X1 U615 ( .A1(n549), .A2(n560), .ZN(n551) );
  XNOR2_X1 U616 ( .A(KEYINPUT116), .B(KEYINPUT117), .ZN(n550) );
  XNOR2_X1 U617 ( .A(n551), .B(n550), .ZN(n552) );
  XNOR2_X1 U618 ( .A(G141GAT), .B(n552), .ZN(G1344GAT) );
  XOR2_X1 U619 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n554) );
  XNOR2_X1 U620 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n553) );
  XNOR2_X1 U621 ( .A(n554), .B(n553), .ZN(n556) );
  NOR2_X1 U622 ( .A1(n456), .A2(n560), .ZN(n555) );
  XOR2_X1 U623 ( .A(n556), .B(n555), .Z(G1345GAT) );
  NOR2_X1 U624 ( .A1(n557), .A2(n560), .ZN(n559) );
  XNOR2_X1 U625 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n558) );
  XNOR2_X1 U626 ( .A(n559), .B(n558), .ZN(G1346GAT) );
  NOR2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n562) );
  XOR2_X1 U628 ( .A(G162GAT), .B(n562), .Z(G1347GAT) );
  NAND2_X1 U629 ( .A1(n576), .A2(n569), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n563), .B(G169GAT), .ZN(G1348GAT) );
  NAND2_X1 U631 ( .A1(n569), .A2(n564), .ZN(n566) );
  XOR2_X1 U632 ( .A(KEYINPUT123), .B(KEYINPUT57), .Z(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n568) );
  XOR2_X1 U634 ( .A(G176GAT), .B(KEYINPUT56), .Z(n567) );
  XNOR2_X1 U635 ( .A(n568), .B(n567), .ZN(G1349GAT) );
  NAND2_X1 U636 ( .A1(n585), .A2(n569), .ZN(n570) );
  XNOR2_X1 U637 ( .A(n570), .B(G183GAT), .ZN(G1350GAT) );
  XOR2_X1 U638 ( .A(G197GAT), .B(KEYINPUT125), .Z(n578) );
  AND2_X1 U639 ( .A1(n572), .A2(n571), .ZN(n573) );
  NAND2_X1 U640 ( .A1(n574), .A2(n573), .ZN(n575) );
  XOR2_X1 U641 ( .A(KEYINPUT124), .B(n575), .Z(n588) );
  NAND2_X1 U642 ( .A1(n588), .A2(n576), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n580) );
  XOR2_X1 U644 ( .A(KEYINPUT59), .B(KEYINPUT60), .Z(n579) );
  XNOR2_X1 U645 ( .A(n580), .B(n579), .ZN(G1352GAT) );
  XOR2_X1 U646 ( .A(KEYINPUT61), .B(KEYINPUT126), .Z(n583) );
  NAND2_X1 U647 ( .A1(n588), .A2(n581), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(G204GAT), .B(n584), .ZN(G1353GAT) );
  NAND2_X1 U650 ( .A1(n588), .A2(n585), .ZN(n586) );
  XNOR2_X1 U651 ( .A(n586), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U652 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n590) );
  NAND2_X1 U653 ( .A1(n588), .A2(n587), .ZN(n589) );
  XNOR2_X1 U654 ( .A(n590), .B(n589), .ZN(n591) );
  XNOR2_X1 U655 ( .A(G218GAT), .B(n591), .ZN(G1355GAT) );
endmodule

