//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 1 0 0 0 0 1 0 1 1 0 0 1 0 0 0 0 1 1 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 0 1 1 0 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n447, new_n451, new_n452, new_n453, new_n454, new_n457,
    new_n458, new_n459, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n534,
    new_n535, new_n536, new_n537, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n548, new_n550, new_n551, new_n552,
    new_n554, new_n555, new_n556, new_n557, new_n558, new_n559, new_n560,
    new_n561, new_n562, new_n563, new_n564, new_n567, new_n568, new_n569,
    new_n570, new_n572, new_n573, new_n574, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n603, new_n604, new_n607, new_n609, new_n610, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n656, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n826, new_n827, new_n828, new_n829, new_n830, new_n831,
    new_n832, new_n833, new_n834, new_n835, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1111, new_n1112,
    new_n1113, new_n1114;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  XOR2_X1   g006(.A(KEYINPUT65), .B(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XOR2_X1   g015(.A(KEYINPUT66), .B(G57), .Z(G237));
  XNOR2_X1  g016(.A(KEYINPUT67), .B(G108), .ZN(G238));
  NAND4_X1  g017(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g018(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g019(.A(G452), .Z(G391));
  AND2_X1   g020(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XOR2_X1   g022(.A(new_n447), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g023(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g024(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g025(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n451));
  XOR2_X1   g026(.A(new_n451), .B(KEYINPUT2), .Z(new_n452));
  NOR4_X1   g027(.A1(G237), .A2(G238), .A3(G235), .A4(G236), .ZN(new_n453));
  NAND2_X1  g028(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g029(.A(new_n454), .ZN(G325));
  XOR2_X1   g030(.A(new_n454), .B(KEYINPUT68), .Z(G261));
  INV_X1    g031(.A(G567), .ZN(new_n457));
  NOR2_X1   g032(.A1(new_n453), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n452), .ZN(new_n459));
  AOI21_X1  g034(.A(new_n458), .B1(new_n459), .B2(G2106), .ZN(G319));
  NAND2_X1  g035(.A1(G113), .A2(G2104), .ZN(new_n461));
  INV_X1    g036(.A(KEYINPUT3), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(G125), .ZN(new_n467));
  OAI21_X1  g042(.A(new_n461), .B1(new_n466), .B2(new_n467), .ZN(new_n468));
  NOR2_X1   g043(.A1(new_n464), .A2(G2105), .ZN(new_n469));
  AOI22_X1  g044(.A1(new_n468), .A2(G2105), .B1(G101), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  OAI21_X1  g046(.A(new_n471), .B1(new_n462), .B2(G2104), .ZN(new_n472));
  NAND2_X1  g047(.A1(new_n472), .A2(new_n463), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  NAND3_X1  g049(.A1(new_n471), .A2(new_n462), .A3(G2104), .ZN(new_n475));
  NAND4_X1  g050(.A1(new_n473), .A2(G137), .A3(new_n474), .A4(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n470), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n480));
  AOI21_X1  g055(.A(KEYINPUT69), .B1(new_n464), .B2(KEYINPUT3), .ZN(new_n481));
  NOR2_X1   g056(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n474), .B(new_n475), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  INV_X1    g058(.A(G136), .ZN(new_n484));
  OAI21_X1  g059(.A(new_n480), .B1(new_n483), .B2(new_n484), .ZN(new_n485));
  OAI211_X1 g060(.A(G2105), .B(new_n475), .C1(new_n481), .C2(new_n482), .ZN(new_n486));
  INV_X1    g061(.A(new_n486), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n485), .B1(G124), .B2(new_n487), .ZN(G162));
  INV_X1    g063(.A(G138), .ZN(new_n489));
  OAI21_X1  g064(.A(KEYINPUT4), .B1(new_n483), .B2(new_n489), .ZN(new_n490));
  INV_X1    g065(.A(KEYINPUT4), .ZN(new_n491));
  NOR2_X1   g066(.A1(new_n489), .A2(G2105), .ZN(new_n492));
  AND4_X1   g067(.A1(new_n491), .A2(new_n492), .A3(new_n463), .A4(new_n465), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(new_n494));
  NAND2_X1  g069(.A1(new_n490), .A2(new_n494), .ZN(new_n495));
  INV_X1    g070(.A(G126), .ZN(new_n496));
  OAI21_X1  g071(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n474), .A2(G114), .ZN(new_n498));
  OAI22_X1  g073(.A1(new_n486), .A2(new_n496), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(new_n499), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n495), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(new_n501), .ZN(G164));
  INV_X1    g077(.A(KEYINPUT70), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n503), .A2(KEYINPUT6), .A3(G651), .ZN(new_n504));
  AOI21_X1  g079(.A(KEYINPUT6), .B1(new_n503), .B2(G651), .ZN(new_n505));
  NOR2_X1   g080(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g081(.A(G543), .ZN(new_n507));
  NOR2_X1   g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n508), .A2(G50), .ZN(new_n509));
  INV_X1    g084(.A(G88), .ZN(new_n510));
  INV_X1    g085(.A(new_n506), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n507), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n513), .A2(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(new_n515), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n509), .B1(new_n510), .B2(new_n517), .ZN(new_n518));
  AOI22_X1  g093(.A1(new_n516), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n519));
  INV_X1    g094(.A(G651), .ZN(new_n520));
  NOR2_X1   g095(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OR2_X1    g096(.A1(new_n518), .A2(new_n521), .ZN(G303));
  INV_X1    g097(.A(G303), .ZN(G166));
  XNOR2_X1  g098(.A(KEYINPUT71), .B(KEYINPUT7), .ZN(new_n524));
  XNOR2_X1  g099(.A(new_n524), .B(KEYINPUT72), .ZN(new_n525));
  NAND3_X1  g100(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n526));
  XNOR2_X1  g101(.A(new_n525), .B(new_n526), .ZN(new_n527));
  NOR2_X1   g102(.A1(new_n506), .A2(new_n515), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n528), .A2(G89), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n508), .A2(G51), .ZN(new_n530));
  NAND3_X1  g105(.A1(new_n516), .A2(G63), .A3(G651), .ZN(new_n531));
  NAND3_X1  g106(.A1(new_n529), .A2(new_n530), .A3(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n527), .A2(new_n532), .ZN(G168));
  AOI22_X1  g108(.A1(new_n516), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n534));
  INV_X1    g109(.A(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n535), .A2(G651), .B1(G52), .B2(new_n508), .ZN(new_n536));
  NAND2_X1  g111(.A1(new_n528), .A2(G90), .ZN(new_n537));
  NAND2_X1  g112(.A1(new_n536), .A2(new_n537), .ZN(G301));
  INV_X1    g113(.A(G301), .ZN(G171));
  NAND2_X1  g114(.A1(G68), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G56), .ZN(new_n541));
  OAI21_X1  g116(.A(new_n540), .B1(new_n515), .B2(new_n541), .ZN(new_n542));
  AOI22_X1  g117(.A1(new_n508), .A2(G43), .B1(G651), .B2(new_n542), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n528), .A2(G81), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(new_n545), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n546), .A2(G860), .ZN(G153));
  AND3_X1   g122(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G36), .ZN(G176));
  NAND2_X1  g124(.A1(G1), .A2(G3), .ZN(new_n550));
  XNOR2_X1  g125(.A(new_n550), .B(KEYINPUT8), .ZN(new_n551));
  NAND2_X1  g126(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT73), .ZN(G188));
  AND3_X1   g128(.A1(new_n508), .A2(KEYINPUT9), .A3(G53), .ZN(new_n554));
  AOI21_X1  g129(.A(KEYINPUT9), .B1(new_n508), .B2(G53), .ZN(new_n555));
  NOR2_X1   g130(.A1(new_n554), .A2(new_n555), .ZN(new_n556));
  NAND2_X1  g131(.A1(G78), .A2(G543), .ZN(new_n557));
  XNOR2_X1  g132(.A(new_n515), .B(KEYINPUT74), .ZN(new_n558));
  XNOR2_X1  g133(.A(KEYINPUT75), .B(G65), .ZN(new_n559));
  OAI21_X1  g134(.A(new_n557), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n560), .A2(G651), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n528), .A2(G91), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n556), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT76), .ZN(new_n564));
  INV_X1    g139(.A(new_n564), .ZN(G299));
  INV_X1    g140(.A(G168), .ZN(G286));
  NAND2_X1  g141(.A1(new_n508), .A2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n528), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n516), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n570));
  XNOR2_X1  g145(.A(new_n570), .B(KEYINPUT77), .ZN(G288));
  INV_X1    g146(.A(KEYINPUT78), .ZN(new_n572));
  INV_X1    g147(.A(G86), .ZN(new_n573));
  OAI21_X1  g148(.A(new_n572), .B1(new_n517), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n528), .A2(KEYINPUT78), .A3(G86), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g151(.A1(G73), .A2(G543), .ZN(new_n577));
  INV_X1    g152(.A(G61), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n515), .B2(new_n578), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n508), .A2(G48), .B1(G651), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g155(.A1(new_n576), .A2(new_n580), .ZN(G305));
  AOI22_X1  g156(.A1(new_n516), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n582));
  NOR2_X1   g157(.A1(new_n582), .A2(new_n520), .ZN(new_n583));
  XNOR2_X1  g158(.A(new_n583), .B(KEYINPUT79), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n508), .A2(G47), .ZN(new_n585));
  INV_X1    g160(.A(G85), .ZN(new_n586));
  OAI21_X1  g161(.A(new_n585), .B1(new_n586), .B2(new_n517), .ZN(new_n587));
  AND2_X1   g162(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n588));
  NOR2_X1   g163(.A1(new_n587), .A2(KEYINPUT80), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n584), .B1(new_n588), .B2(new_n589), .ZN(G290));
  NAND2_X1  g165(.A1(G301), .A2(G868), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n528), .A2(G92), .ZN(new_n592));
  XOR2_X1   g167(.A(new_n592), .B(KEYINPUT10), .Z(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n558), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n508), .A2(G54), .ZN(new_n598));
  NAND3_X1  g173(.A1(new_n593), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  INV_X1    g174(.A(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G284));
  OAI21_X1  g176(.A(new_n591), .B1(new_n600), .B2(G868), .ZN(G321));
  NAND2_X1  g177(.A1(G286), .A2(G868), .ZN(new_n603));
  XOR2_X1   g178(.A(new_n564), .B(KEYINPUT81), .Z(new_n604));
  OAI21_X1  g179(.A(new_n603), .B1(new_n604), .B2(G868), .ZN(G297));
  XNOR2_X1  g180(.A(G297), .B(KEYINPUT82), .ZN(G280));
  XOR2_X1   g181(.A(KEYINPUT83), .B(G559), .Z(new_n607));
  OAI21_X1  g182(.A(new_n600), .B1(G860), .B2(new_n607), .ZN(G148));
  NAND2_X1  g183(.A1(new_n600), .A2(new_n607), .ZN(new_n609));
  NAND2_X1  g184(.A1(new_n609), .A2(G868), .ZN(new_n610));
  OAI21_X1  g185(.A(new_n610), .B1(G868), .B2(new_n546), .ZN(G323));
  XNOR2_X1  g186(.A(G323), .B(KEYINPUT11), .ZN(G282));
  OR2_X1    g187(.A1(G99), .A2(G2105), .ZN(new_n613));
  OAI211_X1 g188(.A(new_n613), .B(G2104), .C1(G111), .C2(new_n474), .ZN(new_n614));
  INV_X1    g189(.A(G135), .ZN(new_n615));
  OAI21_X1  g190(.A(new_n614), .B1(new_n483), .B2(new_n615), .ZN(new_n616));
  AOI21_X1  g191(.A(new_n616), .B1(G123), .B2(new_n487), .ZN(new_n617));
  XNOR2_X1  g192(.A(new_n617), .B(G2096), .ZN(new_n618));
  INV_X1    g193(.A(new_n466), .ZN(new_n619));
  NAND2_X1  g194(.A1(new_n619), .A2(new_n469), .ZN(new_n620));
  XOR2_X1   g195(.A(KEYINPUT84), .B(KEYINPUT12), .Z(new_n621));
  XNOR2_X1  g196(.A(new_n620), .B(new_n621), .ZN(new_n622));
  XNOR2_X1  g197(.A(KEYINPUT13), .B(G2100), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n622), .B(new_n623), .ZN(new_n624));
  NAND2_X1  g199(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  XOR2_X1   g200(.A(new_n625), .B(KEYINPUT85), .Z(G156));
  XOR2_X1   g201(.A(KEYINPUT88), .B(G2438), .Z(new_n627));
  XNOR2_X1  g202(.A(G2427), .B(G2430), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n627), .B(new_n628), .ZN(new_n629));
  XOR2_X1   g204(.A(KEYINPUT15), .B(G2435), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n629), .B(new_n630), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(KEYINPUT14), .ZN(new_n632));
  XNOR2_X1  g207(.A(G2443), .B(G2446), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n632), .B(new_n633), .ZN(new_n634));
  XNOR2_X1  g209(.A(G2451), .B(G2454), .ZN(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT87), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT86), .B(KEYINPUT16), .ZN(new_n637));
  XNOR2_X1  g212(.A(new_n636), .B(new_n637), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n634), .B(new_n638), .ZN(new_n639));
  XNOR2_X1  g214(.A(G1341), .B(G1348), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n641), .A2(G14), .ZN(new_n642));
  INV_X1    g217(.A(new_n642), .ZN(G401));
  XOR2_X1   g218(.A(G2072), .B(G2078), .Z(new_n644));
  XOR2_X1   g219(.A(G2067), .B(G2678), .Z(new_n645));
  INV_X1    g220(.A(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2084), .B(G2090), .Z(new_n647));
  NAND2_X1  g222(.A1(new_n646), .A2(new_n647), .ZN(new_n648));
  AOI21_X1  g223(.A(new_n644), .B1(new_n648), .B2(KEYINPUT18), .ZN(new_n649));
  XNOR2_X1  g224(.A(new_n649), .B(G2096), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(G2100), .ZN(new_n651));
  AND2_X1   g226(.A1(new_n648), .A2(KEYINPUT17), .ZN(new_n652));
  OR2_X1    g227(.A1(new_n646), .A2(new_n647), .ZN(new_n653));
  AOI21_X1  g228(.A(KEYINPUT18), .B1(new_n652), .B2(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(new_n651), .B(new_n654), .Z(G227));
  XNOR2_X1  g230(.A(G1971), .B(G1976), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT19), .ZN(new_n657));
  XOR2_X1   g232(.A(G1956), .B(G2474), .Z(new_n658));
  XOR2_X1   g233(.A(G1961), .B(G1966), .Z(new_n659));
  NAND2_X1  g234(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n660), .ZN(new_n661));
  NOR2_X1   g236(.A1(new_n658), .A2(new_n659), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI22_X1  g238(.A1(new_n661), .A2(KEYINPUT20), .B1(new_n657), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(KEYINPUT20), .B2(new_n661), .ZN(new_n665));
  NAND3_X1  g240(.A1(new_n663), .A2(new_n657), .A3(new_n660), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g242(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n668));
  INV_X1    g243(.A(G1981), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n668), .B(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(G1991), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(G1996), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n667), .B(new_n672), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT89), .B(G1986), .ZN(new_n674));
  XOR2_X1   g249(.A(new_n673), .B(new_n674), .Z(G229));
  INV_X1    g250(.A(G16), .ZN(new_n676));
  NAND2_X1  g251(.A1(new_n676), .A2(G22), .ZN(new_n677));
  OAI21_X1  g252(.A(new_n677), .B1(G166), .B2(new_n676), .ZN(new_n678));
  INV_X1    g253(.A(G1971), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND2_X1   g255(.A1(new_n676), .A2(G6), .ZN(new_n681));
  AOI21_X1  g256(.A(new_n681), .B1(G305), .B2(G16), .ZN(new_n682));
  XNOR2_X1  g257(.A(KEYINPUT32), .B(G1981), .ZN(new_n683));
  XNOR2_X1  g258(.A(new_n682), .B(new_n683), .ZN(new_n684));
  INV_X1    g259(.A(G1976), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n676), .A2(G23), .ZN(new_n686));
  INV_X1    g261(.A(new_n570), .ZN(new_n687));
  OAI21_X1  g262(.A(new_n686), .B1(new_n687), .B2(new_n676), .ZN(new_n688));
  AND2_X1   g263(.A1(new_n688), .A2(KEYINPUT33), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n688), .A2(KEYINPUT33), .ZN(new_n690));
  OAI21_X1  g265(.A(new_n685), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OR3_X1    g266(.A1(new_n689), .A2(new_n690), .A3(new_n685), .ZN(new_n692));
  NAND4_X1  g267(.A1(new_n680), .A2(new_n684), .A3(new_n691), .A4(new_n692), .ZN(new_n693));
  OR2_X1    g268(.A1(new_n693), .A2(KEYINPUT34), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G24), .ZN(new_n695));
  XNOR2_X1  g270(.A(G290), .B(KEYINPUT90), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT91), .B(G1986), .Z(new_n698));
  INV_X1    g273(.A(new_n698), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n697), .B(new_n699), .ZN(new_n700));
  AOI21_X1  g275(.A(KEYINPUT92), .B1(new_n693), .B2(KEYINPUT34), .ZN(new_n701));
  INV_X1    g276(.A(G29), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n702), .A2(G25), .ZN(new_n703));
  OR2_X1    g278(.A1(G95), .A2(G2105), .ZN(new_n704));
  OAI211_X1 g279(.A(new_n704), .B(G2104), .C1(G107), .C2(new_n474), .ZN(new_n705));
  INV_X1    g280(.A(G131), .ZN(new_n706));
  OAI21_X1  g281(.A(new_n705), .B1(new_n483), .B2(new_n706), .ZN(new_n707));
  AOI21_X1  g282(.A(new_n707), .B1(G119), .B2(new_n487), .ZN(new_n708));
  OAI21_X1  g283(.A(new_n703), .B1(new_n708), .B2(new_n702), .ZN(new_n709));
  XNOR2_X1  g284(.A(KEYINPUT35), .B(G1991), .ZN(new_n710));
  INV_X1    g285(.A(new_n710), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n709), .B(new_n711), .ZN(new_n712));
  NAND4_X1  g287(.A1(new_n694), .A2(new_n700), .A3(new_n701), .A4(new_n712), .ZN(new_n713));
  XNOR2_X1  g288(.A(new_n713), .B(KEYINPUT36), .ZN(new_n714));
  XNOR2_X1  g289(.A(KEYINPUT31), .B(G11), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n676), .A2(KEYINPUT23), .A3(G20), .ZN(new_n716));
  INV_X1    g291(.A(KEYINPUT23), .ZN(new_n717));
  INV_X1    g292(.A(G20), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n717), .B1(new_n718), .B2(G16), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n716), .B(new_n719), .C1(new_n564), .C2(new_n676), .ZN(new_n720));
  XNOR2_X1  g295(.A(KEYINPUT97), .B(G1956), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  NAND2_X1  g297(.A1(new_n487), .A2(G129), .ZN(new_n723));
  NAND4_X1  g298(.A1(new_n473), .A2(G141), .A3(new_n474), .A4(new_n475), .ZN(new_n724));
  NAND2_X1  g299(.A1(new_n469), .A2(G105), .ZN(new_n725));
  NAND3_X1  g300(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n726));
  XOR2_X1   g301(.A(new_n726), .B(KEYINPUT26), .Z(new_n727));
  NAND4_X1  g302(.A1(new_n723), .A2(new_n724), .A3(new_n725), .A4(new_n727), .ZN(new_n728));
  OR2_X1    g303(.A1(new_n728), .A2(new_n702), .ZN(new_n729));
  NOR2_X1   g304(.A1(G29), .A2(G32), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(KEYINPUT95), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g306(.A(new_n731), .B1(KEYINPUT95), .B2(new_n729), .ZN(new_n732));
  XOR2_X1   g307(.A(KEYINPUT27), .B(G1996), .Z(new_n733));
  XNOR2_X1  g308(.A(new_n732), .B(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(new_n734), .ZN(new_n735));
  NOR2_X1   g310(.A1(new_n722), .A2(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n702), .A2(G27), .ZN(new_n737));
  OAI21_X1  g312(.A(new_n737), .B1(G164), .B2(new_n702), .ZN(new_n738));
  INV_X1    g313(.A(G2078), .ZN(new_n739));
  XNOR2_X1  g314(.A(new_n738), .B(new_n739), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n702), .A2(G35), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G162), .B2(new_n702), .ZN(new_n742));
  XOR2_X1   g317(.A(new_n742), .B(KEYINPUT29), .Z(new_n743));
  INV_X1    g318(.A(G2090), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NOR2_X1   g320(.A1(G16), .A2(G21), .ZN(new_n746));
  AOI21_X1  g321(.A(new_n746), .B1(G168), .B2(G16), .ZN(new_n747));
  NOR2_X1   g322(.A1(new_n747), .A2(G1966), .ZN(new_n748));
  INV_X1    g323(.A(KEYINPUT30), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n749), .A2(G28), .ZN(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(KEYINPUT96), .ZN(new_n751));
  OAI211_X1 g326(.A(new_n751), .B(new_n702), .C1(new_n749), .C2(G28), .ZN(new_n752));
  INV_X1    g327(.A(new_n747), .ZN(new_n753));
  INV_X1    g328(.A(G1966), .ZN(new_n754));
  OAI21_X1  g329(.A(new_n752), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g330(.A(G2072), .ZN(new_n756));
  OR2_X1    g331(.A1(G29), .A2(G33), .ZN(new_n757));
  AOI22_X1  g332(.A1(new_n619), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n474), .ZN(new_n759));
  INV_X1    g334(.A(G139), .ZN(new_n760));
  NOR2_X1   g335(.A1(new_n483), .A2(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n469), .A2(G103), .ZN(new_n762));
  XNOR2_X1  g337(.A(new_n762), .B(KEYINPUT25), .ZN(new_n763));
  OR3_X1    g338(.A1(new_n759), .A2(new_n761), .A3(new_n763), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n757), .B1(new_n764), .B2(new_n702), .ZN(new_n765));
  AOI211_X1 g340(.A(new_n748), .B(new_n755), .C1(new_n756), .C2(new_n765), .ZN(new_n766));
  NAND4_X1  g341(.A1(new_n736), .A2(new_n740), .A3(new_n745), .A4(new_n766), .ZN(new_n767));
  NAND2_X1  g342(.A1(G171), .A2(G16), .ZN(new_n768));
  OAI21_X1  g343(.A(new_n768), .B1(G5), .B2(G16), .ZN(new_n769));
  INV_X1    g344(.A(G1961), .ZN(new_n770));
  AND2_X1   g345(.A1(new_n676), .A2(G19), .ZN(new_n771));
  AOI21_X1  g346(.A(new_n771), .B1(new_n545), .B2(G16), .ZN(new_n772));
  INV_X1    g347(.A(new_n772), .ZN(new_n773));
  AOI22_X1  g348(.A1(new_n769), .A2(new_n770), .B1(new_n773), .B2(G1341), .ZN(new_n774));
  OAI21_X1  g349(.A(new_n774), .B1(G1341), .B2(new_n773), .ZN(new_n775));
  NAND2_X1  g350(.A1(KEYINPUT24), .A2(G34), .ZN(new_n776));
  INV_X1    g351(.A(new_n776), .ZN(new_n777));
  NOR2_X1   g352(.A1(KEYINPUT24), .A2(G34), .ZN(new_n778));
  NOR3_X1   g353(.A1(new_n777), .A2(new_n778), .A3(G29), .ZN(new_n779));
  AOI21_X1  g354(.A(new_n779), .B1(new_n477), .B2(G29), .ZN(new_n780));
  INV_X1    g355(.A(G2084), .ZN(new_n781));
  NAND2_X1  g356(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  INV_X1    g357(.A(G2067), .ZN(new_n783));
  XNOR2_X1  g358(.A(KEYINPUT94), .B(KEYINPUT28), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n702), .A2(G26), .ZN(new_n785));
  XNOR2_X1  g360(.A(new_n784), .B(new_n785), .ZN(new_n786));
  OR2_X1    g361(.A1(G104), .A2(G2105), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n787), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n788));
  INV_X1    g363(.A(G140), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n483), .B2(new_n789), .ZN(new_n790));
  AOI21_X1  g365(.A(new_n790), .B1(G128), .B2(new_n487), .ZN(new_n791));
  INV_X1    g366(.A(new_n791), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n786), .B1(new_n792), .B2(G29), .ZN(new_n793));
  OAI221_X1 g368(.A(new_n782), .B1(new_n783), .B2(new_n793), .C1(new_n769), .C2(new_n770), .ZN(new_n794));
  NOR2_X1   g369(.A1(new_n775), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g370(.A(new_n795), .B1(new_n781), .B2(new_n780), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n793), .A2(new_n783), .ZN(new_n797));
  OAI21_X1  g372(.A(new_n797), .B1(new_n765), .B2(new_n756), .ZN(new_n798));
  NOR2_X1   g373(.A1(new_n743), .A2(new_n744), .ZN(new_n799));
  NOR4_X1   g374(.A1(new_n767), .A2(new_n796), .A3(new_n798), .A4(new_n799), .ZN(new_n800));
  AND3_X1   g375(.A1(new_n714), .A2(new_n715), .A3(new_n800), .ZN(new_n801));
  NAND2_X1  g376(.A1(new_n600), .A2(G16), .ZN(new_n802));
  OAI21_X1  g377(.A(new_n802), .B1(G4), .B2(G16), .ZN(new_n803));
  XNOR2_X1  g378(.A(KEYINPUT93), .B(G1348), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n803), .B(new_n804), .ZN(new_n805));
  INV_X1    g380(.A(new_n805), .ZN(new_n806));
  NAND2_X1  g381(.A1(new_n617), .A2(G29), .ZN(new_n807));
  NAND4_X1  g382(.A1(new_n801), .A2(KEYINPUT98), .A3(new_n806), .A4(new_n807), .ZN(new_n808));
  INV_X1    g383(.A(KEYINPUT98), .ZN(new_n809));
  NAND4_X1  g384(.A1(new_n714), .A2(new_n800), .A3(new_n807), .A4(new_n715), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n809), .B1(new_n810), .B2(new_n805), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n808), .A2(new_n811), .ZN(G311));
  NAND3_X1  g387(.A1(new_n801), .A2(new_n806), .A3(new_n807), .ZN(G150));
  NAND2_X1  g388(.A1(new_n528), .A2(G93), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n508), .A2(G55), .ZN(new_n815));
  AOI22_X1  g390(.A1(new_n516), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n816));
  OAI211_X1 g391(.A(new_n814), .B(new_n815), .C1(new_n520), .C2(new_n816), .ZN(new_n817));
  NAND2_X1  g392(.A1(new_n817), .A2(G860), .ZN(new_n818));
  XOR2_X1   g393(.A(new_n818), .B(KEYINPUT37), .Z(new_n819));
  NAND2_X1  g394(.A1(new_n600), .A2(G559), .ZN(new_n820));
  XNOR2_X1  g395(.A(new_n820), .B(KEYINPUT38), .ZN(new_n821));
  XOR2_X1   g396(.A(new_n817), .B(new_n545), .Z(new_n822));
  XNOR2_X1  g397(.A(new_n822), .B(KEYINPUT39), .ZN(new_n823));
  XNOR2_X1  g398(.A(new_n821), .B(new_n823), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n819), .B1(new_n824), .B2(G860), .ZN(G145));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n501), .B(new_n728), .ZN(new_n827));
  OR2_X1    g402(.A1(new_n827), .A2(new_n791), .ZN(new_n828));
  NAND2_X1  g403(.A1(new_n827), .A2(new_n791), .ZN(new_n829));
  NAND3_X1  g404(.A1(new_n828), .A2(new_n764), .A3(new_n829), .ZN(new_n830));
  XOR2_X1   g405(.A(new_n830), .B(KEYINPUT100), .Z(new_n831));
  XOR2_X1   g406(.A(new_n708), .B(new_n622), .Z(new_n832));
  INV_X1    g407(.A(G142), .ZN(new_n833));
  OAI21_X1  g408(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n834));
  NOR2_X1   g409(.A1(new_n474), .A2(G118), .ZN(new_n835));
  OAI22_X1  g410(.A1(new_n483), .A2(new_n833), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  AOI21_X1  g411(.A(new_n836), .B1(G130), .B2(new_n487), .ZN(new_n837));
  XNOR2_X1  g412(.A(new_n832), .B(new_n837), .ZN(new_n838));
  AOI21_X1  g413(.A(new_n764), .B1(new_n828), .B2(new_n829), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n839), .B(KEYINPUT99), .ZN(new_n840));
  AND3_X1   g415(.A1(new_n831), .A2(new_n838), .A3(new_n840), .ZN(new_n841));
  AOI21_X1  g416(.A(new_n838), .B1(new_n831), .B2(new_n840), .ZN(new_n842));
  OAI21_X1  g417(.A(new_n826), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  XNOR2_X1  g418(.A(G160), .B(new_n617), .ZN(new_n844));
  XOR2_X1   g419(.A(new_n844), .B(G162), .Z(new_n845));
  INV_X1    g420(.A(new_n845), .ZN(new_n846));
  OAI211_X1 g421(.A(new_n843), .B(new_n846), .C1(new_n826), .C2(new_n842), .ZN(new_n847));
  INV_X1    g422(.A(G37), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n845), .B1(new_n841), .B2(new_n842), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n847), .A2(new_n848), .A3(new_n849), .ZN(new_n850));
  XNOR2_X1  g425(.A(new_n850), .B(KEYINPUT40), .ZN(G395));
  NOR2_X1   g426(.A1(new_n817), .A2(G868), .ZN(new_n852));
  XNOR2_X1  g427(.A(new_n609), .B(new_n822), .ZN(new_n853));
  INV_X1    g428(.A(new_n853), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n564), .A2(new_n599), .ZN(new_n855));
  INV_X1    g430(.A(new_n855), .ZN(new_n856));
  NOR2_X1   g431(.A1(new_n564), .A2(new_n599), .ZN(new_n857));
  OAI21_X1  g432(.A(KEYINPUT102), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  NOR2_X1   g433(.A1(new_n857), .A2(KEYINPUT102), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n854), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(KEYINPUT102), .ZN(new_n862));
  NAND2_X1  g437(.A1(G299), .A2(new_n600), .ZN(new_n863));
  AOI21_X1  g438(.A(new_n862), .B1(new_n863), .B2(new_n855), .ZN(new_n864));
  OAI21_X1  g439(.A(KEYINPUT41), .B1(new_n864), .B2(new_n859), .ZN(new_n865));
  INV_X1    g440(.A(KEYINPUT41), .ZN(new_n866));
  NAND3_X1  g441(.A1(new_n863), .A2(new_n866), .A3(new_n855), .ZN(new_n867));
  AND2_X1   g442(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  XNOR2_X1  g443(.A(G303), .B(G305), .ZN(new_n869));
  XNOR2_X1  g444(.A(new_n869), .B(KEYINPUT103), .ZN(new_n870));
  XNOR2_X1  g445(.A(G290), .B(new_n687), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n870), .B(new_n871), .ZN(new_n872));
  XNOR2_X1  g447(.A(new_n872), .B(KEYINPUT42), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT104), .ZN(new_n874));
  OAI221_X1 g449(.A(new_n861), .B1(new_n854), .B2(new_n868), .C1(new_n873), .C2(new_n874), .ZN(new_n875));
  AND2_X1   g450(.A1(new_n873), .A2(new_n874), .ZN(new_n876));
  XNOR2_X1  g451(.A(new_n875), .B(new_n876), .ZN(new_n877));
  AOI21_X1  g452(.A(new_n852), .B1(new_n877), .B2(G868), .ZN(G295));
  AOI21_X1  g453(.A(new_n852), .B1(new_n877), .B2(G868), .ZN(G331));
  INV_X1    g454(.A(new_n872), .ZN(new_n880));
  XNOR2_X1  g455(.A(G168), .B(G301), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n822), .ZN(new_n882));
  INV_X1    g457(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n865), .B2(new_n867), .ZN(new_n884));
  NOR3_X1   g459(.A1(new_n864), .A2(new_n859), .A3(new_n882), .ZN(new_n885));
  OAI21_X1  g460(.A(new_n880), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  OAI211_X1 g461(.A(new_n858), .B(new_n860), .C1(new_n883), .C2(new_n866), .ZN(new_n887));
  OAI211_X1 g462(.A(new_n882), .B(KEYINPUT41), .C1(new_n857), .C2(new_n856), .ZN(new_n888));
  NAND3_X1  g463(.A1(new_n872), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n889), .A2(KEYINPUT105), .ZN(new_n890));
  INV_X1    g465(.A(KEYINPUT105), .ZN(new_n891));
  NAND4_X1  g466(.A1(new_n872), .A2(new_n887), .A3(new_n891), .A4(new_n888), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n886), .A2(new_n848), .A3(new_n890), .A4(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n893), .A2(KEYINPUT43), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT106), .ZN(new_n895));
  NAND2_X1  g470(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  OR3_X1    g471(.A1(new_n884), .A2(new_n880), .A3(new_n885), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT43), .ZN(new_n898));
  NAND4_X1  g473(.A1(new_n897), .A2(new_n898), .A3(new_n848), .A4(new_n886), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n893), .A2(KEYINPUT106), .A3(KEYINPUT43), .ZN(new_n900));
  NAND4_X1  g475(.A1(new_n896), .A2(KEYINPUT44), .A3(new_n899), .A4(new_n900), .ZN(new_n901));
  NAND2_X1  g476(.A1(new_n893), .A2(new_n898), .ZN(new_n902));
  NAND4_X1  g477(.A1(new_n897), .A2(KEYINPUT43), .A3(new_n848), .A4(new_n886), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  OAI21_X1  g479(.A(new_n901), .B1(KEYINPUT44), .B2(new_n904), .ZN(G397));
  INV_X1    g480(.A(G1384), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n473), .A2(G138), .A3(new_n474), .A4(new_n475), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n493), .B1(new_n907), .B2(KEYINPUT4), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n906), .B1(new_n908), .B2(new_n499), .ZN(new_n909));
  INV_X1    g484(.A(KEYINPUT45), .ZN(new_n910));
  NAND2_X1  g485(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n470), .A2(G40), .A3(new_n476), .ZN(new_n912));
  NOR2_X1   g487(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND3_X1   g488(.A1(new_n913), .A2(G1996), .A3(new_n728), .ZN(new_n914));
  OR3_X1    g489(.A1(new_n911), .A2(G1996), .A3(new_n912), .ZN(new_n915));
  NOR2_X1   g490(.A1(new_n915), .A2(new_n728), .ZN(new_n916));
  XOR2_X1   g491(.A(new_n916), .B(KEYINPUT107), .Z(new_n917));
  XNOR2_X1  g492(.A(new_n791), .B(new_n783), .ZN(new_n918));
  AOI211_X1 g493(.A(new_n914), .B(new_n917), .C1(new_n913), .C2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(new_n708), .B(new_n711), .ZN(new_n920));
  NAND2_X1  g495(.A1(new_n913), .A2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n919), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(G290), .B(G1986), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n913), .B2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n909), .A2(KEYINPUT50), .ZN(new_n925));
  INV_X1    g500(.A(new_n912), .ZN(new_n926));
  INV_X1    g501(.A(KEYINPUT50), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(new_n906), .C1(new_n908), .C2(new_n499), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n925), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n929), .A2(KEYINPUT117), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT117), .ZN(new_n931));
  NAND4_X1  g506(.A1(new_n925), .A2(new_n931), .A3(new_n926), .A4(new_n928), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g508(.A(G1348), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n909), .A2(new_n912), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n936), .A2(new_n783), .ZN(new_n937));
  NAND3_X1  g512(.A1(new_n935), .A2(KEYINPUT60), .A3(new_n937), .ZN(new_n938));
  INV_X1    g513(.A(KEYINPUT119), .ZN(new_n939));
  NAND2_X1  g514(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  NAND4_X1  g515(.A1(new_n935), .A2(KEYINPUT119), .A3(KEYINPUT60), .A4(new_n937), .ZN(new_n941));
  NAND3_X1  g516(.A1(new_n940), .A2(new_n600), .A3(new_n941), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n935), .A2(new_n937), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT60), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n938), .A2(new_n939), .A3(new_n599), .ZN(new_n946));
  NAND3_X1  g521(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  NAND3_X1  g522(.A1(new_n501), .A2(KEYINPUT45), .A3(new_n906), .ZN(new_n948));
  NAND3_X1  g523(.A1(new_n948), .A2(new_n911), .A3(new_n926), .ZN(new_n949));
  XNOR2_X1  g524(.A(KEYINPUT58), .B(G1341), .ZN(new_n950));
  OAI22_X1  g525(.A1(new_n949), .A2(G1996), .B1(new_n936), .B2(new_n950), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT118), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n952), .A2(KEYINPUT59), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n546), .A3(new_n953), .ZN(new_n954));
  OR2_X1    g529(.A1(new_n952), .A2(KEYINPUT59), .ZN(new_n955));
  XNOR2_X1  g530(.A(new_n954), .B(new_n955), .ZN(new_n956));
  INV_X1    g531(.A(KEYINPUT61), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT57), .ZN(new_n958));
  XNOR2_X1  g533(.A(new_n563), .B(new_n958), .ZN(new_n959));
  INV_X1    g534(.A(new_n949), .ZN(new_n960));
  XNOR2_X1  g535(.A(KEYINPUT56), .B(G2072), .ZN(new_n961));
  NAND2_X1  g536(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(G1956), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n929), .A2(new_n963), .ZN(new_n964));
  NAND3_X1  g539(.A1(new_n959), .A2(new_n962), .A3(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(new_n965), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n959), .B1(new_n962), .B2(new_n964), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n957), .B1(new_n966), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n962), .A2(new_n964), .ZN(new_n969));
  INV_X1    g544(.A(new_n959), .ZN(new_n970));
  NAND2_X1  g545(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n971), .A2(KEYINPUT61), .A3(new_n965), .ZN(new_n972));
  AND3_X1   g547(.A1(new_n956), .A2(new_n968), .A3(new_n972), .ZN(new_n973));
  NAND2_X1  g548(.A1(new_n947), .A2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n943), .A2(new_n600), .A3(new_n965), .ZN(new_n975));
  NAND3_X1  g550(.A1(new_n974), .A2(new_n975), .A3(new_n971), .ZN(new_n976));
  NAND2_X1  g551(.A1(new_n976), .A2(KEYINPUT120), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n933), .A2(new_n770), .ZN(new_n978));
  NAND3_X1  g553(.A1(new_n960), .A2(KEYINPUT53), .A3(new_n739), .ZN(new_n979));
  NAND2_X1  g554(.A1(new_n949), .A2(KEYINPUT108), .ZN(new_n980));
  INV_X1    g555(.A(KEYINPUT108), .ZN(new_n981));
  NAND4_X1  g556(.A1(new_n948), .A2(new_n911), .A3(new_n981), .A4(new_n926), .ZN(new_n982));
  NAND3_X1  g557(.A1(new_n980), .A2(new_n739), .A3(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT124), .ZN(new_n984));
  INV_X1    g559(.A(KEYINPUT53), .ZN(new_n985));
  AND3_X1   g560(.A1(new_n983), .A2(new_n984), .A3(new_n985), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n983), .B2(new_n985), .ZN(new_n987));
  OAI211_X1 g562(.A(new_n978), .B(new_n979), .C1(new_n986), .C2(new_n987), .ZN(new_n988));
  NOR2_X1   g563(.A1(new_n988), .A2(G171), .ZN(new_n989));
  INV_X1    g564(.A(new_n989), .ZN(new_n990));
  NAND2_X1  g565(.A1(new_n988), .A2(G171), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT125), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT54), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n990), .B(new_n991), .C1(new_n992), .C2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(new_n991), .ZN(new_n995));
  OAI211_X1 g570(.A(KEYINPUT125), .B(KEYINPUT54), .C1(new_n995), .C2(new_n989), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n994), .A2(new_n996), .ZN(new_n997));
  XNOR2_X1  g572(.A(KEYINPUT114), .B(G86), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n580), .B1(new_n517), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(G1981), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT113), .ZN(new_n1001));
  INV_X1    g576(.A(G305), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n1001), .B1(new_n1002), .B2(new_n669), .ZN(new_n1003));
  NOR3_X1   g578(.A1(G305), .A2(KEYINPUT113), .A3(G1981), .ZN(new_n1004));
  OAI21_X1  g579(.A(new_n1000), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  INV_X1    g580(.A(KEYINPUT49), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(G8), .ZN(new_n1008));
  NOR2_X1   g583(.A1(new_n936), .A2(new_n1008), .ZN(new_n1009));
  OAI211_X1 g584(.A(KEYINPUT49), .B(new_n1000), .C1(new_n1003), .C2(new_n1004), .ZN(new_n1010));
  NAND3_X1  g585(.A1(new_n1007), .A2(new_n1009), .A3(new_n1010), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n687), .A2(KEYINPUT112), .A3(G1976), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n1009), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g588(.A(KEYINPUT112), .B1(new_n687), .B2(G1976), .ZN(new_n1014));
  OAI21_X1  g589(.A(KEYINPUT52), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  NOR2_X1   g590(.A1(new_n1013), .A2(new_n1014), .ZN(new_n1016));
  AOI21_X1  g591(.A(KEYINPUT52), .B1(G288), .B2(new_n685), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AND3_X1   g593(.A1(new_n1011), .A2(new_n1015), .A3(new_n1018), .ZN(new_n1019));
  XNOR2_X1  g594(.A(KEYINPUT109), .B(G1971), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n1020), .B1(new_n980), .B2(new_n982), .ZN(new_n1021));
  INV_X1    g596(.A(new_n929), .ZN(new_n1022));
  XNOR2_X1  g597(.A(KEYINPUT110), .B(G2090), .ZN(new_n1023));
  NAND2_X1  g598(.A1(new_n1022), .A2(new_n1023), .ZN(new_n1024));
  INV_X1    g599(.A(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT111), .ZN(new_n1026));
  OR3_X1    g601(.A1(new_n1021), .A2(new_n1025), .A3(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(G303), .A2(G8), .ZN(new_n1028));
  XNOR2_X1  g603(.A(new_n1028), .B(KEYINPUT55), .ZN(new_n1029));
  INV_X1    g604(.A(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1026), .B1(new_n1021), .B2(new_n1025), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1027), .A2(G8), .A3(new_n1030), .A4(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT115), .ZN(new_n1033));
  OAI21_X1  g608(.A(new_n1023), .B1(new_n929), .B2(new_n1033), .ZN(new_n1034));
  AOI21_X1  g609(.A(new_n1034), .B1(new_n1033), .B2(new_n929), .ZN(new_n1035));
  OAI21_X1  g610(.A(G8), .B1(new_n1035), .B2(new_n1021), .ZN(new_n1036));
  NAND2_X1  g611(.A1(new_n1036), .A2(new_n1029), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n992), .A2(new_n993), .ZN(new_n1038));
  NAND4_X1  g613(.A1(new_n1019), .A2(new_n1032), .A3(new_n1037), .A4(new_n1038), .ZN(new_n1039));
  INV_X1    g614(.A(KEYINPUT123), .ZN(new_n1040));
  NOR2_X1   g615(.A1(G168), .A2(new_n1008), .ZN(new_n1041));
  INV_X1    g616(.A(new_n1041), .ZN(new_n1042));
  NAND4_X1  g617(.A1(new_n925), .A2(new_n781), .A3(new_n926), .A4(new_n928), .ZN(new_n1043));
  XNOR2_X1  g618(.A(new_n1043), .B(KEYINPUT116), .ZN(new_n1044));
  NAND2_X1  g619(.A1(new_n949), .A2(new_n754), .ZN(new_n1045));
  AOI21_X1  g620(.A(new_n1008), .B1(new_n1044), .B2(new_n1045), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT122), .ZN(new_n1047));
  OAI21_X1  g622(.A(new_n1042), .B1(new_n1046), .B2(new_n1047), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n925), .A2(new_n928), .ZN(new_n1049));
  NAND4_X1  g624(.A1(new_n1049), .A2(KEYINPUT116), .A3(new_n781), .A4(new_n926), .ZN(new_n1050));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n1051));
  NAND2_X1  g626(.A1(new_n1043), .A2(new_n1051), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1050), .A2(new_n1045), .A3(new_n1052), .ZN(new_n1053));
  NAND3_X1  g628(.A1(new_n1053), .A2(new_n1047), .A3(G8), .ZN(new_n1054));
  INV_X1    g629(.A(KEYINPUT51), .ZN(new_n1055));
  NAND2_X1  g630(.A1(new_n1054), .A2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n1040), .B1(new_n1048), .B2(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1053), .A2(G8), .ZN(new_n1058));
  AOI21_X1  g633(.A(new_n1041), .B1(new_n1058), .B2(KEYINPUT122), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1059), .A2(KEYINPUT123), .A3(new_n1055), .A4(new_n1054), .ZN(new_n1060));
  INV_X1    g635(.A(KEYINPUT121), .ZN(new_n1061));
  NAND3_X1  g636(.A1(new_n1044), .A2(new_n1061), .A3(new_n1045), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1053), .A2(KEYINPUT121), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1062), .A2(new_n1063), .ZN(new_n1064));
  OAI211_X1 g639(.A(KEYINPUT51), .B(G8), .C1(new_n1064), .C2(G286), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1057), .A2(new_n1060), .A3(new_n1065), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1041), .ZN(new_n1067));
  AOI21_X1  g642(.A(new_n1039), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT120), .ZN(new_n1069));
  NAND4_X1  g644(.A1(new_n974), .A2(new_n1069), .A3(new_n975), .A4(new_n971), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n977), .A2(new_n997), .A3(new_n1068), .A4(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(new_n1019), .ZN(new_n1072));
  NOR2_X1   g647(.A1(new_n1072), .A2(new_n1032), .ZN(new_n1073));
  AND2_X1   g648(.A1(new_n1007), .A2(new_n1010), .ZN(new_n1074));
  OR2_X1    g649(.A1(G288), .A2(G1976), .ZN(new_n1075));
  OAI22_X1  g650(.A1(new_n1074), .A2(new_n1075), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1076));
  AND2_X1   g651(.A1(new_n1076), .A2(new_n1009), .ZN(new_n1077));
  INV_X1    g652(.A(KEYINPUT63), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1019), .A2(new_n1032), .A3(new_n1037), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1046), .A2(G168), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1078), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NAND3_X1  g656(.A1(new_n1027), .A2(G8), .A3(new_n1031), .ZN(new_n1082));
  AOI21_X1  g657(.A(new_n1078), .B1(new_n1082), .B2(new_n1029), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1080), .ZN(new_n1084));
  NAND4_X1  g659(.A1(new_n1083), .A2(new_n1032), .A3(new_n1019), .A4(new_n1084), .ZN(new_n1085));
  AOI211_X1 g660(.A(new_n1073), .B(new_n1077), .C1(new_n1081), .C2(new_n1085), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1071), .A2(new_n1086), .ZN(new_n1087));
  INV_X1    g662(.A(KEYINPUT62), .ZN(new_n1088));
  NAND3_X1  g663(.A1(new_n1066), .A2(new_n1088), .A3(new_n1067), .ZN(new_n1089));
  NOR2_X1   g664(.A1(new_n1079), .A2(new_n991), .ZN(new_n1090));
  AND3_X1   g665(.A1(new_n1089), .A2(KEYINPUT126), .A3(new_n1090), .ZN(new_n1091));
  AOI21_X1  g666(.A(KEYINPUT126), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1093));
  NOR3_X1   g668(.A1(new_n1091), .A2(new_n1092), .A3(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n924), .B1(new_n1087), .B2(new_n1094), .ZN(new_n1095));
  OAI21_X1  g670(.A(new_n913), .B1(new_n918), .B2(new_n728), .ZN(new_n1096));
  XNOR2_X1  g671(.A(new_n1096), .B(KEYINPUT127), .ZN(new_n1097));
  XNOR2_X1  g672(.A(new_n915), .B(KEYINPUT46), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1097), .A2(new_n1098), .ZN(new_n1099));
  XOR2_X1   g674(.A(new_n1099), .B(KEYINPUT47), .Z(new_n1100));
  NAND3_X1  g675(.A1(new_n919), .A2(new_n711), .A3(new_n708), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n791), .A2(new_n783), .ZN(new_n1102));
  AOI211_X1 g677(.A(new_n912), .B(new_n911), .C1(new_n1101), .C2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(new_n922), .ZN(new_n1104));
  NOR2_X1   g679(.A1(G290), .A2(G1986), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1105), .A2(new_n913), .ZN(new_n1106));
  XNOR2_X1  g681(.A(new_n1106), .B(KEYINPUT48), .ZN(new_n1107));
  AOI211_X1 g682(.A(new_n1100), .B(new_n1103), .C1(new_n1104), .C2(new_n1107), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1095), .A2(new_n1108), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g684(.A(G227), .ZN(new_n1111));
  NAND3_X1  g685(.A1(new_n850), .A2(new_n642), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g686(.A(G229), .ZN(new_n1113));
  NAND4_X1  g687(.A1(new_n902), .A2(G319), .A3(new_n903), .A4(new_n1113), .ZN(new_n1114));
  NOR2_X1   g688(.A1(new_n1112), .A2(new_n1114), .ZN(G308));
  INV_X1    g689(.A(G308), .ZN(G225));
endmodule


