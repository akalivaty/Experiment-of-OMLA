

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U550 ( .A1(n519), .A2(G2105), .ZN(n886) );
  NOR2_X2 U551 ( .A1(n528), .A2(n527), .ZN(G160) );
  NOR2_X1 U552 ( .A1(n804), .A2(n803), .ZN(n805) );
  NOR2_X1 U553 ( .A1(n740), .A2(n766), .ZN(n516) );
  NOR2_X1 U554 ( .A1(G651), .A2(G543), .ZN(n636) );
  NOR2_X1 U555 ( .A1(G651), .A2(n623), .ZN(n635) );
  INV_X1 U556 ( .A(G2104), .ZN(n519) );
  NAND2_X1 U557 ( .A1(G101), .A2(n886), .ZN(n517) );
  XNOR2_X1 U558 ( .A(n517), .B(KEYINPUT65), .ZN(n518) );
  XNOR2_X1 U559 ( .A(n518), .B(KEYINPUT23), .ZN(n521) );
  INV_X1 U560 ( .A(G2105), .ZN(n522) );
  NOR2_X1 U561 ( .A1(n519), .A2(n522), .ZN(n878) );
  NAND2_X1 U562 ( .A1(n878), .A2(G113), .ZN(n520) );
  NAND2_X1 U563 ( .A1(n521), .A2(n520), .ZN(n528) );
  NOR2_X1 U564 ( .A1(G2104), .A2(n522), .ZN(n879) );
  NAND2_X1 U565 ( .A1(n879), .A2(G125), .ZN(n526) );
  NOR2_X1 U566 ( .A1(G2104), .A2(G2105), .ZN(n523) );
  XOR2_X1 U567 ( .A(KEYINPUT17), .B(n523), .Z(n524) );
  XNOR2_X2 U568 ( .A(n524), .B(KEYINPUT66), .ZN(n883) );
  NAND2_X1 U569 ( .A1(G137), .A2(n883), .ZN(n525) );
  NAND2_X1 U570 ( .A1(n526), .A2(n525), .ZN(n527) );
  AND2_X1 U571 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U572 ( .A(G57), .ZN(G237) );
  INV_X1 U573 ( .A(G132), .ZN(G219) );
  INV_X1 U574 ( .A(G82), .ZN(G220) );
  NAND2_X1 U575 ( .A1(G88), .A2(n636), .ZN(n530) );
  XOR2_X1 U576 ( .A(KEYINPUT0), .B(G543), .Z(n623) );
  INV_X1 U577 ( .A(G651), .ZN(n531) );
  NOR2_X1 U578 ( .A1(n623), .A2(n531), .ZN(n633) );
  NAND2_X1 U579 ( .A1(G75), .A2(n633), .ZN(n529) );
  NAND2_X1 U580 ( .A1(n530), .A2(n529), .ZN(n536) );
  NOR2_X1 U581 ( .A1(G543), .A2(n531), .ZN(n532) );
  XOR2_X1 U582 ( .A(KEYINPUT1), .B(n532), .Z(n639) );
  NAND2_X1 U583 ( .A1(G62), .A2(n639), .ZN(n534) );
  NAND2_X1 U584 ( .A1(G50), .A2(n635), .ZN(n533) );
  NAND2_X1 U585 ( .A1(n534), .A2(n533), .ZN(n535) );
  NOR2_X1 U586 ( .A1(n536), .A2(n535), .ZN(G166) );
  NAND2_X1 U587 ( .A1(G76), .A2(n633), .ZN(n540) );
  XOR2_X1 U588 ( .A(KEYINPUT73), .B(KEYINPUT4), .Z(n538) );
  NAND2_X1 U589 ( .A1(G89), .A2(n636), .ZN(n537) );
  XNOR2_X1 U590 ( .A(n538), .B(n537), .ZN(n539) );
  NAND2_X1 U591 ( .A1(n540), .A2(n539), .ZN(n541) );
  XNOR2_X1 U592 ( .A(n541), .B(KEYINPUT5), .ZN(n542) );
  XNOR2_X1 U593 ( .A(KEYINPUT74), .B(n542), .ZN(n547) );
  NAND2_X1 U594 ( .A1(G63), .A2(n639), .ZN(n544) );
  NAND2_X1 U595 ( .A1(G51), .A2(n635), .ZN(n543) );
  NAND2_X1 U596 ( .A1(n544), .A2(n543), .ZN(n545) );
  XOR2_X1 U597 ( .A(KEYINPUT6), .B(n545), .Z(n546) );
  NAND2_X1 U598 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U599 ( .A(KEYINPUT7), .B(n548), .ZN(G168) );
  XNOR2_X1 U600 ( .A(G168), .B(KEYINPUT8), .ZN(n549) );
  XNOR2_X1 U601 ( .A(n549), .B(KEYINPUT75), .ZN(G286) );
  NAND2_X1 U602 ( .A1(G102), .A2(n886), .ZN(n551) );
  NAND2_X1 U603 ( .A1(G138), .A2(n883), .ZN(n550) );
  NAND2_X1 U604 ( .A1(n551), .A2(n550), .ZN(n555) );
  NAND2_X1 U605 ( .A1(G114), .A2(n878), .ZN(n553) );
  NAND2_X1 U606 ( .A1(G126), .A2(n879), .ZN(n552) );
  NAND2_X1 U607 ( .A1(n553), .A2(n552), .ZN(n554) );
  NOR2_X1 U608 ( .A1(n555), .A2(n554), .ZN(G164) );
  NAND2_X1 U609 ( .A1(G7), .A2(G661), .ZN(n556) );
  XNOR2_X1 U610 ( .A(n556), .B(KEYINPUT10), .ZN(G223) );
  INV_X1 U611 ( .A(G223), .ZN(n827) );
  NAND2_X1 U612 ( .A1(n827), .A2(G567), .ZN(n557) );
  XOR2_X1 U613 ( .A(KEYINPUT11), .B(n557), .Z(G234) );
  NAND2_X1 U614 ( .A1(G81), .A2(n636), .ZN(n558) );
  XNOR2_X1 U615 ( .A(n558), .B(KEYINPUT12), .ZN(n559) );
  XNOR2_X1 U616 ( .A(n559), .B(KEYINPUT68), .ZN(n561) );
  NAND2_X1 U617 ( .A1(G68), .A2(n633), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U619 ( .A(KEYINPUT13), .B(n562), .ZN(n568) );
  NAND2_X1 U620 ( .A1(G56), .A2(n639), .ZN(n563) );
  XOR2_X1 U621 ( .A(KEYINPUT14), .B(n563), .Z(n566) );
  NAND2_X1 U622 ( .A1(G43), .A2(n635), .ZN(n564) );
  XNOR2_X1 U623 ( .A(KEYINPUT69), .B(n564), .ZN(n565) );
  NOR2_X1 U624 ( .A1(n566), .A2(n565), .ZN(n567) );
  NAND2_X1 U625 ( .A1(n568), .A2(n567), .ZN(n972) );
  INV_X1 U626 ( .A(n972), .ZN(n649) );
  NAND2_X1 U627 ( .A1(n649), .A2(G860), .ZN(G153) );
  NAND2_X1 U628 ( .A1(G90), .A2(n636), .ZN(n570) );
  NAND2_X1 U629 ( .A1(G77), .A2(n633), .ZN(n569) );
  NAND2_X1 U630 ( .A1(n570), .A2(n569), .ZN(n571) );
  XNOR2_X1 U631 ( .A(KEYINPUT9), .B(n571), .ZN(n575) );
  NAND2_X1 U632 ( .A1(G64), .A2(n639), .ZN(n573) );
  NAND2_X1 U633 ( .A1(G52), .A2(n635), .ZN(n572) );
  AND2_X1 U634 ( .A1(n573), .A2(n572), .ZN(n574) );
  NAND2_X1 U635 ( .A1(n575), .A2(n574), .ZN(G301) );
  NAND2_X1 U636 ( .A1(G301), .A2(G868), .ZN(n576) );
  XNOR2_X1 U637 ( .A(n576), .B(KEYINPUT70), .ZN(n586) );
  NAND2_X1 U638 ( .A1(G92), .A2(n636), .ZN(n578) );
  NAND2_X1 U639 ( .A1(G79), .A2(n633), .ZN(n577) );
  NAND2_X1 U640 ( .A1(n578), .A2(n577), .ZN(n582) );
  NAND2_X1 U641 ( .A1(G66), .A2(n639), .ZN(n580) );
  NAND2_X1 U642 ( .A1(G54), .A2(n635), .ZN(n579) );
  NAND2_X1 U643 ( .A1(n580), .A2(n579), .ZN(n581) );
  NOR2_X1 U644 ( .A1(n582), .A2(n581), .ZN(n584) );
  XNOR2_X1 U645 ( .A(KEYINPUT71), .B(KEYINPUT15), .ZN(n583) );
  XNOR2_X1 U646 ( .A(n584), .B(n583), .ZN(n985) );
  OR2_X1 U647 ( .A1(G868), .A2(n985), .ZN(n585) );
  NAND2_X1 U648 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U649 ( .A(KEYINPUT72), .B(n587), .ZN(G284) );
  NAND2_X1 U650 ( .A1(G65), .A2(n639), .ZN(n589) );
  NAND2_X1 U651 ( .A1(G53), .A2(n635), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n593) );
  NAND2_X1 U653 ( .A1(G91), .A2(n636), .ZN(n591) );
  NAND2_X1 U654 ( .A1(G78), .A2(n633), .ZN(n590) );
  NAND2_X1 U655 ( .A1(n591), .A2(n590), .ZN(n592) );
  NOR2_X1 U656 ( .A1(n593), .A2(n592), .ZN(n983) );
  INV_X1 U657 ( .A(n983), .ZN(G299) );
  INV_X1 U658 ( .A(G868), .ZN(n656) );
  NOR2_X1 U659 ( .A1(G286), .A2(n656), .ZN(n595) );
  NOR2_X1 U660 ( .A1(G868), .A2(G299), .ZN(n594) );
  NOR2_X1 U661 ( .A1(n595), .A2(n594), .ZN(G297) );
  INV_X1 U662 ( .A(G860), .ZN(n596) );
  NAND2_X1 U663 ( .A1(n596), .A2(G559), .ZN(n597) );
  NAND2_X1 U664 ( .A1(n597), .A2(n985), .ZN(n598) );
  XNOR2_X1 U665 ( .A(n598), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U666 ( .A1(G868), .A2(n972), .ZN(n601) );
  NAND2_X1 U667 ( .A1(G868), .A2(n985), .ZN(n599) );
  NOR2_X1 U668 ( .A1(G559), .A2(n599), .ZN(n600) );
  NOR2_X1 U669 ( .A1(n601), .A2(n600), .ZN(G282) );
  NAND2_X1 U670 ( .A1(G123), .A2(n879), .ZN(n602) );
  XNOR2_X1 U671 ( .A(n602), .B(KEYINPUT18), .ZN(n604) );
  NAND2_X1 U672 ( .A1(n878), .A2(G111), .ZN(n603) );
  NAND2_X1 U673 ( .A1(n604), .A2(n603), .ZN(n608) );
  NAND2_X1 U674 ( .A1(G99), .A2(n886), .ZN(n606) );
  NAND2_X1 U675 ( .A1(G135), .A2(n883), .ZN(n605) );
  NAND2_X1 U676 ( .A1(n606), .A2(n605), .ZN(n607) );
  NOR2_X1 U677 ( .A1(n608), .A2(n607), .ZN(n954) );
  XNOR2_X1 U678 ( .A(G2096), .B(n954), .ZN(n610) );
  INV_X1 U679 ( .A(G2100), .ZN(n609) );
  NAND2_X1 U680 ( .A1(n610), .A2(n609), .ZN(G156) );
  NAND2_X1 U681 ( .A1(n985), .A2(G559), .ZN(n652) );
  XNOR2_X1 U682 ( .A(n972), .B(n652), .ZN(n611) );
  NOR2_X1 U683 ( .A1(n611), .A2(G860), .ZN(n619) );
  NAND2_X1 U684 ( .A1(G67), .A2(n639), .ZN(n613) );
  NAND2_X1 U685 ( .A1(G55), .A2(n635), .ZN(n612) );
  NAND2_X1 U686 ( .A1(n613), .A2(n612), .ZN(n614) );
  XNOR2_X1 U687 ( .A(KEYINPUT76), .B(n614), .ZN(n618) );
  NAND2_X1 U688 ( .A1(G93), .A2(n636), .ZN(n616) );
  NAND2_X1 U689 ( .A1(G80), .A2(n633), .ZN(n615) );
  NAND2_X1 U690 ( .A1(n616), .A2(n615), .ZN(n617) );
  OR2_X1 U691 ( .A1(n618), .A2(n617), .ZN(n657) );
  XOR2_X1 U692 ( .A(n619), .B(n657), .Z(G145) );
  NAND2_X1 U693 ( .A1(G49), .A2(n635), .ZN(n621) );
  NAND2_X1 U694 ( .A1(G74), .A2(G651), .ZN(n620) );
  NAND2_X1 U695 ( .A1(n621), .A2(n620), .ZN(n622) );
  NOR2_X1 U696 ( .A1(n639), .A2(n622), .ZN(n625) );
  NAND2_X1 U697 ( .A1(n623), .A2(G87), .ZN(n624) );
  NAND2_X1 U698 ( .A1(n625), .A2(n624), .ZN(G288) );
  NAND2_X1 U699 ( .A1(G60), .A2(n639), .ZN(n627) );
  NAND2_X1 U700 ( .A1(G72), .A2(n633), .ZN(n626) );
  NAND2_X1 U701 ( .A1(n627), .A2(n626), .ZN(n630) );
  NAND2_X1 U702 ( .A1(G85), .A2(n636), .ZN(n628) );
  XNOR2_X1 U703 ( .A(KEYINPUT67), .B(n628), .ZN(n629) );
  NOR2_X1 U704 ( .A1(n630), .A2(n629), .ZN(n632) );
  NAND2_X1 U705 ( .A1(n635), .A2(G47), .ZN(n631) );
  NAND2_X1 U706 ( .A1(n632), .A2(n631), .ZN(G290) );
  NAND2_X1 U707 ( .A1(G73), .A2(n633), .ZN(n634) );
  XNOR2_X1 U708 ( .A(n634), .B(KEYINPUT2), .ZN(n644) );
  NAND2_X1 U709 ( .A1(G48), .A2(n635), .ZN(n638) );
  NAND2_X1 U710 ( .A1(G86), .A2(n636), .ZN(n637) );
  NAND2_X1 U711 ( .A1(n638), .A2(n637), .ZN(n642) );
  NAND2_X1 U712 ( .A1(G61), .A2(n639), .ZN(n640) );
  XNOR2_X1 U713 ( .A(KEYINPUT77), .B(n640), .ZN(n641) );
  NOR2_X1 U714 ( .A1(n642), .A2(n641), .ZN(n643) );
  NAND2_X1 U715 ( .A1(n644), .A2(n643), .ZN(G305) );
  XNOR2_X1 U716 ( .A(G290), .B(KEYINPUT19), .ZN(n646) );
  XNOR2_X1 U717 ( .A(n983), .B(G166), .ZN(n645) );
  XNOR2_X1 U718 ( .A(n646), .B(n645), .ZN(n647) );
  XOR2_X1 U719 ( .A(n647), .B(G305), .Z(n648) );
  XNOR2_X1 U720 ( .A(G288), .B(n648), .ZN(n651) );
  XOR2_X1 U721 ( .A(n657), .B(n649), .Z(n650) );
  XNOR2_X1 U722 ( .A(n651), .B(n650), .ZN(n899) );
  XNOR2_X1 U723 ( .A(n899), .B(KEYINPUT78), .ZN(n653) );
  XNOR2_X1 U724 ( .A(n653), .B(n652), .ZN(n654) );
  NAND2_X1 U725 ( .A1(n654), .A2(G868), .ZN(n655) );
  XOR2_X1 U726 ( .A(KEYINPUT79), .B(n655), .Z(n659) );
  NAND2_X1 U727 ( .A1(n657), .A2(n656), .ZN(n658) );
  NAND2_X1 U728 ( .A1(n659), .A2(n658), .ZN(G295) );
  NAND2_X1 U729 ( .A1(G2084), .A2(G2078), .ZN(n660) );
  XOR2_X1 U730 ( .A(KEYINPUT20), .B(n660), .Z(n661) );
  NAND2_X1 U731 ( .A1(n661), .A2(G2090), .ZN(n662) );
  XNOR2_X1 U732 ( .A(n662), .B(KEYINPUT80), .ZN(n663) );
  XNOR2_X1 U733 ( .A(KEYINPUT21), .B(n663), .ZN(n664) );
  NAND2_X1 U734 ( .A1(G2072), .A2(n664), .ZN(G158) );
  XNOR2_X1 U735 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U736 ( .A1(G220), .A2(G219), .ZN(n665) );
  XNOR2_X1 U737 ( .A(KEYINPUT22), .B(n665), .ZN(n666) );
  NAND2_X1 U738 ( .A1(n666), .A2(G96), .ZN(n667) );
  NOR2_X1 U739 ( .A1(n667), .A2(G218), .ZN(n668) );
  XNOR2_X1 U740 ( .A(n668), .B(KEYINPUT81), .ZN(n832) );
  NAND2_X1 U741 ( .A1(n832), .A2(G2106), .ZN(n673) );
  NAND2_X1 U742 ( .A1(G69), .A2(G120), .ZN(n669) );
  NOR2_X1 U743 ( .A1(G237), .A2(n669), .ZN(n670) );
  NAND2_X1 U744 ( .A1(G108), .A2(n670), .ZN(n831) );
  NAND2_X1 U745 ( .A1(G567), .A2(n831), .ZN(n671) );
  XNOR2_X1 U746 ( .A(KEYINPUT82), .B(n671), .ZN(n672) );
  NAND2_X1 U747 ( .A1(n673), .A2(n672), .ZN(n833) );
  NAND2_X1 U748 ( .A1(G661), .A2(G483), .ZN(n674) );
  NOR2_X1 U749 ( .A1(n833), .A2(n674), .ZN(n675) );
  XOR2_X1 U750 ( .A(KEYINPUT83), .B(n675), .Z(n830) );
  NAND2_X1 U751 ( .A1(n830), .A2(G36), .ZN(G176) );
  INV_X1 U752 ( .A(G166), .ZN(G303) );
  INV_X1 U753 ( .A(G301), .ZN(G171) );
  NAND2_X1 U754 ( .A1(G160), .A2(G40), .ZN(n783) );
  INV_X1 U755 ( .A(n783), .ZN(n676) );
  NOR2_X1 U756 ( .A1(G164), .A2(G1384), .ZN(n782) );
  NAND2_X1 U757 ( .A1(n676), .A2(n782), .ZN(n677) );
  XNOR2_X1 U758 ( .A(n677), .B(KEYINPUT64), .ZN(n678) );
  INV_X1 U759 ( .A(n678), .ZN(n704) );
  INV_X1 U760 ( .A(n704), .ZN(n719) );
  NOR2_X1 U761 ( .A1(n719), .A2(G2084), .ZN(n736) );
  NAND2_X1 U762 ( .A1(n678), .A2(G8), .ZN(n766) );
  NOR2_X1 U763 ( .A1(n766), .A2(G1966), .ZN(n679) );
  XNOR2_X1 U764 ( .A(n679), .B(KEYINPUT91), .ZN(n735) );
  NAND2_X1 U765 ( .A1(G8), .A2(n735), .ZN(n680) );
  NOR2_X1 U766 ( .A1(n736), .A2(n680), .ZN(n681) );
  XOR2_X1 U767 ( .A(KEYINPUT30), .B(n681), .Z(n682) );
  NOR2_X1 U768 ( .A1(G168), .A2(n682), .ZN(n686) );
  XNOR2_X1 U769 ( .A(KEYINPUT25), .B(G2078), .ZN(n921) );
  NAND2_X1 U770 ( .A1(n704), .A2(n921), .ZN(n684) );
  INV_X1 U771 ( .A(G1961), .ZN(n1010) );
  NAND2_X1 U772 ( .A1(n719), .A2(n1010), .ZN(n683) );
  NAND2_X1 U773 ( .A1(n684), .A2(n683), .ZN(n689) );
  NOR2_X1 U774 ( .A1(G171), .A2(n689), .ZN(n685) );
  NOR2_X1 U775 ( .A1(n686), .A2(n685), .ZN(n687) );
  XOR2_X1 U776 ( .A(n687), .B(KEYINPUT96), .Z(n688) );
  XNOR2_X1 U777 ( .A(n688), .B(KEYINPUT31), .ZN(n732) );
  NAND2_X1 U778 ( .A1(n689), .A2(G171), .ZN(n717) );
  NAND2_X1 U779 ( .A1(G2072), .A2(n704), .ZN(n690) );
  XOR2_X1 U780 ( .A(KEYINPUT27), .B(n690), .Z(n692) );
  NAND2_X1 U781 ( .A1(n719), .A2(G1956), .ZN(n691) );
  NAND2_X1 U782 ( .A1(n692), .A2(n691), .ZN(n693) );
  XOR2_X1 U783 ( .A(KEYINPUT92), .B(n693), .Z(n696) );
  NOR2_X1 U784 ( .A1(n983), .A2(n696), .ZN(n695) );
  XNOR2_X1 U785 ( .A(KEYINPUT93), .B(KEYINPUT28), .ZN(n694) );
  XNOR2_X1 U786 ( .A(n695), .B(n694), .ZN(n714) );
  NAND2_X1 U787 ( .A1(n983), .A2(n696), .ZN(n712) );
  AND2_X1 U788 ( .A1(n704), .A2(G1996), .ZN(n698) );
  XOR2_X1 U789 ( .A(KEYINPUT26), .B(KEYINPUT94), .Z(n697) );
  XNOR2_X1 U790 ( .A(n698), .B(n697), .ZN(n700) );
  NAND2_X1 U791 ( .A1(n719), .A2(G1341), .ZN(n699) );
  NAND2_X1 U792 ( .A1(n700), .A2(n699), .ZN(n701) );
  NOR2_X1 U793 ( .A1(n972), .A2(n701), .ZN(n703) );
  NOR2_X1 U794 ( .A1(n703), .A2(n985), .ZN(n702) );
  XNOR2_X1 U795 ( .A(n702), .B(KEYINPUT95), .ZN(n710) );
  NAND2_X1 U796 ( .A1(n703), .A2(n985), .ZN(n708) );
  NOR2_X1 U797 ( .A1(n719), .A2(G2067), .ZN(n706) );
  NOR2_X1 U798 ( .A1(G1348), .A2(n704), .ZN(n705) );
  NOR2_X1 U799 ( .A1(n706), .A2(n705), .ZN(n707) );
  NAND2_X1 U800 ( .A1(n708), .A2(n707), .ZN(n709) );
  NAND2_X1 U801 ( .A1(n710), .A2(n709), .ZN(n711) );
  NAND2_X1 U802 ( .A1(n712), .A2(n711), .ZN(n713) );
  NAND2_X1 U803 ( .A1(n714), .A2(n713), .ZN(n715) );
  XOR2_X1 U804 ( .A(KEYINPUT29), .B(n715), .Z(n716) );
  NAND2_X1 U805 ( .A1(n717), .A2(n716), .ZN(n733) );
  INV_X1 U806 ( .A(G8), .ZN(n724) );
  NOR2_X1 U807 ( .A1(G1971), .A2(n766), .ZN(n718) );
  XNOR2_X1 U808 ( .A(KEYINPUT97), .B(n718), .ZN(n722) );
  NOR2_X1 U809 ( .A1(n719), .A2(G2090), .ZN(n720) );
  NOR2_X1 U810 ( .A1(G166), .A2(n720), .ZN(n721) );
  NAND2_X1 U811 ( .A1(n722), .A2(n721), .ZN(n723) );
  OR2_X1 U812 ( .A1(n724), .A2(n723), .ZN(n726) );
  AND2_X1 U813 ( .A1(n733), .A2(n726), .ZN(n725) );
  NAND2_X1 U814 ( .A1(n732), .A2(n725), .ZN(n730) );
  INV_X1 U815 ( .A(n726), .ZN(n728) );
  AND2_X1 U816 ( .A1(G286), .A2(G8), .ZN(n727) );
  OR2_X1 U817 ( .A1(n728), .A2(n727), .ZN(n729) );
  NAND2_X1 U818 ( .A1(n730), .A2(n729), .ZN(n731) );
  XNOR2_X1 U819 ( .A(n731), .B(KEYINPUT32), .ZN(n756) );
  XOR2_X1 U820 ( .A(G1981), .B(G305), .Z(n979) );
  AND2_X1 U821 ( .A1(n756), .A2(n979), .ZN(n745) );
  NAND2_X1 U822 ( .A1(n733), .A2(n732), .ZN(n734) );
  AND2_X1 U823 ( .A1(n735), .A2(n734), .ZN(n738) );
  NAND2_X1 U824 ( .A1(G8), .A2(n736), .ZN(n737) );
  NAND2_X1 U825 ( .A1(n738), .A2(n737), .ZN(n757) );
  NAND2_X1 U826 ( .A1(G288), .A2(G1976), .ZN(n739) );
  XNOR2_X1 U827 ( .A(n739), .B(KEYINPUT98), .ZN(n978) );
  INV_X1 U828 ( .A(n978), .ZN(n740) );
  NOR2_X1 U829 ( .A1(KEYINPUT33), .A2(n516), .ZN(n743) );
  NOR2_X1 U830 ( .A1(G1976), .A2(G288), .ZN(n748) );
  NAND2_X1 U831 ( .A1(n748), .A2(KEYINPUT33), .ZN(n741) );
  NOR2_X1 U832 ( .A1(n741), .A2(n766), .ZN(n742) );
  NOR2_X1 U833 ( .A1(n743), .A2(n742), .ZN(n746) );
  AND2_X1 U834 ( .A1(n757), .A2(n746), .ZN(n744) );
  NAND2_X1 U835 ( .A1(n745), .A2(n744), .ZN(n755) );
  INV_X1 U836 ( .A(n979), .ZN(n753) );
  INV_X1 U837 ( .A(n746), .ZN(n751) );
  NOR2_X1 U838 ( .A1(G1971), .A2(G303), .ZN(n747) );
  NOR2_X1 U839 ( .A1(n748), .A2(n747), .ZN(n976) );
  INV_X1 U840 ( .A(KEYINPUT33), .ZN(n749) );
  AND2_X1 U841 ( .A1(n976), .A2(n749), .ZN(n750) );
  OR2_X1 U842 ( .A1(n751), .A2(n750), .ZN(n752) );
  OR2_X1 U843 ( .A1(n753), .A2(n752), .ZN(n754) );
  NAND2_X1 U844 ( .A1(n755), .A2(n754), .ZN(n771) );
  NAND2_X1 U845 ( .A1(n757), .A2(n756), .ZN(n765) );
  NAND2_X1 U846 ( .A1(G8), .A2(G166), .ZN(n758) );
  NOR2_X1 U847 ( .A1(G2090), .A2(n758), .ZN(n759) );
  XNOR2_X1 U848 ( .A(n759), .B(KEYINPUT99), .ZN(n763) );
  NOR2_X1 U849 ( .A1(G1981), .A2(G305), .ZN(n760) );
  XOR2_X1 U850 ( .A(n760), .B(KEYINPUT24), .Z(n761) );
  NOR2_X1 U851 ( .A1(n766), .A2(n761), .ZN(n767) );
  INV_X1 U852 ( .A(n767), .ZN(n762) );
  AND2_X1 U853 ( .A1(n763), .A2(n762), .ZN(n764) );
  NAND2_X1 U854 ( .A1(n765), .A2(n764), .ZN(n769) );
  OR2_X1 U855 ( .A1(n767), .A2(n766), .ZN(n768) );
  AND2_X1 U856 ( .A1(n769), .A2(n768), .ZN(n770) );
  NOR2_X1 U857 ( .A1(n771), .A2(n770), .ZN(n804) );
  XNOR2_X1 U858 ( .A(G2067), .B(KEYINPUT37), .ZN(n820) );
  NAND2_X1 U859 ( .A1(G104), .A2(n886), .ZN(n773) );
  NAND2_X1 U860 ( .A1(G140), .A2(n883), .ZN(n772) );
  NAND2_X1 U861 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U862 ( .A(KEYINPUT34), .B(n774), .ZN(n779) );
  NAND2_X1 U863 ( .A1(G116), .A2(n878), .ZN(n776) );
  NAND2_X1 U864 ( .A1(G128), .A2(n879), .ZN(n775) );
  NAND2_X1 U865 ( .A1(n776), .A2(n775), .ZN(n777) );
  XOR2_X1 U866 ( .A(n777), .B(KEYINPUT35), .Z(n778) );
  NOR2_X1 U867 ( .A1(n779), .A2(n778), .ZN(n780) );
  XOR2_X1 U868 ( .A(KEYINPUT36), .B(n780), .Z(n781) );
  XNOR2_X1 U869 ( .A(KEYINPUT87), .B(n781), .ZN(n895) );
  NOR2_X1 U870 ( .A1(n820), .A2(n895), .ZN(n959) );
  NOR2_X1 U871 ( .A1(n783), .A2(n782), .ZN(n784) );
  XNOR2_X1 U872 ( .A(n784), .B(KEYINPUT85), .ZN(n807) );
  INV_X1 U873 ( .A(n807), .ZN(n822) );
  NAND2_X1 U874 ( .A1(n959), .A2(n822), .ZN(n819) );
  NAND2_X1 U875 ( .A1(G105), .A2(n886), .ZN(n785) );
  XNOR2_X1 U876 ( .A(n785), .B(KEYINPUT38), .ZN(n792) );
  NAND2_X1 U877 ( .A1(n879), .A2(G129), .ZN(n787) );
  NAND2_X1 U878 ( .A1(G141), .A2(n883), .ZN(n786) );
  NAND2_X1 U879 ( .A1(n787), .A2(n786), .ZN(n790) );
  NAND2_X1 U880 ( .A1(n878), .A2(G117), .ZN(n788) );
  XOR2_X1 U881 ( .A(KEYINPUT90), .B(n788), .Z(n789) );
  NOR2_X1 U882 ( .A1(n790), .A2(n789), .ZN(n791) );
  NAND2_X1 U883 ( .A1(n792), .A2(n791), .ZN(n890) );
  NAND2_X1 U884 ( .A1(G1996), .A2(n890), .ZN(n802) );
  NAND2_X1 U885 ( .A1(n879), .A2(G119), .ZN(n793) );
  XNOR2_X1 U886 ( .A(n793), .B(KEYINPUT88), .ZN(n795) );
  NAND2_X1 U887 ( .A1(G107), .A2(n878), .ZN(n794) );
  NAND2_X1 U888 ( .A1(n795), .A2(n794), .ZN(n796) );
  XNOR2_X1 U889 ( .A(KEYINPUT89), .B(n796), .ZN(n800) );
  NAND2_X1 U890 ( .A1(n883), .A2(G131), .ZN(n798) );
  NAND2_X1 U891 ( .A1(G95), .A2(n886), .ZN(n797) );
  AND2_X1 U892 ( .A1(n798), .A2(n797), .ZN(n799) );
  NAND2_X1 U893 ( .A1(n800), .A2(n799), .ZN(n867) );
  NAND2_X1 U894 ( .A1(G1991), .A2(n867), .ZN(n801) );
  NAND2_X1 U895 ( .A1(n802), .A2(n801), .ZN(n955) );
  NAND2_X1 U896 ( .A1(n822), .A2(n955), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n819), .A2(n811), .ZN(n803) );
  XNOR2_X1 U898 ( .A(n805), .B(KEYINPUT100), .ZN(n810) );
  XOR2_X1 U899 ( .A(KEYINPUT84), .B(G1986), .Z(n806) );
  XNOR2_X1 U900 ( .A(G290), .B(n806), .ZN(n975) );
  NOR2_X1 U901 ( .A1(n807), .A2(n975), .ZN(n808) );
  XOR2_X1 U902 ( .A(KEYINPUT86), .B(n808), .Z(n809) );
  NAND2_X1 U903 ( .A1(n810), .A2(n809), .ZN(n825) );
  NOR2_X1 U904 ( .A1(G1996), .A2(n890), .ZN(n948) );
  INV_X1 U905 ( .A(n811), .ZN(n814) );
  NOR2_X1 U906 ( .A1(G1986), .A2(G290), .ZN(n812) );
  NOR2_X1 U907 ( .A1(G1991), .A2(n867), .ZN(n956) );
  NOR2_X1 U908 ( .A1(n812), .A2(n956), .ZN(n813) );
  NOR2_X1 U909 ( .A1(n814), .A2(n813), .ZN(n815) );
  NOR2_X1 U910 ( .A1(n948), .A2(n815), .ZN(n816) );
  XOR2_X1 U911 ( .A(n816), .B(KEYINPUT39), .Z(n817) );
  XNOR2_X1 U912 ( .A(KEYINPUT101), .B(n817), .ZN(n818) );
  NAND2_X1 U913 ( .A1(n819), .A2(n818), .ZN(n821) );
  NAND2_X1 U914 ( .A1(n820), .A2(n895), .ZN(n945) );
  NAND2_X1 U915 ( .A1(n821), .A2(n945), .ZN(n823) );
  NAND2_X1 U916 ( .A1(n823), .A2(n822), .ZN(n824) );
  NAND2_X1 U917 ( .A1(n825), .A2(n824), .ZN(n826) );
  XNOR2_X1 U918 ( .A(n826), .B(KEYINPUT40), .ZN(G329) );
  NAND2_X1 U919 ( .A1(G2106), .A2(n827), .ZN(G217) );
  AND2_X1 U920 ( .A1(G15), .A2(G2), .ZN(n828) );
  NAND2_X1 U921 ( .A1(G661), .A2(n828), .ZN(G259) );
  NAND2_X1 U922 ( .A1(G3), .A2(G1), .ZN(n829) );
  NAND2_X1 U923 ( .A1(n830), .A2(n829), .ZN(G188) );
  INV_X1 U925 ( .A(G120), .ZN(G236) );
  INV_X1 U926 ( .A(G96), .ZN(G221) );
  INV_X1 U927 ( .A(G69), .ZN(G235) );
  NOR2_X1 U928 ( .A1(n832), .A2(n831), .ZN(G325) );
  INV_X1 U929 ( .A(G325), .ZN(G261) );
  INV_X1 U930 ( .A(n833), .ZN(G319) );
  XOR2_X1 U931 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n835) );
  XNOR2_X1 U932 ( .A(KEYINPUT104), .B(G2096), .ZN(n834) );
  XNOR2_X1 U933 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U934 ( .A(n836), .B(KEYINPUT105), .Z(n838) );
  XNOR2_X1 U935 ( .A(G2078), .B(G2072), .ZN(n837) );
  XNOR2_X1 U936 ( .A(n838), .B(n837), .ZN(n842) );
  XOR2_X1 U937 ( .A(G2100), .B(G2090), .Z(n840) );
  XNOR2_X1 U938 ( .A(G2084), .B(G2067), .ZN(n839) );
  XNOR2_X1 U939 ( .A(n840), .B(n839), .ZN(n841) );
  XOR2_X1 U940 ( .A(n842), .B(n841), .Z(n844) );
  XNOR2_X1 U941 ( .A(G2678), .B(KEYINPUT43), .ZN(n843) );
  XNOR2_X1 U942 ( .A(n844), .B(n843), .ZN(G227) );
  XOR2_X1 U943 ( .A(G1981), .B(G1971), .Z(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1956), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n847), .B(G2474), .Z(n849) );
  XNOR2_X1 U947 ( .A(G1996), .B(G1991), .ZN(n848) );
  XNOR2_X1 U948 ( .A(n849), .B(n848), .ZN(n853) );
  XOR2_X1 U949 ( .A(KEYINPUT41), .B(G1986), .Z(n851) );
  XNOR2_X1 U950 ( .A(G1961), .B(G1976), .ZN(n850) );
  XNOR2_X1 U951 ( .A(n851), .B(n850), .ZN(n852) );
  XNOR2_X1 U952 ( .A(n853), .B(n852), .ZN(G229) );
  NAND2_X1 U953 ( .A1(G100), .A2(n886), .ZN(n854) );
  XNOR2_X1 U954 ( .A(n854), .B(KEYINPUT108), .ZN(n857) );
  NAND2_X1 U955 ( .A1(n883), .A2(G136), .ZN(n855) );
  XOR2_X1 U956 ( .A(KEYINPUT107), .B(n855), .Z(n856) );
  NAND2_X1 U957 ( .A1(n857), .A2(n856), .ZN(n862) );
  NAND2_X1 U958 ( .A1(G124), .A2(n879), .ZN(n858) );
  XNOR2_X1 U959 ( .A(n858), .B(KEYINPUT44), .ZN(n860) );
  NAND2_X1 U960 ( .A1(n878), .A2(G112), .ZN(n859) );
  NAND2_X1 U961 ( .A1(n860), .A2(n859), .ZN(n861) );
  NOR2_X1 U962 ( .A1(n862), .A2(n861), .ZN(G162) );
  XOR2_X1 U963 ( .A(KEYINPUT46), .B(KEYINPUT48), .Z(n864) );
  XNOR2_X1 U964 ( .A(G162), .B(KEYINPUT111), .ZN(n863) );
  XNOR2_X1 U965 ( .A(n864), .B(n863), .ZN(n865) );
  XNOR2_X1 U966 ( .A(G164), .B(n865), .ZN(n894) );
  XOR2_X1 U967 ( .A(G160), .B(n954), .Z(n866) );
  XNOR2_X1 U968 ( .A(n867), .B(n866), .ZN(n877) );
  NAND2_X1 U969 ( .A1(G106), .A2(n886), .ZN(n869) );
  NAND2_X1 U970 ( .A1(G142), .A2(n883), .ZN(n868) );
  NAND2_X1 U971 ( .A1(n869), .A2(n868), .ZN(n870) );
  XNOR2_X1 U972 ( .A(n870), .B(KEYINPUT45), .ZN(n872) );
  NAND2_X1 U973 ( .A1(G118), .A2(n878), .ZN(n871) );
  NAND2_X1 U974 ( .A1(n872), .A2(n871), .ZN(n875) );
  NAND2_X1 U975 ( .A1(G130), .A2(n879), .ZN(n873) );
  XNOR2_X1 U976 ( .A(KEYINPUT109), .B(n873), .ZN(n874) );
  NOR2_X1 U977 ( .A1(n875), .A2(n874), .ZN(n876) );
  XNOR2_X1 U978 ( .A(n877), .B(n876), .ZN(n892) );
  NAND2_X1 U979 ( .A1(G115), .A2(n878), .ZN(n881) );
  NAND2_X1 U980 ( .A1(G127), .A2(n879), .ZN(n880) );
  NAND2_X1 U981 ( .A1(n881), .A2(n880), .ZN(n882) );
  XNOR2_X1 U982 ( .A(n882), .B(KEYINPUT47), .ZN(n885) );
  NAND2_X1 U983 ( .A1(G139), .A2(n883), .ZN(n884) );
  NAND2_X1 U984 ( .A1(n885), .A2(n884), .ZN(n889) );
  NAND2_X1 U985 ( .A1(n886), .A2(G103), .ZN(n887) );
  XOR2_X1 U986 ( .A(KEYINPUT110), .B(n887), .Z(n888) );
  NOR2_X1 U987 ( .A1(n889), .A2(n888), .ZN(n941) );
  XNOR2_X1 U988 ( .A(n890), .B(n941), .ZN(n891) );
  XNOR2_X1 U989 ( .A(n892), .B(n891), .ZN(n893) );
  XNOR2_X1 U990 ( .A(n894), .B(n893), .ZN(n896) );
  XOR2_X1 U991 ( .A(n896), .B(n895), .Z(n897) );
  NOR2_X1 U992 ( .A1(G37), .A2(n897), .ZN(G395) );
  XOR2_X1 U993 ( .A(n985), .B(G286), .Z(n898) );
  XNOR2_X1 U994 ( .A(n899), .B(n898), .ZN(n900) );
  XNOR2_X1 U995 ( .A(n900), .B(G171), .ZN(n901) );
  NOR2_X1 U996 ( .A1(G37), .A2(n901), .ZN(G397) );
  XNOR2_X1 U997 ( .A(G2427), .B(KEYINPUT102), .ZN(n911) );
  XOR2_X1 U998 ( .A(G2430), .B(G2446), .Z(n903) );
  XNOR2_X1 U999 ( .A(G2435), .B(G2438), .ZN(n902) );
  XNOR2_X1 U1000 ( .A(n903), .B(n902), .ZN(n907) );
  XOR2_X1 U1001 ( .A(G2454), .B(KEYINPUT103), .Z(n905) );
  XNOR2_X1 U1002 ( .A(G1348), .B(G1341), .ZN(n904) );
  XNOR2_X1 U1003 ( .A(n905), .B(n904), .ZN(n906) );
  XOR2_X1 U1004 ( .A(n907), .B(n906), .Z(n909) );
  XNOR2_X1 U1005 ( .A(G2451), .B(G2443), .ZN(n908) );
  XNOR2_X1 U1006 ( .A(n909), .B(n908), .ZN(n910) );
  XNOR2_X1 U1007 ( .A(n911), .B(n910), .ZN(n912) );
  NAND2_X1 U1008 ( .A1(n912), .A2(G14), .ZN(n918) );
  NAND2_X1 U1009 ( .A1(G319), .A2(n918), .ZN(n915) );
  NOR2_X1 U1010 ( .A1(G227), .A2(G229), .ZN(n913) );
  XNOR2_X1 U1011 ( .A(KEYINPUT49), .B(n913), .ZN(n914) );
  NOR2_X1 U1012 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1013 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1014 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1015 ( .A(G225), .ZN(G308) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G1991), .B(G25), .Z(n919) );
  NAND2_X1 U1019 ( .A1(G28), .A2(n919), .ZN(n920) );
  XNOR2_X1 U1020 ( .A(KEYINPUT117), .B(n920), .ZN(n931) );
  XNOR2_X1 U1021 ( .A(G27), .B(n921), .ZN(n925) );
  XNOR2_X1 U1022 ( .A(G1996), .B(G32), .ZN(n923) );
  XNOR2_X1 U1023 ( .A(G33), .B(G2072), .ZN(n922) );
  NOR2_X1 U1024 ( .A1(n923), .A2(n922), .ZN(n924) );
  NAND2_X1 U1025 ( .A1(n925), .A2(n924), .ZN(n928) );
  XNOR2_X1 U1026 ( .A(KEYINPUT118), .B(G2067), .ZN(n926) );
  XNOR2_X1 U1027 ( .A(G26), .B(n926), .ZN(n927) );
  NOR2_X1 U1028 ( .A1(n928), .A2(n927), .ZN(n929) );
  XOR2_X1 U1029 ( .A(KEYINPUT119), .B(n929), .Z(n930) );
  NAND2_X1 U1030 ( .A1(n931), .A2(n930), .ZN(n932) );
  XNOR2_X1 U1031 ( .A(n932), .B(KEYINPUT53), .ZN(n935) );
  XOR2_X1 U1032 ( .A(G2084), .B(G34), .Z(n933) );
  XNOR2_X1 U1033 ( .A(KEYINPUT54), .B(n933), .ZN(n934) );
  NAND2_X1 U1034 ( .A1(n935), .A2(n934), .ZN(n938) );
  XNOR2_X1 U1035 ( .A(KEYINPUT116), .B(G2090), .ZN(n936) );
  XNOR2_X1 U1036 ( .A(G35), .B(n936), .ZN(n937) );
  NOR2_X1 U1037 ( .A1(n938), .A2(n937), .ZN(n939) );
  XOR2_X1 U1038 ( .A(KEYINPUT55), .B(n939), .Z(n940) );
  NOR2_X1 U1039 ( .A1(G29), .A2(n940), .ZN(n970) );
  XOR2_X1 U1040 ( .A(G2072), .B(n941), .Z(n943) );
  XOR2_X1 U1041 ( .A(G164), .B(G2078), .Z(n942) );
  NOR2_X1 U1042 ( .A1(n943), .A2(n942), .ZN(n944) );
  XNOR2_X1 U1043 ( .A(n944), .B(KEYINPUT50), .ZN(n946) );
  NAND2_X1 U1044 ( .A1(n946), .A2(n945), .ZN(n952) );
  XOR2_X1 U1045 ( .A(G2090), .B(G162), .Z(n947) );
  NOR2_X1 U1046 ( .A1(n948), .A2(n947), .ZN(n949) );
  XOR2_X1 U1047 ( .A(KEYINPUT112), .B(n949), .Z(n950) );
  XOR2_X1 U1048 ( .A(KEYINPUT51), .B(n950), .Z(n951) );
  NOR2_X1 U1049 ( .A1(n952), .A2(n951), .ZN(n962) );
  XOR2_X1 U1050 ( .A(G2084), .B(G160), .Z(n953) );
  NOR2_X1 U1051 ( .A1(n954), .A2(n953), .ZN(n958) );
  NOR2_X1 U1052 ( .A1(n956), .A2(n955), .ZN(n957) );
  NAND2_X1 U1053 ( .A1(n958), .A2(n957), .ZN(n960) );
  NOR2_X1 U1054 ( .A1(n960), .A2(n959), .ZN(n961) );
  NAND2_X1 U1055 ( .A1(n962), .A2(n961), .ZN(n963) );
  XNOR2_X1 U1056 ( .A(KEYINPUT52), .B(n963), .ZN(n964) );
  XOR2_X1 U1057 ( .A(KEYINPUT113), .B(n964), .Z(n965) );
  NOR2_X1 U1058 ( .A1(KEYINPUT55), .A2(n965), .ZN(n966) );
  XOR2_X1 U1059 ( .A(KEYINPUT114), .B(n966), .Z(n967) );
  NAND2_X1 U1060 ( .A1(n967), .A2(G29), .ZN(n968) );
  XNOR2_X1 U1061 ( .A(KEYINPUT115), .B(n968), .ZN(n969) );
  NOR2_X1 U1062 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1063 ( .A1(G11), .A2(n971), .ZN(n1029) );
  XNOR2_X1 U1064 ( .A(G16), .B(KEYINPUT56), .ZN(n997) );
  XNOR2_X1 U1065 ( .A(G301), .B(G1961), .ZN(n974) );
  XNOR2_X1 U1066 ( .A(n972), .B(G1341), .ZN(n973) );
  NOR2_X1 U1067 ( .A1(n974), .A2(n973), .ZN(n995) );
  AND2_X1 U1068 ( .A1(n976), .A2(n975), .ZN(n977) );
  NAND2_X1 U1069 ( .A1(n978), .A2(n977), .ZN(n993) );
  XNOR2_X1 U1070 ( .A(G1966), .B(G168), .ZN(n980) );
  NAND2_X1 U1071 ( .A1(n980), .A2(n979), .ZN(n981) );
  XNOR2_X1 U1072 ( .A(n981), .B(KEYINPUT120), .ZN(n982) );
  XNOR2_X1 U1073 ( .A(KEYINPUT57), .B(n982), .ZN(n991) );
  XNOR2_X1 U1074 ( .A(n983), .B(G1956), .ZN(n984) );
  XNOR2_X1 U1075 ( .A(n984), .B(KEYINPUT121), .ZN(n989) );
  XNOR2_X1 U1076 ( .A(G1348), .B(n985), .ZN(n987) );
  NAND2_X1 U1077 ( .A1(G1971), .A2(G303), .ZN(n986) );
  NAND2_X1 U1078 ( .A1(n987), .A2(n986), .ZN(n988) );
  NOR2_X1 U1079 ( .A1(n989), .A2(n988), .ZN(n990) );
  NAND2_X1 U1080 ( .A1(n991), .A2(n990), .ZN(n992) );
  NOR2_X1 U1081 ( .A1(n993), .A2(n992), .ZN(n994) );
  NAND2_X1 U1082 ( .A1(n995), .A2(n994), .ZN(n996) );
  NAND2_X1 U1083 ( .A1(n997), .A2(n996), .ZN(n1026) );
  INV_X1 U1084 ( .A(G16), .ZN(n1024) );
  XOR2_X1 U1085 ( .A(G1348), .B(KEYINPUT59), .Z(n998) );
  XNOR2_X1 U1086 ( .A(G4), .B(n998), .ZN(n1005) );
  XOR2_X1 U1087 ( .A(G1341), .B(G19), .Z(n1002) );
  XNOR2_X1 U1088 ( .A(G1956), .B(G20), .ZN(n1000) );
  XNOR2_X1 U1089 ( .A(G1981), .B(G6), .ZN(n999) );
  NOR2_X1 U1090 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  NAND2_X1 U1091 ( .A1(n1002), .A2(n1001), .ZN(n1003) );
  XOR2_X1 U1092 ( .A(KEYINPUT123), .B(n1003), .Z(n1004) );
  NOR2_X1 U1093 ( .A1(n1005), .A2(n1004), .ZN(n1006) );
  XOR2_X1 U1094 ( .A(KEYINPUT60), .B(n1006), .Z(n1008) );
  XNOR2_X1 U1095 ( .A(G1966), .B(G21), .ZN(n1007) );
  NOR2_X1 U1096 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  XNOR2_X1 U1097 ( .A(n1009), .B(KEYINPUT124), .ZN(n1013) );
  XNOR2_X1 U1098 ( .A(G5), .B(KEYINPUT122), .ZN(n1011) );
  XNOR2_X1 U1099 ( .A(n1011), .B(n1010), .ZN(n1012) );
  NAND2_X1 U1100 ( .A1(n1013), .A2(n1012), .ZN(n1021) );
  XNOR2_X1 U1101 ( .A(G1976), .B(G23), .ZN(n1015) );
  XNOR2_X1 U1102 ( .A(G1986), .B(G24), .ZN(n1014) );
  NOR2_X1 U1103 ( .A1(n1015), .A2(n1014), .ZN(n1018) );
  XNOR2_X1 U1104 ( .A(G1971), .B(KEYINPUT125), .ZN(n1016) );
  XNOR2_X1 U1105 ( .A(n1016), .B(G22), .ZN(n1017) );
  NAND2_X1 U1106 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  XNOR2_X1 U1107 ( .A(KEYINPUT58), .B(n1019), .ZN(n1020) );
  NOR2_X1 U1108 ( .A1(n1021), .A2(n1020), .ZN(n1022) );
  XNOR2_X1 U1109 ( .A(KEYINPUT61), .B(n1022), .ZN(n1023) );
  NAND2_X1 U1110 ( .A1(n1024), .A2(n1023), .ZN(n1025) );
  NAND2_X1 U1111 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1112 ( .A(n1027), .B(KEYINPUT126), .ZN(n1028) );
  NOR2_X1 U1113 ( .A1(n1029), .A2(n1028), .ZN(n1030) );
  XOR2_X1 U1114 ( .A(n1030), .B(KEYINPUT62), .Z(n1031) );
  XNOR2_X1 U1115 ( .A(KEYINPUT127), .B(n1031), .ZN(G311) );
  INV_X1 U1116 ( .A(G311), .ZN(G150) );
endmodule

