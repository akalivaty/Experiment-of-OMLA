//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 1 1 0 1 0 1 1 1 1 1 0 0 1 1 1 0 1 1 0 0 1 0 0 0 1 0 1 0 0 1 0 1 0 0 1 1 1 0 1 0 0 1 1 1 0 0 0 1 0 0 0 1 0 0 0 1 1 0 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:22 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n230, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1225, new_n1226, new_n1227, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1233, new_n1234, new_n1235, new_n1236,
    new_n1237, new_n1239, new_n1240, new_n1241, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1299,
    new_n1300, new_n1301, new_n1302, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309;
  INV_X1    g0000(.A(G50), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  NOR2_X1   g0004(.A1(new_n204), .A2(G77), .ZN(G353));
  OAI21_X1  g0005(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0006(.A(G1), .ZN(new_n207));
  INV_X1    g0007(.A(G20), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  INV_X1    g0009(.A(new_n209), .ZN(new_n210));
  NOR2_X1   g0010(.A1(new_n210), .A2(G13), .ZN(new_n211));
  OAI211_X1 g0011(.A(new_n211), .B(G250), .C1(G257), .C2(G264), .ZN(new_n212));
  XOR2_X1   g0012(.A(KEYINPUT64), .B(KEYINPUT0), .Z(new_n213));
  XNOR2_X1  g0013(.A(new_n212), .B(new_n213), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n202), .A2(new_n203), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n215), .A2(G50), .ZN(new_n216));
  NAND2_X1  g0016(.A1(G1), .A2(G13), .ZN(new_n217));
  OR3_X1    g0017(.A1(new_n216), .A2(new_n208), .A3(new_n217), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G68), .A2(G238), .B1(G77), .B2(G244), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n220));
  NAND2_X1  g0020(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  XOR2_X1   g0021(.A(new_n221), .B(KEYINPUT65), .Z(new_n222));
  AOI22_X1  g0022(.A1(G58), .A2(G232), .B1(G107), .B2(G264), .ZN(new_n223));
  XNOR2_X1  g0023(.A(new_n223), .B(KEYINPUT66), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G87), .A2(G250), .B1(G97), .B2(G257), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n210), .B1(new_n222), .B2(new_n226), .ZN(new_n227));
  OAI211_X1 g0027(.A(new_n214), .B(new_n218), .C1(new_n227), .C2(KEYINPUT1), .ZN(new_n228));
  AOI21_X1  g0028(.A(new_n228), .B1(KEYINPUT1), .B2(new_n227), .ZN(G361));
  XNOR2_X1  g0029(.A(G238), .B(G244), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(G232), .ZN(new_n231));
  XNOR2_X1  g0031(.A(KEYINPUT2), .B(G226), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(G264), .B(G270), .Z(new_n234));
  XNOR2_X1  g0034(.A(G250), .B(G257), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n233), .B(new_n236), .ZN(G358));
  XNOR2_X1  g0037(.A(G87), .B(G97), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(KEYINPUT67), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G107), .B(G116), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(G58), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G68), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(new_n241), .B(new_n244), .Z(G351));
  NAND3_X1  g0045(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(new_n217), .ZN(new_n247));
  INV_X1    g0047(.A(new_n247), .ZN(new_n248));
  XNOR2_X1  g0048(.A(KEYINPUT15), .B(G87), .ZN(new_n249));
  INV_X1    g0049(.A(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  OAI21_X1  g0051(.A(KEYINPUT68), .B1(new_n251), .B2(G20), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT68), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(new_n208), .A3(G33), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n252), .A2(new_n254), .ZN(new_n255));
  AOI22_X1  g0055(.A1(new_n250), .A2(new_n255), .B1(G20), .B2(G77), .ZN(new_n256));
  XNOR2_X1  g0056(.A(KEYINPUT8), .B(G58), .ZN(new_n257));
  INV_X1    g0057(.A(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(KEYINPUT70), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n259), .A2(new_n208), .A3(new_n251), .ZN(new_n260));
  OAI21_X1  g0060(.A(KEYINPUT70), .B1(G20), .B2(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n258), .A2(new_n262), .ZN(new_n263));
  AOI21_X1  g0063(.A(new_n248), .B1(new_n256), .B2(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(G13), .ZN(new_n265));
  NOR3_X1   g0065(.A1(new_n265), .A2(new_n208), .A3(G1), .ZN(new_n266));
  NOR2_X1   g0066(.A1(new_n266), .A2(new_n247), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n208), .A2(G1), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  NAND3_X1  g0069(.A1(new_n267), .A2(G77), .A3(new_n269), .ZN(new_n270));
  INV_X1    g0070(.A(new_n266), .ZN(new_n271));
  OAI21_X1  g0071(.A(new_n270), .B1(G77), .B2(new_n271), .ZN(new_n272));
  NOR2_X1   g0072(.A1(new_n264), .A2(new_n272), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n217), .B1(G33), .B2(G41), .ZN(new_n274));
  INV_X1    g0074(.A(G274), .ZN(new_n275));
  OAI21_X1  g0075(.A(new_n207), .B1(G41), .B2(G45), .ZN(new_n276));
  NOR3_X1   g0076(.A1(new_n274), .A2(new_n275), .A3(new_n276), .ZN(new_n277));
  INV_X1    g0077(.A(G41), .ZN(new_n278));
  OAI211_X1 g0078(.A(G1), .B(G13), .C1(new_n251), .C2(new_n278), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n279), .A2(new_n276), .ZN(new_n280));
  INV_X1    g0080(.A(new_n280), .ZN(new_n281));
  AOI21_X1  g0081(.A(new_n277), .B1(G244), .B2(new_n281), .ZN(new_n282));
  AND2_X1   g0082(.A1(KEYINPUT3), .A2(G33), .ZN(new_n283));
  NOR2_X1   g0083(.A1(KEYINPUT3), .A2(G33), .ZN(new_n284));
  NOR2_X1   g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g0085(.A(G1698), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  AOI22_X1  g0087(.A1(new_n287), .A2(G238), .B1(G107), .B2(new_n285), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT3), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(new_n251), .ZN(new_n290));
  NAND2_X1  g0090(.A1(KEYINPUT3), .A2(G33), .ZN(new_n291));
  NAND2_X1  g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  NAND3_X1  g0092(.A1(new_n292), .A2(G232), .A3(new_n286), .ZN(new_n293));
  AND2_X1   g0093(.A1(new_n288), .A2(new_n293), .ZN(new_n294));
  OAI21_X1  g0094(.A(new_n282), .B1(new_n294), .B2(new_n279), .ZN(new_n295));
  INV_X1    g0095(.A(G169), .ZN(new_n296));
  AOI21_X1  g0096(.A(new_n273), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(G179), .B2(new_n295), .ZN(new_n298));
  NAND2_X1  g0098(.A1(new_n295), .A2(G200), .ZN(new_n299));
  INV_X1    g0099(.A(G190), .ZN(new_n300));
  OAI211_X1 g0100(.A(new_n299), .B(new_n273), .C1(new_n300), .C2(new_n295), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n298), .A2(new_n301), .ZN(new_n302));
  XNOR2_X1  g0102(.A(new_n302), .B(KEYINPUT72), .ZN(new_n303));
  OAI21_X1  g0103(.A(KEYINPUT75), .B1(new_n283), .B2(new_n284), .ZN(new_n304));
  INV_X1    g0104(.A(KEYINPUT75), .ZN(new_n305));
  NAND3_X1  g0105(.A1(new_n290), .A2(new_n305), .A3(new_n291), .ZN(new_n306));
  NAND3_X1  g0106(.A1(new_n304), .A2(new_n306), .A3(new_n208), .ZN(new_n307));
  INV_X1    g0107(.A(KEYINPUT7), .ZN(new_n308));
  AND2_X1   g0108(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND4_X1  g0109(.A1(new_n290), .A2(KEYINPUT7), .A3(new_n208), .A4(new_n291), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n310), .A2(KEYINPUT76), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT76), .ZN(new_n312));
  NAND4_X1  g0112(.A1(new_n285), .A2(new_n312), .A3(KEYINPUT7), .A4(new_n208), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n311), .A2(new_n313), .ZN(new_n314));
  OAI21_X1  g0114(.A(G68), .B1(new_n309), .B2(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n262), .A2(G159), .ZN(new_n316));
  NAND2_X1  g0116(.A1(G58), .A2(G68), .ZN(new_n317));
  AOI21_X1  g0117(.A(new_n208), .B1(new_n215), .B2(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n319), .A3(KEYINPUT77), .ZN(new_n320));
  INV_X1    g0120(.A(KEYINPUT77), .ZN(new_n321));
  INV_X1    g0121(.A(G159), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n260), .B2(new_n261), .ZN(new_n323));
  OAI21_X1  g0123(.A(new_n321), .B1(new_n323), .B2(new_n318), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n320), .A2(KEYINPUT78), .A3(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(KEYINPUT78), .B1(new_n320), .B2(new_n324), .ZN(new_n327));
  OAI211_X1 g0127(.A(new_n315), .B(KEYINPUT16), .C1(new_n326), .C2(new_n327), .ZN(new_n328));
  XOR2_X1   g0128(.A(KEYINPUT79), .B(KEYINPUT16), .Z(new_n329));
  NAND3_X1  g0129(.A1(new_n290), .A2(new_n208), .A3(new_n291), .ZN(new_n330));
  NAND2_X1  g0130(.A1(new_n330), .A2(new_n308), .ZN(new_n331));
  NAND3_X1  g0131(.A1(new_n331), .A2(KEYINPUT80), .A3(new_n310), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT80), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n330), .A2(new_n333), .A3(new_n308), .ZN(new_n334));
  AND3_X1   g0134(.A1(new_n332), .A2(G68), .A3(new_n334), .ZN(new_n335));
  NAND2_X1  g0135(.A1(new_n320), .A2(new_n324), .ZN(new_n336));
  OAI21_X1  g0136(.A(new_n329), .B1(new_n335), .B2(new_n336), .ZN(new_n337));
  NAND3_X1  g0137(.A1(new_n328), .A2(new_n247), .A3(new_n337), .ZN(new_n338));
  NOR2_X1   g0138(.A1(new_n257), .A2(new_n268), .ZN(new_n339));
  AOI211_X1 g0139(.A(new_n247), .B(new_n266), .C1(new_n339), .C2(KEYINPUT81), .ZN(new_n340));
  NOR2_X1   g0140(.A1(new_n339), .A2(KEYINPUT81), .ZN(new_n341));
  INV_X1    g0141(.A(new_n341), .ZN(new_n342));
  AOI22_X1  g0142(.A1(new_n340), .A2(new_n342), .B1(new_n257), .B2(new_n266), .ZN(new_n343));
  AND2_X1   g0143(.A1(new_n338), .A2(new_n343), .ZN(new_n344));
  OR2_X1    g0144(.A1(new_n286), .A2(G226), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n292), .B(new_n345), .C1(G223), .C2(G1698), .ZN(new_n346));
  NAND2_X1  g0146(.A1(G33), .A2(G87), .ZN(new_n347));
  AOI21_X1  g0147(.A(new_n279), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(G232), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n279), .A2(G274), .ZN(new_n350));
  OAI22_X1  g0150(.A1(new_n349), .A2(new_n280), .B1(new_n350), .B2(new_n276), .ZN(new_n351));
  INV_X1    g0151(.A(G179), .ZN(new_n352));
  NOR3_X1   g0152(.A1(new_n348), .A2(new_n351), .A3(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  OAI21_X1  g0154(.A(G169), .B1(new_n348), .B2(new_n351), .ZN(new_n355));
  AOI21_X1  g0155(.A(KEYINPUT82), .B1(new_n354), .B2(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n354), .A2(KEYINPUT82), .A3(new_n355), .ZN(new_n358));
  NAND2_X1  g0158(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(KEYINPUT18), .B1(new_n344), .B2(new_n359), .ZN(new_n360));
  NOR2_X1   g0160(.A1(new_n348), .A2(new_n351), .ZN(new_n361));
  INV_X1    g0161(.A(G200), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n363), .B1(G190), .B2(new_n361), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n344), .A2(KEYINPUT17), .A3(new_n364), .ZN(new_n365));
  NAND3_X1  g0165(.A1(new_n338), .A2(new_n364), .A3(new_n343), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT17), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  INV_X1    g0168(.A(new_n358), .ZN(new_n369));
  NOR2_X1   g0169(.A1(new_n369), .A2(new_n356), .ZN(new_n370));
  NAND2_X1  g0170(.A1(new_n338), .A2(new_n343), .ZN(new_n371));
  INV_X1    g0171(.A(KEYINPUT18), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n370), .A2(new_n371), .A3(new_n372), .ZN(new_n373));
  NAND4_X1  g0173(.A1(new_n360), .A2(new_n365), .A3(new_n368), .A4(new_n373), .ZN(new_n374));
  XNOR2_X1  g0174(.A(new_n255), .B(KEYINPUT69), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n375), .A2(G77), .ZN(new_n376));
  AOI22_X1  g0176(.A1(new_n262), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n248), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g0178(.A1(new_n378), .A2(KEYINPUT11), .ZN(new_n379));
  NAND3_X1  g0179(.A1(new_n267), .A2(G68), .A3(new_n269), .ZN(new_n380));
  NOR3_X1   g0180(.A1(new_n271), .A2(KEYINPUT12), .A3(G68), .ZN(new_n381));
  INV_X1    g0181(.A(KEYINPUT12), .ZN(new_n382));
  AOI21_X1  g0182(.A(new_n382), .B1(new_n266), .B2(new_n203), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n380), .B1(new_n381), .B2(new_n383), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n384), .B1(new_n378), .B2(KEYINPUT11), .ZN(new_n385));
  NAND2_X1  g0185(.A1(new_n379), .A2(new_n385), .ZN(new_n386));
  NAND3_X1  g0186(.A1(new_n292), .A2(G232), .A3(G1698), .ZN(new_n387));
  NAND3_X1  g0187(.A1(new_n292), .A2(G226), .A3(new_n286), .ZN(new_n388));
  INV_X1    g0188(.A(G97), .ZN(new_n389));
  NOR2_X1   g0189(.A1(new_n251), .A2(new_n389), .ZN(new_n390));
  INV_X1    g0190(.A(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n387), .A2(new_n388), .A3(new_n391), .ZN(new_n392));
  NAND2_X1  g0192(.A1(new_n392), .A2(new_n274), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n277), .B1(G238), .B2(new_n281), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n395), .A2(KEYINPUT13), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT13), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n393), .A2(new_n397), .A3(new_n394), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n396), .A2(G179), .A3(new_n398), .ZN(new_n399));
  NAND2_X1  g0199(.A1(KEYINPUT74), .A2(G169), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n400), .B1(new_n396), .B2(new_n398), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT14), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n399), .B1(new_n401), .B2(new_n402), .ZN(new_n403));
  INV_X1    g0203(.A(new_n400), .ZN(new_n404));
  INV_X1    g0204(.A(new_n398), .ZN(new_n405));
  AOI21_X1  g0205(.A(new_n397), .B1(new_n393), .B2(new_n394), .ZN(new_n406));
  OAI211_X1 g0206(.A(new_n402), .B(new_n404), .C1(new_n405), .C2(new_n406), .ZN(new_n407));
  INV_X1    g0207(.A(new_n407), .ZN(new_n408));
  OAI21_X1  g0208(.A(new_n386), .B1(new_n403), .B2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  OAI21_X1  g0210(.A(G200), .B1(new_n405), .B2(new_n406), .ZN(new_n411));
  NAND3_X1  g0211(.A1(new_n396), .A2(G190), .A3(new_n398), .ZN(new_n412));
  NAND4_X1  g0212(.A1(new_n379), .A2(new_n411), .A3(new_n385), .A4(new_n412), .ZN(new_n413));
  INV_X1    g0213(.A(new_n413), .ZN(new_n414));
  NOR4_X1   g0214(.A1(new_n303), .A2(new_n374), .A3(new_n410), .A4(new_n414), .ZN(new_n415));
  AOI22_X1  g0215(.A1(new_n287), .A2(G223), .B1(G77), .B2(new_n285), .ZN(new_n416));
  NOR2_X1   g0216(.A1(new_n285), .A2(G1698), .ZN(new_n417));
  NAND2_X1  g0217(.A1(new_n417), .A2(G222), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n416), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g0219(.A1(new_n419), .A2(new_n274), .ZN(new_n420));
  AOI21_X1  g0220(.A(new_n277), .B1(G226), .B2(new_n281), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n420), .A2(new_n421), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n422), .A2(G200), .ZN(new_n423));
  NAND3_X1  g0223(.A1(new_n420), .A2(G190), .A3(new_n421), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  INV_X1    g0225(.A(new_n425), .ZN(new_n426));
  AOI22_X1  g0226(.A1(new_n375), .A2(new_n258), .B1(G150), .B2(new_n262), .ZN(new_n427));
  INV_X1    g0227(.A(KEYINPUT71), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n427), .A2(new_n428), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n204), .A2(G20), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  NOR2_X1   g0231(.A1(new_n427), .A2(new_n428), .ZN(new_n432));
  OAI21_X1  g0232(.A(new_n247), .B1(new_n431), .B2(new_n432), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT9), .ZN(new_n434));
  NOR2_X1   g0234(.A1(new_n268), .A2(new_n201), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n267), .A2(new_n435), .B1(new_n201), .B2(new_n266), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n436), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n434), .B1(new_n433), .B2(new_n436), .ZN(new_n439));
  OAI21_X1  g0239(.A(new_n426), .B1(new_n438), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n433), .A2(new_n436), .ZN(new_n441));
  NAND2_X1  g0241(.A1(new_n441), .A2(KEYINPUT9), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(new_n437), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT10), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT73), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n423), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g0246(.A1(new_n422), .A2(KEYINPUT73), .A3(G200), .ZN(new_n447));
  AND4_X1   g0247(.A1(new_n444), .A2(new_n446), .A3(new_n447), .A4(new_n424), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n440), .A2(KEYINPUT10), .B1(new_n443), .B2(new_n448), .ZN(new_n449));
  NOR2_X1   g0249(.A1(new_n422), .A2(G179), .ZN(new_n450));
  AOI21_X1  g0250(.A(new_n450), .B1(new_n296), .B2(new_n422), .ZN(new_n451));
  NAND2_X1  g0251(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n452), .ZN(new_n453));
  NOR2_X1   g0253(.A1(new_n449), .A2(new_n453), .ZN(new_n454));
  AND2_X1   g0254(.A1(new_n415), .A2(new_n454), .ZN(new_n455));
  NOR2_X1   g0255(.A1(new_n271), .A2(G97), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n207), .A2(G33), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n267), .A2(new_n457), .ZN(new_n458));
  INV_X1    g0258(.A(new_n458), .ZN(new_n459));
  AOI21_X1  g0259(.A(new_n456), .B1(new_n459), .B2(G97), .ZN(new_n460));
  INV_X1    g0260(.A(KEYINPUT83), .ZN(new_n461));
  NAND3_X1  g0261(.A1(new_n332), .A2(G107), .A3(new_n334), .ZN(new_n462));
  INV_X1    g0262(.A(KEYINPUT6), .ZN(new_n463));
  INV_X1    g0263(.A(G107), .ZN(new_n464));
  NOR2_X1   g0264(.A1(new_n389), .A2(new_n464), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n463), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n464), .A2(KEYINPUT6), .A3(G97), .ZN(new_n468));
  NAND2_X1  g0268(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  AOI22_X1  g0269(.A1(new_n469), .A2(G20), .B1(G77), .B2(new_n262), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n462), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n461), .B1(new_n471), .B2(new_n247), .ZN(new_n472));
  AOI211_X1 g0272(.A(KEYINPUT83), .B(new_n248), .C1(new_n462), .C2(new_n470), .ZN(new_n473));
  OAI21_X1  g0273(.A(new_n460), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n207), .A2(G45), .ZN(new_n475));
  INV_X1    g0275(.A(new_n475), .ZN(new_n476));
  XNOR2_X1  g0276(.A(KEYINPUT5), .B(G41), .ZN(new_n477));
  AOI21_X1  g0277(.A(new_n274), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(G257), .ZN(new_n479));
  AND2_X1   g0279(.A1(new_n477), .A2(new_n476), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n274), .A2(new_n275), .ZN(new_n481));
  NAND2_X1  g0281(.A1(new_n480), .A2(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n479), .A2(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n417), .A2(KEYINPUT4), .A3(G244), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n292), .A2(G244), .A3(new_n286), .ZN(new_n485));
  INV_X1    g0285(.A(KEYINPUT4), .ZN(new_n486));
  NAND2_X1  g0286(.A1(new_n485), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(G33), .A2(G283), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n292), .A2(G250), .A3(G1698), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n484), .A2(new_n487), .A3(new_n488), .A4(new_n489), .ZN(new_n490));
  AOI21_X1  g0290(.A(new_n483), .B1(new_n490), .B2(new_n274), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n491), .A2(new_n362), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n488), .B(new_n489), .C1(new_n485), .C2(new_n486), .ZN(new_n493));
  AOI21_X1  g0293(.A(KEYINPUT4), .B1(new_n417), .B2(G244), .ZN(new_n494));
  OAI21_X1  g0294(.A(new_n274), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  AND2_X1   g0295(.A1(new_n479), .A2(new_n482), .ZN(new_n496));
  NAND2_X1  g0296(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n497), .A2(new_n300), .ZN(new_n498));
  NOR3_X1   g0298(.A1(new_n474), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(KEYINPUT84), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n474), .A2(new_n500), .ZN(new_n501));
  OAI211_X1 g0301(.A(KEYINPUT84), .B(new_n460), .C1(new_n472), .C2(new_n473), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n501), .A2(new_n502), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n491), .A2(G179), .ZN(new_n504));
  NAND2_X1  g0304(.A1(new_n497), .A2(G169), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n499), .B1(new_n503), .B2(new_n506), .ZN(new_n507));
  NAND3_X1  g0307(.A1(new_n292), .A2(G257), .A3(G1698), .ZN(new_n508));
  NAND2_X1  g0308(.A1(G33), .A2(G294), .ZN(new_n509));
  OAI211_X1 g0309(.A(G250), .B(new_n286), .C1(new_n283), .C2(new_n284), .ZN(new_n510));
  NAND3_X1  g0310(.A1(new_n508), .A2(new_n509), .A3(new_n510), .ZN(new_n511));
  AOI22_X1  g0311(.A1(new_n511), .A2(new_n274), .B1(G264), .B2(new_n478), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n512), .A2(new_n482), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n296), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n512), .A2(new_n352), .A3(new_n482), .ZN(new_n515));
  NAND3_X1  g0315(.A1(new_n292), .A2(new_n208), .A3(G87), .ZN(new_n516));
  NOR2_X1   g0316(.A1(KEYINPUT87), .A2(KEYINPUT22), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  XOR2_X1   g0318(.A(KEYINPUT87), .B(KEYINPUT22), .Z(new_n519));
  NAND4_X1  g0319(.A1(new_n519), .A2(new_n208), .A3(G87), .A4(new_n292), .ZN(new_n520));
  INV_X1    g0320(.A(G116), .ZN(new_n521));
  NOR3_X1   g0321(.A1(new_n251), .A2(new_n521), .A3(G20), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT88), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n523), .B1(new_n208), .B2(G107), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n524), .A2(KEYINPUT23), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT23), .ZN(new_n526));
  OAI211_X1 g0326(.A(new_n523), .B(new_n526), .C1(new_n208), .C2(G107), .ZN(new_n527));
  AOI21_X1  g0327(.A(new_n522), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND3_X1  g0328(.A1(new_n518), .A2(new_n520), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g0329(.A1(new_n529), .A2(KEYINPUT24), .ZN(new_n530));
  INV_X1    g0330(.A(KEYINPUT24), .ZN(new_n531));
  NAND4_X1  g0331(.A1(new_n518), .A2(new_n528), .A3(new_n520), .A4(new_n531), .ZN(new_n532));
  AOI21_X1  g0332(.A(new_n248), .B1(new_n530), .B2(new_n532), .ZN(new_n533));
  AND3_X1   g0333(.A1(new_n266), .A2(KEYINPUT25), .A3(new_n464), .ZN(new_n534));
  AOI21_X1  g0334(.A(KEYINPUT25), .B1(new_n266), .B2(new_n464), .ZN(new_n535));
  OAI22_X1  g0335(.A1(new_n458), .A2(new_n464), .B1(new_n534), .B2(new_n535), .ZN(new_n536));
  OAI211_X1 g0336(.A(new_n514), .B(new_n515), .C1(new_n533), .C2(new_n536), .ZN(new_n537));
  NOR2_X1   g0337(.A1(new_n533), .A2(new_n536), .ZN(new_n538));
  AND3_X1   g0338(.A1(new_n512), .A2(G190), .A3(new_n482), .ZN(new_n539));
  AOI21_X1  g0339(.A(new_n362), .B1(new_n512), .B2(new_n482), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n538), .A2(new_n541), .A3(KEYINPUT89), .ZN(new_n542));
  AOI21_X1  g0342(.A(KEYINPUT89), .B1(new_n538), .B2(new_n541), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n537), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n292), .A2(G238), .A3(new_n286), .ZN(new_n545));
  NAND3_X1  g0345(.A1(new_n292), .A2(G244), .A3(G1698), .ZN(new_n546));
  NAND2_X1  g0346(.A1(G33), .A2(G116), .ZN(new_n547));
  NAND3_X1  g0347(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n548), .A2(new_n274), .ZN(new_n549));
  NAND2_X1  g0349(.A1(new_n475), .A2(G250), .ZN(new_n550));
  OAI21_X1  g0350(.A(KEYINPUT85), .B1(new_n274), .B2(new_n550), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n279), .A2(G274), .A3(new_n476), .ZN(new_n552));
  INV_X1    g0352(.A(KEYINPUT85), .ZN(new_n553));
  NAND4_X1  g0353(.A1(new_n279), .A2(new_n553), .A3(G250), .A4(new_n475), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n551), .A2(new_n552), .A3(new_n554), .ZN(new_n555));
  INV_X1    g0355(.A(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n549), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n557), .A2(G200), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n292), .A2(new_n208), .A3(G68), .ZN(new_n559));
  AOI21_X1  g0359(.A(new_n389), .B1(new_n252), .B2(new_n254), .ZN(new_n560));
  XNOR2_X1  g0360(.A(KEYINPUT86), .B(KEYINPUT19), .ZN(new_n561));
  AOI21_X1  g0361(.A(G20), .B1(new_n561), .B2(new_n390), .ZN(new_n562));
  NOR3_X1   g0362(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n563));
  OAI221_X1 g0363(.A(new_n559), .B1(new_n560), .B2(new_n561), .C1(new_n562), .C2(new_n563), .ZN(new_n564));
  AOI22_X1  g0364(.A1(new_n564), .A2(new_n247), .B1(new_n266), .B2(new_n249), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n459), .A2(G87), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n549), .A2(new_n556), .A3(G190), .ZN(new_n567));
  NAND4_X1  g0367(.A1(new_n558), .A2(new_n565), .A3(new_n566), .A4(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n557), .A2(new_n296), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n555), .B1(new_n274), .B2(new_n548), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n352), .ZN(new_n571));
  NOR2_X1   g0371(.A1(new_n562), .A2(new_n563), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n559), .B1(new_n560), .B2(new_n561), .ZN(new_n573));
  OAI21_X1  g0373(.A(new_n247), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n459), .A2(new_n250), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n249), .A2(new_n266), .ZN(new_n576));
  NAND3_X1  g0376(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n569), .A2(new_n571), .A3(new_n577), .ZN(new_n578));
  NAND2_X1  g0378(.A1(new_n568), .A2(new_n578), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  NAND3_X1  g0380(.A1(new_n292), .A2(G264), .A3(G1698), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n292), .A2(G257), .A3(new_n286), .ZN(new_n582));
  NAND2_X1  g0382(.A1(new_n285), .A2(G303), .ZN(new_n583));
  NAND3_X1  g0383(.A1(new_n581), .A2(new_n582), .A3(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n584), .A2(new_n274), .ZN(new_n585));
  AOI22_X1  g0385(.A1(new_n478), .A2(G270), .B1(new_n480), .B2(new_n481), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n267), .A2(G116), .A3(new_n457), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n266), .A2(new_n521), .ZN(new_n589));
  AOI22_X1  g0389(.A1(new_n246), .A2(new_n217), .B1(G20), .B2(new_n521), .ZN(new_n590));
  OAI211_X1 g0390(.A(new_n488), .B(new_n208), .C1(G33), .C2(new_n389), .ZN(new_n591));
  AND3_X1   g0391(.A1(new_n590), .A2(KEYINPUT20), .A3(new_n591), .ZN(new_n592));
  AOI21_X1  g0392(.A(KEYINPUT20), .B1(new_n590), .B2(new_n591), .ZN(new_n593));
  OAI211_X1 g0393(.A(new_n588), .B(new_n589), .C1(new_n592), .C2(new_n593), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n587), .A2(G169), .A3(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT21), .ZN(new_n596));
  NAND2_X1  g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n594), .A2(G179), .A3(new_n585), .A4(new_n586), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n587), .A2(KEYINPUT21), .A3(G169), .A4(new_n594), .ZN(new_n599));
  AND3_X1   g0399(.A1(new_n597), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  AOI21_X1  g0400(.A(new_n594), .B1(new_n587), .B2(G200), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n601), .B1(new_n300), .B2(new_n587), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n580), .A2(new_n600), .A3(new_n602), .ZN(new_n603));
  NOR2_X1   g0403(.A1(new_n544), .A2(new_n603), .ZN(new_n604));
  AND3_X1   g0404(.A1(new_n455), .A2(new_n507), .A3(new_n604), .ZN(G372));
  OAI21_X1  g0405(.A(new_n409), .B1(new_n414), .B2(new_n298), .ZN(new_n606));
  NAND3_X1  g0406(.A1(new_n606), .A2(new_n368), .A3(new_n365), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n354), .A2(new_n355), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n371), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g0409(.A1(new_n609), .A2(KEYINPUT18), .ZN(new_n610));
  NAND3_X1  g0410(.A1(new_n371), .A2(new_n372), .A3(new_n608), .ZN(new_n611));
  AND2_X1   g0411(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n607), .A2(new_n612), .ZN(new_n613));
  OAI21_X1  g0413(.A(new_n448), .B1(new_n438), .B2(new_n439), .ZN(new_n614));
  AOI21_X1  g0414(.A(new_n425), .B1(new_n442), .B2(new_n437), .ZN(new_n615));
  OAI21_X1  g0415(.A(new_n614), .B1(new_n615), .B2(new_n444), .ZN(new_n616));
  AOI21_X1  g0416(.A(new_n453), .B1(new_n613), .B2(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n455), .ZN(new_n618));
  NAND3_X1  g0418(.A1(new_n574), .A2(new_n566), .A3(new_n576), .ZN(new_n619));
  NAND2_X1  g0419(.A1(new_n619), .A2(KEYINPUT91), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT91), .ZN(new_n621));
  NAND4_X1  g0421(.A1(new_n574), .A2(new_n566), .A3(new_n621), .A4(new_n576), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n620), .A2(new_n622), .ZN(new_n623));
  INV_X1    g0423(.A(new_n567), .ZN(new_n624));
  INV_X1    g0424(.A(KEYINPUT90), .ZN(new_n625));
  AND3_X1   g0425(.A1(new_n548), .A2(new_n625), .A3(new_n274), .ZN(new_n626));
  AOI21_X1  g0426(.A(new_n625), .B1(new_n548), .B2(new_n274), .ZN(new_n627));
  OAI21_X1  g0427(.A(new_n556), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n624), .B1(new_n628), .B2(G200), .ZN(new_n629));
  AND2_X1   g0429(.A1(new_n571), .A2(new_n577), .ZN(new_n630));
  NAND2_X1  g0430(.A1(new_n628), .A2(new_n296), .ZN(new_n631));
  AOI22_X1  g0431(.A1(new_n623), .A2(new_n629), .B1(new_n630), .B2(new_n631), .ZN(new_n632));
  AND2_X1   g0432(.A1(new_n599), .A2(new_n598), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n537), .A2(new_n633), .A3(new_n597), .ZN(new_n634));
  OAI211_X1 g0434(.A(new_n632), .B(new_n634), .C1(new_n542), .C2(new_n543), .ZN(new_n635));
  INV_X1    g0435(.A(new_n635), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n636), .A2(new_n507), .B1(new_n630), .B2(new_n631), .ZN(new_n637));
  AND2_X1   g0437(.A1(new_n474), .A2(new_n506), .ZN(new_n638));
  INV_X1    g0438(.A(KEYINPUT26), .ZN(new_n639));
  AND3_X1   g0439(.A1(new_n638), .A2(new_n632), .A3(new_n639), .ZN(new_n640));
  NAND2_X1  g0440(.A1(new_n471), .A2(new_n247), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n641), .A2(KEYINPUT83), .ZN(new_n642));
  NAND3_X1  g0442(.A1(new_n471), .A2(new_n461), .A3(new_n247), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  AOI21_X1  g0444(.A(KEYINPUT84), .B1(new_n644), .B2(new_n460), .ZN(new_n645));
  INV_X1    g0445(.A(new_n502), .ZN(new_n646));
  OAI211_X1 g0446(.A(new_n506), .B(new_n580), .C1(new_n645), .C2(new_n646), .ZN(new_n647));
  AOI21_X1  g0447(.A(new_n640), .B1(KEYINPUT26), .B2(new_n647), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n637), .A2(new_n648), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(new_n617), .B1(new_n618), .B2(new_n650), .ZN(G369));
  NAND2_X1  g0451(.A1(new_n633), .A2(new_n597), .ZN(new_n652));
  NAND3_X1  g0452(.A1(new_n207), .A2(new_n208), .A3(G13), .ZN(new_n653));
  OR2_X1    g0453(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n654));
  NAND2_X1  g0454(.A1(new_n653), .A2(KEYINPUT27), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n654), .A2(G213), .A3(new_n655), .ZN(new_n656));
  INV_X1    g0456(.A(G343), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  AND2_X1   g0458(.A1(new_n594), .A2(new_n658), .ZN(new_n659));
  NAND2_X1  g0459(.A1(new_n652), .A2(new_n659), .ZN(new_n660));
  NAND2_X1  g0460(.A1(new_n600), .A2(new_n602), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n660), .B1(new_n661), .B2(new_n659), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n662), .A2(G330), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT92), .Z(new_n664));
  INV_X1    g0464(.A(new_n658), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n537), .A2(new_n665), .ZN(new_n666));
  XNOR2_X1  g0466(.A(new_n666), .B(KEYINPUT93), .ZN(new_n667));
  OAI221_X1 g0467(.A(new_n537), .B1(new_n538), .B2(new_n665), .C1(new_n542), .C2(new_n543), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  NOR2_X1   g0470(.A1(new_n600), .A2(new_n658), .ZN(new_n671));
  INV_X1    g0471(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n667), .B2(new_n668), .ZN(new_n673));
  INV_X1    g0473(.A(new_n537), .ZN(new_n674));
  AOI21_X1  g0474(.A(new_n673), .B1(new_n674), .B2(new_n665), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n670), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g0476(.A(new_n676), .B(KEYINPUT94), .Z(G399));
  INV_X1    g0477(.A(new_n211), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n678), .A2(G41), .ZN(new_n679));
  INV_X1    g0479(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n563), .A2(new_n521), .ZN(new_n681));
  XOR2_X1   g0481(.A(new_n681), .B(KEYINPUT95), .Z(new_n682));
  NAND3_X1  g0482(.A1(new_n680), .A2(G1), .A3(new_n682), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n683), .B1(new_n216), .B2(new_n680), .ZN(new_n684));
  XNOR2_X1  g0484(.A(new_n684), .B(KEYINPUT28), .ZN(new_n685));
  INV_X1    g0485(.A(G330), .ZN(new_n686));
  AND2_X1   g0486(.A1(new_n570), .A2(new_n512), .ZN(new_n687));
  INV_X1    g0487(.A(KEYINPUT96), .ZN(new_n688));
  OAI21_X1  g0488(.A(new_n688), .B1(new_n587), .B2(new_n352), .ZN(new_n689));
  NAND4_X1  g0489(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT96), .A4(G179), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n687), .A2(new_n689), .A3(new_n491), .A4(new_n690), .ZN(new_n691));
  INV_X1    g0491(.A(KEYINPUT30), .ZN(new_n692));
  NAND2_X1  g0492(.A1(new_n692), .A2(KEYINPUT97), .ZN(new_n693));
  INV_X1    g0493(.A(new_n693), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g0495(.A1(new_n491), .A2(new_n512), .A3(new_n570), .ZN(new_n696));
  NAND4_X1  g0496(.A1(new_n696), .A2(new_n693), .A3(new_n690), .A4(new_n689), .ZN(new_n697));
  AOI21_X1  g0497(.A(G179), .B1(new_n585), .B2(new_n586), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n628), .A2(new_n497), .A3(new_n513), .A4(new_n698), .ZN(new_n699));
  NAND3_X1  g0499(.A1(new_n695), .A2(new_n697), .A3(new_n699), .ZN(new_n700));
  AND3_X1   g0500(.A1(new_n700), .A2(KEYINPUT31), .A3(new_n658), .ZN(new_n701));
  AOI21_X1  g0501(.A(KEYINPUT31), .B1(new_n700), .B2(new_n658), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n604), .A2(new_n507), .A3(new_n665), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n686), .B1(new_n703), .B2(new_n704), .ZN(new_n705));
  AOI21_X1  g0505(.A(new_n658), .B1(new_n637), .B2(new_n648), .ZN(new_n706));
  OR2_X1    g0506(.A1(new_n706), .A2(KEYINPUT29), .ZN(new_n707));
  AND2_X1   g0507(.A1(new_n504), .A2(new_n505), .ZN(new_n708));
  AOI211_X1 g0508(.A(new_n708), .B(new_n579), .C1(new_n501), .C2(new_n502), .ZN(new_n709));
  OAI21_X1  g0509(.A(KEYINPUT98), .B1(new_n709), .B2(KEYINPUT26), .ZN(new_n710));
  NAND3_X1  g0510(.A1(new_n638), .A2(new_n632), .A3(KEYINPUT26), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT98), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n647), .A2(new_n712), .A3(new_n639), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n711), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g0514(.A(new_n658), .B1(new_n714), .B2(new_n637), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(KEYINPUT29), .ZN(new_n716));
  AOI21_X1  g0516(.A(new_n705), .B1(new_n707), .B2(new_n716), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n685), .B1(new_n717), .B2(G1), .ZN(G364));
  NOR2_X1   g0518(.A1(new_n265), .A2(G20), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n207), .B1(new_n719), .B2(G45), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n679), .A2(new_n721), .ZN(new_n722));
  INV_X1    g0522(.A(new_n722), .ZN(new_n723));
  OAI21_X1  g0523(.A(new_n723), .B1(new_n662), .B2(G330), .ZN(new_n724));
  NOR2_X1   g0524(.A1(G13), .A2(G33), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g0526(.A1(new_n726), .A2(G20), .ZN(new_n727));
  INV_X1    g0527(.A(new_n727), .ZN(new_n728));
  NOR2_X1   g0528(.A1(new_n662), .A2(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n217), .B1(G20), .B2(new_n296), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n727), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT100), .Z(new_n732));
  NOR2_X1   g0532(.A1(new_n678), .A2(new_n285), .ZN(new_n733));
  AOI22_X1  g0533(.A1(new_n733), .A2(G355), .B1(new_n521), .B2(new_n678), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n304), .A2(new_n306), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n678), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g0536(.A(new_n736), .B1(G45), .B2(new_n216), .ZN(new_n737));
  INV_X1    g0537(.A(G45), .ZN(new_n738));
  NOR2_X1   g0538(.A1(new_n244), .A2(new_n738), .ZN(new_n739));
  OAI21_X1  g0539(.A(new_n734), .B1(new_n737), .B2(new_n739), .ZN(new_n740));
  AOI21_X1  g0540(.A(new_n732), .B1(new_n740), .B2(KEYINPUT99), .ZN(new_n741));
  OAI21_X1  g0541(.A(new_n741), .B1(KEYINPUT99), .B2(new_n740), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n208), .A2(G179), .ZN(new_n743));
  NOR2_X1   g0543(.A1(G190), .A2(G200), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(KEYINPUT32), .B1(new_n745), .B2(new_n322), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n208), .A2(new_n352), .ZN(new_n747));
  NAND2_X1  g0547(.A1(new_n747), .A2(G200), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n748), .A2(new_n300), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n748), .A2(G190), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  OAI221_X1 g0552(.A(new_n746), .B1(new_n750), .B2(new_n201), .C1(new_n203), .C2(new_n752), .ZN(new_n753));
  NOR3_X1   g0553(.A1(new_n300), .A2(G179), .A3(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(new_n208), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NAND3_X1  g0556(.A1(new_n743), .A2(G190), .A3(G200), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI22_X1  g0558(.A1(new_n756), .A2(G97), .B1(new_n758), .B2(G87), .ZN(new_n759));
  NAND3_X1  g0559(.A1(new_n743), .A2(new_n300), .A3(G200), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(G107), .ZN(new_n762));
  INV_X1    g0562(.A(new_n745), .ZN(new_n763));
  NAND2_X1  g0563(.A1(new_n763), .A2(G159), .ZN(new_n764));
  OAI211_X1 g0564(.A(new_n759), .B(new_n762), .C1(KEYINPUT32), .C2(new_n764), .ZN(new_n765));
  NAND2_X1  g0565(.A1(new_n747), .A2(new_n744), .ZN(new_n766));
  INV_X1    g0566(.A(G77), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n747), .A2(G190), .A3(new_n362), .ZN(new_n768));
  OAI221_X1 g0568(.A(new_n292), .B1(new_n766), .B2(new_n767), .C1(new_n202), .C2(new_n768), .ZN(new_n769));
  NOR3_X1   g0569(.A1(new_n753), .A2(new_n765), .A3(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(new_n768), .ZN(new_n771));
  AOI22_X1  g0571(.A1(new_n771), .A2(G322), .B1(new_n763), .B2(G329), .ZN(new_n772));
  INV_X1    g0572(.A(G311), .ZN(new_n773));
  OAI211_X1 g0573(.A(new_n772), .B(new_n285), .C1(new_n773), .C2(new_n766), .ZN(new_n774));
  INV_X1    g0574(.A(G317), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n776));
  OR2_X1    g0576(.A1(new_n775), .A2(KEYINPUT33), .ZN(new_n777));
  NAND3_X1  g0577(.A1(new_n751), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g0578(.A1(new_n749), .A2(G326), .ZN(new_n779));
  INV_X1    g0579(.A(G294), .ZN(new_n780));
  OAI211_X1 g0580(.A(new_n778), .B(new_n779), .C1(new_n780), .C2(new_n755), .ZN(new_n781));
  INV_X1    g0581(.A(G283), .ZN(new_n782));
  INV_X1    g0582(.A(G303), .ZN(new_n783));
  OAI22_X1  g0583(.A1(new_n782), .A2(new_n760), .B1(new_n757), .B2(new_n783), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n774), .A2(new_n781), .A3(new_n784), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n730), .B1(new_n770), .B2(new_n785), .ZN(new_n786));
  NAND3_X1  g0586(.A1(new_n742), .A2(new_n722), .A3(new_n786), .ZN(new_n787));
  OAI22_X1  g0587(.A1(new_n664), .A2(new_n724), .B1(new_n729), .B2(new_n787), .ZN(G396));
  NOR2_X1   g0588(.A1(new_n298), .A2(new_n658), .ZN(new_n789));
  OAI21_X1  g0589(.A(new_n301), .B1(new_n273), .B2(new_n665), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n789), .B1(new_n790), .B2(new_n298), .ZN(new_n791));
  OR2_X1    g0591(.A1(new_n706), .A2(new_n791), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n649), .A2(new_n665), .A3(new_n791), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  NAND2_X1  g0594(.A1(new_n703), .A2(new_n704), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n794), .B1(new_n686), .B2(new_n796), .ZN(new_n797));
  NAND3_X1  g0597(.A1(new_n792), .A2(new_n705), .A3(new_n793), .ZN(new_n798));
  NAND3_X1  g0598(.A1(new_n797), .A2(new_n723), .A3(new_n798), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n730), .A2(new_n725), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n723), .B1(new_n767), .B2(new_n800), .ZN(new_n801));
  INV_X1    g0601(.A(G87), .ZN(new_n802));
  OAI22_X1  g0602(.A1(new_n750), .A2(new_n783), .B1(new_n760), .B2(new_n802), .ZN(new_n803));
  AOI21_X1  g0603(.A(new_n803), .B1(G107), .B2(new_n758), .ZN(new_n804));
  OAI22_X1  g0604(.A1(new_n768), .A2(new_n780), .B1(new_n745), .B2(new_n773), .ZN(new_n805));
  INV_X1    g0605(.A(new_n766), .ZN(new_n806));
  AOI211_X1 g0606(.A(new_n292), .B(new_n805), .C1(G116), .C2(new_n806), .ZN(new_n807));
  AOI22_X1  g0607(.A1(G97), .A2(new_n756), .B1(new_n751), .B2(G283), .ZN(new_n808));
  NAND3_X1  g0608(.A1(new_n804), .A2(new_n807), .A3(new_n808), .ZN(new_n809));
  AOI22_X1  g0609(.A1(new_n771), .A2(G143), .B1(new_n806), .B2(G159), .ZN(new_n810));
  INV_X1    g0610(.A(G137), .ZN(new_n811));
  INV_X1    g0611(.A(G150), .ZN(new_n812));
  OAI221_X1 g0612(.A(new_n810), .B1(new_n750), .B2(new_n811), .C1(new_n812), .C2(new_n752), .ZN(new_n813));
  INV_X1    g0613(.A(KEYINPUT34), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  INV_X1    g0615(.A(new_n735), .ZN(new_n816));
  AOI21_X1  g0616(.A(new_n816), .B1(G132), .B2(new_n763), .ZN(new_n817));
  NOR2_X1   g0617(.A1(new_n757), .A2(new_n201), .ZN(new_n818));
  NOR2_X1   g0618(.A1(new_n760), .A2(new_n203), .ZN(new_n819));
  AOI211_X1 g0619(.A(new_n818), .B(new_n819), .C1(G58), .C2(new_n756), .ZN(new_n820));
  NAND3_X1  g0620(.A1(new_n815), .A2(new_n817), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n813), .A2(new_n814), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n809), .B1(new_n821), .B2(new_n822), .ZN(new_n823));
  INV_X1    g0623(.A(KEYINPUT101), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n730), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n823), .A2(new_n824), .ZN(new_n827));
  OAI221_X1 g0627(.A(new_n801), .B1(new_n826), .B2(new_n827), .C1(new_n791), .C2(new_n726), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n799), .A2(new_n828), .ZN(new_n829));
  XOR2_X1   g0629(.A(new_n829), .B(KEYINPUT102), .Z(new_n830));
  INV_X1    g0630(.A(new_n830), .ZN(G384));
  NOR2_X1   g0631(.A1(new_n719), .A2(new_n207), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n386), .A2(new_n658), .ZN(new_n833));
  NAND3_X1  g0633(.A1(new_n409), .A2(new_n413), .A3(new_n833), .ZN(new_n834));
  OAI211_X1 g0634(.A(new_n386), .B(new_n658), .C1(new_n403), .C2(new_n408), .ZN(new_n835));
  NAND2_X1  g0635(.A1(new_n834), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n836), .A2(new_n791), .ZN(new_n837));
  AOI21_X1  g0637(.A(new_n837), .B1(new_n704), .B2(new_n703), .ZN(new_n838));
  INV_X1    g0638(.A(new_n343), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT78), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n336), .A2(new_n840), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n307), .A2(new_n308), .ZN(new_n842));
  NAND3_X1  g0642(.A1(new_n842), .A2(new_n311), .A3(new_n313), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n841), .A2(new_n325), .B1(new_n843), .B2(G68), .ZN(new_n844));
  AOI21_X1  g0644(.A(new_n248), .B1(new_n844), .B2(KEYINPUT16), .ZN(new_n845));
  OAI21_X1  g0645(.A(new_n315), .B1(new_n326), .B2(new_n327), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(new_n329), .ZN(new_n847));
  AOI21_X1  g0647(.A(new_n839), .B1(new_n845), .B2(new_n847), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n366), .B1(new_n848), .B2(new_n656), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n845), .A2(new_n847), .ZN(new_n850));
  AOI22_X1  g0650(.A1(new_n850), .A2(new_n343), .B1(new_n355), .B2(new_n354), .ZN(new_n851));
  OAI21_X1  g0651(.A(KEYINPUT37), .B1(new_n849), .B2(new_n851), .ZN(new_n852));
  XOR2_X1   g0652(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n853));
  AOI21_X1  g0653(.A(new_n853), .B1(new_n370), .B2(new_n371), .ZN(new_n854));
  INV_X1    g0654(.A(new_n656), .ZN(new_n855));
  AOI21_X1  g0655(.A(KEYINPUT105), .B1(new_n371), .B2(new_n855), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT105), .ZN(new_n857));
  AOI211_X1 g0657(.A(new_n857), .B(new_n656), .C1(new_n338), .C2(new_n343), .ZN(new_n858));
  OAI211_X1 g0658(.A(new_n366), .B(new_n854), .C1(new_n856), .C2(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n852), .A2(new_n859), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n848), .A2(new_n656), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n374), .A2(new_n861), .ZN(new_n862));
  AND3_X1   g0662(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n863));
  AOI21_X1  g0663(.A(KEYINPUT38), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  OAI21_X1  g0664(.A(new_n838), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT40), .ZN(new_n866));
  AOI211_X1 g0666(.A(new_n866), .B(new_n837), .C1(new_n704), .C2(new_n703), .ZN(new_n867));
  NAND3_X1  g0667(.A1(new_n860), .A2(new_n862), .A3(KEYINPUT38), .ZN(new_n868));
  OAI211_X1 g0668(.A(new_n366), .B(new_n609), .C1(new_n856), .C2(new_n858), .ZN(new_n869));
  NAND2_X1  g0669(.A1(new_n869), .A2(new_n853), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n856), .A2(new_n858), .ZN(new_n871));
  NAND4_X1  g0671(.A1(new_n610), .A2(new_n365), .A3(new_n368), .A4(new_n611), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n870), .A2(new_n859), .B1(new_n871), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n868), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n874));
  AOI22_X1  g0674(.A1(new_n865), .A2(new_n866), .B1(new_n867), .B2(new_n874), .ZN(new_n875));
  XOR2_X1   g0675(.A(new_n875), .B(KEYINPUT107), .Z(new_n876));
  OR3_X1    g0676(.A1(new_n876), .A2(new_n618), .A3(new_n796), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n876), .B1(new_n618), .B2(new_n796), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n877), .A2(G330), .A3(new_n878), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n612), .A2(new_n855), .ZN(new_n880));
  INV_X1    g0680(.A(new_n836), .ZN(new_n881));
  XNOR2_X1  g0681(.A(new_n789), .B(KEYINPUT104), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  AOI21_X1  g0683(.A(new_n881), .B1(new_n793), .B2(new_n883), .ZN(new_n884));
  INV_X1    g0684(.A(new_n864), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n885), .A2(new_n868), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n880), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT39), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n874), .A2(new_n888), .ZN(new_n889));
  NOR2_X1   g0689(.A1(new_n409), .A2(new_n658), .ZN(new_n890));
  NAND3_X1  g0690(.A1(new_n885), .A2(KEYINPUT39), .A3(new_n868), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n889), .A2(new_n890), .A3(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n887), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n707), .A2(new_n455), .A3(new_n716), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n617), .ZN(new_n895));
  XNOR2_X1  g0695(.A(new_n893), .B(new_n895), .ZN(new_n896));
  AOI21_X1  g0696(.A(new_n832), .B1(new_n879), .B2(new_n896), .ZN(new_n897));
  OAI21_X1  g0697(.A(new_n897), .B1(new_n896), .B2(new_n879), .ZN(new_n898));
  NOR3_X1   g0698(.A1(new_n217), .A2(new_n208), .A3(new_n521), .ZN(new_n899));
  XOR2_X1   g0699(.A(new_n469), .B(KEYINPUT103), .Z(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT35), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g0703(.A(new_n903), .B1(new_n902), .B2(new_n901), .ZN(new_n904));
  XOR2_X1   g0704(.A(new_n904), .B(KEYINPUT36), .Z(new_n905));
  NAND2_X1  g0705(.A1(new_n317), .A2(G77), .ZN(new_n906));
  OAI22_X1  g0706(.A1(new_n216), .A2(new_n906), .B1(G50), .B2(new_n203), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n907), .A2(G1), .A3(new_n265), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n898), .A2(new_n905), .A3(new_n908), .ZN(G367));
  NAND2_X1  g0709(.A1(new_n474), .A2(new_n658), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n507), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n638), .A2(new_n658), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n673), .ZN(new_n914));
  XOR2_X1   g0714(.A(new_n914), .B(KEYINPUT42), .Z(new_n915));
  AOI22_X1  g0715(.A1(new_n913), .A2(new_n674), .B1(new_n506), .B2(new_n503), .ZN(new_n916));
  OR2_X1    g0716(.A1(new_n916), .A2(new_n658), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NAND3_X1  g0718(.A1(new_n620), .A2(new_n622), .A3(new_n658), .ZN(new_n919));
  NAND2_X1  g0719(.A1(new_n632), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g0720(.A1(new_n630), .A2(new_n631), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n920), .B1(new_n921), .B2(new_n919), .ZN(new_n922));
  XNOR2_X1  g0722(.A(KEYINPUT108), .B(KEYINPUT43), .ZN(new_n923));
  NOR2_X1   g0723(.A1(new_n922), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g0724(.A(new_n924), .B1(KEYINPUT43), .B2(new_n922), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n918), .A2(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT109), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n926), .A2(new_n927), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n915), .A2(new_n917), .A3(new_n924), .ZN(new_n929));
  NAND3_X1  g0729(.A1(new_n918), .A2(KEYINPUT109), .A3(new_n925), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n928), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  INV_X1    g0731(.A(new_n913), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n931), .B1(new_n670), .B2(new_n932), .ZN(new_n933));
  NOR2_X1   g0733(.A1(new_n670), .A2(new_n932), .ZN(new_n934));
  NAND4_X1  g0734(.A1(new_n928), .A2(new_n934), .A3(new_n929), .A4(new_n930), .ZN(new_n935));
  XOR2_X1   g0735(.A(new_n679), .B(KEYINPUT41), .Z(new_n936));
  NOR2_X1   g0736(.A1(new_n675), .A2(new_n913), .ZN(new_n937));
  XNOR2_X1  g0737(.A(new_n937), .B(KEYINPUT44), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n675), .A2(new_n913), .ZN(new_n939));
  INV_X1    g0739(.A(KEYINPUT45), .ZN(new_n940));
  XNOR2_X1  g0740(.A(new_n939), .B(new_n940), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n938), .A2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n670), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n942), .A2(new_n943), .ZN(new_n944));
  NAND3_X1  g0744(.A1(new_n667), .A2(new_n668), .A3(new_n672), .ZN(new_n945));
  INV_X1    g0745(.A(KEYINPUT110), .ZN(new_n946));
  NAND2_X1  g0746(.A1(new_n945), .A2(new_n946), .ZN(new_n947));
  NAND2_X1  g0747(.A1(new_n669), .A2(new_n671), .ZN(new_n948));
  XNOR2_X1  g0748(.A(new_n947), .B(new_n948), .ZN(new_n949));
  INV_X1    g0749(.A(KEYINPUT111), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n949), .A2(new_n950), .A3(new_n664), .ZN(new_n951));
  XNOR2_X1  g0751(.A(new_n664), .B(new_n950), .ZN(new_n952));
  OAI21_X1  g0752(.A(new_n951), .B1(new_n952), .B2(new_n949), .ZN(new_n953));
  NAND3_X1  g0753(.A1(new_n938), .A2(new_n670), .A3(new_n941), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n944), .A2(new_n717), .A3(new_n953), .A4(new_n954), .ZN(new_n955));
  AOI21_X1  g0755(.A(new_n936), .B1(new_n955), .B2(new_n717), .ZN(new_n956));
  OAI211_X1 g0756(.A(new_n933), .B(new_n935), .C1(new_n956), .C2(new_n721), .ZN(new_n957));
  INV_X1    g0757(.A(new_n732), .ZN(new_n958));
  OAI21_X1  g0758(.A(new_n958), .B1(new_n211), .B2(new_n249), .ZN(new_n959));
  NOR3_X1   g0759(.A1(new_n236), .A2(new_n678), .A3(new_n735), .ZN(new_n960));
  OAI21_X1  g0760(.A(new_n722), .B1(new_n959), .B2(new_n960), .ZN(new_n961));
  OAI22_X1  g0761(.A1(new_n768), .A2(new_n783), .B1(new_n745), .B2(new_n775), .ZN(new_n962));
  OAI21_X1  g0762(.A(new_n816), .B1(new_n389), .B2(new_n760), .ZN(new_n963));
  AOI211_X1 g0763(.A(new_n962), .B(new_n963), .C1(G283), .C2(new_n806), .ZN(new_n964));
  AOI21_X1  g0764(.A(KEYINPUT112), .B1(new_n758), .B2(G116), .ZN(new_n965));
  XNOR2_X1  g0765(.A(new_n965), .B(KEYINPUT46), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n780), .A2(new_n752), .B1(new_n750), .B2(new_n773), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G107), .B2(new_n756), .ZN(new_n968));
  NAND3_X1  g0768(.A1(new_n964), .A2(new_n966), .A3(new_n968), .ZN(new_n969));
  INV_X1    g0769(.A(KEYINPUT113), .ZN(new_n970));
  OR2_X1    g0770(.A1(new_n969), .A2(new_n970), .ZN(new_n971));
  NOR2_X1   g0771(.A1(new_n760), .A2(new_n767), .ZN(new_n972));
  NOR2_X1   g0772(.A1(new_n972), .A2(new_n285), .ZN(new_n973));
  XOR2_X1   g0773(.A(new_n973), .B(KEYINPUT114), .Z(new_n974));
  OAI22_X1  g0774(.A1(new_n766), .A2(new_n201), .B1(new_n745), .B2(new_n811), .ZN(new_n975));
  AOI21_X1  g0775(.A(new_n975), .B1(G150), .B2(new_n771), .ZN(new_n976));
  AOI22_X1  g0776(.A1(G143), .A2(new_n749), .B1(new_n751), .B2(G159), .ZN(new_n977));
  AOI22_X1  g0777(.A1(new_n756), .A2(G68), .B1(new_n758), .B2(G58), .ZN(new_n978));
  NAND4_X1  g0778(.A1(new_n974), .A2(new_n976), .A3(new_n977), .A4(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n969), .A2(new_n970), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n971), .A2(new_n979), .A3(new_n980), .ZN(new_n981));
  XNOR2_X1  g0781(.A(new_n981), .B(KEYINPUT47), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n961), .B1(new_n982), .B2(new_n730), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n728), .B2(new_n922), .ZN(new_n984));
  NAND2_X1  g0784(.A1(new_n957), .A2(new_n984), .ZN(G387));
  NAND3_X1  g0785(.A1(new_n667), .A2(new_n668), .A3(new_n727), .ZN(new_n986));
  OAI21_X1  g0786(.A(new_n736), .B1(new_n233), .B2(new_n738), .ZN(new_n987));
  INV_X1    g0787(.A(new_n733), .ZN(new_n988));
  OAI21_X1  g0788(.A(new_n987), .B1(new_n682), .B2(new_n988), .ZN(new_n989));
  OR3_X1    g0789(.A1(new_n257), .A2(KEYINPUT50), .A3(G50), .ZN(new_n990));
  OAI21_X1  g0790(.A(KEYINPUT50), .B1(new_n257), .B2(G50), .ZN(new_n991));
  AOI21_X1  g0791(.A(G45), .B1(G68), .B2(G77), .ZN(new_n992));
  NAND4_X1  g0792(.A1(new_n682), .A2(new_n990), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  AOI22_X1  g0793(.A1(new_n989), .A2(new_n993), .B1(new_n464), .B2(new_n678), .ZN(new_n994));
  OAI21_X1  g0794(.A(new_n722), .B1(new_n994), .B2(new_n732), .ZN(new_n995));
  NOR2_X1   g0795(.A1(new_n757), .A2(new_n767), .ZN(new_n996));
  OAI21_X1  g0796(.A(new_n735), .B1(new_n812), .B2(new_n745), .ZN(new_n997));
  AOI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(G97), .C2(new_n761), .ZN(new_n998));
  XOR2_X1   g0798(.A(new_n998), .B(KEYINPUT115), .Z(new_n999));
  NOR2_X1   g0799(.A1(new_n755), .A2(new_n249), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(new_n771), .A2(G50), .B1(new_n806), .B2(G68), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n1001), .B1(new_n257), .B2(new_n752), .ZN(new_n1002));
  AOI211_X1 g0802(.A(new_n1000), .B(new_n1002), .C1(G159), .C2(new_n749), .ZN(new_n1003));
  NAND2_X1  g0803(.A1(new_n999), .A2(new_n1003), .ZN(new_n1004));
  AOI22_X1  g0804(.A1(new_n771), .A2(G317), .B1(new_n806), .B2(G303), .ZN(new_n1005));
  NAND2_X1  g0805(.A1(new_n749), .A2(G322), .ZN(new_n1006));
  OAI211_X1 g0806(.A(new_n1005), .B(new_n1006), .C1(new_n773), .C2(new_n752), .ZN(new_n1007));
  INV_X1    g0807(.A(KEYINPUT48), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  OAI221_X1 g0809(.A(new_n1009), .B1(new_n782), .B2(new_n755), .C1(new_n780), .C2(new_n757), .ZN(new_n1010));
  NOR2_X1   g0810(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1011));
  NOR2_X1   g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n760), .A2(new_n521), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n735), .B(new_n1014), .C1(G326), .C2(new_n763), .ZN(new_n1015));
  NAND2_X1  g0815(.A1(new_n1013), .A2(new_n1015), .ZN(new_n1016));
  NOR2_X1   g0816(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n1004), .B1(new_n1016), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n995), .B1(new_n1018), .B2(new_n730), .ZN(new_n1019));
  AOI22_X1  g0819(.A1(new_n953), .A2(new_n721), .B1(new_n986), .B2(new_n1019), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n953), .A2(new_n717), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n679), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n953), .A2(new_n717), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1020), .B1(new_n1022), .B2(new_n1023), .ZN(G393));
  INV_X1    g0824(.A(new_n954), .ZN(new_n1025));
  AOI21_X1  g0825(.A(new_n670), .B1(new_n938), .B2(new_n941), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1021), .B1(new_n1025), .B2(new_n1026), .ZN(new_n1027));
  NAND3_X1  g0827(.A1(new_n1027), .A2(new_n955), .A3(new_n679), .ZN(new_n1028));
  AND2_X1   g0828(.A1(new_n241), .A2(new_n736), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n958), .B1(new_n389), .B2(new_n211), .ZN(new_n1030));
  OAI22_X1  g0830(.A1(new_n750), .A2(new_n812), .B1(new_n322), .B2(new_n768), .ZN(new_n1031));
  XOR2_X1   g0831(.A(new_n1031), .B(KEYINPUT51), .Z(new_n1032));
  NOR2_X1   g0832(.A1(new_n755), .A2(new_n767), .ZN(new_n1033));
  OAI22_X1  g0833(.A1(new_n203), .A2(new_n757), .B1(new_n760), .B2(new_n802), .ZN(new_n1034));
  AOI211_X1 g0834(.A(new_n1033), .B(new_n1034), .C1(G50), .C2(new_n751), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(new_n258), .A2(new_n806), .B1(new_n763), .B2(G143), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n1035), .A2(new_n735), .A3(new_n1036), .ZN(new_n1037));
  AOI22_X1  g0837(.A1(G317), .A2(new_n749), .B1(new_n771), .B2(G311), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  OAI21_X1  g0839(.A(new_n762), .B1(new_n752), .B2(new_n783), .ZN(new_n1040));
  AOI21_X1  g0840(.A(new_n292), .B1(new_n763), .B2(G322), .ZN(new_n1041));
  OAI21_X1  g0841(.A(new_n1041), .B1(new_n780), .B2(new_n766), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n755), .A2(new_n521), .B1(new_n757), .B2(new_n782), .ZN(new_n1043));
  OR3_X1    g0843(.A1(new_n1040), .A2(new_n1042), .A3(new_n1043), .ZN(new_n1044));
  OAI22_X1  g0844(.A1(new_n1032), .A2(new_n1037), .B1(new_n1039), .B2(new_n1044), .ZN(new_n1045));
  XNOR2_X1  g0845(.A(new_n1045), .B(KEYINPUT116), .ZN(new_n1046));
  INV_X1    g0846(.A(new_n730), .ZN(new_n1047));
  OAI221_X1 g0847(.A(new_n722), .B1(new_n1029), .B2(new_n1030), .C1(new_n1046), .C2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n932), .B2(new_n727), .ZN(new_n1049));
  NOR2_X1   g0849(.A1(new_n1025), .A2(new_n1026), .ZN(new_n1050));
  AOI21_X1  g0850(.A(new_n1049), .B1(new_n1050), .B2(new_n721), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1028), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1052), .A2(KEYINPUT117), .ZN(new_n1053));
  INV_X1    g0853(.A(KEYINPUT117), .ZN(new_n1054));
  NAND3_X1  g0854(.A1(new_n1028), .A2(new_n1051), .A3(new_n1054), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1053), .A2(new_n1055), .ZN(G390));
  AOI21_X1  g0856(.A(new_n726), .B1(new_n889), .B2(new_n891), .ZN(new_n1057));
  INV_X1    g0857(.A(new_n800), .ZN(new_n1058));
  AOI22_X1  g0858(.A1(G97), .A2(new_n806), .B1(new_n763), .B2(G294), .ZN(new_n1059));
  OAI211_X1 g0859(.A(new_n1059), .B(new_n285), .C1(new_n521), .C2(new_n768), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n819), .B(new_n1060), .C1(G87), .C2(new_n758), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n752), .A2(new_n464), .ZN(new_n1062));
  AOI211_X1 g0862(.A(new_n1033), .B(new_n1062), .C1(G283), .C2(new_n749), .ZN(new_n1063));
  NOR2_X1   g0863(.A1(new_n757), .A2(new_n812), .ZN(new_n1064));
  XNOR2_X1  g0864(.A(new_n1064), .B(KEYINPUT53), .ZN(new_n1065));
  OAI22_X1  g0865(.A1(new_n752), .A2(new_n811), .B1(new_n760), .B2(new_n201), .ZN(new_n1066));
  INV_X1    g0866(.A(G128), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n750), .A2(new_n1067), .B1(new_n322), .B2(new_n755), .ZN(new_n1068));
  INV_X1    g0868(.A(G125), .ZN(new_n1069));
  OAI21_X1  g0869(.A(new_n292), .B1(new_n745), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g0870(.A(G132), .ZN(new_n1071));
  XNOR2_X1  g0871(.A(KEYINPUT54), .B(G143), .ZN(new_n1072));
  OAI22_X1  g0872(.A1(new_n768), .A2(new_n1071), .B1(new_n766), .B2(new_n1072), .ZN(new_n1073));
  NOR4_X1   g0873(.A1(new_n1066), .A2(new_n1068), .A3(new_n1070), .A4(new_n1073), .ZN(new_n1074));
  AOI22_X1  g0874(.A1(new_n1061), .A2(new_n1063), .B1(new_n1065), .B2(new_n1074), .ZN(new_n1075));
  OAI221_X1 g0875(.A(new_n722), .B1(new_n258), .B2(new_n1058), .C1(new_n1075), .C2(new_n1047), .ZN(new_n1076));
  NOR2_X1   g0876(.A1(new_n1057), .A2(new_n1076), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n889), .A2(new_n891), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n890), .ZN(new_n1079));
  AOI21_X1  g0879(.A(new_n882), .B1(new_n706), .B2(new_n791), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n1079), .B1(new_n1080), .B2(new_n881), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n1078), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n791), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n658), .B(new_n1083), .C1(new_n714), .C2(new_n637), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n836), .B1(new_n1084), .B2(new_n882), .ZN(new_n1085));
  INV_X1    g0885(.A(KEYINPUT38), .ZN(new_n1086));
  INV_X1    g0886(.A(new_n856), .ZN(new_n1087));
  INV_X1    g0887(.A(new_n858), .ZN(new_n1088));
  AOI22_X1  g0888(.A1(new_n1087), .A2(new_n1088), .B1(new_n344), .B2(new_n364), .ZN(new_n1089));
  AOI22_X1  g0889(.A1(new_n1089), .A2(new_n854), .B1(new_n869), .B2(new_n853), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n872), .A2(new_n871), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1086), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1093));
  AOI21_X1  g0893(.A(new_n890), .B1(new_n1093), .B2(new_n868), .ZN(new_n1094));
  AOI21_X1  g0894(.A(KEYINPUT118), .B1(new_n1085), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g0895(.A1(new_n713), .A2(new_n711), .ZN(new_n1096));
  AOI21_X1  g0896(.A(new_n712), .B1(new_n647), .B2(new_n639), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n637), .B1(new_n1096), .B2(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1098), .A2(new_n665), .A3(new_n791), .ZN(new_n1099));
  AOI21_X1  g0899(.A(new_n881), .B1(new_n1099), .B2(new_n883), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n870), .A2(new_n859), .ZN(new_n1101));
  AOI21_X1  g0901(.A(KEYINPUT38), .B1(new_n1101), .B2(new_n1091), .ZN(new_n1102));
  OAI21_X1  g0902(.A(new_n1079), .B1(new_n1102), .B2(new_n863), .ZN(new_n1103));
  INV_X1    g0903(.A(KEYINPUT118), .ZN(new_n1104));
  NOR3_X1   g0904(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .ZN(new_n1105));
  OAI21_X1  g0905(.A(new_n1082), .B1(new_n1095), .B2(new_n1105), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n705), .A2(new_n791), .A3(new_n836), .ZN(new_n1107));
  NOR2_X1   g0907(.A1(new_n1107), .A2(KEYINPUT119), .ZN(new_n1108));
  INV_X1    g0908(.A(new_n1108), .ZN(new_n1109));
  NAND2_X1  g0909(.A1(new_n1106), .A2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1104), .B1(new_n1100), .B2(new_n1103), .ZN(new_n1111));
  AOI21_X1  g0911(.A(new_n882), .B1(new_n715), .B2(new_n791), .ZN(new_n1112));
  OAI211_X1 g0912(.A(new_n1094), .B(KEYINPUT118), .C1(new_n1112), .C2(new_n881), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1111), .A2(new_n1113), .ZN(new_n1114));
  NAND3_X1  g0914(.A1(new_n1114), .A2(new_n1082), .A3(new_n1108), .ZN(new_n1115));
  NAND2_X1  g0915(.A1(new_n1110), .A2(new_n1115), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n1077), .B1(new_n1116), .B2(new_n721), .ZN(new_n1117));
  INV_X1    g0917(.A(new_n1117), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n455), .A2(new_n705), .ZN(new_n1119));
  NAND3_X1  g0919(.A1(new_n894), .A2(new_n617), .A3(new_n1119), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n705), .A2(new_n791), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1122), .A2(new_n881), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1123), .A2(new_n1107), .ZN(new_n1124));
  INV_X1    g0924(.A(new_n1080), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n1124), .A2(new_n1125), .ZN(new_n1126));
  NAND3_X1  g0926(.A1(new_n1112), .A2(new_n1123), .A3(new_n1107), .ZN(new_n1127));
  NAND2_X1  g0927(.A1(new_n1126), .A2(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1121), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(new_n1129), .ZN(new_n1130));
  AOI221_X4 g0930(.A(new_n1109), .B1(new_n1078), .B2(new_n1081), .C1(new_n1111), .C2(new_n1113), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1108), .B1(new_n1114), .B2(new_n1082), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  NAND3_X1  g0933(.A1(new_n1110), .A2(new_n1115), .A3(new_n1129), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1133), .A2(new_n1134), .A3(new_n679), .ZN(new_n1135));
  INV_X1    g0935(.A(KEYINPUT120), .ZN(new_n1136));
  NAND2_X1  g0936(.A1(new_n1135), .A2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g0937(.A1(new_n1133), .A2(new_n1134), .A3(KEYINPUT120), .A4(new_n679), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1118), .B1(new_n1137), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(new_n1139), .ZN(G378));
  XNOR2_X1  g0940(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1141));
  INV_X1    g0941(.A(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n656), .B1(new_n433), .B2(new_n436), .ZN(new_n1143));
  NOR3_X1   g0943(.A1(new_n449), .A2(new_n453), .A3(new_n1143), .ZN(new_n1144));
  INV_X1    g0944(.A(new_n1143), .ZN(new_n1145));
  AOI21_X1  g0945(.A(new_n1145), .B1(new_n616), .B2(new_n452), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1142), .B1(new_n1144), .B2(new_n1146), .ZN(new_n1147));
  OAI21_X1  g0947(.A(new_n1143), .B1(new_n449), .B2(new_n453), .ZN(new_n1148));
  NAND3_X1  g0948(.A1(new_n616), .A2(new_n452), .A3(new_n1145), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n1148), .A2(new_n1149), .A3(new_n1141), .ZN(new_n1150));
  NAND2_X1  g0950(.A1(new_n1147), .A2(new_n1150), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND2_X1  g0952(.A1(new_n1152), .A2(new_n725), .ZN(new_n1153));
  OAI21_X1  g0953(.A(new_n722), .B1(G50), .B2(new_n1058), .ZN(new_n1154));
  NOR2_X1   g0954(.A1(new_n735), .A2(G41), .ZN(new_n1155));
  AOI211_X1 g0955(.A(G50), .B(new_n1155), .C1(new_n251), .C2(new_n278), .ZN(new_n1156));
  AOI22_X1  g0956(.A1(new_n771), .A2(G107), .B1(new_n763), .B2(G283), .ZN(new_n1157));
  OAI21_X1  g0957(.A(new_n1157), .B1(new_n249), .B2(new_n766), .ZN(new_n1158));
  AOI211_X1 g0958(.A(new_n996), .B(new_n1158), .C1(G68), .C2(new_n756), .ZN(new_n1159));
  NOR2_X1   g0959(.A1(new_n760), .A2(new_n202), .ZN(new_n1160));
  NOR2_X1   g0960(.A1(new_n752), .A2(new_n389), .ZN(new_n1161));
  AOI211_X1 g0961(.A(new_n1160), .B(new_n1161), .C1(G116), .C2(new_n749), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1159), .A2(new_n1162), .A3(new_n1155), .ZN(new_n1163));
  INV_X1    g0963(.A(KEYINPUT58), .ZN(new_n1164));
  AOI21_X1  g0964(.A(new_n1156), .B1(new_n1163), .B2(new_n1164), .ZN(new_n1165));
  AOI211_X1 g0965(.A(G33), .B(G41), .C1(new_n763), .C2(G124), .ZN(new_n1166));
  OAI22_X1  g0966(.A1(new_n768), .A2(new_n1067), .B1(new_n757), .B2(new_n1072), .ZN(new_n1167));
  XNOR2_X1  g0967(.A(new_n1167), .B(KEYINPUT121), .ZN(new_n1168));
  OAI22_X1  g0968(.A1(new_n750), .A2(new_n1069), .B1(new_n766), .B2(new_n811), .ZN(new_n1169));
  OAI22_X1  g0969(.A1(new_n752), .A2(new_n1071), .B1(new_n812), .B2(new_n755), .ZN(new_n1170));
  NOR3_X1   g0970(.A1(new_n1168), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT59), .ZN(new_n1172));
  OAI221_X1 g0972(.A(new_n1166), .B1(new_n322), .B2(new_n760), .C1(new_n1171), .C2(new_n1172), .ZN(new_n1173));
  AND2_X1   g0973(.A1(new_n1171), .A2(new_n1172), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1165), .B1(new_n1164), .B2(new_n1163), .C1(new_n1173), .C2(new_n1174), .ZN(new_n1175));
  AOI21_X1  g0975(.A(new_n1154), .B1(new_n1175), .B2(new_n730), .ZN(new_n1176));
  NAND2_X1  g0976(.A1(new_n1153), .A2(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n865), .A2(new_n866), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n867), .A2(new_n874), .ZN(new_n1179));
  AND4_X1   g0979(.A1(G330), .A2(new_n1178), .A3(new_n1179), .A4(new_n1151), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n1151), .B1(new_n875), .B2(G330), .ZN(new_n1181));
  OAI21_X1  g0981(.A(new_n893), .B1(new_n1180), .B2(new_n1181), .ZN(new_n1182));
  AND2_X1   g0982(.A1(new_n887), .A2(new_n892), .ZN(new_n1183));
  NAND3_X1  g0983(.A1(new_n1178), .A2(G330), .A3(new_n1179), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n1184), .A2(new_n1152), .ZN(new_n1185));
  NAND3_X1  g0985(.A1(new_n875), .A2(G330), .A3(new_n1151), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1183), .A2(new_n1185), .A3(new_n1186), .ZN(new_n1187));
  NAND2_X1  g0987(.A1(new_n1182), .A2(new_n1187), .ZN(new_n1188));
  INV_X1    g0988(.A(new_n1188), .ZN(new_n1189));
  OAI211_X1 g0989(.A(KEYINPUT122), .B(new_n1177), .C1(new_n1189), .C2(new_n720), .ZN(new_n1190));
  INV_X1    g0990(.A(KEYINPUT122), .ZN(new_n1191));
  AOI21_X1  g0991(.A(new_n720), .B1(new_n1182), .B2(new_n1187), .ZN(new_n1192));
  INV_X1    g0992(.A(new_n1177), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1191), .B1(new_n1192), .B2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1190), .A2(new_n1194), .ZN(new_n1195));
  AOI21_X1  g0995(.A(new_n1120), .B1(new_n1116), .B2(new_n1128), .ZN(new_n1196));
  INV_X1    g0996(.A(KEYINPUT123), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n1182), .A2(new_n1187), .A3(new_n1197), .ZN(new_n1198));
  NAND4_X1  g0998(.A1(new_n1183), .A2(new_n1185), .A3(KEYINPUT123), .A4(new_n1186), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1199), .ZN(new_n1200));
  OAI21_X1  g1000(.A(new_n679), .B1(new_n1196), .B2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1133), .A2(new_n1121), .ZN(new_n1202));
  AOI21_X1  g1002(.A(KEYINPUT57), .B1(new_n1202), .B2(new_n1188), .ZN(new_n1203));
  OAI21_X1  g1003(.A(new_n1195), .B1(new_n1201), .B2(new_n1203), .ZN(G375));
  INV_X1    g1004(.A(new_n1128), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1205), .A2(new_n1120), .ZN(new_n1206));
  INV_X1    g1006(.A(new_n936), .ZN(new_n1207));
  NAND3_X1  g1007(.A1(new_n1206), .A2(new_n1207), .A3(new_n1129), .ZN(new_n1208));
  AOI22_X1  g1008(.A1(new_n749), .A2(G132), .B1(new_n758), .B2(G159), .ZN(new_n1209));
  OAI221_X1 g1009(.A(new_n1209), .B1(new_n201), .B2(new_n755), .C1(new_n752), .C2(new_n1072), .ZN(new_n1210));
  AOI22_X1  g1010(.A1(new_n771), .A2(G137), .B1(new_n763), .B2(G128), .ZN(new_n1211));
  OAI21_X1  g1011(.A(new_n1211), .B1(new_n812), .B2(new_n766), .ZN(new_n1212));
  NOR4_X1   g1012(.A1(new_n1210), .A2(new_n816), .A3(new_n1160), .A4(new_n1212), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(G116), .A2(new_n751), .B1(new_n749), .B2(G294), .ZN(new_n1214));
  OAI21_X1  g1014(.A(new_n1214), .B1(new_n389), .B2(new_n757), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n292), .B1(new_n763), .B2(G303), .ZN(new_n1216));
  OAI221_X1 g1016(.A(new_n1216), .B1(new_n464), .B2(new_n766), .C1(new_n782), .C2(new_n768), .ZN(new_n1217));
  NOR4_X1   g1017(.A1(new_n1215), .A2(new_n1217), .A3(new_n972), .A4(new_n1000), .ZN(new_n1218));
  OAI21_X1  g1018(.A(new_n730), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n723), .B1(new_n203), .B2(new_n800), .ZN(new_n1220));
  OAI211_X1 g1020(.A(new_n1219), .B(new_n1220), .C1(new_n836), .C2(new_n726), .ZN(new_n1221));
  OAI21_X1  g1021(.A(new_n1221), .B1(new_n1205), .B2(new_n720), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1222), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1208), .A2(new_n1223), .ZN(G381));
  OR2_X1    g1024(.A1(G393), .A2(G396), .ZN(new_n1225));
  OR4_X1    g1025(.A1(G384), .A2(G387), .A3(G381), .A4(new_n1225), .ZN(new_n1226));
  NOR2_X1   g1026(.A1(new_n1226), .A2(G390), .ZN(new_n1227));
  AND3_X1   g1027(.A1(new_n1198), .A2(KEYINPUT57), .A3(new_n1199), .ZN(new_n1228));
  AOI21_X1  g1028(.A(new_n680), .B1(new_n1228), .B2(new_n1202), .ZN(new_n1229));
  INV_X1    g1029(.A(KEYINPUT57), .ZN(new_n1230));
  OAI21_X1  g1030(.A(new_n1230), .B1(new_n1196), .B2(new_n1189), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n1229), .A2(new_n1231), .B1(new_n1194), .B2(new_n1190), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1135), .A2(new_n1117), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(KEYINPUT124), .ZN(new_n1234));
  INV_X1    g1034(.A(KEYINPUT124), .ZN(new_n1235));
  NAND3_X1  g1035(.A1(new_n1135), .A2(new_n1117), .A3(new_n1235), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1234), .A2(new_n1236), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1227), .A2(new_n1232), .A3(new_n1237), .ZN(G407));
  NAND2_X1  g1038(.A1(new_n657), .A2(G213), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1232), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(G407), .A2(G213), .A3(new_n1241), .ZN(G409));
  NAND2_X1  g1042(.A1(new_n1206), .A2(KEYINPUT125), .ZN(new_n1243));
  INV_X1    g1043(.A(KEYINPUT60), .ZN(new_n1244));
  NAND2_X1  g1044(.A1(new_n1243), .A2(new_n1244), .ZN(new_n1245));
  NAND3_X1  g1045(.A1(new_n1206), .A2(KEYINPUT125), .A3(KEYINPUT60), .ZN(new_n1246));
  NAND2_X1  g1046(.A1(new_n1245), .A2(new_n1246), .ZN(new_n1247));
  NOR2_X1   g1047(.A1(new_n1130), .A2(new_n680), .ZN(new_n1248));
  NAND2_X1  g1048(.A1(new_n1247), .A2(new_n1248), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1249), .A2(new_n830), .A3(new_n1223), .ZN(new_n1250));
  NAND2_X1  g1050(.A1(new_n1129), .A2(new_n679), .ZN(new_n1251));
  AOI21_X1  g1051(.A(new_n1251), .B1(new_n1245), .B2(new_n1246), .ZN(new_n1252));
  OAI21_X1  g1052(.A(G384), .B1(new_n1252), .B2(new_n1222), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1250), .A2(new_n1253), .ZN(new_n1254));
  NOR2_X1   g1054(.A1(G375), .A2(new_n1139), .ZN(new_n1255));
  NAND3_X1  g1055(.A1(new_n1202), .A2(new_n1207), .A3(new_n1188), .ZN(new_n1256));
  NAND3_X1  g1056(.A1(new_n1198), .A2(new_n721), .A3(new_n1199), .ZN(new_n1257));
  AND2_X1   g1057(.A1(new_n1257), .A2(new_n1177), .ZN(new_n1258));
  AOI22_X1  g1058(.A1(new_n1234), .A2(new_n1236), .B1(new_n1256), .B2(new_n1258), .ZN(new_n1259));
  OAI211_X1 g1059(.A(new_n1239), .B(new_n1254), .C1(new_n1255), .C2(new_n1259), .ZN(new_n1260));
  NAND2_X1  g1060(.A1(new_n1260), .A2(KEYINPUT62), .ZN(new_n1261));
  INV_X1    g1061(.A(KEYINPUT61), .ZN(new_n1262));
  AND2_X1   g1062(.A1(new_n1240), .A2(G2897), .ZN(new_n1263));
  AND3_X1   g1063(.A1(new_n1250), .A2(new_n1253), .A3(new_n1263), .ZN(new_n1264));
  AOI21_X1  g1064(.A(new_n1263), .B1(new_n1250), .B2(new_n1253), .ZN(new_n1265));
  NOR2_X1   g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NAND2_X1  g1066(.A1(new_n1258), .A2(new_n1256), .ZN(new_n1267));
  AOI22_X1  g1067(.A1(G378), .A2(new_n1232), .B1(new_n1237), .B2(new_n1267), .ZN(new_n1268));
  OAI21_X1  g1068(.A(new_n1266), .B1(new_n1268), .B2(new_n1240), .ZN(new_n1269));
  INV_X1    g1069(.A(new_n1236), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1235), .B1(new_n1135), .B2(new_n1117), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n1267), .B1(new_n1270), .B2(new_n1271), .ZN(new_n1272));
  OAI21_X1  g1072(.A(new_n1272), .B1(new_n1139), .B2(G375), .ZN(new_n1273));
  INV_X1    g1073(.A(KEYINPUT62), .ZN(new_n1274));
  NAND4_X1  g1074(.A1(new_n1273), .A2(new_n1274), .A3(new_n1239), .A4(new_n1254), .ZN(new_n1275));
  NAND4_X1  g1075(.A1(new_n1261), .A2(new_n1262), .A3(new_n1269), .A4(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(G393), .A2(G396), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1225), .A2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1278), .A2(KEYINPUT126), .ZN(new_n1279));
  INV_X1    g1079(.A(KEYINPUT126), .ZN(new_n1280));
  AOI21_X1  g1080(.A(new_n1280), .B1(new_n1225), .B2(new_n1277), .ZN(new_n1281));
  NOR2_X1   g1081(.A1(new_n1279), .A2(new_n1281), .ZN(new_n1282));
  NAND3_X1  g1082(.A1(G390), .A2(new_n957), .A3(new_n984), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(G387), .A2(new_n1055), .A3(new_n1053), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1282), .A2(new_n1283), .A3(new_n1284), .ZN(new_n1285));
  AND2_X1   g1085(.A1(new_n1283), .A2(new_n1284), .ZN(new_n1286));
  INV_X1    g1086(.A(new_n1281), .ZN(new_n1287));
  OAI21_X1  g1087(.A(new_n1285), .B1(new_n1286), .B2(new_n1287), .ZN(new_n1288));
  NAND2_X1  g1088(.A1(new_n1276), .A2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1273), .A2(new_n1239), .ZN(new_n1290));
  AOI21_X1  g1090(.A(KEYINPUT61), .B1(new_n1290), .B2(new_n1266), .ZN(new_n1291));
  INV_X1    g1091(.A(KEYINPUT63), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1260), .A2(new_n1292), .ZN(new_n1293));
  AOI21_X1  g1093(.A(new_n1287), .B1(new_n1283), .B2(new_n1284), .ZN(new_n1294));
  AOI21_X1  g1094(.A(new_n1294), .B1(new_n1286), .B2(new_n1282), .ZN(new_n1295));
  NAND4_X1  g1095(.A1(new_n1273), .A2(KEYINPUT63), .A3(new_n1239), .A4(new_n1254), .ZN(new_n1296));
  NAND4_X1  g1096(.A1(new_n1291), .A2(new_n1293), .A3(new_n1295), .A4(new_n1296), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1289), .A2(new_n1297), .ZN(G405));
  NAND2_X1  g1098(.A1(new_n1254), .A2(KEYINPUT127), .ZN(new_n1299));
  NAND2_X1  g1099(.A1(G378), .A2(new_n1232), .ZN(new_n1300));
  NAND2_X1  g1100(.A1(new_n1237), .A2(G375), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NOR2_X1   g1102(.A1(new_n1295), .A2(new_n1302), .ZN(new_n1303));
  INV_X1    g1103(.A(new_n1302), .ZN(new_n1304));
  NOR2_X1   g1104(.A1(new_n1288), .A2(new_n1304), .ZN(new_n1305));
  OAI21_X1  g1105(.A(new_n1299), .B1(new_n1303), .B2(new_n1305), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1295), .A2(new_n1302), .ZN(new_n1307));
  NAND2_X1  g1107(.A1(new_n1288), .A2(new_n1304), .ZN(new_n1308));
  NAND4_X1  g1108(.A1(new_n1307), .A2(new_n1308), .A3(KEYINPUT127), .A4(new_n1254), .ZN(new_n1309));
  NAND2_X1  g1109(.A1(new_n1306), .A2(new_n1309), .ZN(G402));
endmodule


