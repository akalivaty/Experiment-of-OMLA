//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 1 0 1 0 1 0 0 0 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 0 0 1 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:01 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n610, new_n611, new_n612, new_n613,
    new_n614, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n621, new_n622, new_n623, new_n624, new_n625, new_n626, new_n627,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n733, new_n734, new_n735, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n745, new_n746, new_n747,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n755, new_n756, new_n757, new_n758, new_n759, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n782, new_n783, new_n784, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n802, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n811, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n836, new_n837, new_n838,
    new_n839, new_n840, new_n841, new_n842, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n945,
    new_n946, new_n947, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n971, new_n972, new_n974, new_n975, new_n976,
    new_n977, new_n979, new_n980, new_n981, new_n982, new_n983, new_n984,
    new_n985, new_n986, new_n987, new_n988, new_n989, new_n990, new_n991,
    new_n992, new_n993, new_n994, new_n995, new_n996, new_n998, new_n999,
    new_n1000, new_n1002, new_n1003, new_n1004, new_n1005, new_n1006,
    new_n1007, new_n1008, new_n1009, new_n1010, new_n1011, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1019, new_n1020, new_n1021, new_n1022, new_n1023, new_n1024,
    new_n1025, new_n1026, new_n1027, new_n1028, new_n1029, new_n1030,
    new_n1031, new_n1032, new_n1033, new_n1034, new_n1035, new_n1036,
    new_n1037, new_n1038, new_n1039, new_n1041, new_n1042, new_n1043,
    new_n1044, new_n1045, new_n1046, new_n1047, new_n1048, new_n1049,
    new_n1050, new_n1051, new_n1052, new_n1053;
  NOR2_X1   g000(.A1(G237), .A2(G953), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(G210), .ZN(new_n188));
  XNOR2_X1  g002(.A(new_n188), .B(KEYINPUT27), .ZN(new_n189));
  XNOR2_X1  g003(.A(KEYINPUT26), .B(G101), .ZN(new_n190));
  XNOR2_X1  g004(.A(new_n189), .B(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(new_n191), .ZN(new_n192));
  XOR2_X1   g006(.A(KEYINPUT2), .B(G113), .Z(new_n193));
  XNOR2_X1  g007(.A(G116), .B(G119), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n193), .A2(new_n194), .ZN(new_n195));
  INV_X1    g009(.A(G119), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n196), .A2(G116), .ZN(new_n197));
  INV_X1    g011(.A(G116), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n198), .A2(G119), .ZN(new_n199));
  NAND2_X1  g013(.A1(new_n197), .A2(new_n199), .ZN(new_n200));
  XNOR2_X1  g014(.A(KEYINPUT2), .B(G113), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n200), .A2(new_n201), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n195), .A2(new_n202), .ZN(new_n203));
  INV_X1    g017(.A(new_n203), .ZN(new_n204));
  INV_X1    g018(.A(G146), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n205), .A2(G143), .ZN(new_n206));
  AND2_X1   g020(.A1(KEYINPUT65), .A2(G146), .ZN(new_n207));
  NOR2_X1   g021(.A1(KEYINPUT65), .A2(G146), .ZN(new_n208));
  NOR2_X1   g022(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  OAI21_X1  g023(.A(new_n206), .B1(new_n209), .B2(G143), .ZN(new_n210));
  NAND2_X1  g024(.A1(KEYINPUT0), .A2(G128), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT64), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT64), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n213), .A2(KEYINPUT0), .A3(G128), .ZN(new_n214));
  OR2_X1    g028(.A1(KEYINPUT0), .A2(G128), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n212), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(new_n216), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n210), .A2(new_n217), .ZN(new_n218));
  INV_X1    g032(.A(KEYINPUT65), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n219), .A2(new_n205), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT65), .A2(G146), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G143), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(G143), .ZN(new_n223));
  NAND2_X1  g037(.A1(new_n223), .A2(G146), .ZN(new_n224));
  NAND4_X1  g038(.A1(new_n222), .A2(KEYINPUT0), .A3(G128), .A4(new_n224), .ZN(new_n225));
  INV_X1    g039(.A(KEYINPUT66), .ZN(new_n226));
  INV_X1    g040(.A(G134), .ZN(new_n227));
  OAI22_X1  g041(.A1(new_n226), .A2(KEYINPUT11), .B1(new_n227), .B2(G137), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G137), .ZN(new_n230));
  NAND4_X1  g044(.A1(new_n229), .A2(new_n230), .A3(KEYINPUT66), .A4(G134), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n228), .A2(new_n231), .ZN(new_n232));
  INV_X1    g046(.A(G131), .ZN(new_n233));
  OAI22_X1  g047(.A1(KEYINPUT66), .A2(new_n229), .B1(new_n230), .B2(G134), .ZN(new_n234));
  INV_X1    g048(.A(new_n234), .ZN(new_n235));
  AND3_X1   g049(.A1(new_n232), .A2(new_n233), .A3(new_n235), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n233), .B1(new_n232), .B2(new_n235), .ZN(new_n237));
  OAI211_X1 g051(.A(new_n218), .B(new_n225), .C1(new_n236), .C2(new_n237), .ZN(new_n238));
  INV_X1    g052(.A(G128), .ZN(new_n239));
  NOR2_X1   g053(.A1(new_n239), .A2(KEYINPUT1), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n222), .A2(new_n224), .A3(new_n240), .ZN(new_n241));
  AOI21_X1  g055(.A(new_n239), .B1(new_n222), .B2(KEYINPUT1), .ZN(new_n242));
  INV_X1    g056(.A(new_n206), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n220), .A2(new_n221), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n243), .B1(new_n244), .B2(new_n223), .ZN(new_n245));
  OAI21_X1  g059(.A(new_n241), .B1(new_n242), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n230), .A2(G134), .ZN(new_n247));
  NAND2_X1  g061(.A1(new_n227), .A2(G137), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n233), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n234), .B1(new_n228), .B2(new_n231), .ZN(new_n250));
  AOI21_X1  g064(.A(new_n249), .B1(new_n250), .B2(new_n233), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n246), .A2(new_n251), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n238), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n253), .A2(KEYINPUT30), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  NAND3_X1  g069(.A1(new_n238), .A2(new_n252), .A3(new_n255), .ZN(new_n256));
  AOI21_X1  g070(.A(new_n204), .B1(new_n254), .B2(new_n256), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT67), .ZN(new_n258));
  NOR2_X1   g072(.A1(new_n193), .A2(new_n194), .ZN(new_n259));
  NOR2_X1   g073(.A1(new_n200), .A2(new_n201), .ZN(new_n260));
  OAI21_X1  g074(.A(new_n258), .B1(new_n259), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g075(.A1(new_n195), .A2(KEYINPUT67), .A3(new_n202), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  AND3_X1   g077(.A1(new_n238), .A2(new_n252), .A3(new_n263), .ZN(new_n264));
  OAI21_X1  g078(.A(new_n192), .B1(new_n257), .B2(new_n264), .ZN(new_n265));
  AOI21_X1  g079(.A(new_n204), .B1(new_n238), .B2(new_n252), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n266), .B1(new_n264), .B2(KEYINPUT28), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n238), .A2(new_n252), .A3(new_n263), .ZN(new_n268));
  INV_X1    g082(.A(KEYINPUT28), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  NAND4_X1  g084(.A1(new_n267), .A2(KEYINPUT69), .A3(new_n191), .A4(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n253), .A2(new_n203), .ZN(new_n272));
  NAND4_X1  g086(.A1(new_n238), .A2(new_n252), .A3(new_n263), .A4(KEYINPUT28), .ZN(new_n273));
  NAND4_X1  g087(.A1(new_n270), .A2(new_n272), .A3(new_n191), .A4(new_n273), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT69), .ZN(new_n275));
  NAND2_X1  g089(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  INV_X1    g090(.A(KEYINPUT29), .ZN(new_n277));
  NAND4_X1  g091(.A1(new_n265), .A2(new_n271), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n278), .A2(KEYINPUT70), .ZN(new_n279));
  INV_X1    g093(.A(new_n263), .ZN(new_n280));
  NAND2_X1  g094(.A1(new_n253), .A2(new_n280), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n281), .A2(KEYINPUT71), .A3(new_n268), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  NAND4_X1  g097(.A1(new_n238), .A2(new_n252), .A3(new_n263), .A4(new_n283), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n282), .A2(KEYINPUT28), .A3(new_n284), .ZN(new_n285));
  AND3_X1   g099(.A1(new_n268), .A2(KEYINPUT72), .A3(new_n269), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT72), .B1(new_n268), .B2(new_n269), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NOR2_X1   g102(.A1(new_n192), .A2(new_n277), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n285), .A2(new_n288), .A3(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(G902), .ZN(new_n291));
  AND2_X1   g105(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g106(.A1(new_n238), .A2(new_n252), .A3(new_n255), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n255), .B1(new_n238), .B2(new_n252), .ZN(new_n294));
  OAI21_X1  g108(.A(new_n203), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n268), .ZN(new_n296));
  AOI21_X1  g110(.A(KEYINPUT29), .B1(new_n296), .B2(new_n192), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT70), .ZN(new_n298));
  NAND4_X1  g112(.A1(new_n297), .A2(new_n298), .A3(new_n276), .A4(new_n271), .ZN(new_n299));
  NAND3_X1  g113(.A1(new_n279), .A2(new_n292), .A3(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G472), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n295), .A2(new_n191), .A3(new_n268), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT31), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n295), .A2(KEYINPUT31), .A3(new_n191), .A4(new_n268), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n267), .A2(new_n270), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n307), .A2(new_n192), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NOR2_X1   g123(.A1(G472), .A2(G902), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n309), .A2(KEYINPUT32), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(KEYINPUT68), .B(KEYINPUT32), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n304), .A2(new_n305), .B1(new_n192), .B2(new_n307), .ZN(new_n313));
  INV_X1    g127(.A(new_n310), .ZN(new_n314));
  OAI21_X1  g128(.A(new_n312), .B1(new_n313), .B2(new_n314), .ZN(new_n315));
  NAND3_X1  g129(.A1(new_n301), .A2(new_n311), .A3(new_n315), .ZN(new_n316));
  OAI21_X1  g130(.A(G214), .B1(G237), .B2(G902), .ZN(new_n317));
  OAI21_X1  g131(.A(new_n225), .B1(new_n245), .B2(new_n216), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n318), .A2(G125), .ZN(new_n319));
  INV_X1    g133(.A(G125), .ZN(new_n320));
  OAI211_X1 g134(.A(new_n320), .B(new_n241), .C1(new_n242), .C2(new_n245), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n319), .A2(new_n321), .ZN(new_n322));
  INV_X1    g136(.A(G224), .ZN(new_n323));
  OR3_X1    g137(.A1(new_n323), .A2(KEYINPUT83), .A3(G953), .ZN(new_n324));
  OAI21_X1  g138(.A(KEYINPUT83), .B1(new_n323), .B2(G953), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n324), .A2(new_n325), .ZN(new_n326));
  XNOR2_X1  g140(.A(new_n326), .B(KEYINPUT84), .ZN(new_n327));
  XNOR2_X1  g141(.A(new_n322), .B(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(new_n328), .ZN(new_n329));
  INV_X1    g143(.A(G113), .ZN(new_n330));
  AND2_X1   g144(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n331));
  NOR2_X1   g145(.A1(KEYINPUT80), .A2(KEYINPUT5), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g147(.A(new_n197), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n330), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  XNOR2_X1  g149(.A(KEYINPUT80), .B(KEYINPUT5), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n194), .A2(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n335), .A2(new_n337), .ZN(new_n338));
  INV_X1    g152(.A(G104), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n339), .A2(KEYINPUT3), .ZN(new_n340));
  OR2_X1    g154(.A1(KEYINPUT78), .A2(G107), .ZN(new_n341));
  NAND2_X1  g155(.A1(KEYINPUT78), .A2(G107), .ZN(new_n342));
  NAND3_X1  g156(.A1(new_n340), .A2(new_n341), .A3(new_n342), .ZN(new_n343));
  INV_X1    g157(.A(G107), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT3), .ZN(new_n345));
  OAI21_X1  g159(.A(new_n344), .B1(new_n345), .B2(G104), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n345), .A2(G104), .ZN(new_n347));
  NAND2_X1  g161(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(G101), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n343), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g164(.A(new_n349), .B1(G104), .B2(G107), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n341), .A2(new_n342), .ZN(new_n352));
  OAI21_X1  g166(.A(new_n351), .B1(new_n352), .B2(G104), .ZN(new_n353));
  NAND4_X1  g167(.A1(new_n338), .A2(new_n195), .A3(new_n350), .A4(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n350), .A2(KEYINPUT4), .ZN(new_n355));
  AOI21_X1  g169(.A(new_n349), .B1(new_n343), .B2(new_n348), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT4), .ZN(new_n358));
  AND2_X1   g172(.A1(KEYINPUT78), .A2(G107), .ZN(new_n359));
  NOR2_X1   g173(.A1(KEYINPUT78), .A2(G107), .ZN(new_n360));
  NOR3_X1   g174(.A1(new_n347), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  AOI21_X1  g175(.A(G107), .B1(new_n339), .B2(KEYINPUT3), .ZN(new_n362));
  NOR2_X1   g176(.A1(new_n362), .A2(new_n340), .ZN(new_n363));
  OAI211_X1 g177(.A(new_n358), .B(G101), .C1(new_n361), .C2(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n364), .A2(new_n203), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n354), .B1(new_n357), .B2(new_n365), .ZN(new_n366));
  XNOR2_X1  g180(.A(G110), .B(G122), .ZN(new_n367));
  INV_X1    g181(.A(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n366), .A2(new_n368), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT82), .B(KEYINPUT6), .ZN(new_n370));
  NOR2_X1   g184(.A1(new_n369), .A2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n371), .ZN(new_n372));
  AOI22_X1  g186(.A1(new_n356), .A2(new_n358), .B1(new_n202), .B2(new_n195), .ZN(new_n373));
  OAI21_X1  g187(.A(G101), .B1(new_n361), .B2(new_n363), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n374), .A2(KEYINPUT4), .A3(new_n350), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n350), .A2(new_n353), .ZN(new_n376));
  AOI21_X1  g190(.A(new_n260), .B1(new_n335), .B2(new_n337), .ZN(new_n377));
  AOI22_X1  g191(.A1(new_n373), .A2(new_n375), .B1(new_n376), .B2(new_n377), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n378), .A2(new_n367), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n369), .A2(new_n379), .A3(KEYINPUT81), .A4(KEYINPUT6), .ZN(new_n380));
  INV_X1    g194(.A(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT6), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n382), .B1(new_n366), .B2(new_n368), .ZN(new_n383));
  AOI21_X1  g197(.A(KEYINPUT81), .B1(new_n383), .B2(new_n379), .ZN(new_n384));
  OAI211_X1 g198(.A(new_n329), .B(new_n372), .C1(new_n381), .C2(new_n384), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n373), .A2(new_n375), .ZN(new_n386));
  AND3_X1   g200(.A1(new_n386), .A2(new_n354), .A3(new_n367), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n324), .A2(KEYINPUT7), .A3(new_n325), .ZN(new_n388));
  INV_X1    g202(.A(new_n388), .ZN(new_n389));
  INV_X1    g203(.A(new_n321), .ZN(new_n390));
  AOI21_X1  g204(.A(new_n320), .B1(new_n218), .B2(new_n225), .ZN(new_n391));
  OAI21_X1  g205(.A(new_n389), .B1(new_n390), .B2(new_n391), .ZN(new_n392));
  NAND3_X1  g206(.A1(new_n319), .A2(new_n321), .A3(new_n388), .ZN(new_n393));
  INV_X1    g207(.A(new_n335), .ZN(new_n394));
  AND2_X1   g208(.A1(new_n194), .A2(KEYINPUT5), .ZN(new_n395));
  OAI21_X1  g209(.A(new_n195), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n376), .ZN(new_n397));
  XOR2_X1   g211(.A(new_n367), .B(KEYINPUT8), .Z(new_n398));
  NAND2_X1  g212(.A1(new_n350), .A2(new_n353), .ZN(new_n399));
  AOI21_X1  g213(.A(new_n398), .B1(new_n377), .B2(new_n399), .ZN(new_n400));
  AOI22_X1  g214(.A1(new_n392), .A2(new_n393), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  AOI21_X1  g215(.A(new_n387), .B1(new_n401), .B2(KEYINPUT85), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n400), .A2(new_n397), .ZN(new_n403));
  INV_X1    g217(.A(new_n393), .ZN(new_n404));
  AOI21_X1  g218(.A(new_n388), .B1(new_n319), .B2(new_n321), .ZN(new_n405));
  OAI21_X1  g219(.A(new_n403), .B1(new_n404), .B2(new_n405), .ZN(new_n406));
  INV_X1    g220(.A(KEYINPUT85), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  AOI21_X1  g222(.A(G902), .B1(new_n402), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g223(.A(G210), .B1(G237), .B2(G902), .ZN(new_n410));
  AND3_X1   g224(.A1(new_n385), .A2(new_n409), .A3(new_n410), .ZN(new_n411));
  AOI21_X1  g225(.A(new_n410), .B1(new_n385), .B2(new_n409), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n317), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(G140), .ZN(new_n414));
  NAND2_X1  g228(.A1(new_n414), .A2(G125), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n320), .A2(G140), .ZN(new_n416));
  NAND4_X1  g230(.A1(new_n220), .A2(new_n415), .A3(new_n416), .A4(new_n221), .ZN(new_n417));
  XNOR2_X1  g231(.A(G125), .B(G140), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n417), .B1(new_n205), .B2(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(KEYINPUT18), .A2(G131), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  AND3_X1   g235(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n422));
  AOI21_X1  g236(.A(G143), .B1(new_n187), .B2(G214), .ZN(new_n423));
  OAI21_X1  g237(.A(new_n421), .B1(new_n422), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g238(.A1(new_n187), .A2(G214), .ZN(new_n425));
  NAND2_X1  g239(.A1(new_n425), .A2(new_n223), .ZN(new_n426));
  NAND3_X1  g240(.A1(new_n187), .A2(G143), .A3(G214), .ZN(new_n427));
  NAND3_X1  g241(.A1(new_n426), .A2(new_n427), .A3(new_n420), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n419), .A2(new_n424), .A3(new_n428), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n429), .A2(KEYINPUT87), .ZN(new_n430));
  INV_X1    g244(.A(KEYINPUT87), .ZN(new_n431));
  NAND4_X1  g245(.A1(new_n419), .A2(new_n424), .A3(new_n428), .A4(new_n431), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n430), .A2(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n415), .A2(new_n416), .ZN(new_n434));
  INV_X1    g248(.A(KEYINPUT19), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n434), .A2(new_n435), .ZN(new_n436));
  NAND2_X1  g250(.A1(new_n418), .A2(KEYINPUT19), .ZN(new_n437));
  AOI21_X1  g251(.A(new_n244), .B1(new_n436), .B2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n415), .A2(new_n416), .A3(KEYINPUT16), .ZN(new_n439));
  OR3_X1    g253(.A1(new_n320), .A2(KEYINPUT16), .A3(G140), .ZN(new_n440));
  AND3_X1   g254(.A1(new_n439), .A2(G146), .A3(new_n440), .ZN(new_n441));
  NOR2_X1   g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  OAI21_X1  g256(.A(G131), .B1(new_n422), .B2(new_n423), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n426), .A2(new_n233), .A3(new_n427), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n442), .A2(new_n445), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n433), .A2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT90), .ZN(new_n448));
  XNOR2_X1  g262(.A(G113), .B(G122), .ZN(new_n449));
  XNOR2_X1  g263(.A(new_n449), .B(KEYINPUT89), .ZN(new_n450));
  XOR2_X1   g264(.A(KEYINPUT88), .B(G104), .Z(new_n451));
  XNOR2_X1  g265(.A(new_n450), .B(new_n451), .ZN(new_n452));
  INV_X1    g266(.A(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n447), .A2(new_n448), .A3(new_n453), .ZN(new_n454));
  AOI22_X1  g268(.A1(new_n430), .A2(new_n432), .B1(new_n442), .B2(new_n445), .ZN(new_n455));
  OAI21_X1  g269(.A(KEYINPUT90), .B1(new_n455), .B2(new_n452), .ZN(new_n456));
  AOI21_X1  g270(.A(G146), .B1(new_n439), .B2(new_n440), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n441), .A2(new_n457), .ZN(new_n458));
  OAI211_X1 g272(.A(KEYINPUT17), .B(G131), .C1(new_n422), .C2(new_n423), .ZN(new_n459));
  OAI211_X1 g273(.A(new_n458), .B(new_n459), .C1(KEYINPUT17), .C2(new_n445), .ZN(new_n460));
  NAND3_X1  g274(.A1(new_n433), .A2(new_n452), .A3(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n454), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NOR2_X1   g276(.A1(G475), .A2(G902), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  XOR2_X1   g278(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n465));
  INV_X1    g279(.A(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n464), .A2(new_n466), .ZN(new_n467));
  OAI21_X1  g281(.A(new_n467), .B1(KEYINPUT20), .B2(new_n464), .ZN(new_n468));
  INV_X1    g282(.A(G122), .ZN(new_n469));
  AOI21_X1  g283(.A(KEYINPUT14), .B1(new_n469), .B2(G116), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(G116), .ZN(new_n471));
  OAI21_X1  g285(.A(KEYINPUT91), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT91), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n198), .A2(G122), .ZN(new_n474));
  NOR2_X1   g288(.A1(new_n198), .A2(G122), .ZN(new_n475));
  OAI211_X1 g289(.A(new_n473), .B(new_n474), .C1(new_n475), .C2(KEYINPUT14), .ZN(new_n476));
  OR2_X1    g290(.A1(new_n474), .A2(KEYINPUT14), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n472), .A2(new_n476), .A3(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n478), .A2(G107), .ZN(new_n479));
  INV_X1    g293(.A(KEYINPUT92), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n478), .A2(KEYINPUT92), .A3(G107), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n223), .A2(G128), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n239), .A2(G143), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n485), .A2(G134), .ZN(new_n486));
  NAND3_X1  g300(.A1(new_n483), .A2(new_n484), .A3(new_n227), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n469), .A2(G116), .ZN(new_n489));
  NAND4_X1  g303(.A1(new_n341), .A2(new_n489), .A3(new_n474), .A4(new_n342), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(new_n491), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n481), .A2(new_n482), .A3(new_n492), .ZN(new_n493));
  OAI21_X1  g307(.A(new_n352), .B1(new_n475), .B2(new_n471), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n494), .A2(new_n490), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT13), .ZN(new_n496));
  NAND2_X1  g310(.A1(new_n483), .A2(new_n496), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n484), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n483), .A2(new_n496), .ZN(new_n499));
  OAI21_X1  g313(.A(G134), .B1(new_n498), .B2(new_n499), .ZN(new_n500));
  AND3_X1   g314(.A1(new_n495), .A2(new_n500), .A3(new_n487), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  XNOR2_X1  g316(.A(KEYINPUT9), .B(G234), .ZN(new_n503));
  INV_X1    g317(.A(G217), .ZN(new_n504));
  OR3_X1    g318(.A1(new_n503), .A2(new_n504), .A3(G953), .ZN(new_n505));
  INV_X1    g319(.A(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n493), .A2(new_n502), .A3(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(new_n506), .B1(new_n493), .B2(new_n502), .ZN(new_n509));
  OAI211_X1 g323(.A(KEYINPUT93), .B(new_n291), .C1(new_n508), .C2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(G478), .ZN(new_n511));
  NOR2_X1   g325(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g327(.A1(new_n493), .A2(new_n502), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n514), .A2(new_n505), .ZN(new_n515));
  NAND2_X1  g329(.A1(new_n515), .A2(new_n507), .ZN(new_n516));
  INV_X1    g330(.A(new_n512), .ZN(new_n517));
  NAND4_X1  g331(.A1(new_n516), .A2(KEYINPUT93), .A3(new_n291), .A4(new_n517), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  INV_X1    g334(.A(G475), .ZN(new_n521));
  NAND2_X1  g335(.A1(new_n433), .A2(new_n460), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n522), .A2(new_n453), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n523), .A2(new_n461), .ZN(new_n524));
  AOI21_X1  g338(.A(new_n521), .B1(new_n524), .B2(new_n291), .ZN(new_n525));
  INV_X1    g339(.A(new_n525), .ZN(new_n526));
  NAND2_X1  g340(.A1(G234), .A2(G237), .ZN(new_n527));
  INV_X1    g341(.A(G953), .ZN(new_n528));
  AND3_X1   g342(.A1(new_n527), .A2(G952), .A3(new_n528), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n527), .A2(G902), .A3(G953), .ZN(new_n530));
  XNOR2_X1  g344(.A(KEYINPUT21), .B(G898), .ZN(new_n531));
  AOI21_X1  g345(.A(new_n529), .B1(new_n530), .B2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n532), .ZN(new_n533));
  NAND4_X1  g347(.A1(new_n468), .A2(new_n520), .A3(new_n526), .A4(new_n533), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n413), .A2(new_n534), .ZN(new_n535));
  INV_X1    g349(.A(KEYINPUT24), .ZN(new_n536));
  NOR2_X1   g350(.A1(new_n536), .A2(G110), .ZN(new_n537));
  INV_X1    g351(.A(G110), .ZN(new_n538));
  NOR2_X1   g352(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n539));
  OAI21_X1  g353(.A(KEYINPUT73), .B1(new_n537), .B2(new_n539), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n538), .A2(KEYINPUT24), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n536), .A2(G110), .ZN(new_n542));
  INV_X1    g356(.A(KEYINPUT73), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n540), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n196), .A2(G128), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n239), .A2(G119), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g362(.A(KEYINPUT23), .ZN(new_n549));
  OAI21_X1  g363(.A(new_n549), .B1(new_n196), .B2(G128), .ZN(new_n550));
  NAND3_X1  g364(.A1(new_n239), .A2(KEYINPUT23), .A3(G119), .ZN(new_n551));
  AND3_X1   g365(.A1(new_n550), .A2(new_n546), .A3(new_n551), .ZN(new_n552));
  AOI22_X1  g366(.A1(new_n545), .A2(new_n548), .B1(new_n538), .B2(new_n552), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n439), .A2(new_n440), .A3(G146), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(new_n417), .ZN(new_n555));
  OAI21_X1  g369(.A(KEYINPUT75), .B1(new_n553), .B2(new_n555), .ZN(new_n556));
  AND3_X1   g370(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n557));
  AOI21_X1  g371(.A(new_n543), .B1(new_n541), .B2(new_n542), .ZN(new_n558));
  NOR2_X1   g372(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(new_n548), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n550), .A2(new_n546), .A3(new_n551), .ZN(new_n561));
  OAI22_X1  g375(.A1(new_n559), .A2(new_n560), .B1(G110), .B2(new_n561), .ZN(new_n562));
  INV_X1    g376(.A(new_n555), .ZN(new_n563));
  INV_X1    g377(.A(KEYINPUT75), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n562), .A2(new_n563), .A3(new_n564), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n556), .A2(new_n565), .ZN(new_n566));
  NAND3_X1  g380(.A1(new_n540), .A2(new_n560), .A3(new_n544), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n561), .A2(G110), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  OAI21_X1  g383(.A(KEYINPUT74), .B1(new_n458), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n439), .A2(new_n440), .ZN(new_n571));
  NAND2_X1  g385(.A1(new_n571), .A2(new_n205), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n572), .A2(new_n554), .ZN(new_n573));
  INV_X1    g387(.A(KEYINPUT74), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n573), .A2(new_n574), .A3(new_n567), .A4(new_n568), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n528), .A2(G221), .A3(G234), .ZN(new_n577));
  XNOR2_X1  g391(.A(new_n577), .B(KEYINPUT76), .ZN(new_n578));
  XNOR2_X1  g392(.A(KEYINPUT22), .B(G137), .ZN(new_n579));
  XNOR2_X1  g393(.A(new_n578), .B(new_n579), .ZN(new_n580));
  AND3_X1   g394(.A1(new_n566), .A2(new_n576), .A3(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n580), .B1(new_n566), .B2(new_n576), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  INV_X1    g397(.A(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n504), .B1(G234), .B2(new_n291), .ZN(new_n585));
  NOR2_X1   g399(.A1(new_n585), .A2(G902), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NOR2_X1   g401(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n583), .A2(KEYINPUT25), .A3(new_n291), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n566), .A2(new_n576), .ZN(new_n590));
  INV_X1    g404(.A(new_n580), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n566), .A2(new_n576), .A3(new_n580), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n592), .A2(new_n291), .A3(new_n593), .ZN(new_n594));
  INV_X1    g408(.A(KEYINPUT25), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n594), .A2(new_n595), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n589), .A2(new_n596), .ZN(new_n597));
  AOI21_X1  g411(.A(new_n588), .B1(new_n597), .B2(new_n585), .ZN(new_n598));
  NAND4_X1  g412(.A1(new_n375), .A2(new_n218), .A3(new_n225), .A4(new_n364), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT10), .ZN(new_n600));
  INV_X1    g414(.A(new_n241), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n206), .A2(KEYINPUT1), .ZN(new_n602));
  AOI22_X1  g416(.A1(new_n222), .A2(new_n224), .B1(new_n602), .B2(G128), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g418(.A(new_n600), .B1(new_n604), .B2(new_n399), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n376), .A2(new_n246), .A3(KEYINPUT10), .ZN(new_n606));
  NOR2_X1   g420(.A1(new_n236), .A2(new_n237), .ZN(new_n607));
  NAND4_X1  g421(.A1(new_n599), .A2(new_n605), .A3(new_n606), .A4(new_n607), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n528), .A2(G227), .ZN(new_n609));
  XNOR2_X1  g423(.A(new_n609), .B(KEYINPUT77), .ZN(new_n610));
  XNOR2_X1  g424(.A(G110), .B(G140), .ZN(new_n611));
  XOR2_X1   g425(.A(new_n610), .B(new_n611), .Z(new_n612));
  AND2_X1   g426(.A1(new_n608), .A2(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n599), .A2(new_n605), .A3(new_n606), .ZN(new_n614));
  INV_X1    g428(.A(new_n607), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n614), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n613), .A2(new_n616), .ZN(new_n617));
  INV_X1    g431(.A(new_n608), .ZN(new_n618));
  OAI21_X1  g432(.A(KEYINPUT79), .B1(new_n376), .B2(new_n246), .ZN(new_n619));
  AND2_X1   g433(.A1(new_n222), .A2(KEYINPUT1), .ZN(new_n620));
  OAI21_X1  g434(.A(new_n210), .B1(new_n620), .B2(new_n239), .ZN(new_n621));
  INV_X1    g435(.A(KEYINPUT79), .ZN(new_n622));
  NAND4_X1  g436(.A1(new_n621), .A2(new_n399), .A3(new_n622), .A4(new_n241), .ZN(new_n623));
  OAI21_X1  g437(.A(new_n376), .B1(new_n601), .B2(new_n603), .ZN(new_n624));
  NAND3_X1  g438(.A1(new_n619), .A2(new_n623), .A3(new_n624), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n625), .A2(new_n615), .ZN(new_n626));
  INV_X1    g440(.A(KEYINPUT12), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND3_X1  g442(.A1(new_n625), .A2(KEYINPUT12), .A3(new_n615), .ZN(new_n629));
  AOI21_X1  g443(.A(new_n618), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  OAI211_X1 g444(.A(G469), .B(new_n617), .C1(new_n630), .C2(new_n612), .ZN(new_n631));
  INV_X1    g445(.A(G469), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n608), .A2(new_n612), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n633), .B1(new_n628), .B2(new_n629), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n612), .B1(new_n616), .B2(new_n608), .ZN(new_n635));
  OAI211_X1 g449(.A(new_n632), .B(new_n291), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  NAND2_X1  g450(.A1(G469), .A2(G902), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n631), .A2(new_n636), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g452(.A(G221), .B1(new_n503), .B2(G902), .ZN(new_n639));
  NAND2_X1  g453(.A1(new_n638), .A2(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n640), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n316), .A2(new_n535), .A3(new_n598), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G101), .ZN(G3));
  OAI21_X1  g457(.A(G472), .B1(new_n313), .B2(G902), .ZN(new_n644));
  NAND2_X1  g458(.A1(new_n309), .A2(new_n310), .ZN(new_n645));
  AND3_X1   g459(.A1(new_n644), .A2(new_n645), .A3(new_n598), .ZN(new_n646));
  INV_X1    g460(.A(new_n317), .ZN(new_n647));
  INV_X1    g461(.A(new_n410), .ZN(new_n648));
  INV_X1    g462(.A(KEYINPUT81), .ZN(new_n649));
  OAI21_X1  g463(.A(KEYINPUT6), .B1(new_n378), .B2(new_n367), .ZN(new_n650));
  OAI21_X1  g464(.A(new_n649), .B1(new_n650), .B2(new_n387), .ZN(new_n651));
  AOI211_X1 g465(.A(new_n328), .B(new_n371), .C1(new_n651), .C2(new_n380), .ZN(new_n652));
  OAI211_X1 g466(.A(KEYINPUT85), .B(new_n403), .C1(new_n404), .C2(new_n405), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n653), .A2(new_n379), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n401), .A2(KEYINPUT85), .ZN(new_n655));
  OAI21_X1  g469(.A(new_n291), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  OAI21_X1  g470(.A(new_n648), .B1(new_n652), .B2(new_n656), .ZN(new_n657));
  NAND3_X1  g471(.A1(new_n385), .A2(new_n409), .A3(new_n410), .ZN(new_n658));
  AOI211_X1 g472(.A(new_n532), .B(new_n647), .C1(new_n657), .C2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(KEYINPUT20), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n462), .A2(new_n660), .A3(new_n463), .ZN(new_n661));
  AOI21_X1  g475(.A(new_n465), .B1(new_n462), .B2(new_n463), .ZN(new_n662));
  OAI21_X1  g476(.A(new_n526), .B1(new_n661), .B2(new_n662), .ZN(new_n663));
  OAI21_X1  g477(.A(KEYINPUT33), .B1(new_n506), .B2(KEYINPUT94), .ZN(new_n664));
  OAI21_X1  g478(.A(new_n664), .B1(new_n508), .B2(new_n509), .ZN(new_n665));
  INV_X1    g479(.A(new_n664), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n515), .A2(new_n507), .A3(new_n666), .ZN(new_n667));
  AOI21_X1  g481(.A(new_n511), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI211_X1 g482(.A(new_n511), .B(new_n291), .C1(new_n508), .C2(new_n509), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n511), .A2(new_n291), .ZN(new_n670));
  INV_X1    g484(.A(new_n670), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n669), .A2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  NAND2_X1  g487(.A1(new_n663), .A2(new_n673), .ZN(new_n674));
  INV_X1    g488(.A(new_n674), .ZN(new_n675));
  NAND4_X1  g489(.A1(new_n646), .A2(new_n641), .A3(new_n659), .A4(new_n675), .ZN(new_n676));
  XOR2_X1   g490(.A(KEYINPUT34), .B(G104), .Z(new_n677));
  XNOR2_X1  g491(.A(new_n676), .B(new_n677), .ZN(G6));
  AND2_X1   g492(.A1(new_n646), .A2(new_n641), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n647), .B1(new_n657), .B2(new_n658), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n462), .A2(new_n465), .A3(new_n463), .ZN(new_n681));
  NAND2_X1  g495(.A1(new_n467), .A2(new_n681), .ZN(new_n682));
  AOI21_X1  g496(.A(new_n525), .B1(new_n513), .B2(new_n518), .ZN(new_n683));
  AND3_X1   g497(.A1(new_n682), .A2(new_n683), .A3(new_n533), .ZN(new_n684));
  AND2_X1   g498(.A1(new_n680), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g499(.A1(new_n679), .A2(new_n685), .ZN(new_n686));
  XOR2_X1   g500(.A(KEYINPUT35), .B(G107), .Z(new_n687));
  XNOR2_X1  g501(.A(new_n686), .B(new_n687), .ZN(G9));
  AOI21_X1  g502(.A(KEYINPUT25), .B1(new_n583), .B2(new_n291), .ZN(new_n689));
  NOR4_X1   g503(.A1(new_n581), .A2(new_n582), .A3(new_n595), .A4(G902), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n585), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  NOR2_X1   g505(.A1(new_n591), .A2(KEYINPUT36), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n590), .B(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n586), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n691), .A2(new_n694), .ZN(new_n695));
  AND3_X1   g509(.A1(new_n644), .A2(new_n695), .A3(new_n645), .ZN(new_n696));
  NAND3_X1  g510(.A1(new_n535), .A2(new_n696), .A3(new_n641), .ZN(new_n697));
  XNOR2_X1  g511(.A(KEYINPUT37), .B(G110), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(KEYINPUT96), .ZN(new_n699));
  XOR2_X1   g513(.A(new_n699), .B(KEYINPUT95), .Z(new_n700));
  XNOR2_X1  g514(.A(new_n697), .B(new_n700), .ZN(G12));
  AOI22_X1  g515(.A1(new_n597), .A2(new_n585), .B1(new_n586), .B2(new_n693), .ZN(new_n702));
  NOR2_X1   g516(.A1(new_n413), .A2(new_n702), .ZN(new_n703));
  INV_X1    g517(.A(G900), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n529), .B1(new_n530), .B2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n705), .ZN(new_n706));
  AND3_X1   g520(.A1(new_n682), .A2(new_n683), .A3(new_n706), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n316), .A2(new_n641), .A3(new_n703), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G128), .ZN(G30));
  INV_X1    g523(.A(KEYINPUT97), .ZN(new_n710));
  OAI21_X1  g524(.A(new_n710), .B1(new_n411), .B2(new_n412), .ZN(new_n711));
  NAND3_X1  g525(.A1(new_n657), .A2(KEYINPUT97), .A3(new_n658), .ZN(new_n712));
  XNOR2_X1  g526(.A(KEYINPUT98), .B(KEYINPUT38), .ZN(new_n713));
  AND3_X1   g527(.A1(new_n711), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n713), .B1(new_n711), .B2(new_n712), .ZN(new_n715));
  OR2_X1    g529(.A1(new_n714), .A2(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n663), .A2(new_n519), .ZN(new_n717));
  NOR3_X1   g531(.A1(new_n717), .A2(new_n695), .A3(new_n647), .ZN(new_n718));
  NAND2_X1  g532(.A1(new_n296), .A2(new_n191), .ZN(new_n719));
  AND2_X1   g533(.A1(new_n282), .A2(new_n284), .ZN(new_n720));
  OAI211_X1 g534(.A(new_n719), .B(new_n291), .C1(new_n191), .C2(new_n720), .ZN(new_n721));
  AND3_X1   g535(.A1(new_n721), .A2(KEYINPUT99), .A3(G472), .ZN(new_n722));
  AOI21_X1  g536(.A(KEYINPUT99), .B1(new_n721), .B2(G472), .ZN(new_n723));
  OAI211_X1 g537(.A(new_n311), .B(new_n315), .C1(new_n722), .C2(new_n723), .ZN(new_n724));
  XOR2_X1   g538(.A(new_n705), .B(KEYINPUT39), .Z(new_n725));
  INV_X1    g539(.A(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n640), .A2(new_n726), .ZN(new_n727));
  INV_X1    g541(.A(KEYINPUT40), .ZN(new_n728));
  OAI211_X1 g542(.A(new_n718), .B(new_n724), .C1(new_n727), .C2(new_n728), .ZN(new_n729));
  NOR3_X1   g543(.A1(new_n640), .A2(KEYINPUT40), .A3(new_n726), .ZN(new_n730));
  NOR3_X1   g544(.A1(new_n716), .A2(new_n729), .A3(new_n730), .ZN(new_n731));
  XNOR2_X1  g545(.A(new_n731), .B(new_n223), .ZN(G45));
  NAND3_X1  g546(.A1(new_n663), .A2(new_n673), .A3(new_n706), .ZN(new_n733));
  NOR3_X1   g547(.A1(new_n413), .A2(new_n733), .A3(new_n702), .ZN(new_n734));
  NAND3_X1  g548(.A1(new_n734), .A2(new_n316), .A3(new_n641), .ZN(new_n735));
  XNOR2_X1  g549(.A(new_n735), .B(G146), .ZN(G48));
  NOR2_X1   g550(.A1(new_n634), .A2(new_n635), .ZN(new_n737));
  OAI21_X1  g551(.A(G469), .B1(new_n737), .B2(G902), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n738), .A2(new_n639), .A3(new_n636), .ZN(new_n739));
  INV_X1    g553(.A(new_n598), .ZN(new_n740));
  NOR2_X1   g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  NAND4_X1  g555(.A1(new_n316), .A2(new_n675), .A3(new_n741), .A4(new_n659), .ZN(new_n742));
  XNOR2_X1  g556(.A(KEYINPUT41), .B(G113), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n742), .B(new_n743), .ZN(G15));
  INV_X1    g558(.A(G472), .ZN(new_n745));
  NAND2_X1  g559(.A1(new_n290), .A2(new_n291), .ZN(new_n746));
  AOI21_X1  g560(.A(new_n746), .B1(KEYINPUT70), .B2(new_n278), .ZN(new_n747));
  AOI21_X1  g561(.A(new_n745), .B1(new_n747), .B2(new_n299), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n311), .A2(new_n315), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  AND3_X1   g564(.A1(new_n625), .A2(KEYINPUT12), .A3(new_n615), .ZN(new_n751));
  AOI21_X1  g565(.A(KEYINPUT12), .B1(new_n625), .B2(new_n615), .ZN(new_n752));
  OAI21_X1  g566(.A(new_n613), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(new_n616), .A2(new_n608), .ZN(new_n754));
  INV_X1    g568(.A(new_n612), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n753), .A2(new_n756), .ZN(new_n757));
  AOI21_X1  g571(.A(new_n632), .B1(new_n757), .B2(new_n291), .ZN(new_n758));
  AOI211_X1 g572(.A(G469), .B(G902), .C1(new_n753), .C2(new_n756), .ZN(new_n759));
  INV_X1    g573(.A(new_n639), .ZN(new_n760));
  NOR3_X1   g574(.A1(new_n758), .A2(new_n759), .A3(new_n760), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n761), .A2(new_n680), .A3(new_n684), .A4(new_n598), .ZN(new_n762));
  OAI21_X1  g576(.A(KEYINPUT100), .B1(new_n750), .B2(new_n762), .ZN(new_n763));
  INV_X1    g577(.A(KEYINPUT100), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n316), .A2(new_n685), .A3(new_n764), .A4(new_n741), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n763), .A2(new_n765), .ZN(new_n766));
  XNOR2_X1  g580(.A(new_n766), .B(G116), .ZN(G18));
  INV_X1    g581(.A(KEYINPUT101), .ZN(new_n768));
  OAI21_X1  g582(.A(new_n768), .B1(new_n413), .B2(new_n739), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n761), .A2(new_n680), .A3(KEYINPUT101), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n534), .A2(new_n702), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n769), .A2(new_n316), .A3(new_n770), .A4(new_n771), .ZN(new_n772));
  XOR2_X1   g586(.A(KEYINPUT102), .B(G119), .Z(new_n773));
  XNOR2_X1  g587(.A(new_n772), .B(new_n773), .ZN(G21));
  AND2_X1   g588(.A1(new_n304), .A2(new_n305), .ZN(new_n775));
  AOI21_X1  g589(.A(new_n191), .B1(new_n285), .B2(new_n288), .ZN(new_n776));
  OAI21_X1  g590(.A(new_n310), .B1(new_n775), .B2(new_n776), .ZN(new_n777));
  AND3_X1   g591(.A1(new_n644), .A2(new_n777), .A3(new_n598), .ZN(new_n778));
  NOR2_X1   g592(.A1(new_n717), .A2(new_n532), .ZN(new_n779));
  NAND4_X1  g593(.A1(new_n778), .A2(new_n680), .A3(new_n761), .A4(new_n779), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(G122), .ZN(G24));
  INV_X1    g595(.A(new_n733), .ZN(new_n782));
  AND3_X1   g596(.A1(new_n644), .A2(new_n695), .A3(new_n777), .ZN(new_n783));
  NAND4_X1  g597(.A1(new_n769), .A2(new_n770), .A3(new_n782), .A4(new_n783), .ZN(new_n784));
  XNOR2_X1  g598(.A(new_n784), .B(G125), .ZN(G27));
  XOR2_X1   g599(.A(new_n637), .B(KEYINPUT103), .Z(new_n786));
  NAND3_X1  g600(.A1(new_n631), .A2(new_n636), .A3(new_n786), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n787), .A2(new_n639), .ZN(new_n788));
  NAND3_X1  g602(.A1(new_n657), .A2(new_n317), .A3(new_n658), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n788), .A2(new_n789), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n316), .A2(new_n790), .A3(new_n598), .A4(new_n782), .ZN(new_n791));
  XOR2_X1   g605(.A(KEYINPUT104), .B(KEYINPUT42), .Z(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT32), .B1(new_n309), .B2(new_n310), .ZN(new_n794));
  INV_X1    g608(.A(KEYINPUT32), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n313), .A2(new_n795), .A3(new_n314), .ZN(new_n796));
  NOR2_X1   g610(.A1(new_n794), .A2(new_n796), .ZN(new_n797));
  AOI21_X1  g611(.A(new_n740), .B1(new_n797), .B2(new_n301), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n798), .A2(KEYINPUT42), .A3(new_n782), .A4(new_n790), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g614(.A(new_n800), .B(G131), .ZN(G33));
  NAND4_X1  g615(.A1(new_n316), .A2(new_n790), .A3(new_n598), .A4(new_n707), .ZN(new_n802));
  XNOR2_X1  g616(.A(new_n802), .B(G134), .ZN(G36));
  OR2_X1    g617(.A1(new_n668), .A2(new_n672), .ZN(new_n804));
  NOR2_X1   g618(.A1(new_n804), .A2(new_n663), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT43), .ZN(new_n806));
  AOI21_X1  g620(.A(new_n702), .B1(new_n645), .B2(new_n644), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n806), .A2(KEYINPUT44), .A3(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(new_n789), .ZN(new_n809));
  AND3_X1   g623(.A1(new_n808), .A2(KEYINPUT107), .A3(new_n809), .ZN(new_n810));
  AOI21_X1  g624(.A(KEYINPUT107), .B1(new_n808), .B2(new_n809), .ZN(new_n811));
  AND2_X1   g625(.A1(new_n806), .A2(new_n807), .ZN(new_n812));
  OAI22_X1  g626(.A1(new_n810), .A2(new_n811), .B1(KEYINPUT44), .B2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(new_n786), .ZN(new_n814));
  OAI21_X1  g628(.A(new_n617), .B1(new_n630), .B2(new_n612), .ZN(new_n815));
  INV_X1    g629(.A(KEYINPUT45), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n815), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n817), .A2(G469), .ZN(new_n818));
  NOR2_X1   g632(.A1(new_n815), .A2(new_n816), .ZN(new_n819));
  OR3_X1    g633(.A1(new_n818), .A2(KEYINPUT105), .A3(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(KEYINPUT105), .B1(new_n818), .B2(new_n819), .ZN(new_n821));
  AOI21_X1  g635(.A(new_n814), .B1(new_n820), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g636(.A(new_n636), .B1(new_n822), .B2(KEYINPUT46), .ZN(new_n823));
  INV_X1    g637(.A(KEYINPUT46), .ZN(new_n824));
  AOI211_X1 g638(.A(new_n824), .B(new_n814), .C1(new_n820), .C2(new_n821), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n639), .B1(new_n823), .B2(new_n825), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT106), .B1(new_n826), .B2(new_n726), .ZN(new_n827));
  AND2_X1   g641(.A1(new_n820), .A2(new_n821), .ZN(new_n828));
  OAI21_X1  g642(.A(new_n824), .B1(new_n828), .B2(new_n814), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n822), .A2(KEYINPUT46), .ZN(new_n830));
  NAND3_X1  g644(.A1(new_n829), .A2(new_n636), .A3(new_n830), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT106), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n831), .A2(new_n832), .A3(new_n639), .A4(new_n725), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n813), .B1(new_n827), .B2(new_n833), .ZN(new_n834));
  XNOR2_X1  g648(.A(new_n834), .B(new_n230), .ZN(G39));
  NOR4_X1   g649(.A1(new_n316), .A2(new_n598), .A3(new_n733), .A4(new_n789), .ZN(new_n836));
  INV_X1    g650(.A(new_n836), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n831), .A2(KEYINPUT47), .A3(new_n639), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT47), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n826), .A2(new_n839), .ZN(new_n840));
  AOI21_X1  g654(.A(new_n837), .B1(new_n838), .B2(new_n840), .ZN(new_n841));
  XOR2_X1   g655(.A(KEYINPUT108), .B(G140), .Z(new_n842));
  XNOR2_X1  g656(.A(new_n841), .B(new_n842), .ZN(G42));
  NOR3_X1   g657(.A1(new_n740), .A2(new_n760), .A3(new_n647), .ZN(new_n844));
  INV_X1    g658(.A(KEYINPUT49), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n758), .A2(new_n759), .ZN(new_n846));
  OAI211_X1 g660(.A(new_n844), .B(new_n805), .C1(new_n845), .C2(new_n846), .ZN(new_n847));
  AOI21_X1  g661(.A(new_n847), .B1(new_n845), .B2(new_n846), .ZN(new_n848));
  INV_X1    g662(.A(new_n724), .ZN(new_n849));
  NAND3_X1  g663(.A1(new_n848), .A2(new_n849), .A3(new_n716), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n739), .A2(new_n789), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n598), .A3(new_n529), .A4(new_n851), .ZN(new_n852));
  XOR2_X1   g666(.A(new_n852), .B(KEYINPUT114), .Z(new_n853));
  AND2_X1   g667(.A1(new_n853), .A2(new_n675), .ZN(new_n854));
  NAND3_X1  g668(.A1(new_n806), .A2(new_n529), .A3(new_n851), .ZN(new_n855));
  INV_X1    g669(.A(new_n798), .ZN(new_n856));
  NOR2_X1   g670(.A1(new_n855), .A2(new_n856), .ZN(new_n857));
  XNOR2_X1  g671(.A(new_n857), .B(KEYINPUT48), .ZN(new_n858));
  NAND3_X1  g672(.A1(new_n806), .A2(new_n529), .A3(new_n778), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n769), .A2(new_n770), .ZN(new_n860));
  OAI211_X1 g674(.A(G952), .B(new_n528), .C1(new_n859), .C2(new_n860), .ZN(new_n861));
  NOR3_X1   g675(.A1(new_n854), .A2(new_n858), .A3(new_n861), .ZN(new_n862));
  XOR2_X1   g676(.A(new_n862), .B(KEYINPUT115), .Z(new_n863));
  INV_X1    g677(.A(new_n859), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n864), .A2(new_n647), .A3(new_n716), .A4(new_n761), .ZN(new_n865));
  INV_X1    g679(.A(KEYINPUT113), .ZN(new_n866));
  OR3_X1    g680(.A1(new_n865), .A2(new_n866), .A3(KEYINPUT50), .ZN(new_n867));
  NAND4_X1  g681(.A1(new_n853), .A2(new_n468), .A3(new_n526), .A4(new_n804), .ZN(new_n868));
  NAND4_X1  g682(.A1(new_n806), .A2(new_n529), .A3(new_n783), .A4(new_n851), .ZN(new_n869));
  XNOR2_X1  g683(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n865), .A2(new_n870), .ZN(new_n871));
  NAND4_X1  g685(.A1(new_n867), .A2(new_n868), .A3(new_n869), .A4(new_n871), .ZN(new_n872));
  INV_X1    g686(.A(new_n846), .ZN(new_n873));
  OAI211_X1 g687(.A(new_n838), .B(new_n840), .C1(new_n639), .C2(new_n873), .ZN(new_n874));
  NOR2_X1   g688(.A1(new_n859), .A2(new_n789), .ZN(new_n875));
  AOI21_X1  g689(.A(new_n872), .B1(new_n874), .B2(new_n875), .ZN(new_n876));
  OAI21_X1  g690(.A(new_n863), .B1(new_n876), .B2(KEYINPUT51), .ZN(new_n877));
  NOR2_X1   g691(.A1(new_n413), .A2(new_n717), .ZN(new_n878));
  INV_X1    g692(.A(new_n788), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n695), .A2(new_n705), .ZN(new_n880));
  NAND4_X1  g694(.A1(new_n878), .A2(new_n724), .A3(new_n879), .A4(new_n880), .ZN(new_n881));
  NAND4_X1  g695(.A1(new_n708), .A2(new_n784), .A3(new_n735), .A4(new_n881), .ZN(new_n882));
  NAND2_X1  g696(.A1(new_n882), .A2(KEYINPUT52), .ZN(new_n883));
  AND2_X1   g697(.A1(new_n311), .A2(new_n315), .ZN(new_n884));
  AOI21_X1  g698(.A(new_n640), .B1(new_n884), .B2(new_n301), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n703), .C1(new_n707), .C2(new_n782), .ZN(new_n886));
  INV_X1    g700(.A(KEYINPUT52), .ZN(new_n887));
  NAND4_X1  g701(.A1(new_n886), .A2(new_n887), .A3(new_n784), .A4(new_n881), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n883), .A2(new_n888), .ZN(new_n889));
  AND3_X1   g703(.A1(new_n772), .A2(new_n642), .A3(new_n742), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n468), .A2(new_n683), .ZN(new_n891));
  INV_X1    g705(.A(new_n891), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n659), .A2(new_n892), .ZN(new_n893));
  INV_X1    g707(.A(KEYINPUT109), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND3_X1  g709(.A1(new_n659), .A2(KEYINPUT109), .A3(new_n892), .ZN(new_n896));
  NAND3_X1  g710(.A1(new_n895), .A2(new_n679), .A3(new_n896), .ZN(new_n897));
  AND3_X1   g711(.A1(new_n780), .A2(new_n697), .A3(new_n676), .ZN(new_n898));
  NAND4_X1  g712(.A1(new_n890), .A2(new_n766), .A3(new_n897), .A4(new_n898), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT110), .ZN(new_n900));
  INV_X1    g714(.A(new_n681), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n901), .A2(new_n662), .ZN(new_n902));
  INV_X1    g716(.A(new_n461), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n452), .B1(new_n433), .B2(new_n460), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n291), .B1(new_n903), .B2(new_n904), .ZN(new_n905));
  AOI21_X1  g719(.A(new_n705), .B1(new_n905), .B2(G475), .ZN(new_n906));
  NAND3_X1  g720(.A1(new_n513), .A2(new_n906), .A3(new_n518), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n900), .B1(new_n902), .B2(new_n907), .ZN(new_n908));
  NAND4_X1  g722(.A1(new_n520), .A2(new_n682), .A3(KEYINPUT110), .A4(new_n906), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n789), .A2(new_n702), .ZN(new_n911));
  NAND4_X1  g725(.A1(new_n885), .A2(KEYINPUT111), .A3(new_n910), .A4(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(KEYINPUT111), .ZN(new_n913));
  OAI21_X1  g727(.A(new_n641), .B1(new_n748), .B2(new_n749), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n911), .A2(new_n910), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n912), .A2(new_n916), .ZN(new_n917));
  NAND3_X1  g731(.A1(new_n790), .A2(new_n783), .A3(new_n782), .ZN(new_n918));
  AND2_X1   g732(.A1(new_n802), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g733(.A1(new_n800), .A2(new_n917), .A3(new_n919), .ZN(new_n920));
  NOR3_X1   g734(.A1(new_n889), .A2(new_n899), .A3(new_n920), .ZN(new_n921));
  XNOR2_X1  g735(.A(KEYINPUT112), .B(KEYINPUT53), .ZN(new_n922));
  INV_X1    g736(.A(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n921), .A2(new_n923), .ZN(new_n924));
  OAI21_X1  g738(.A(new_n924), .B1(KEYINPUT53), .B2(new_n921), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n925), .A2(KEYINPUT54), .ZN(new_n926));
  AND2_X1   g740(.A1(new_n883), .A2(new_n888), .ZN(new_n927));
  NAND3_X1  g741(.A1(new_n898), .A2(new_n766), .A3(new_n897), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n772), .A2(new_n642), .A3(new_n742), .ZN(new_n929));
  NOR2_X1   g743(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  AND3_X1   g744(.A1(new_n800), .A2(new_n917), .A3(new_n919), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n927), .A2(KEYINPUT53), .A3(new_n930), .A4(new_n931), .ZN(new_n932));
  OAI21_X1  g746(.A(new_n932), .B1(new_n921), .B2(new_n923), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n926), .B1(KEYINPUT54), .B2(new_n933), .ZN(new_n934));
  AND2_X1   g748(.A1(new_n876), .A2(KEYINPUT51), .ZN(new_n935));
  NOR3_X1   g749(.A1(new_n877), .A2(new_n934), .A3(new_n935), .ZN(new_n936));
  NOR2_X1   g750(.A1(G952), .A2(G953), .ZN(new_n937));
  OAI21_X1  g751(.A(new_n850), .B1(new_n936), .B2(new_n937), .ZN(G75));
  OAI21_X1  g752(.A(new_n372), .B1(new_n381), .B2(new_n384), .ZN(new_n939));
  NAND2_X1  g753(.A1(new_n939), .A2(new_n328), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n940), .A2(new_n385), .ZN(new_n941));
  XNOR2_X1  g755(.A(KEYINPUT116), .B(KEYINPUT55), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n941), .B(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  NAND2_X1  g758(.A1(new_n930), .A2(new_n931), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n922), .B1(new_n945), .B2(new_n889), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n291), .B1(new_n946), .B2(new_n932), .ZN(new_n947));
  AND2_X1   g761(.A1(new_n947), .A2(G210), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n944), .B1(new_n948), .B2(KEYINPUT56), .ZN(new_n949));
  NOR2_X1   g763(.A1(new_n528), .A2(G952), .ZN(new_n950));
  INV_X1    g764(.A(new_n950), .ZN(new_n951));
  NAND2_X1  g765(.A1(new_n949), .A2(new_n951), .ZN(new_n952));
  NOR2_X1   g766(.A1(new_n948), .A2(KEYINPUT117), .ZN(new_n953));
  NAND3_X1  g767(.A1(new_n947), .A2(KEYINPUT117), .A3(G210), .ZN(new_n954));
  NOR2_X1   g768(.A1(new_n944), .A2(KEYINPUT56), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n954), .A2(new_n955), .ZN(new_n956));
  NOR2_X1   g770(.A1(new_n953), .A2(new_n956), .ZN(new_n957));
  OAI21_X1  g771(.A(KEYINPUT118), .B1(new_n952), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g772(.A1(new_n954), .A2(new_n955), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n959), .B1(KEYINPUT117), .B2(new_n948), .ZN(new_n960));
  INV_X1    g774(.A(KEYINPUT118), .ZN(new_n961));
  NAND4_X1  g775(.A1(new_n960), .A2(new_n949), .A3(new_n961), .A4(new_n951), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n958), .A2(new_n962), .ZN(G51));
  XNOR2_X1  g777(.A(new_n933), .B(KEYINPUT54), .ZN(new_n964));
  XNOR2_X1  g778(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n965));
  XNOR2_X1  g779(.A(new_n786), .B(new_n965), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n964), .A2(new_n966), .ZN(new_n967));
  NAND2_X1  g781(.A1(new_n967), .A2(new_n757), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n947), .A2(new_n828), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n950), .B1(new_n968), .B2(new_n969), .ZN(G54));
  AND3_X1   g784(.A1(new_n947), .A2(KEYINPUT58), .A3(G475), .ZN(new_n971));
  OAI21_X1  g785(.A(new_n951), .B1(new_n971), .B2(new_n462), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n972), .B1(new_n462), .B2(new_n971), .ZN(G60));
  AND2_X1   g787(.A1(new_n665), .A2(new_n667), .ZN(new_n974));
  XOR2_X1   g788(.A(new_n670), .B(KEYINPUT59), .Z(new_n975));
  AOI21_X1  g789(.A(new_n974), .B1(new_n934), .B2(new_n975), .ZN(new_n976));
  AND3_X1   g790(.A1(new_n964), .A2(new_n974), .A3(new_n975), .ZN(new_n977));
  NOR3_X1   g791(.A1(new_n976), .A2(new_n977), .A3(new_n950), .ZN(G63));
  NAND2_X1  g792(.A1(G217), .A2(G902), .ZN(new_n979));
  XNOR2_X1  g793(.A(new_n979), .B(KEYINPUT60), .ZN(new_n980));
  INV_X1    g794(.A(new_n980), .ZN(new_n981));
  AOI21_X1  g795(.A(new_n583), .B1(new_n933), .B2(new_n981), .ZN(new_n982));
  NOR2_X1   g796(.A1(new_n982), .A2(new_n950), .ZN(new_n983));
  NAND3_X1  g797(.A1(new_n933), .A2(new_n693), .A3(new_n981), .ZN(new_n984));
  NAND3_X1  g798(.A1(new_n983), .A2(KEYINPUT61), .A3(new_n984), .ZN(new_n985));
  INV_X1    g799(.A(KEYINPUT121), .ZN(new_n986));
  OAI21_X1  g800(.A(new_n986), .B1(new_n982), .B2(new_n950), .ZN(new_n987));
  AOI21_X1  g801(.A(new_n980), .B1(new_n946), .B2(new_n932), .ZN(new_n988));
  OAI211_X1 g802(.A(KEYINPUT121), .B(new_n951), .C1(new_n988), .C2(new_n583), .ZN(new_n989));
  INV_X1    g803(.A(KEYINPUT120), .ZN(new_n990));
  NAND2_X1  g804(.A1(new_n984), .A2(new_n990), .ZN(new_n991));
  NAND3_X1  g805(.A1(new_n988), .A2(KEYINPUT120), .A3(new_n693), .ZN(new_n992));
  NAND4_X1  g806(.A1(new_n987), .A2(new_n989), .A3(new_n991), .A4(new_n992), .ZN(new_n993));
  INV_X1    g807(.A(KEYINPUT61), .ZN(new_n994));
  AND3_X1   g808(.A1(new_n993), .A2(KEYINPUT122), .A3(new_n994), .ZN(new_n995));
  AOI21_X1  g809(.A(KEYINPUT122), .B1(new_n993), .B2(new_n994), .ZN(new_n996));
  OAI21_X1  g810(.A(new_n985), .B1(new_n995), .B2(new_n996), .ZN(G66));
  OAI21_X1  g811(.A(G953), .B1(new_n531), .B2(new_n323), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n930), .B2(G953), .ZN(new_n999));
  OAI21_X1  g813(.A(new_n939), .B1(G898), .B2(new_n528), .ZN(new_n1000));
  XNOR2_X1  g814(.A(new_n999), .B(new_n1000), .ZN(G69));
  AOI21_X1  g815(.A(new_n528), .B1(G227), .B2(G900), .ZN(new_n1002));
  AND2_X1   g816(.A1(new_n1002), .A2(KEYINPUT126), .ZN(new_n1003));
  INV_X1    g817(.A(KEYINPUT124), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n834), .A2(new_n841), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n886), .A2(new_n784), .ZN(new_n1006));
  INV_X1    g820(.A(KEYINPUT62), .ZN(new_n1007));
  OR3_X1    g821(.A1(new_n731), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  OAI21_X1  g822(.A(new_n1007), .B1(new_n731), .B2(new_n1006), .ZN(new_n1009));
  NAND2_X1  g823(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  AOI21_X1  g824(.A(new_n789), .B1(new_n674), .B2(new_n891), .ZN(new_n1011));
  NAND4_X1  g825(.A1(new_n316), .A2(new_n1011), .A3(new_n727), .A4(new_n598), .ZN(new_n1012));
  AND2_X1   g826(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1013));
  AOI21_X1  g827(.A(G953), .B1(new_n1005), .B2(new_n1013), .ZN(new_n1014));
  NOR2_X1   g828(.A1(new_n293), .A2(new_n294), .ZN(new_n1015));
  NAND2_X1  g829(.A1(new_n436), .A2(new_n437), .ZN(new_n1016));
  XNOR2_X1  g830(.A(new_n1015), .B(new_n1016), .ZN(new_n1017));
  XOR2_X1   g831(.A(new_n1017), .B(KEYINPUT123), .Z(new_n1018));
  OAI21_X1  g832(.A(new_n1004), .B1(new_n1014), .B2(new_n1018), .ZN(new_n1019));
  INV_X1    g833(.A(new_n1018), .ZN(new_n1020));
  NAND2_X1  g834(.A1(new_n1010), .A2(new_n1012), .ZN(new_n1021));
  NOR3_X1   g835(.A1(new_n1021), .A2(new_n834), .A3(new_n841), .ZN(new_n1022));
  OAI211_X1 g836(.A(KEYINPUT124), .B(new_n1020), .C1(new_n1022), .C2(G953), .ZN(new_n1023));
  AOI21_X1  g837(.A(new_n1003), .B1(new_n1019), .B2(new_n1023), .ZN(new_n1024));
  OR2_X1    g838(.A1(new_n1002), .A2(KEYINPUT126), .ZN(new_n1025));
  INV_X1    g839(.A(new_n1006), .ZN(new_n1026));
  NAND3_X1  g840(.A1(new_n1026), .A2(new_n800), .A3(new_n802), .ZN(new_n1027));
  NAND2_X1  g841(.A1(new_n827), .A2(new_n833), .ZN(new_n1028));
  AND2_X1   g842(.A1(new_n798), .A2(new_n878), .ZN(new_n1029));
  AOI21_X1  g843(.A(new_n1027), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  NAND2_X1  g844(.A1(new_n1005), .A2(new_n1030), .ZN(new_n1031));
  INV_X1    g845(.A(KEYINPUT125), .ZN(new_n1032));
  NAND2_X1  g846(.A1(new_n1031), .A2(new_n1032), .ZN(new_n1033));
  NAND3_X1  g847(.A1(new_n1005), .A2(KEYINPUT125), .A3(new_n1030), .ZN(new_n1034));
  NAND3_X1  g848(.A1(new_n1033), .A2(new_n528), .A3(new_n1034), .ZN(new_n1035));
  AOI21_X1  g849(.A(new_n1017), .B1(G900), .B2(G953), .ZN(new_n1036));
  NAND2_X1  g850(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  AND3_X1   g851(.A1(new_n1024), .A2(new_n1025), .A3(new_n1037), .ZN(new_n1038));
  AOI21_X1  g852(.A(new_n1025), .B1(new_n1024), .B2(new_n1037), .ZN(new_n1039));
  NOR2_X1   g853(.A1(new_n1038), .A2(new_n1039), .ZN(G72));
  INV_X1    g854(.A(KEYINPUT127), .ZN(new_n1041));
  NAND2_X1  g855(.A1(new_n302), .A2(new_n1041), .ZN(new_n1042));
  XOR2_X1   g856(.A(new_n1042), .B(new_n265), .Z(new_n1043));
  NAND2_X1  g857(.A1(G472), .A2(G902), .ZN(new_n1044));
  XOR2_X1   g858(.A(new_n1044), .B(KEYINPUT63), .Z(new_n1045));
  INV_X1    g859(.A(new_n1045), .ZN(new_n1046));
  NOR2_X1   g860(.A1(new_n1043), .A2(new_n1046), .ZN(new_n1047));
  AOI21_X1  g861(.A(new_n950), .B1(new_n925), .B2(new_n1047), .ZN(new_n1048));
  AOI21_X1  g862(.A(new_n1046), .B1(new_n1022), .B2(new_n930), .ZN(new_n1049));
  OAI21_X1  g863(.A(new_n1048), .B1(new_n1049), .B2(new_n719), .ZN(new_n1050));
  NAND3_X1  g864(.A1(new_n1033), .A2(new_n930), .A3(new_n1034), .ZN(new_n1051));
  NAND2_X1  g865(.A1(new_n1051), .A2(new_n1045), .ZN(new_n1052));
  NOR2_X1   g866(.A1(new_n296), .A2(new_n191), .ZN(new_n1053));
  AOI21_X1  g867(.A(new_n1050), .B1(new_n1052), .B2(new_n1053), .ZN(G57));
endmodule


