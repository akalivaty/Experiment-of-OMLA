//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 0 0 0 1 1 1 0 1 0 1 0 1 0 1 1 1 0 0 0 0 1 1 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 1 1 0 1 0 1 1 0 1 1 0 1 0 0 0 0 1 0 0 1 0 1 1 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:38:32 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n231,
    new_n232, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n240, new_n241, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1033,
    new_n1034, new_n1035, new_n1036, new_n1037, new_n1038, new_n1039,
    new_n1040, new_n1041, new_n1042, new_n1043, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1060, new_n1061, new_n1062, new_n1063, new_n1064,
    new_n1065, new_n1066, new_n1067, new_n1068, new_n1069, new_n1070,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1209, new_n1210, new_n1211,
    new_n1212, new_n1213, new_n1214, new_n1215, new_n1216, new_n1217,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1228, new_n1229, new_n1230,
    new_n1231, new_n1232, new_n1234, new_n1235, new_n1236, new_n1237,
    new_n1238, new_n1239, new_n1240, new_n1241, new_n1242, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1302, new_n1303, new_n1304,
    new_n1305, new_n1306, new_n1307, new_n1308, new_n1309, new_n1310,
    new_n1312, new_n1313, new_n1314, new_n1315, new_n1316, new_n1317,
    new_n1318;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(G50), .ZN(new_n202));
  NAND2_X1  g0002(.A1(new_n201), .A2(new_n202), .ZN(new_n203));
  NOR2_X1   g0003(.A1(new_n203), .A2(G77), .ZN(G353));
  OAI21_X1  g0004(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0005(.A(G1), .ZN(new_n206));
  INV_X1    g0006(.A(G20), .ZN(new_n207));
  NOR2_X1   g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  INV_X1    g0008(.A(new_n208), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n209), .A2(G13), .ZN(new_n210));
  OAI211_X1 g0010(.A(new_n210), .B(G250), .C1(G257), .C2(G264), .ZN(new_n211));
  XNOR2_X1  g0011(.A(new_n211), .B(KEYINPUT0), .ZN(new_n212));
  NAND3_X1  g0012(.A1(G1), .A2(G13), .A3(G20), .ZN(new_n213));
  INV_X1    g0013(.A(new_n201), .ZN(new_n214));
  NAND2_X1  g0014(.A1(new_n214), .A2(G50), .ZN(new_n215));
  AOI22_X1  g0015(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n216));
  INV_X1    g0016(.A(G68), .ZN(new_n217));
  INV_X1    g0017(.A(G238), .ZN(new_n218));
  INV_X1    g0018(.A(G87), .ZN(new_n219));
  INV_X1    g0019(.A(G250), .ZN(new_n220));
  OAI221_X1 g0020(.A(new_n216), .B1(new_n217), .B2(new_n218), .C1(new_n219), .C2(new_n220), .ZN(new_n221));
  AOI22_X1  g0021(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n222));
  INV_X1    g0022(.A(G77), .ZN(new_n223));
  INV_X1    g0023(.A(G244), .ZN(new_n224));
  INV_X1    g0024(.A(G107), .ZN(new_n225));
  INV_X1    g0025(.A(G264), .ZN(new_n226));
  OAI221_X1 g0026(.A(new_n222), .B1(new_n223), .B2(new_n224), .C1(new_n225), .C2(new_n226), .ZN(new_n227));
  OAI21_X1  g0027(.A(new_n209), .B1(new_n221), .B2(new_n227), .ZN(new_n228));
  OAI221_X1 g0028(.A(new_n212), .B1(new_n213), .B2(new_n215), .C1(KEYINPUT1), .C2(new_n228), .ZN(new_n229));
  AOI21_X1  g0029(.A(new_n229), .B1(KEYINPUT1), .B2(new_n228), .ZN(G361));
  XNOR2_X1  g0030(.A(G238), .B(G244), .ZN(new_n231));
  INV_X1    g0031(.A(G232), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(KEYINPUT2), .B(G226), .Z(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(G264), .B(G270), .Z(new_n236));
  XNOR2_X1  g0036(.A(G250), .B(G257), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n235), .B(new_n238), .ZN(G358));
  XNOR2_X1  g0039(.A(G68), .B(G77), .ZN(new_n240));
  INV_X1    g0040(.A(G58), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(KEYINPUT64), .B(G50), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XOR2_X1   g0044(.A(G87), .B(G97), .Z(new_n245));
  XOR2_X1   g0045(.A(G107), .B(G116), .Z(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XNOR2_X1  g0047(.A(new_n244), .B(new_n247), .ZN(G351));
  NOR2_X1   g0048(.A1(G20), .A2(G33), .ZN(new_n249));
  AOI22_X1  g0049(.A1(new_n203), .A2(G20), .B1(G150), .B2(new_n249), .ZN(new_n250));
  NAND2_X1  g0050(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n251));
  NAND2_X1  g0051(.A1(KEYINPUT68), .A2(G58), .ZN(new_n252));
  OAI211_X1 g0052(.A(new_n251), .B(KEYINPUT8), .C1(KEYINPUT67), .C2(new_n252), .ZN(new_n253));
  OR2_X1    g0053(.A1(new_n252), .A2(KEYINPUT8), .ZN(new_n254));
  NAND2_X1  g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  INV_X1    g0055(.A(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G33), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n257), .A2(G20), .ZN(new_n258));
  INV_X1    g0058(.A(new_n258), .ZN(new_n259));
  OAI21_X1  g0059(.A(new_n250), .B1(new_n256), .B2(new_n259), .ZN(new_n260));
  NAND3_X1  g0060(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G1), .A2(G13), .ZN(new_n262));
  NAND2_X1  g0062(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND3_X1  g0064(.A1(new_n206), .A2(G13), .A3(G20), .ZN(new_n265));
  NOR2_X1   g0065(.A1(new_n265), .A2(G50), .ZN(new_n266));
  AOI21_X1  g0066(.A(new_n263), .B1(new_n206), .B2(G20), .ZN(new_n267));
  AOI21_X1  g0067(.A(new_n266), .B1(new_n267), .B2(G50), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n264), .A2(new_n268), .ZN(new_n269));
  XOR2_X1   g0069(.A(new_n269), .B(KEYINPUT9), .Z(new_n270));
  AND2_X1   g0070(.A1(KEYINPUT3), .A2(G33), .ZN(new_n271));
  NOR2_X1   g0071(.A1(KEYINPUT3), .A2(G33), .ZN(new_n272));
  NOR3_X1   g0072(.A1(new_n271), .A2(new_n272), .A3(KEYINPUT66), .ZN(new_n273));
  INV_X1    g0073(.A(KEYINPUT66), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT3), .ZN(new_n275));
  NAND2_X1  g0075(.A1(new_n275), .A2(new_n257), .ZN(new_n276));
  NAND2_X1  g0076(.A1(KEYINPUT3), .A2(G33), .ZN(new_n277));
  AOI21_X1  g0077(.A(new_n274), .B1(new_n276), .B2(new_n277), .ZN(new_n278));
  NOR2_X1   g0078(.A1(new_n273), .A2(new_n278), .ZN(new_n279));
  INV_X1    g0079(.A(G1698), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n279), .A2(G222), .A3(new_n280), .ZN(new_n281));
  NAND3_X1  g0081(.A1(new_n279), .A2(G223), .A3(G1698), .ZN(new_n282));
  OAI211_X1 g0082(.A(new_n281), .B(new_n282), .C1(new_n223), .C2(new_n279), .ZN(new_n283));
  AOI21_X1  g0083(.A(new_n262), .B1(G33), .B2(G41), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  OAI21_X1  g0085(.A(new_n206), .B1(G41), .B2(G45), .ZN(new_n286));
  INV_X1    g0086(.A(G274), .ZN(new_n287));
  NOR2_X1   g0087(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  INV_X1    g0088(.A(KEYINPUT65), .ZN(new_n289));
  INV_X1    g0089(.A(G41), .ZN(new_n290));
  OAI211_X1 g0090(.A(G1), .B(G13), .C1(new_n257), .C2(new_n290), .ZN(new_n291));
  AOI21_X1  g0091(.A(new_n289), .B1(new_n291), .B2(new_n286), .ZN(new_n292));
  INV_X1    g0092(.A(new_n292), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n291), .A2(new_n289), .A3(new_n286), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  AOI21_X1  g0095(.A(new_n288), .B1(new_n295), .B2(G226), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n285), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(G200), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G190), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n297), .A2(new_n301), .ZN(new_n302));
  NOR3_X1   g0102(.A1(new_n270), .A2(new_n300), .A3(new_n302), .ZN(new_n303));
  INV_X1    g0103(.A(KEYINPUT10), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n303), .B(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(KEYINPUT72), .ZN(new_n306));
  INV_X1    g0106(.A(new_n294), .ZN(new_n307));
  OAI21_X1  g0107(.A(new_n306), .B1(new_n307), .B2(new_n292), .ZN(new_n308));
  NAND3_X1  g0108(.A1(new_n293), .A2(KEYINPUT72), .A3(new_n294), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n308), .A2(new_n309), .A3(G238), .ZN(new_n310));
  INV_X1    g0110(.A(KEYINPUT13), .ZN(new_n311));
  OAI21_X1  g0111(.A(KEYINPUT66), .B1(new_n271), .B2(new_n272), .ZN(new_n312));
  NAND3_X1  g0112(.A1(new_n276), .A2(new_n274), .A3(new_n277), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n312), .A2(new_n313), .ZN(new_n314));
  NAND2_X1  g0114(.A1(new_n232), .A2(G1698), .ZN(new_n315));
  OAI21_X1  g0115(.A(new_n315), .B1(G226), .B2(G1698), .ZN(new_n316));
  INV_X1    g0116(.A(G97), .ZN(new_n317));
  OAI22_X1  g0117(.A1(new_n314), .A2(new_n316), .B1(new_n257), .B2(new_n317), .ZN(new_n318));
  AOI21_X1  g0118(.A(new_n288), .B1(new_n318), .B2(new_n284), .ZN(new_n319));
  AND3_X1   g0119(.A1(new_n310), .A2(new_n311), .A3(new_n319), .ZN(new_n320));
  AOI21_X1  g0120(.A(new_n311), .B1(new_n310), .B2(new_n319), .ZN(new_n321));
  NOR3_X1   g0121(.A1(new_n320), .A2(new_n321), .A3(new_n301), .ZN(new_n322));
  NAND2_X1  g0122(.A1(new_n310), .A2(new_n319), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n323), .A2(KEYINPUT13), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n310), .A2(new_n311), .A3(new_n319), .ZN(new_n325));
  AOI21_X1  g0125(.A(new_n299), .B1(new_n324), .B2(new_n325), .ZN(new_n326));
  OAI22_X1  g0126(.A1(new_n259), .A2(new_n223), .B1(new_n207), .B2(G68), .ZN(new_n327));
  INV_X1    g0127(.A(new_n249), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n328), .A2(new_n202), .ZN(new_n329));
  OAI21_X1  g0129(.A(new_n263), .B1(new_n327), .B2(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT11), .ZN(new_n331));
  AND2_X1   g0131(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n330), .A2(new_n331), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n267), .A2(G68), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT12), .ZN(new_n335));
  INV_X1    g0135(.A(new_n265), .ZN(new_n336));
  AOI21_X1  g0136(.A(new_n335), .B1(new_n336), .B2(new_n217), .ZN(new_n337));
  NOR3_X1   g0137(.A1(new_n265), .A2(KEYINPUT12), .A3(G68), .ZN(new_n338));
  OAI21_X1  g0138(.A(new_n334), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  NOR3_X1   g0139(.A1(new_n332), .A2(new_n333), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n340), .ZN(new_n341));
  NOR3_X1   g0141(.A1(new_n322), .A2(new_n326), .A3(new_n341), .ZN(new_n342));
  OAI21_X1  g0142(.A(G169), .B1(new_n320), .B2(new_n321), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n343), .A2(KEYINPUT14), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT14), .ZN(new_n345));
  OAI211_X1 g0145(.A(new_n345), .B(G169), .C1(new_n320), .C2(new_n321), .ZN(new_n346));
  NAND3_X1  g0146(.A1(new_n324), .A2(G179), .A3(new_n325), .ZN(new_n347));
  NAND3_X1  g0147(.A1(new_n344), .A2(new_n346), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n342), .B1(new_n348), .B2(new_n341), .ZN(new_n349));
  INV_X1    g0149(.A(G169), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n297), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(new_n269), .ZN(new_n352));
  INV_X1    g0152(.A(G179), .ZN(new_n353));
  AOI21_X1  g0153(.A(new_n352), .B1(new_n353), .B2(new_n298), .ZN(new_n354));
  INV_X1    g0154(.A(new_n354), .ZN(new_n355));
  NAND3_X1  g0155(.A1(new_n305), .A2(new_n349), .A3(new_n355), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT67), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G58), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n251), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g0159(.A(new_n214), .B1(new_n359), .B2(new_n217), .ZN(new_n360));
  AOI22_X1  g0160(.A1(new_n360), .A2(G20), .B1(G159), .B2(new_n249), .ZN(new_n361));
  NAND3_X1  g0161(.A1(new_n276), .A2(new_n207), .A3(new_n277), .ZN(new_n362));
  INV_X1    g0162(.A(KEYINPUT73), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT7), .ZN(new_n364));
  AND3_X1   g0164(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  AOI21_X1  g0165(.A(new_n363), .B1(new_n362), .B2(new_n364), .ZN(new_n366));
  NOR2_X1   g0166(.A1(new_n362), .A2(new_n364), .ZN(new_n367));
  NOR3_X1   g0167(.A1(new_n365), .A2(new_n366), .A3(new_n367), .ZN(new_n368));
  OAI211_X1 g0168(.A(KEYINPUT16), .B(new_n361), .C1(new_n368), .C2(new_n217), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n251), .A2(new_n358), .ZN(new_n370));
  AOI21_X1  g0170(.A(new_n201), .B1(new_n370), .B2(G68), .ZN(new_n371));
  INV_X1    g0171(.A(G159), .ZN(new_n372));
  OAI22_X1  g0172(.A1(new_n371), .A2(new_n207), .B1(new_n372), .B2(new_n328), .ZN(new_n373));
  NOR3_X1   g0173(.A1(new_n271), .A2(new_n272), .A3(G20), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n374), .A2(KEYINPUT7), .ZN(new_n375));
  AOI21_X1  g0175(.A(G20), .B1(new_n312), .B2(new_n313), .ZN(new_n376));
  OAI21_X1  g0176(.A(new_n375), .B1(new_n376), .B2(KEYINPUT7), .ZN(new_n377));
  AOI21_X1  g0177(.A(new_n373), .B1(new_n377), .B2(G68), .ZN(new_n378));
  OAI211_X1 g0178(.A(new_n369), .B(new_n263), .C1(KEYINPUT16), .C2(new_n378), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n256), .A2(new_n336), .ZN(new_n380));
  NAND2_X1  g0180(.A1(new_n255), .A2(new_n267), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  INV_X1    g0182(.A(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n276), .A2(new_n277), .ZN(new_n384));
  OR2_X1    g0184(.A1(new_n280), .A2(G226), .ZN(new_n385));
  OAI211_X1 g0185(.A(new_n384), .B(new_n385), .C1(G223), .C2(G1698), .ZN(new_n386));
  NAND2_X1  g0186(.A1(G33), .A2(G87), .ZN(new_n387));
  AOI21_X1  g0187(.A(new_n291), .B1(new_n386), .B2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(new_n288), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n291), .A2(new_n286), .ZN(new_n390));
  OAI21_X1  g0190(.A(new_n389), .B1(new_n390), .B2(new_n232), .ZN(new_n391));
  NOR3_X1   g0191(.A1(new_n388), .A2(new_n301), .A3(new_n391), .ZN(new_n392));
  OR2_X1    g0192(.A1(new_n388), .A2(new_n391), .ZN(new_n393));
  AOI21_X1  g0193(.A(new_n392), .B1(new_n393), .B2(G200), .ZN(new_n394));
  NAND4_X1  g0194(.A1(new_n379), .A2(KEYINPUT74), .A3(new_n383), .A4(new_n394), .ZN(new_n395));
  XNOR2_X1  g0195(.A(new_n395), .B(KEYINPUT17), .ZN(new_n396));
  INV_X1    g0196(.A(new_n263), .ZN(new_n397));
  OAI21_X1  g0197(.A(KEYINPUT73), .B1(new_n374), .B2(KEYINPUT7), .ZN(new_n398));
  NAND3_X1  g0198(.A1(new_n362), .A2(new_n363), .A3(new_n364), .ZN(new_n399));
  NAND3_X1  g0199(.A1(new_n398), .A2(new_n375), .A3(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n373), .B1(new_n400), .B2(G68), .ZN(new_n401));
  AOI21_X1  g0201(.A(new_n397), .B1(new_n401), .B2(KEYINPUT16), .ZN(new_n402));
  OAI21_X1  g0202(.A(new_n207), .B1(new_n273), .B2(new_n278), .ZN(new_n403));
  AOI21_X1  g0203(.A(new_n367), .B1(new_n403), .B2(new_n364), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n361), .B1(new_n404), .B2(new_n217), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT16), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n382), .B1(new_n402), .B2(new_n407), .ZN(new_n408));
  NOR3_X1   g0208(.A1(new_n388), .A2(new_n353), .A3(new_n391), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n409), .B1(new_n393), .B2(G169), .ZN(new_n410));
  OAI21_X1  g0210(.A(KEYINPUT18), .B1(new_n408), .B2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n369), .A2(new_n263), .ZN(new_n412));
  NOR2_X1   g0212(.A1(new_n378), .A2(KEYINPUT16), .ZN(new_n413));
  OAI21_X1  g0213(.A(new_n383), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g0214(.A(KEYINPUT18), .ZN(new_n415));
  INV_X1    g0215(.A(new_n410), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n414), .A2(new_n415), .A3(new_n416), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n396), .A2(new_n411), .A3(new_n417), .ZN(new_n418));
  INV_X1    g0218(.A(KEYINPUT71), .ZN(new_n419));
  NAND4_X1  g0219(.A1(new_n312), .A2(new_n313), .A3(G232), .A4(new_n280), .ZN(new_n420));
  INV_X1    g0220(.A(KEYINPUT69), .ZN(new_n421));
  XNOR2_X1  g0221(.A(new_n420), .B(new_n421), .ZN(new_n422));
  OAI21_X1  g0222(.A(G107), .B1(new_n273), .B2(new_n278), .ZN(new_n423));
  NAND4_X1  g0223(.A1(new_n312), .A2(new_n313), .A3(G238), .A4(G1698), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n423), .A2(new_n424), .ZN(new_n425));
  OAI21_X1  g0225(.A(new_n284), .B1(new_n422), .B2(new_n425), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n288), .B1(new_n295), .B2(G244), .ZN(new_n427));
  AOI21_X1  g0227(.A(G169), .B1(new_n426), .B2(new_n427), .ZN(new_n428));
  NAND2_X1  g0228(.A1(new_n267), .A2(G77), .ZN(new_n429));
  NAND2_X1  g0229(.A1(new_n336), .A2(new_n223), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  XNOR2_X1  g0231(.A(KEYINPUT8), .B(G58), .ZN(new_n432));
  INV_X1    g0232(.A(new_n432), .ZN(new_n433));
  AOI22_X1  g0233(.A1(new_n433), .A2(new_n249), .B1(G20), .B2(G77), .ZN(new_n434));
  XNOR2_X1  g0234(.A(KEYINPUT15), .B(G87), .ZN(new_n435));
  XNOR2_X1  g0235(.A(new_n435), .B(KEYINPUT70), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n434), .B1(new_n436), .B2(new_n259), .ZN(new_n437));
  AOI21_X1  g0237(.A(new_n431), .B1(new_n437), .B2(new_n263), .ZN(new_n438));
  OAI21_X1  g0238(.A(new_n419), .B1(new_n428), .B2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n279), .A2(new_n421), .A3(G232), .A4(new_n280), .ZN(new_n440));
  NAND2_X1  g0240(.A1(new_n420), .A2(KEYINPUT69), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n425), .B1(new_n440), .B2(new_n441), .ZN(new_n442));
  OAI21_X1  g0242(.A(new_n427), .B1(new_n442), .B2(new_n291), .ZN(new_n443));
  AOI21_X1  g0243(.A(new_n438), .B1(new_n443), .B2(new_n350), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT71), .ZN(new_n445));
  INV_X1    g0245(.A(new_n427), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n440), .A2(new_n441), .ZN(new_n447));
  INV_X1    g0247(.A(new_n425), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n446), .B1(new_n449), .B2(new_n284), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n450), .A2(new_n353), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n439), .A2(new_n445), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(new_n438), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n443), .B2(G200), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n454), .B1(new_n301), .B2(new_n443), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n356), .A2(new_n418), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(new_n457), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n265), .A2(G97), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n206), .A2(G33), .ZN(new_n460));
  NAND3_X1  g0260(.A1(new_n397), .A2(new_n265), .A3(new_n460), .ZN(new_n461));
  INV_X1    g0261(.A(new_n461), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n462), .B2(G97), .ZN(new_n463));
  NOR2_X1   g0263(.A1(KEYINPUT75), .A2(KEYINPUT6), .ZN(new_n464));
  AND2_X1   g0264(.A1(G97), .A2(G107), .ZN(new_n465));
  NOR2_X1   g0265(.A1(G97), .A2(G107), .ZN(new_n466));
  OAI21_X1  g0266(.A(new_n464), .B1(new_n465), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n317), .A2(KEYINPUT6), .ZN(new_n468));
  OAI21_X1  g0268(.A(new_n468), .B1(KEYINPUT75), .B2(KEYINPUT6), .ZN(new_n469));
  XNOR2_X1  g0269(.A(G97), .B(G107), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n467), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n471), .A2(G20), .ZN(new_n472));
  NAND2_X1  g0272(.A1(new_n249), .A2(G77), .ZN(new_n473));
  NAND2_X1  g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n474), .B1(G107), .B2(new_n377), .ZN(new_n475));
  OAI21_X1  g0275(.A(new_n463), .B1(new_n475), .B2(new_n397), .ZN(new_n476));
  OAI211_X1 g0276(.A(G244), .B(new_n280), .C1(new_n271), .C2(new_n272), .ZN(new_n477));
  INV_X1    g0277(.A(KEYINPUT4), .ZN(new_n478));
  AOI22_X1  g0278(.A1(new_n477), .A2(new_n478), .B1(G33), .B2(G283), .ZN(new_n479));
  NAND4_X1  g0279(.A1(new_n312), .A2(new_n313), .A3(G250), .A4(G1698), .ZN(new_n480));
  NOR2_X1   g0280(.A1(new_n478), .A2(new_n224), .ZN(new_n481));
  NAND4_X1  g0281(.A1(new_n312), .A2(new_n313), .A3(new_n280), .A4(new_n481), .ZN(new_n482));
  NAND3_X1  g0282(.A1(new_n479), .A2(new_n480), .A3(new_n482), .ZN(new_n483));
  INV_X1    g0283(.A(KEYINPUT76), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NAND4_X1  g0285(.A1(new_n479), .A2(new_n480), .A3(new_n482), .A4(KEYINPUT76), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(new_n486), .A3(new_n284), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n206), .A2(G45), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT5), .A2(G41), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  NAND2_X1  g0290(.A1(KEYINPUT5), .A2(G41), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n488), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND3_X1  g0292(.A1(new_n492), .A2(G274), .A3(new_n291), .ZN(new_n493));
  INV_X1    g0293(.A(G45), .ZN(new_n494));
  NOR2_X1   g0294(.A1(new_n494), .A2(G1), .ZN(new_n495));
  INV_X1    g0295(.A(new_n491), .ZN(new_n496));
  OAI21_X1  g0296(.A(new_n495), .B1(new_n496), .B2(new_n489), .ZN(new_n497));
  NAND3_X1  g0297(.A1(new_n497), .A2(G257), .A3(new_n291), .ZN(new_n498));
  NAND2_X1  g0298(.A1(new_n493), .A2(new_n498), .ZN(new_n499));
  INV_X1    g0299(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g0300(.A1(new_n487), .A2(new_n353), .A3(new_n500), .ZN(new_n501));
  AOI21_X1  g0301(.A(new_n291), .B1(new_n483), .B2(new_n484), .ZN(new_n502));
  AOI21_X1  g0302(.A(new_n499), .B1(new_n502), .B2(new_n486), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n476), .B(new_n501), .C1(G169), .C2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n487), .A2(G190), .A3(new_n500), .ZN(new_n505));
  INV_X1    g0305(.A(new_n463), .ZN(new_n506));
  AOI22_X1  g0306(.A1(new_n471), .A2(G20), .B1(G77), .B2(new_n249), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n404), .B2(new_n225), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n506), .B1(new_n508), .B2(new_n263), .ZN(new_n509));
  OAI211_X1 g0309(.A(new_n505), .B(new_n509), .C1(new_n299), .C2(new_n503), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n218), .A2(new_n280), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n224), .A2(G1698), .ZN(new_n512));
  OAI211_X1 g0312(.A(new_n511), .B(new_n512), .C1(new_n271), .C2(new_n272), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G116), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n291), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n488), .A2(G250), .ZN(new_n516));
  OAI22_X1  g0316(.A1(new_n284), .A2(new_n516), .B1(new_n287), .B2(new_n488), .ZN(new_n517));
  OR4_X1    g0317(.A1(KEYINPUT78), .A2(new_n515), .A3(new_n301), .A4(new_n517), .ZN(new_n518));
  NOR2_X1   g0318(.A1(new_n495), .A2(new_n220), .ZN(new_n519));
  AOI22_X1  g0319(.A1(new_n519), .A2(new_n291), .B1(G274), .B2(new_n495), .ZN(new_n520));
  NOR2_X1   g0320(.A1(G238), .A2(G1698), .ZN(new_n521));
  AOI21_X1  g0321(.A(new_n521), .B1(new_n224), .B2(G1698), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n522), .A2(new_n384), .B1(G33), .B2(G116), .ZN(new_n523));
  OAI21_X1  g0323(.A(new_n520), .B1(new_n523), .B2(new_n291), .ZN(new_n524));
  OAI21_X1  g0324(.A(KEYINPUT78), .B1(new_n524), .B2(new_n301), .ZN(new_n525));
  AOI22_X1  g0325(.A1(new_n518), .A2(new_n525), .B1(G200), .B2(new_n524), .ZN(new_n526));
  NAND3_X1  g0326(.A1(new_n384), .A2(new_n207), .A3(G68), .ZN(new_n527));
  NAND2_X1  g0327(.A1(new_n527), .A2(KEYINPUT77), .ZN(new_n528));
  INV_X1    g0328(.A(KEYINPUT19), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n258), .A2(new_n529), .A3(G97), .ZN(new_n530));
  AOI21_X1  g0330(.A(G20), .B1(G33), .B2(G97), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n219), .B2(new_n466), .ZN(new_n532));
  OAI21_X1  g0332(.A(new_n530), .B1(new_n532), .B2(new_n529), .ZN(new_n533));
  INV_X1    g0333(.A(KEYINPUT77), .ZN(new_n534));
  NAND4_X1  g0334(.A1(new_n384), .A2(new_n534), .A3(new_n207), .A4(G68), .ZN(new_n535));
  NAND3_X1  g0335(.A1(new_n528), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n536), .A2(new_n263), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n436), .A2(new_n336), .ZN(new_n538));
  NAND2_X1  g0338(.A1(new_n462), .A2(G87), .ZN(new_n539));
  AND3_X1   g0339(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  NOR2_X1   g0340(.A1(new_n524), .A2(G179), .ZN(new_n541));
  AOI21_X1  g0341(.A(new_n541), .B1(new_n350), .B2(new_n524), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n537), .B(new_n538), .C1(new_n461), .C2(new_n436), .ZN(new_n543));
  AOI22_X1  g0343(.A1(new_n526), .A2(new_n540), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n504), .A2(new_n510), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(G116), .ZN(new_n546));
  NAND2_X1  g0346(.A1(new_n336), .A2(new_n546), .ZN(new_n547));
  NAND4_X1  g0347(.A1(new_n397), .A2(G116), .A3(new_n265), .A4(new_n460), .ZN(new_n548));
  AOI22_X1  g0348(.A1(new_n261), .A2(new_n262), .B1(G20), .B2(new_n546), .ZN(new_n549));
  NAND2_X1  g0349(.A1(G33), .A2(G283), .ZN(new_n550));
  OAI211_X1 g0350(.A(new_n550), .B(new_n207), .C1(G33), .C2(new_n317), .ZN(new_n551));
  AND3_X1   g0351(.A1(new_n549), .A2(KEYINPUT20), .A3(new_n551), .ZN(new_n552));
  AOI21_X1  g0352(.A(KEYINPUT20), .B1(new_n549), .B2(new_n551), .ZN(new_n553));
  OAI211_X1 g0353(.A(new_n547), .B(new_n548), .C1(new_n552), .C2(new_n553), .ZN(new_n554));
  OAI21_X1  g0354(.A(G303), .B1(new_n273), .B2(new_n278), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n226), .A2(G1698), .ZN(new_n556));
  OAI221_X1 g0356(.A(new_n556), .B1(G257), .B2(G1698), .C1(new_n271), .C2(new_n272), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n291), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND3_X1  g0358(.A1(new_n497), .A2(G270), .A3(new_n291), .ZN(new_n559));
  NAND2_X1  g0359(.A1(new_n493), .A2(new_n559), .ZN(new_n560));
  OAI211_X1 g0360(.A(new_n554), .B(G169), .C1(new_n558), .C2(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(KEYINPUT21), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(new_n560), .ZN(new_n564));
  INV_X1    g0364(.A(G303), .ZN(new_n565));
  AOI21_X1  g0365(.A(new_n565), .B1(new_n312), .B2(new_n313), .ZN(new_n566));
  INV_X1    g0366(.A(new_n557), .ZN(new_n567));
  OAI21_X1  g0367(.A(new_n284), .B1(new_n566), .B2(new_n567), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n564), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n569), .A2(KEYINPUT21), .A3(G169), .A4(new_n554), .ZN(new_n570));
  NOR2_X1   g0370(.A1(new_n558), .A2(new_n560), .ZN(new_n571));
  NAND3_X1  g0371(.A1(new_n571), .A2(G179), .A3(new_n554), .ZN(new_n572));
  AND3_X1   g0372(.A1(new_n563), .A2(new_n570), .A3(new_n572), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n497), .A2(G264), .A3(new_n291), .ZN(new_n574));
  MUX2_X1   g0374(.A(G250), .B(G257), .S(G1698), .Z(new_n575));
  AOI22_X1  g0375(.A1(new_n575), .A2(new_n384), .B1(G33), .B2(G294), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n493), .B(new_n574), .C1(new_n576), .C2(new_n291), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(G179), .ZN(new_n578));
  AOI21_X1  g0378(.A(new_n578), .B1(new_n350), .B2(new_n577), .ZN(new_n579));
  OAI211_X1 g0379(.A(new_n207), .B(G87), .C1(new_n271), .C2(new_n272), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(KEYINPUT22), .ZN(new_n581));
  OR3_X1    g0381(.A1(new_n219), .A2(KEYINPUT22), .A3(G20), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n581), .B1(new_n314), .B2(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n225), .A2(G20), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n584), .A2(KEYINPUT79), .A3(KEYINPUT23), .ZN(new_n585));
  INV_X1    g0385(.A(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n207), .A2(G33), .A3(G116), .ZN(new_n587));
  OAI21_X1  g0387(.A(new_n587), .B1(new_n584), .B2(KEYINPUT23), .ZN(new_n588));
  AOI21_X1  g0388(.A(KEYINPUT79), .B1(new_n584), .B2(KEYINPUT23), .ZN(new_n589));
  NOR3_X1   g0389(.A1(new_n586), .A2(new_n588), .A3(new_n589), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n583), .A2(new_n590), .ZN(new_n591));
  NAND2_X1  g0391(.A1(new_n591), .A2(KEYINPUT24), .ZN(new_n592));
  INV_X1    g0392(.A(KEYINPUT24), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n583), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  AOI21_X1  g0394(.A(new_n397), .B1(new_n592), .B2(new_n594), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT25), .ZN(new_n596));
  NOR3_X1   g0396(.A1(new_n265), .A2(new_n596), .A3(G107), .ZN(new_n597));
  INV_X1    g0397(.A(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(new_n596), .B1(new_n265), .B2(G107), .ZN(new_n599));
  AOI22_X1  g0399(.A1(new_n462), .A2(G107), .B1(new_n598), .B2(new_n599), .ZN(new_n600));
  INV_X1    g0400(.A(new_n600), .ZN(new_n601));
  OAI21_X1  g0401(.A(new_n579), .B1(new_n595), .B2(new_n601), .ZN(new_n602));
  AND3_X1   g0402(.A1(new_n583), .A2(new_n590), .A3(new_n593), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n593), .B1(new_n583), .B2(new_n590), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n263), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n575), .A2(new_n384), .ZN(new_n606));
  NAND2_X1  g0406(.A1(G33), .A2(G294), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n606), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g0408(.A1(new_n608), .A2(new_n284), .ZN(new_n609));
  NAND4_X1  g0409(.A1(new_n609), .A2(G190), .A3(new_n493), .A4(new_n574), .ZN(new_n610));
  NAND2_X1  g0410(.A1(new_n577), .A2(G200), .ZN(new_n611));
  NAND4_X1  g0411(.A1(new_n605), .A2(new_n600), .A3(new_n610), .A4(new_n611), .ZN(new_n612));
  NAND3_X1  g0412(.A1(new_n564), .A2(new_n568), .A3(G190), .ZN(new_n613));
  INV_X1    g0413(.A(new_n554), .ZN(new_n614));
  OAI211_X1 g0414(.A(new_n613), .B(new_n614), .C1(new_n571), .C2(new_n299), .ZN(new_n615));
  NAND4_X1  g0415(.A1(new_n573), .A2(new_n602), .A3(new_n612), .A4(new_n615), .ZN(new_n616));
  NOR3_X1   g0416(.A1(new_n458), .A2(new_n545), .A3(new_n616), .ZN(G372));
  NAND2_X1  g0417(.A1(new_n577), .A2(new_n350), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(G179), .B2(new_n577), .ZN(new_n619));
  AOI21_X1  g0419(.A(new_n619), .B1(new_n605), .B2(new_n600), .ZN(new_n620));
  XNOR2_X1  g0420(.A(new_n620), .B(KEYINPUT80), .ZN(new_n621));
  INV_X1    g0421(.A(new_n573), .ZN(new_n622));
  NOR2_X1   g0422(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AND2_X1   g0423(.A1(new_n504), .A2(new_n510), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n624), .A2(new_n544), .A3(new_n612), .ZN(new_n625));
  NOR2_X1   g0425(.A1(new_n623), .A2(new_n625), .ZN(new_n626));
  INV_X1    g0426(.A(new_n504), .ZN(new_n627));
  NAND2_X1  g0427(.A1(new_n627), .A2(new_n544), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n628), .A2(KEYINPUT26), .ZN(new_n629));
  NAND2_X1  g0429(.A1(new_n542), .A2(new_n543), .ZN(new_n630));
  XNOR2_X1  g0430(.A(KEYINPUT81), .B(KEYINPUT26), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n627), .A2(new_n544), .A3(new_n631), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n629), .A2(new_n630), .A3(new_n632), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n457), .B1(new_n626), .B2(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n348), .A2(new_n341), .ZN(new_n635));
  OAI21_X1  g0435(.A(new_n635), .B1(new_n452), .B2(new_n342), .ZN(new_n636));
  OR2_X1    g0436(.A1(new_n636), .A2(KEYINPUT83), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT17), .ZN(new_n638));
  XNOR2_X1  g0438(.A(new_n395), .B(new_n638), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n636), .B2(KEYINPUT83), .ZN(new_n640));
  AND2_X1   g0440(.A1(new_n637), .A2(new_n640), .ZN(new_n641));
  AND3_X1   g0441(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT82), .ZN(new_n642));
  AOI21_X1  g0442(.A(KEYINPUT82), .B1(new_n411), .B2(new_n417), .ZN(new_n643));
  NOR2_X1   g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g0444(.A(new_n644), .ZN(new_n645));
  OAI21_X1  g0445(.A(new_n305), .B1(new_n641), .B2(new_n645), .ZN(new_n646));
  NAND3_X1  g0446(.A1(new_n634), .A2(new_n355), .A3(new_n646), .ZN(G369));
  INV_X1    g0447(.A(G13), .ZN(new_n648));
  NOR3_X1   g0448(.A1(new_n648), .A2(G1), .A3(G20), .ZN(new_n649));
  INV_X1    g0449(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g0450(.A(G213), .B1(new_n650), .B2(KEYINPUT27), .ZN(new_n651));
  AOI21_X1  g0451(.A(KEYINPUT84), .B1(new_n650), .B2(KEYINPUT27), .ZN(new_n652));
  INV_X1    g0452(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g0453(.A1(new_n650), .A2(KEYINPUT84), .A3(KEYINPUT27), .ZN(new_n654));
  AOI21_X1  g0454(.A(new_n651), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n655), .A2(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n656), .A2(new_n614), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n622), .A2(new_n657), .ZN(new_n658));
  NAND4_X1  g0458(.A1(new_n615), .A2(new_n563), .A3(new_n570), .A4(new_n572), .ZN(new_n659));
  OAI21_X1  g0459(.A(new_n658), .B1(new_n659), .B2(new_n657), .ZN(new_n660));
  XNOR2_X1  g0460(.A(new_n660), .B(KEYINPUT85), .ZN(new_n661));
  NAND2_X1  g0461(.A1(new_n661), .A2(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n656), .ZN(new_n663));
  OAI21_X1  g0463(.A(new_n663), .B1(new_n595), .B2(new_n601), .ZN(new_n664));
  NAND3_X1  g0464(.A1(new_n602), .A2(new_n664), .A3(new_n612), .ZN(new_n665));
  XOR2_X1   g0465(.A(new_n665), .B(KEYINPUT86), .Z(new_n666));
  AOI21_X1  g0466(.A(new_n666), .B1(new_n620), .B2(new_n663), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n662), .A2(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n573), .A2(new_n663), .ZN(new_n669));
  NAND2_X1  g0469(.A1(new_n666), .A2(new_n669), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n621), .A2(new_n656), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OR2_X1    g0472(.A1(new_n668), .A2(new_n672), .ZN(G399));
  INV_X1    g0473(.A(new_n210), .ZN(new_n674));
  NOR2_X1   g0474(.A1(new_n674), .A2(G41), .ZN(new_n675));
  NAND3_X1  g0475(.A1(new_n466), .A2(new_n219), .A3(new_n546), .ZN(new_n676));
  NOR3_X1   g0476(.A1(new_n675), .A2(new_n206), .A3(new_n676), .ZN(new_n677));
  INV_X1    g0477(.A(new_n215), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n677), .B1(new_n678), .B2(new_n675), .ZN(new_n679));
  XOR2_X1   g0479(.A(new_n679), .B(KEYINPUT28), .Z(new_n680));
  INV_X1    g0480(.A(KEYINPUT89), .ZN(new_n681));
  NOR3_X1   g0481(.A1(new_n558), .A2(new_n353), .A3(new_n560), .ZN(new_n682));
  OAI21_X1  g0482(.A(new_n574), .B1(new_n576), .B2(new_n291), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n683), .A2(new_n524), .ZN(new_n684));
  NAND4_X1  g0484(.A1(new_n487), .A2(new_n682), .A3(new_n500), .A4(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(KEYINPUT30), .ZN(new_n686));
  NAND2_X1  g0486(.A1(new_n487), .A2(new_n500), .ZN(new_n687));
  OAI211_X1 g0487(.A(KEYINPUT87), .B(new_n520), .C1(new_n523), .C2(new_n291), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT87), .ZN(new_n689));
  OAI21_X1  g0489(.A(new_n689), .B1(new_n515), .B2(new_n517), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n577), .A2(new_n688), .A3(new_n690), .A4(new_n353), .ZN(new_n691));
  NOR2_X1   g0491(.A1(new_n691), .A2(new_n571), .ZN(new_n692));
  AOI22_X1  g0492(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n692), .ZN(new_n693));
  NAND4_X1  g0493(.A1(new_n503), .A2(KEYINPUT30), .A3(new_n682), .A4(new_n684), .ZN(new_n694));
  AOI21_X1  g0494(.A(new_n656), .B1(new_n693), .B2(new_n694), .ZN(new_n695));
  INV_X1    g0495(.A(new_n695), .ZN(new_n696));
  NOR3_X1   g0496(.A1(new_n545), .A2(new_n616), .A3(new_n663), .ZN(new_n697));
  INV_X1    g0497(.A(KEYINPUT31), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n696), .B1(new_n697), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g0499(.A(KEYINPUT88), .B1(new_n695), .B2(KEYINPUT31), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n686), .ZN(new_n701));
  NAND2_X1  g0501(.A1(new_n687), .A2(new_n692), .ZN(new_n702));
  NAND3_X1  g0502(.A1(new_n701), .A2(new_n694), .A3(new_n702), .ZN(new_n703));
  AND4_X1   g0503(.A1(KEYINPUT88), .A2(new_n703), .A3(KEYINPUT31), .A4(new_n663), .ZN(new_n704));
  NOR2_X1   g0504(.A1(new_n700), .A2(new_n704), .ZN(new_n705));
  NAND2_X1  g0505(.A1(new_n699), .A2(new_n705), .ZN(new_n706));
  AOI21_X1  g0506(.A(new_n681), .B1(new_n706), .B2(G330), .ZN(new_n707));
  INV_X1    g0507(.A(G330), .ZN(new_n708));
  AOI211_X1 g0508(.A(KEYINPUT89), .B(new_n708), .C1(new_n699), .C2(new_n705), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n707), .A2(new_n709), .ZN(new_n710));
  OAI21_X1  g0510(.A(new_n656), .B1(new_n626), .B2(new_n633), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n625), .B1(new_n602), .B2(new_n573), .ZN(new_n714));
  INV_X1    g0514(.A(new_n631), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n628), .A2(new_n715), .ZN(new_n716));
  OAI211_X1 g0516(.A(new_n716), .B(new_n630), .C1(KEYINPUT26), .C2(new_n628), .ZN(new_n717));
  OAI211_X1 g0517(.A(KEYINPUT29), .B(new_n656), .C1(new_n714), .C2(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n713), .A2(new_n718), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n710), .A2(new_n719), .ZN(new_n720));
  INV_X1    g0520(.A(new_n720), .ZN(new_n721));
  OAI21_X1  g0521(.A(new_n680), .B1(new_n721), .B2(G1), .ZN(G364));
  NOR2_X1   g0522(.A1(new_n648), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n206), .B1(new_n723), .B2(G45), .ZN(new_n724));
  INV_X1    g0524(.A(new_n724), .ZN(new_n725));
  OR3_X1    g0525(.A1(new_n675), .A2(KEYINPUT90), .A3(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(KEYINPUT90), .B1(new_n675), .B2(new_n725), .ZN(new_n727));
  NAND2_X1  g0527(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  INV_X1    g0528(.A(new_n728), .ZN(new_n729));
  AOI21_X1  g0529(.A(new_n729), .B1(new_n661), .B2(G330), .ZN(new_n730));
  OAI21_X1  g0530(.A(new_n730), .B1(G330), .B2(new_n661), .ZN(new_n731));
  NOR2_X1   g0531(.A1(new_n674), .A2(new_n314), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G355), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n733), .B1(G116), .B2(new_n210), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n244), .A2(G45), .ZN(new_n735));
  NOR2_X1   g0535(.A1(new_n674), .A2(new_n384), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n737), .B1(new_n494), .B2(new_n678), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n734), .B1(new_n735), .B2(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(G13), .A2(G33), .ZN(new_n740));
  XNOR2_X1  g0540(.A(new_n740), .B(KEYINPUT91), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n741), .A2(G20), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n262), .B1(G20), .B2(new_n350), .ZN(new_n743));
  NOR2_X1   g0543(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  OAI21_X1  g0545(.A(new_n729), .B1(new_n739), .B2(new_n745), .ZN(new_n746));
  OR3_X1    g0546(.A1(new_n207), .A2(KEYINPUT93), .A3(G190), .ZN(new_n747));
  NOR2_X1   g0547(.A1(G179), .A2(G200), .ZN(new_n748));
  OAI21_X1  g0548(.A(KEYINPUT93), .B1(new_n207), .B2(G190), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n747), .A2(new_n748), .A3(new_n749), .ZN(new_n750));
  XNOR2_X1  g0550(.A(KEYINPUT94), .B(G159), .ZN(new_n751));
  NOR2_X1   g0551(.A1(new_n750), .A2(new_n751), .ZN(new_n752));
  XNOR2_X1  g0552(.A(new_n752), .B(KEYINPUT95), .ZN(new_n753));
  OR2_X1    g0553(.A1(new_n753), .A2(KEYINPUT32), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n753), .A2(KEYINPUT32), .ZN(new_n755));
  AOI21_X1  g0555(.A(new_n207), .B1(new_n748), .B2(G190), .ZN(new_n756));
  XNOR2_X1  g0556(.A(new_n756), .B(KEYINPUT96), .ZN(new_n757));
  NAND2_X1  g0557(.A1(new_n757), .A2(G97), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n353), .A2(new_n299), .ZN(new_n759));
  NAND2_X1  g0559(.A1(G20), .A2(G190), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  AND3_X1   g0561(.A1(new_n759), .A2(KEYINPUT92), .A3(new_n761), .ZN(new_n762));
  AOI21_X1  g0562(.A(KEYINPUT92), .B1(new_n759), .B2(new_n761), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n299), .A2(G179), .ZN(new_n765));
  NAND3_X1  g0565(.A1(new_n747), .A2(new_n765), .A3(new_n749), .ZN(new_n766));
  OAI22_X1  g0566(.A1(new_n764), .A2(new_n202), .B1(new_n225), .B2(new_n766), .ZN(new_n767));
  NOR2_X1   g0567(.A1(new_n207), .A2(G190), .ZN(new_n768));
  AND2_X1   g0568(.A1(new_n759), .A2(new_n768), .ZN(new_n769));
  INV_X1    g0569(.A(new_n769), .ZN(new_n770));
  NOR3_X1   g0570(.A1(new_n760), .A2(new_n353), .A3(G200), .ZN(new_n771));
  INV_X1    g0571(.A(new_n771), .ZN(new_n772));
  OAI22_X1  g0572(.A1(new_n770), .A2(new_n217), .B1(new_n359), .B2(new_n772), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n353), .A2(G200), .ZN(new_n774));
  NAND2_X1  g0574(.A1(new_n774), .A2(new_n768), .ZN(new_n775));
  NAND2_X1  g0575(.A1(new_n765), .A2(new_n761), .ZN(new_n776));
  OAI22_X1  g0576(.A1(new_n775), .A2(new_n223), .B1(new_n776), .B2(new_n219), .ZN(new_n777));
  NOR4_X1   g0577(.A1(new_n767), .A2(new_n773), .A3(new_n314), .A4(new_n777), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n754), .A2(new_n755), .A3(new_n758), .A4(new_n778), .ZN(new_n779));
  INV_X1    g0579(.A(G311), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n775), .A2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(G317), .ZN(new_n782));
  AND2_X1   g0582(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n783));
  NOR2_X1   g0583(.A1(new_n782), .A2(KEYINPUT33), .ZN(new_n784));
  NOR3_X1   g0584(.A1(new_n770), .A2(new_n783), .A3(new_n784), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n781), .B(new_n785), .C1(G322), .C2(new_n771), .ZN(new_n786));
  INV_X1    g0586(.A(new_n756), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n279), .B1(G294), .B2(new_n787), .ZN(new_n788));
  INV_X1    g0588(.A(new_n764), .ZN(new_n789));
  INV_X1    g0589(.A(new_n766), .ZN(new_n790));
  AOI22_X1  g0590(.A1(new_n789), .A2(G326), .B1(G283), .B2(new_n790), .ZN(new_n791));
  XNOR2_X1  g0591(.A(new_n776), .B(KEYINPUT97), .ZN(new_n792));
  INV_X1    g0592(.A(new_n750), .ZN(new_n793));
  AOI22_X1  g0593(.A1(new_n792), .A2(G303), .B1(G329), .B2(new_n793), .ZN(new_n794));
  NAND4_X1  g0594(.A1(new_n786), .A2(new_n788), .A3(new_n791), .A4(new_n794), .ZN(new_n795));
  NAND2_X1  g0595(.A1(new_n779), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g0596(.A(new_n746), .B1(new_n796), .B2(new_n743), .ZN(new_n797));
  INV_X1    g0597(.A(new_n742), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n660), .B2(new_n798), .ZN(new_n799));
  AND2_X1   g0599(.A1(new_n731), .A2(new_n799), .ZN(new_n800));
  INV_X1    g0600(.A(new_n800), .ZN(G396));
  NOR2_X1   g0601(.A1(new_n438), .A2(new_n656), .ZN(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(new_n803));
  OAI21_X1  g0603(.A(new_n451), .B1(new_n444), .B2(KEYINPUT71), .ZN(new_n804));
  NOR3_X1   g0604(.A1(new_n428), .A2(new_n419), .A3(new_n438), .ZN(new_n805));
  OAI211_X1 g0605(.A(new_n455), .B(new_n803), .C1(new_n804), .C2(new_n805), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n806), .A2(KEYINPUT99), .ZN(new_n807));
  INV_X1    g0607(.A(KEYINPUT99), .ZN(new_n808));
  NAND4_X1  g0608(.A1(new_n452), .A2(new_n808), .A3(new_n455), .A4(new_n803), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n807), .A2(new_n809), .ZN(new_n810));
  INV_X1    g0610(.A(KEYINPUT100), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n811), .B1(new_n452), .B2(new_n803), .ZN(new_n812));
  INV_X1    g0612(.A(new_n804), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n813), .A2(KEYINPUT100), .A3(new_n445), .A4(new_n802), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n812), .A2(new_n814), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n810), .A2(new_n815), .ZN(new_n816));
  XNOR2_X1  g0616(.A(new_n711), .B(new_n816), .ZN(new_n817));
  INV_X1    g0617(.A(new_n817), .ZN(new_n818));
  AOI21_X1  g0618(.A(new_n729), .B1(new_n818), .B2(new_n710), .ZN(new_n819));
  INV_X1    g0619(.A(new_n819), .ZN(new_n820));
  NOR2_X1   g0620(.A1(new_n818), .A2(new_n710), .ZN(new_n821));
  NOR2_X1   g0621(.A1(new_n816), .A2(new_n741), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n743), .A2(new_n740), .ZN(new_n823));
  INV_X1    g0623(.A(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(G283), .ZN(new_n825));
  OAI221_X1 g0625(.A(new_n314), .B1(new_n546), .B2(new_n775), .C1(new_n770), .C2(new_n825), .ZN(new_n826));
  NAND2_X1  g0626(.A1(new_n790), .A2(G87), .ZN(new_n827));
  INV_X1    g0627(.A(new_n792), .ZN(new_n828));
  OAI221_X1 g0628(.A(new_n827), .B1(new_n565), .B2(new_n764), .C1(new_n828), .C2(new_n225), .ZN(new_n829));
  AOI211_X1 g0629(.A(new_n826), .B(new_n829), .C1(G311), .C2(new_n793), .ZN(new_n830));
  INV_X1    g0630(.A(G294), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n758), .B1(new_n831), .B2(new_n772), .ZN(new_n832));
  XNOR2_X1  g0632(.A(new_n832), .B(KEYINPUT98), .ZN(new_n833));
  NAND2_X1  g0633(.A1(new_n769), .A2(G150), .ZN(new_n834));
  INV_X1    g0634(.A(G143), .ZN(new_n835));
  OAI221_X1 g0635(.A(new_n834), .B1(new_n835), .B2(new_n772), .C1(new_n775), .C2(new_n751), .ZN(new_n836));
  AOI21_X1  g0636(.A(new_n836), .B1(G137), .B2(new_n789), .ZN(new_n837));
  OR2_X1    g0637(.A1(new_n837), .A2(KEYINPUT34), .ZN(new_n838));
  AOI22_X1  g0638(.A1(G68), .A2(new_n790), .B1(new_n793), .B2(G132), .ZN(new_n839));
  INV_X1    g0639(.A(new_n384), .ZN(new_n840));
  AOI21_X1  g0640(.A(new_n840), .B1(new_n787), .B2(new_n370), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n839), .B(new_n841), .C1(new_n202), .C2(new_n828), .ZN(new_n842));
  AOI21_X1  g0642(.A(new_n842), .B1(KEYINPUT34), .B2(new_n837), .ZN(new_n843));
  AOI22_X1  g0643(.A1(new_n830), .A2(new_n833), .B1(new_n838), .B2(new_n843), .ZN(new_n844));
  INV_X1    g0644(.A(new_n743), .ZN(new_n845));
  OAI221_X1 g0645(.A(new_n729), .B1(G77), .B2(new_n824), .C1(new_n844), .C2(new_n845), .ZN(new_n846));
  OAI22_X1  g0646(.A1(new_n820), .A2(new_n821), .B1(new_n822), .B2(new_n846), .ZN(G384));
  AOI211_X1 g0647(.A(new_n546), .B(new_n213), .C1(new_n471), .C2(KEYINPUT35), .ZN(new_n848));
  OAI21_X1  g0648(.A(new_n848), .B1(KEYINPUT35), .B2(new_n471), .ZN(new_n849));
  XNOR2_X1  g0649(.A(new_n849), .B(KEYINPUT36), .ZN(new_n850));
  AOI211_X1 g0650(.A(new_n223), .B(new_n215), .C1(new_n370), .C2(G68), .ZN(new_n851));
  NOR2_X1   g0651(.A1(new_n217), .A2(G50), .ZN(new_n852));
  OAI211_X1 g0652(.A(G1), .B(new_n648), .C1(new_n851), .C2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  XOR2_X1   g0654(.A(new_n854), .B(KEYINPUT101), .Z(new_n855));
  INV_X1    g0655(.A(new_n655), .ZN(new_n856));
  INV_X1    g0656(.A(KEYINPUT103), .ZN(new_n857));
  OR3_X1    g0657(.A1(new_n401), .A2(new_n857), .A3(KEYINPUT16), .ZN(new_n858));
  OAI21_X1  g0658(.A(new_n401), .B1(new_n857), .B2(KEYINPUT16), .ZN(new_n859));
  NAND3_X1  g0659(.A1(new_n858), .A2(new_n263), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g0660(.A(new_n856), .B1(new_n860), .B2(new_n383), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n411), .A2(new_n417), .ZN(new_n862));
  OAI21_X1  g0662(.A(new_n861), .B1(new_n639), .B2(new_n862), .ZN(new_n863));
  AOI22_X1  g0663(.A1(new_n860), .A2(new_n383), .B1(new_n410), .B2(new_n856), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n408), .A2(new_n394), .ZN(new_n865));
  INV_X1    g0665(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g0666(.A(KEYINPUT37), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g0667(.A1(new_n414), .A2(new_n416), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n414), .A2(new_n655), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT37), .ZN(new_n870));
  NAND4_X1  g0670(.A1(new_n868), .A2(new_n869), .A3(new_n865), .A4(new_n870), .ZN(new_n871));
  NAND2_X1  g0671(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND3_X1  g0672(.A1(new_n863), .A2(new_n872), .A3(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(KEYINPUT82), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n862), .A2(new_n874), .ZN(new_n875));
  NAND3_X1  g0675(.A1(new_n411), .A2(new_n417), .A3(KEYINPUT82), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n875), .A2(new_n396), .A3(new_n876), .ZN(new_n877));
  INV_X1    g0677(.A(new_n869), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n868), .A2(new_n869), .A3(new_n865), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n879), .A2(KEYINPUT37), .ZN(new_n880));
  AOI22_X1  g0680(.A1(new_n877), .A2(new_n878), .B1(new_n871), .B2(new_n880), .ZN(new_n881));
  OAI21_X1  g0681(.A(new_n873), .B1(new_n881), .B2(KEYINPUT38), .ZN(new_n882));
  INV_X1    g0682(.A(KEYINPUT39), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n882), .A2(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n863), .A2(new_n872), .ZN(new_n885));
  INV_X1    g0685(.A(KEYINPUT38), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n873), .ZN(new_n888));
  OAI21_X1  g0688(.A(new_n884), .B1(new_n883), .B2(new_n888), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n348), .A2(new_n341), .A3(new_n656), .ZN(new_n890));
  XNOR2_X1  g0690(.A(new_n890), .B(KEYINPUT104), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n889), .A2(new_n891), .ZN(new_n892));
  NOR2_X1   g0692(.A1(new_n452), .A2(new_n663), .ZN(new_n893));
  INV_X1    g0693(.A(new_n893), .ZN(new_n894));
  AOI22_X1  g0694(.A1(new_n807), .A2(new_n809), .B1(new_n812), .B2(new_n814), .ZN(new_n895));
  OAI21_X1  g0695(.A(new_n894), .B1(new_n711), .B2(new_n895), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n341), .A2(new_n663), .ZN(new_n897));
  XNOR2_X1  g0697(.A(new_n897), .B(KEYINPUT102), .ZN(new_n898));
  INV_X1    g0698(.A(new_n897), .ZN(new_n899));
  AOI22_X1  g0699(.A1(new_n349), .A2(new_n898), .B1(new_n348), .B2(new_n899), .ZN(new_n900));
  INV_X1    g0700(.A(new_n900), .ZN(new_n901));
  NAND3_X1  g0701(.A1(new_n896), .A2(new_n888), .A3(new_n901), .ZN(new_n902));
  NAND2_X1  g0702(.A1(new_n645), .A2(new_n856), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n892), .A2(new_n902), .A3(new_n903), .ZN(new_n904));
  NAND3_X1  g0704(.A1(new_n457), .A2(new_n713), .A3(new_n718), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n905), .A2(new_n646), .A3(new_n355), .ZN(new_n906));
  XNOR2_X1  g0706(.A(new_n904), .B(new_n906), .ZN(new_n907));
  INV_X1    g0707(.A(KEYINPUT105), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n882), .A2(KEYINPUT40), .ZN(new_n909));
  NAND3_X1  g0709(.A1(new_n703), .A2(KEYINPUT31), .A3(new_n663), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n699), .A2(new_n910), .ZN(new_n911));
  NAND3_X1  g0711(.A1(new_n901), .A2(new_n911), .A3(new_n816), .ZN(new_n912));
  OAI21_X1  g0712(.A(new_n908), .B1(new_n909), .B2(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n910), .ZN(new_n914));
  NAND2_X1  g0714(.A1(new_n610), .A2(new_n611), .ZN(new_n915));
  NOR3_X1   g0715(.A1(new_n595), .A2(new_n915), .A3(new_n601), .ZN(new_n916));
  NOR3_X1   g0716(.A1(new_n659), .A2(new_n916), .A3(new_n620), .ZN(new_n917));
  NAND4_X1  g0717(.A1(new_n624), .A2(new_n917), .A3(new_n544), .A4(new_n656), .ZN(new_n918));
  NAND2_X1  g0718(.A1(new_n918), .A2(KEYINPUT31), .ZN(new_n919));
  AOI21_X1  g0719(.A(new_n914), .B1(new_n919), .B2(new_n696), .ZN(new_n920));
  NOR3_X1   g0720(.A1(new_n920), .A2(new_n895), .A3(new_n900), .ZN(new_n921));
  NAND4_X1  g0721(.A1(new_n921), .A2(new_n882), .A3(KEYINPUT105), .A4(KEYINPUT40), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n913), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n921), .A2(new_n888), .ZN(new_n924));
  INV_X1    g0724(.A(KEYINPUT40), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  AND2_X1   g0726(.A1(new_n923), .A2(new_n926), .ZN(new_n927));
  NOR2_X1   g0727(.A1(new_n458), .A2(new_n920), .ZN(new_n928));
  AOI21_X1  g0728(.A(new_n708), .B1(new_n927), .B2(new_n928), .ZN(new_n929));
  OAI21_X1  g0729(.A(new_n929), .B1(new_n928), .B2(new_n927), .ZN(new_n930));
  NAND2_X1  g0730(.A1(new_n907), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g0731(.A(new_n931), .B1(new_n206), .B2(new_n723), .ZN(new_n932));
  NOR2_X1   g0732(.A1(new_n907), .A2(new_n930), .ZN(new_n933));
  OAI21_X1  g0733(.A(new_n855), .B1(new_n932), .B2(new_n933), .ZN(G367));
  OAI221_X1 g0734(.A(new_n744), .B1(new_n210), .B2(new_n436), .C1(new_n737), .C2(new_n238), .ZN(new_n935));
  AND2_X1   g0735(.A1(new_n729), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g0736(.A1(new_n540), .A2(new_n656), .ZN(new_n937));
  INV_X1    g0737(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n544), .A2(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(new_n939), .B1(new_n630), .B2(new_n938), .ZN(new_n940));
  NAND3_X1  g0740(.A1(new_n792), .A2(KEYINPUT46), .A3(G116), .ZN(new_n941));
  XOR2_X1   g0741(.A(new_n941), .B(KEYINPUT110), .Z(new_n942));
  INV_X1    g0742(.A(new_n776), .ZN(new_n943));
  AOI21_X1  g0743(.A(KEYINPUT46), .B1(new_n943), .B2(G116), .ZN(new_n944));
  AOI21_X1  g0744(.A(new_n384), .B1(G303), .B2(new_n771), .ZN(new_n945));
  OAI221_X1 g0745(.A(new_n945), .B1(new_n825), .B2(new_n775), .C1(new_n770), .C2(new_n831), .ZN(new_n946));
  AOI211_X1 g0746(.A(new_n944), .B(new_n946), .C1(G107), .C2(new_n787), .ZN(new_n947));
  NOR2_X1   g0747(.A1(new_n750), .A2(new_n782), .ZN(new_n948));
  NOR2_X1   g0748(.A1(new_n766), .A2(new_n317), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n948), .B(new_n949), .C1(new_n789), .C2(G311), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n942), .A2(new_n947), .A3(new_n950), .ZN(new_n951));
  AND2_X1   g0751(.A1(new_n757), .A2(G68), .ZN(new_n952));
  OAI22_X1  g0752(.A1(new_n770), .A2(new_n751), .B1(new_n775), .B2(new_n202), .ZN(new_n953));
  INV_X1    g0753(.A(G150), .ZN(new_n954));
  OAI22_X1  g0754(.A1(new_n772), .A2(new_n954), .B1(new_n359), .B2(new_n776), .ZN(new_n955));
  NOR4_X1   g0755(.A1(new_n952), .A2(new_n314), .A3(new_n953), .A4(new_n955), .ZN(new_n956));
  AOI22_X1  g0756(.A1(G77), .A2(new_n790), .B1(new_n793), .B2(G137), .ZN(new_n957));
  OAI211_X1 g0757(.A(new_n956), .B(new_n957), .C1(new_n835), .C2(new_n764), .ZN(new_n958));
  NAND2_X1  g0758(.A1(new_n951), .A2(new_n958), .ZN(new_n959));
  XOR2_X1   g0759(.A(new_n959), .B(KEYINPUT47), .Z(new_n960));
  OAI221_X1 g0760(.A(new_n936), .B1(new_n798), .B2(new_n940), .C1(new_n960), .C2(new_n845), .ZN(new_n961));
  XOR2_X1   g0761(.A(new_n675), .B(KEYINPUT41), .Z(new_n962));
  OAI21_X1  g0762(.A(new_n624), .B1(new_n509), .B2(new_n656), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n627), .A2(new_n663), .ZN(new_n964));
  NAND2_X1  g0764(.A1(new_n963), .A2(new_n964), .ZN(new_n965));
  INV_X1    g0765(.A(new_n965), .ZN(new_n966));
  NAND2_X1  g0766(.A1(new_n672), .A2(new_n966), .ZN(new_n967));
  XOR2_X1   g0767(.A(new_n967), .B(KEYINPUT44), .Z(new_n968));
  NOR2_X1   g0768(.A1(new_n672), .A2(new_n966), .ZN(new_n969));
  XNOR2_X1  g0769(.A(new_n969), .B(KEYINPUT45), .ZN(new_n970));
  NAND2_X1  g0770(.A1(new_n968), .A2(new_n970), .ZN(new_n971));
  INV_X1    g0771(.A(new_n668), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n971), .B(new_n972), .ZN(new_n973));
  XNOR2_X1  g0773(.A(new_n662), .B(KEYINPUT109), .ZN(new_n974));
  OAI21_X1  g0774(.A(new_n667), .B1(new_n573), .B2(new_n663), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n975), .A2(new_n670), .ZN(new_n976));
  NAND2_X1  g0776(.A1(new_n974), .A2(new_n976), .ZN(new_n977));
  NAND2_X1  g0777(.A1(new_n662), .A2(KEYINPUT109), .ZN(new_n978));
  INV_X1    g0778(.A(new_n978), .ZN(new_n979));
  OAI21_X1  g0779(.A(new_n977), .B1(new_n976), .B2(new_n979), .ZN(new_n980));
  INV_X1    g0780(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n973), .A2(new_n721), .A3(new_n981), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n962), .B1(new_n982), .B2(new_n721), .ZN(new_n983));
  NOR2_X1   g0783(.A1(new_n983), .A2(new_n725), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n940), .A2(KEYINPUT106), .ZN(new_n985));
  NOR2_X1   g0785(.A1(new_n940), .A2(KEYINPUT106), .ZN(new_n986));
  NOR3_X1   g0786(.A1(new_n985), .A2(new_n986), .A3(KEYINPUT43), .ZN(new_n987));
  NAND3_X1  g0787(.A1(new_n965), .A2(new_n666), .A3(new_n669), .ZN(new_n988));
  OR3_X1    g0788(.A1(new_n988), .A2(KEYINPUT107), .A3(KEYINPUT42), .ZN(new_n989));
  OAI21_X1  g0789(.A(KEYINPUT107), .B1(new_n988), .B2(KEYINPUT42), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n988), .A2(KEYINPUT42), .ZN(new_n991));
  OAI21_X1  g0791(.A(new_n504), .B1(new_n963), .B2(new_n602), .ZN(new_n992));
  NAND2_X1  g0792(.A1(new_n992), .A2(new_n656), .ZN(new_n993));
  NAND4_X1  g0793(.A1(new_n989), .A2(new_n990), .A3(new_n991), .A4(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n940), .A2(KEYINPUT43), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n987), .B1(new_n994), .B2(new_n995), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n996), .B1(new_n987), .B2(new_n994), .ZN(new_n997));
  XNOR2_X1  g0797(.A(new_n997), .B(KEYINPUT108), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n972), .A2(new_n966), .ZN(new_n999));
  INV_X1    g0799(.A(new_n999), .ZN(new_n1000));
  XNOR2_X1  g0800(.A(new_n998), .B(new_n1000), .ZN(new_n1001));
  OAI21_X1  g0801(.A(new_n961), .B1(new_n984), .B2(new_n1001), .ZN(G387));
  INV_X1    g0802(.A(new_n775), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n1003), .A2(G303), .B1(new_n769), .B2(G311), .ZN(new_n1004));
  OAI21_X1  g0804(.A(new_n1004), .B1(new_n782), .B2(new_n772), .ZN(new_n1005));
  AOI21_X1  g0805(.A(new_n1005), .B1(new_n789), .B2(G322), .ZN(new_n1006));
  OR2_X1    g0806(.A1(new_n1006), .A2(KEYINPUT48), .ZN(new_n1007));
  NAND2_X1  g0807(.A1(new_n1006), .A2(KEYINPUT48), .ZN(new_n1008));
  AOI22_X1  g0808(.A1(G294), .A2(new_n943), .B1(new_n787), .B2(G283), .ZN(new_n1009));
  NAND3_X1  g0809(.A1(new_n1007), .A2(new_n1008), .A3(new_n1009), .ZN(new_n1010));
  INV_X1    g0810(.A(KEYINPUT49), .ZN(new_n1011));
  OR2_X1    g0811(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1013));
  NOR2_X1   g0813(.A1(new_n766), .A2(new_n546), .ZN(new_n1014));
  AOI211_X1 g0814(.A(new_n384), .B(new_n1014), .C1(G326), .C2(new_n793), .ZN(new_n1015));
  NAND3_X1  g0815(.A1(new_n1012), .A2(new_n1013), .A3(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n772), .A2(new_n202), .B1(new_n775), .B2(new_n217), .ZN(new_n1017));
  OAI21_X1  g0817(.A(new_n384), .B1(new_n776), .B2(new_n223), .ZN(new_n1018));
  NOR3_X1   g0818(.A1(new_n949), .A2(new_n1017), .A3(new_n1018), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n436), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1020), .A2(new_n757), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n789), .A2(G159), .ZN(new_n1022));
  AOI22_X1  g0822(.A1(new_n793), .A2(G150), .B1(new_n255), .B2(new_n769), .ZN(new_n1023));
  NAND4_X1  g0823(.A1(new_n1019), .A2(new_n1021), .A3(new_n1022), .A4(new_n1023), .ZN(new_n1024));
  AOI21_X1  g0824(.A(new_n845), .B1(new_n1016), .B2(new_n1024), .ZN(new_n1025));
  OR2_X1    g0825(.A1(new_n235), .A2(new_n494), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n1026), .A2(new_n736), .B1(new_n676), .B2(new_n732), .ZN(new_n1027));
  INV_X1    g0827(.A(KEYINPUT50), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n433), .B2(new_n202), .ZN(new_n1029));
  NOR3_X1   g0829(.A1(new_n432), .A2(KEYINPUT50), .A3(G50), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n494), .B1(new_n217), .B2(new_n223), .ZN(new_n1031));
  NOR4_X1   g0831(.A1(new_n1029), .A2(new_n1030), .A3(new_n676), .A4(new_n1031), .ZN(new_n1032));
  OAI22_X1  g0832(.A1(new_n1027), .A2(new_n1032), .B1(G107), .B2(new_n210), .ZN(new_n1033));
  AOI211_X1 g0833(.A(new_n728), .B(new_n1025), .C1(new_n744), .C2(new_n1033), .ZN(new_n1034));
  XNOR2_X1  g0834(.A(new_n1034), .B(KEYINPUT111), .ZN(new_n1035));
  NAND2_X1  g0835(.A1(new_n667), .A2(new_n742), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1037));
  XOR2_X1   g0837(.A(new_n1037), .B(KEYINPUT112), .Z(new_n1038));
  AOI21_X1  g0838(.A(new_n1038), .B1(new_n725), .B2(new_n981), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n981), .A2(new_n721), .ZN(new_n1040));
  NAND2_X1  g0840(.A1(new_n980), .A2(new_n720), .ZN(new_n1041));
  XOR2_X1   g0841(.A(new_n675), .B(KEYINPUT113), .Z(new_n1042));
  NAND3_X1  g0842(.A1(new_n1040), .A2(new_n1041), .A3(new_n1042), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1039), .A2(new_n1043), .ZN(G393));
  XNOR2_X1  g0844(.A(new_n971), .B(new_n668), .ZN(new_n1045));
  OR2_X1    g0845(.A1(new_n1045), .A2(KEYINPUT114), .ZN(new_n1046));
  AOI21_X1  g0846(.A(new_n724), .B1(new_n1045), .B2(KEYINPUT114), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n966), .A2(new_n742), .ZN(new_n1048));
  OAI22_X1  g0848(.A1(new_n764), .A2(new_n954), .B1(new_n372), .B2(new_n772), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  NAND2_X1  g0850(.A1(new_n757), .A2(G77), .ZN(new_n1051));
  AOI22_X1  g0851(.A1(new_n433), .A2(new_n1003), .B1(new_n943), .B2(G68), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n840), .B1(new_n769), .B2(G50), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n827), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1054), .B1(G143), .B2(new_n793), .ZN(new_n1055));
  NAND3_X1  g0855(.A1(new_n1050), .A2(new_n1051), .A3(new_n1055), .ZN(new_n1056));
  OAI22_X1  g0856(.A1(new_n764), .A2(new_n782), .B1(new_n780), .B2(new_n772), .ZN(new_n1057));
  XNOR2_X1  g0857(.A(new_n1057), .B(KEYINPUT52), .ZN(new_n1058));
  OAI22_X1  g0858(.A1(new_n770), .A2(new_n565), .B1(new_n776), .B2(new_n825), .ZN(new_n1059));
  OAI21_X1  g0859(.A(new_n314), .B1(new_n546), .B2(new_n756), .ZN(new_n1060));
  AOI211_X1 g0860(.A(new_n1059), .B(new_n1060), .C1(G294), .C2(new_n1003), .ZN(new_n1061));
  AOI22_X1  g0861(.A1(G107), .A2(new_n790), .B1(new_n793), .B2(G322), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1058), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  AOI21_X1  g0863(.A(new_n845), .B1(new_n1056), .B2(new_n1063), .ZN(new_n1064));
  OAI21_X1  g0864(.A(new_n744), .B1(new_n317), .B2(new_n210), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n1065), .B1(new_n247), .B2(new_n736), .ZN(new_n1066));
  NOR3_X1   g0866(.A1(new_n1064), .A2(new_n728), .A3(new_n1066), .ZN(new_n1067));
  AOI22_X1  g0867(.A1(new_n1046), .A2(new_n1047), .B1(new_n1048), .B2(new_n1067), .ZN(new_n1068));
  NAND2_X1  g0868(.A1(new_n1045), .A2(new_n1040), .ZN(new_n1069));
  NAND3_X1  g0869(.A1(new_n982), .A2(new_n1042), .A3(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1068), .A2(new_n1070), .ZN(G390));
  INV_X1    g0871(.A(KEYINPUT116), .ZN(new_n1072));
  AOI21_X1  g0872(.A(new_n708), .B1(new_n699), .B2(new_n910), .ZN(new_n1073));
  OAI21_X1  g0873(.A(new_n816), .B1(new_n1073), .B2(KEYINPUT115), .ZN(new_n1074));
  AOI21_X1  g0874(.A(new_n695), .B1(new_n918), .B2(KEYINPUT31), .ZN(new_n1075));
  OAI21_X1  g0875(.A(G330), .B1(new_n1075), .B2(new_n914), .ZN(new_n1076));
  INV_X1    g0876(.A(KEYINPUT115), .ZN(new_n1077));
  NOR2_X1   g0877(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n1072), .B(new_n900), .C1(new_n1074), .C2(new_n1078), .ZN(new_n1079));
  OAI211_X1 g0879(.A(new_n816), .B(new_n901), .C1(new_n707), .C2(new_n709), .ZN(new_n1080));
  OAI21_X1  g0880(.A(new_n656), .B1(new_n714), .B2(new_n717), .ZN(new_n1081));
  OAI21_X1  g0881(.A(new_n894), .B1(new_n1081), .B2(new_n895), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND3_X1  g0883(.A1(new_n1079), .A2(new_n1080), .A3(new_n1083), .ZN(new_n1084));
  NAND2_X1  g0884(.A1(new_n1073), .A2(KEYINPUT115), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1076), .A2(new_n1077), .ZN(new_n1086));
  NAND3_X1  g0886(.A1(new_n1085), .A2(new_n1086), .A3(new_n816), .ZN(new_n1087));
  AOI21_X1  g0887(.A(new_n1072), .B1(new_n1087), .B2(new_n900), .ZN(new_n1088));
  NOR2_X1   g0888(.A1(new_n912), .A2(new_n708), .ZN(new_n1089));
  OAI21_X1  g0889(.A(new_n816), .B1(new_n707), .B2(new_n709), .ZN(new_n1090));
  AOI21_X1  g0890(.A(new_n1089), .B1(new_n1090), .B2(new_n900), .ZN(new_n1091));
  INV_X1    g0891(.A(new_n896), .ZN(new_n1092));
  OAI22_X1  g0892(.A1(new_n1084), .A2(new_n1088), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n457), .A2(new_n1073), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n905), .A2(new_n646), .A3(new_n1094), .A4(new_n355), .ZN(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  NAND2_X1  g0896(.A1(new_n1093), .A2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g0897(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1098));
  OAI21_X1  g0898(.A(new_n891), .B1(new_n1092), .B2(new_n900), .ZN(new_n1099));
  NAND2_X1  g0899(.A1(new_n1099), .A2(new_n889), .ZN(new_n1100));
  OAI211_X1 g0900(.A(new_n891), .B(new_n882), .C1(new_n1083), .C2(new_n900), .ZN(new_n1101));
  NAND3_X1  g0901(.A1(new_n1100), .A2(new_n1080), .A3(new_n1101), .ZN(new_n1102));
  AND2_X1   g0902(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1103));
  INV_X1    g0903(.A(new_n1089), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1102), .B1(new_n1103), .B2(new_n1104), .ZN(new_n1105));
  INV_X1    g0905(.A(KEYINPUT117), .ZN(new_n1106));
  NAND3_X1  g0906(.A1(new_n1093), .A2(new_n1106), .A3(new_n1096), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1098), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n1104), .B1(new_n1100), .B2(new_n1101), .ZN(new_n1109));
  AOI21_X1  g0909(.A(new_n1109), .B1(new_n1080), .B2(new_n1103), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n900), .B1(new_n1074), .B2(new_n1078), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1111), .A2(KEYINPUT116), .ZN(new_n1112));
  NAND4_X1  g0912(.A1(new_n1112), .A2(new_n1080), .A3(new_n1083), .A4(new_n1079), .ZN(new_n1113));
  INV_X1    g0913(.A(KEYINPUT88), .ZN(new_n1114));
  XNOR2_X1  g0914(.A(new_n910), .B(new_n1114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(G330), .B1(new_n1115), .B2(new_n1075), .ZN(new_n1116));
  NAND2_X1  g0916(.A1(new_n1116), .A2(KEYINPUT89), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n706), .A2(new_n681), .A3(G330), .ZN(new_n1118));
  AOI21_X1  g0918(.A(new_n895), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  OAI21_X1  g0919(.A(new_n1104), .B1(new_n1119), .B2(new_n901), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n896), .ZN(new_n1121));
  AOI211_X1 g0921(.A(KEYINPUT117), .B(new_n1095), .C1(new_n1113), .C2(new_n1121), .ZN(new_n1122));
  AOI21_X1  g0922(.A(new_n1106), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1123));
  OAI21_X1  g0923(.A(new_n1110), .B1(new_n1122), .B2(new_n1123), .ZN(new_n1124));
  NAND3_X1  g0924(.A1(new_n1108), .A2(new_n1124), .A3(new_n1042), .ZN(new_n1125));
  INV_X1    g0925(.A(new_n741), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n889), .A2(new_n1126), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n729), .B1(new_n255), .B2(new_n824), .ZN(new_n1128));
  AOI22_X1  g0928(.A1(new_n792), .A2(G87), .B1(G294), .B2(new_n793), .ZN(new_n1129));
  OAI221_X1 g0929(.A(new_n1129), .B1(new_n217), .B2(new_n766), .C1(new_n825), .C2(new_n764), .ZN(new_n1130));
  OAI22_X1  g0930(.A1(new_n770), .A2(new_n225), .B1(new_n546), .B2(new_n772), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1131), .B1(G97), .B2(new_n1003), .ZN(new_n1132));
  NAND3_X1  g0932(.A1(new_n1132), .A2(new_n314), .A3(new_n1051), .ZN(new_n1133));
  AOI22_X1  g0933(.A1(new_n789), .A2(G128), .B1(G125), .B2(new_n793), .ZN(new_n1134));
  NOR2_X1   g0934(.A1(new_n776), .A2(new_n954), .ZN(new_n1135));
  XNOR2_X1  g0935(.A(new_n1135), .B(KEYINPUT53), .ZN(new_n1136));
  OAI211_X1 g0936(.A(new_n1134), .B(new_n1136), .C1(new_n202), .C2(new_n766), .ZN(new_n1137));
  NAND2_X1  g0937(.A1(new_n757), .A2(G159), .ZN(new_n1138));
  NAND2_X1  g0938(.A1(new_n769), .A2(G137), .ZN(new_n1139));
  XNOR2_X1  g0939(.A(KEYINPUT54), .B(G143), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1140), .ZN(new_n1141));
  AOI22_X1  g0941(.A1(new_n1003), .A2(new_n1141), .B1(G132), .B2(new_n771), .ZN(new_n1142));
  NAND4_X1  g0942(.A1(new_n1138), .A2(new_n279), .A3(new_n1139), .A4(new_n1142), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n1130), .A2(new_n1133), .B1(new_n1137), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g0944(.A(new_n1128), .B1(new_n1144), .B2(new_n743), .ZN(new_n1145));
  AOI22_X1  g0945(.A1(new_n1110), .A2(new_n725), .B1(new_n1127), .B2(new_n1145), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1125), .A2(new_n1146), .ZN(G378));
  AOI21_X1  g0947(.A(new_n869), .B1(new_n644), .B2(new_n396), .ZN(new_n1148));
  AND2_X1   g0948(.A1(new_n880), .A2(new_n871), .ZN(new_n1149));
  OAI21_X1  g0949(.A(new_n886), .B1(new_n1148), .B2(new_n1149), .ZN(new_n1150));
  AOI21_X1  g0950(.A(new_n925), .B1(new_n1150), .B2(new_n873), .ZN(new_n1151));
  AOI21_X1  g0951(.A(KEYINPUT105), .B1(new_n1151), .B2(new_n921), .ZN(new_n1152));
  AND4_X1   g0952(.A1(KEYINPUT105), .A2(new_n921), .A3(new_n882), .A4(KEYINPUT40), .ZN(new_n1153));
  OAI211_X1 g0953(.A(G330), .B(new_n926), .C1(new_n1152), .C2(new_n1153), .ZN(new_n1154));
  INV_X1    g0954(.A(KEYINPUT119), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1154), .A2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n305), .A2(new_n355), .ZN(new_n1157));
  NAND2_X1  g0957(.A1(new_n269), .A2(new_n655), .ZN(new_n1158));
  XNOR2_X1  g0958(.A(new_n1157), .B(new_n1158), .ZN(new_n1159));
  XNOR2_X1  g0959(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1160));
  XOR2_X1   g0960(.A(new_n1159), .B(new_n1160), .Z(new_n1161));
  INV_X1    g0961(.A(new_n1161), .ZN(new_n1162));
  NAND4_X1  g0962(.A1(new_n923), .A2(KEYINPUT119), .A3(G330), .A4(new_n926), .ZN(new_n1163));
  NAND3_X1  g0963(.A1(new_n1156), .A2(new_n1162), .A3(new_n1163), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n927), .A2(KEYINPUT119), .A3(G330), .A4(new_n1161), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(new_n1165), .ZN(new_n1166));
  NAND2_X1  g0966(.A1(new_n1166), .A2(new_n904), .ZN(new_n1167));
  INV_X1    g0967(.A(new_n904), .ZN(new_n1168));
  NAND3_X1  g0968(.A1(new_n1164), .A2(new_n1165), .A3(new_n1168), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1167), .A2(new_n725), .A3(new_n1169), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n728), .B1(new_n202), .B2(new_n823), .ZN(new_n1171));
  AOI22_X1  g0971(.A1(new_n1020), .A2(new_n1003), .B1(new_n793), .B2(G283), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1172), .B1(new_n546), .B2(new_n764), .ZN(new_n1173));
  AOI211_X1 g0973(.A(G41), .B(new_n384), .C1(new_n943), .C2(G77), .ZN(new_n1174));
  OAI221_X1 g0974(.A(new_n1174), .B1(new_n317), .B2(new_n770), .C1(new_n225), .C2(new_n772), .ZN(new_n1175));
  NOR2_X1   g0975(.A1(new_n766), .A2(new_n359), .ZN(new_n1176));
  NOR4_X1   g0976(.A1(new_n1173), .A2(new_n1175), .A3(new_n952), .A4(new_n1176), .ZN(new_n1177));
  OR2_X1    g0977(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1178));
  NAND2_X1  g0978(.A1(new_n1177), .A2(KEYINPUT58), .ZN(new_n1179));
  OAI21_X1  g0979(.A(new_n202), .B1(new_n271), .B2(G41), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1178), .A2(new_n1179), .A3(new_n1180), .ZN(new_n1181));
  AOI211_X1 g0981(.A(G33), .B(G41), .C1(new_n793), .C2(G124), .ZN(new_n1182));
  OAI21_X1  g0982(.A(new_n1182), .B1(new_n766), .B2(new_n751), .ZN(new_n1183));
  XNOR2_X1  g0983(.A(new_n1183), .B(KEYINPUT118), .ZN(new_n1184));
  NAND2_X1  g0984(.A1(new_n789), .A2(G125), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n757), .A2(G150), .ZN(new_n1186));
  AOI22_X1  g0986(.A1(new_n943), .A2(new_n1141), .B1(G128), .B2(new_n771), .ZN(new_n1187));
  AOI22_X1  g0987(.A1(new_n1003), .A2(G137), .B1(new_n769), .B2(G132), .ZN(new_n1188));
  NAND4_X1  g0988(.A1(new_n1185), .A2(new_n1186), .A3(new_n1187), .A4(new_n1188), .ZN(new_n1189));
  XOR2_X1   g0989(.A(new_n1189), .B(KEYINPUT59), .Z(new_n1190));
  AOI21_X1  g0990(.A(new_n1181), .B1(new_n1184), .B2(new_n1190), .ZN(new_n1191));
  OAI221_X1 g0991(.A(new_n1171), .B1(new_n845), .B2(new_n1191), .C1(new_n1162), .C2(new_n741), .ZN(new_n1192));
  AND2_X1   g0992(.A1(new_n1170), .A2(new_n1192), .ZN(new_n1193));
  XNOR2_X1  g0993(.A(new_n1095), .B(KEYINPUT120), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n1124), .A2(new_n1194), .ZN(new_n1195));
  NAND4_X1  g0995(.A1(new_n1195), .A2(KEYINPUT57), .A3(new_n1169), .A4(new_n1167), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1196), .A2(new_n1042), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n1169), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1168), .B1(new_n1164), .B2(new_n1165), .ZN(new_n1199));
  NOR2_X1   g0999(.A1(new_n1198), .A2(new_n1199), .ZN(new_n1200));
  AOI21_X1  g1000(.A(KEYINPUT57), .B1(new_n1200), .B2(new_n1195), .ZN(new_n1201));
  OAI21_X1  g1001(.A(new_n1193), .B1(new_n1197), .B2(new_n1201), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT121), .ZN(new_n1203));
  XNOR2_X1  g1003(.A(new_n1202), .B(new_n1203), .ZN(G375));
  NAND2_X1  g1004(.A1(new_n1093), .A2(new_n725), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n900), .A2(new_n740), .ZN(new_n1206));
  AOI22_X1  g1006(.A1(new_n792), .A2(G97), .B1(G303), .B2(new_n793), .ZN(new_n1207));
  OAI221_X1 g1007(.A(new_n1207), .B1(new_n223), .B2(new_n766), .C1(new_n831), .C2(new_n764), .ZN(new_n1208));
  OAI22_X1  g1008(.A1(new_n770), .A2(new_n546), .B1(new_n825), .B2(new_n772), .ZN(new_n1209));
  AOI21_X1  g1009(.A(new_n1209), .B1(G107), .B2(new_n1003), .ZN(new_n1210));
  NAND3_X1  g1010(.A1(new_n1210), .A2(new_n314), .A3(new_n1021), .ZN(new_n1211));
  AOI22_X1  g1011(.A1(new_n789), .A2(G132), .B1(G128), .B2(new_n793), .ZN(new_n1212));
  OAI21_X1  g1012(.A(new_n1212), .B1(new_n372), .B2(new_n828), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n757), .A2(G50), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1176), .ZN(new_n1215));
  AOI21_X1  g1015(.A(new_n840), .B1(new_n769), .B2(new_n1141), .ZN(new_n1216));
  AOI22_X1  g1016(.A1(new_n1003), .A2(G150), .B1(new_n771), .B2(G137), .ZN(new_n1217));
  NAND4_X1  g1017(.A1(new_n1214), .A2(new_n1215), .A3(new_n1216), .A4(new_n1217), .ZN(new_n1218));
  OAI22_X1  g1018(.A1(new_n1208), .A2(new_n1211), .B1(new_n1213), .B2(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1219), .A2(new_n743), .ZN(new_n1220));
  AOI21_X1  g1020(.A(new_n728), .B1(new_n217), .B2(new_n823), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1206), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1205), .A2(new_n1222), .ZN(new_n1223));
  INV_X1    g1023(.A(new_n1223), .ZN(new_n1224));
  NAND3_X1  g1024(.A1(new_n1113), .A2(new_n1121), .A3(new_n1095), .ZN(new_n1225));
  NAND3_X1  g1025(.A1(new_n1098), .A2(new_n1107), .A3(new_n1225), .ZN(new_n1226));
  OAI21_X1  g1026(.A(new_n1224), .B1(new_n1226), .B2(new_n962), .ZN(G381));
  NOR2_X1   g1027(.A1(G375), .A2(G378), .ZN(new_n1228));
  INV_X1    g1028(.A(G384), .ZN(new_n1229));
  NAND3_X1  g1029(.A1(new_n1068), .A2(new_n1229), .A3(new_n1070), .ZN(new_n1230));
  NAND3_X1  g1030(.A1(new_n1039), .A2(new_n800), .A3(new_n1043), .ZN(new_n1231));
  NOR4_X1   g1031(.A1(G387), .A2(G381), .A3(new_n1230), .A4(new_n1231), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1228), .A2(new_n1232), .ZN(G407));
  INV_X1    g1033(.A(KEYINPUT122), .ZN(new_n1234));
  INV_X1    g1034(.A(G213), .ZN(new_n1235));
  NOR2_X1   g1035(.A1(new_n1235), .A2(G343), .ZN(new_n1236));
  AOI21_X1  g1036(.A(new_n1234), .B1(new_n1228), .B2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(new_n1202), .B(KEYINPUT121), .ZN(new_n1238));
  INV_X1    g1038(.A(G378), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1238), .A2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(new_n1236), .ZN(new_n1241));
  NOR3_X1   g1041(.A1(new_n1240), .A2(KEYINPUT122), .A3(new_n1241), .ZN(new_n1242));
  OAI211_X1 g1042(.A(G213), .B(G407), .C1(new_n1237), .C2(new_n1242), .ZN(G409));
  NAND2_X1  g1043(.A1(new_n1167), .A2(new_n1169), .ZN(new_n1244));
  INV_X1    g1044(.A(new_n1194), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1098), .A2(new_n1107), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1245), .B1(new_n1246), .B2(new_n1110), .ZN(new_n1247));
  NOR3_X1   g1047(.A1(new_n1244), .A2(new_n1247), .A3(new_n962), .ZN(new_n1248));
  NAND4_X1  g1048(.A1(new_n1170), .A2(new_n1125), .A3(new_n1146), .A4(new_n1192), .ZN(new_n1249));
  OAI21_X1  g1049(.A(new_n1241), .B1(new_n1248), .B2(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(new_n1250), .B1(new_n1202), .B2(G378), .ZN(new_n1251));
  INV_X1    g1051(.A(new_n1225), .ZN(new_n1252));
  OAI21_X1  g1052(.A(new_n1042), .B1(new_n1252), .B2(KEYINPUT60), .ZN(new_n1253));
  AOI21_X1  g1053(.A(new_n1253), .B1(new_n1226), .B2(KEYINPUT60), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1229), .B1(new_n1254), .B2(new_n1223), .ZN(new_n1255));
  INV_X1    g1055(.A(KEYINPUT60), .ZN(new_n1256));
  NOR2_X1   g1056(.A1(new_n1122), .A2(new_n1123), .ZN(new_n1257));
  AOI21_X1  g1057(.A(new_n1256), .B1(new_n1257), .B2(new_n1225), .ZN(new_n1258));
  OAI211_X1 g1058(.A(G384), .B(new_n1224), .C1(new_n1258), .C2(new_n1253), .ZN(new_n1259));
  NAND2_X1  g1059(.A1(new_n1255), .A2(new_n1259), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(KEYINPUT62), .B1(new_n1251), .B2(new_n1261), .ZN(new_n1262));
  INV_X1    g1062(.A(KEYINPUT57), .ZN(new_n1263));
  OAI21_X1  g1063(.A(new_n1263), .B1(new_n1244), .B2(new_n1247), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1264), .A2(new_n1042), .A3(new_n1196), .ZN(new_n1265));
  AOI21_X1  g1065(.A(new_n1239), .B1(new_n1265), .B2(new_n1193), .ZN(new_n1266));
  INV_X1    g1066(.A(KEYINPUT62), .ZN(new_n1267));
  NOR4_X1   g1067(.A1(new_n1266), .A2(new_n1267), .A3(new_n1250), .A4(new_n1260), .ZN(new_n1268));
  NOR2_X1   g1068(.A1(new_n1262), .A2(new_n1268), .ZN(new_n1269));
  INV_X1    g1069(.A(KEYINPUT61), .ZN(new_n1270));
  OAI22_X1  g1070(.A1(new_n1266), .A2(new_n1250), .B1(KEYINPUT124), .B2(new_n1260), .ZN(new_n1271));
  NAND2_X1  g1071(.A1(new_n1236), .A2(G2897), .ZN(new_n1272));
  NAND3_X1  g1072(.A1(new_n1260), .A2(KEYINPUT124), .A3(new_n1272), .ZN(new_n1273));
  INV_X1    g1073(.A(new_n1273), .ZN(new_n1274));
  AOI21_X1  g1074(.A(new_n1272), .B1(new_n1260), .B2(KEYINPUT124), .ZN(new_n1275));
  NOR2_X1   g1075(.A1(new_n1274), .A2(new_n1275), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1270), .B1(new_n1271), .B2(new_n1276), .ZN(new_n1277));
  OAI21_X1  g1077(.A(KEYINPUT126), .B1(new_n1269), .B2(new_n1277), .ZN(new_n1278));
  NOR2_X1   g1078(.A1(new_n1260), .A2(KEYINPUT124), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1202), .A2(G378), .ZN(new_n1280));
  INV_X1    g1080(.A(new_n1250), .ZN(new_n1281));
  AOI21_X1  g1081(.A(new_n1279), .B1(new_n1280), .B2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(new_n1275), .ZN(new_n1283));
  NAND2_X1  g1083(.A1(new_n1283), .A2(new_n1273), .ZN(new_n1284));
  AOI21_X1  g1084(.A(KEYINPUT61), .B1(new_n1282), .B2(new_n1284), .ZN(new_n1285));
  INV_X1    g1085(.A(KEYINPUT126), .ZN(new_n1286));
  OAI211_X1 g1086(.A(new_n1285), .B(new_n1286), .C1(new_n1262), .C2(new_n1268), .ZN(new_n1287));
  INV_X1    g1087(.A(new_n1231), .ZN(new_n1288));
  AOI21_X1  g1088(.A(new_n800), .B1(new_n1039), .B2(new_n1043), .ZN(new_n1289));
  OAI211_X1 g1089(.A(new_n1070), .B(new_n1068), .C1(new_n1288), .C2(new_n1289), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1289), .ZN(new_n1291));
  NAND3_X1  g1091(.A1(new_n1291), .A2(G390), .A3(new_n1231), .ZN(new_n1292));
  NAND2_X1  g1092(.A1(new_n1290), .A2(new_n1292), .ZN(new_n1293));
  NAND2_X1  g1093(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1294));
  INV_X1    g1094(.A(new_n1294), .ZN(new_n1295));
  NOR2_X1   g1095(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1296));
  OAI21_X1  g1096(.A(new_n1293), .B1(new_n1295), .B2(new_n1296), .ZN(new_n1297));
  OR2_X1    g1097(.A1(G387), .A2(KEYINPUT125), .ZN(new_n1298));
  NAND4_X1  g1098(.A1(new_n1298), .A2(new_n1294), .A3(new_n1292), .A4(new_n1290), .ZN(new_n1299));
  AND3_X1   g1099(.A1(new_n1297), .A2(new_n1299), .A3(KEYINPUT127), .ZN(new_n1300));
  AOI21_X1  g1100(.A(KEYINPUT127), .B1(new_n1297), .B2(new_n1299), .ZN(new_n1301));
  NOR2_X1   g1101(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1302));
  NAND3_X1  g1102(.A1(new_n1278), .A2(new_n1287), .A3(new_n1302), .ZN(new_n1303));
  NAND3_X1  g1103(.A1(new_n1280), .A2(new_n1261), .A3(new_n1281), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1304), .ZN(new_n1305));
  OR3_X1    g1105(.A1(new_n1305), .A2(KEYINPUT123), .A3(KEYINPUT63), .ZN(new_n1306));
  NAND2_X1  g1106(.A1(new_n1297), .A2(new_n1299), .ZN(new_n1307));
  AOI21_X1  g1107(.A(new_n1307), .B1(KEYINPUT63), .B2(new_n1305), .ZN(new_n1308));
  OAI21_X1  g1108(.A(KEYINPUT123), .B1(new_n1305), .B2(KEYINPUT63), .ZN(new_n1309));
  NAND4_X1  g1109(.A1(new_n1306), .A2(new_n1285), .A3(new_n1308), .A4(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1303), .A2(new_n1310), .ZN(G405));
  OR2_X1    g1111(.A1(new_n1300), .A2(new_n1301), .ZN(new_n1312));
  NOR3_X1   g1112(.A1(new_n1228), .A2(new_n1261), .A3(new_n1266), .ZN(new_n1313));
  AOI21_X1  g1113(.A(new_n1260), .B1(new_n1240), .B2(new_n1280), .ZN(new_n1314));
  OAI21_X1  g1114(.A(new_n1312), .B1(new_n1313), .B2(new_n1314), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n1261), .B1(new_n1228), .B2(new_n1266), .ZN(new_n1316));
  NAND3_X1  g1116(.A1(new_n1240), .A2(new_n1260), .A3(new_n1280), .ZN(new_n1317));
  NAND3_X1  g1117(.A1(new_n1316), .A2(new_n1302), .A3(new_n1317), .ZN(new_n1318));
  NAND2_X1  g1118(.A1(new_n1315), .A2(new_n1318), .ZN(G402));
endmodule


