

module locked_locked_c2670 ( G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, 
        G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, 
        G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, 
        G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, 
        G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, 
        G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, 
        G103, G104, G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, 
        G117, G118, G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, 
        G131, G132, G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, 
        G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, 
        G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, 
        G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, 
        G215, G239, G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, 
        G250, G251, G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, 
        G266, G267, G268, G269, G270, G271, G272, G273, G274, G275, G276, G452, 
        G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341, G1348, 
        G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991, G1996, 
        G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104, G2105, 
        G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454, G2474, 
        G2678, G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, 
        G220, G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, 
        G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, 
        G188, G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, 
        G148, G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, 
        G331, G397, G329, G231, G308, G225, KEYINPUT63, KEYINPUT62, KEYINPUT61, 
        KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, 
        KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49, 
        KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, 
        KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, 
        KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31, 
        KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, 
        KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19, 
        KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, 
        KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, 
        KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, 
        KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, 
        KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, 
        KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, 
        KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, 
        KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, 
        KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, 
        KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, 
        KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87, 
        KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, 
        KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75, 
        KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, 
        KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64 );
  input G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19, G20, G21, G22,
         G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35, G36, G37, G40,
         G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55, G56, G57, G60,
         G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73, G74, G75, G76,
         G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89, G90, G91, G92,
         G93, G94, G95, G96, G99, G100, G101, G102, G103, G104, G105, G106,
         G107, G108, G111, G112, G113, G114, G115, G116, G117, G118, G119,
         G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
         G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177,
         G178, G179, G180, G181, G182, G183, G184, G185, G186, G189, G190,
         G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201,
         G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
         G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246,
         G247, G248, G249, G250, G251, G252, G253, G254, G255, G256, G257,
         G262, G263, G264, G265, G266, G267, G268, G269, G270, G271, G272,
         G273, G274, G275, G276, G452, G483, G543, G559, G567, G651, G661,
         G860, G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971,
         G1976, G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084,
         G2090, G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438,
         G2443, G2446, G2451, G2454, G2474, G2678, KEYINPUT63, KEYINPUT62,
         KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57,
         KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52,
         KEYINPUT51, KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47,
         KEYINPUT46, KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42,
         KEYINPUT41, KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37,
         KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32,
         KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27,
         KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22,
         KEYINPUT21, KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17,
         KEYINPUT16, KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12,
         KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6,
         KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0,
         KEYINPUT127, KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123,
         KEYINPUT122, KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118,
         KEYINPUT117, KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113,
         KEYINPUT112, KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108,
         KEYINPUT107, KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103,
         KEYINPUT102, KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98,
         KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93,
         KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88,
         KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83,
         KEYINPUT82, KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78,
         KEYINPUT77, KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73,
         KEYINPUT72, KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68,
         KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
         G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234,
         G217, G325, G261, G319, G160, G162, G164, G166, G168, G171, G153,
         G176, G188, G299, G301, G286, G303, G288, G305, G290, G284, G321,
         G297, G280, G148, G282, G323, G156, G401, G227, G229, G311, G150,
         G145, G395, G295, G331, G397, G329, G231, G308, G225;
  wire   G1083, G2066, G452, G284, G297, G282, G295, n517, n518, n519, n520,
         n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531,
         n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
         n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
         n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564,
         n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575,
         n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
         n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597,
         n598, n599, n600, n601, n602, n603, n604, n605, n606, n607, n608,
         n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
         n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630,
         n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641,
         n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
         n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663,
         n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674,
         n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
         n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696,
         n697, n698, n699, n700, n701, n702, n703, n704, n705, n706, n707,
         n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718,
         n719, n720, n721, n722, n723, n724, n725, n726, n727, n728, n729,
         n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
         n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, n751,
         n752, n753, n754, n755, n756, n757, n758, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027;
  assign G231 = 1'b0;
  assign G367 = G1083;
  assign G369 = G1083;
  assign G384 = G2066;
  assign G337 = G2066;
  assign G411 = G2066;
  assign G391 = G452;
  assign G409 = G452;
  assign G335 = G452;
  assign G350 = G452;
  assign G321 = G284;
  assign G280 = G297;
  assign G323 = G282;
  assign G331 = G295;

  NOR2_X2 U551 ( .A1(n533), .A2(n534), .ZN(n878) );
  NOR2_X2 U552 ( .A1(G2105), .A2(n533), .ZN(n583) );
  NOR2_X1 U553 ( .A1(G2104), .A2(G2105), .ZN(n529) );
  INV_X1 U554 ( .A(G2104), .ZN(n533) );
  INV_X1 U555 ( .A(G2105), .ZN(n534) );
  NOR2_X2 U556 ( .A1(n591), .A2(n590), .ZN(G160) );
  NOR2_X1 U557 ( .A1(n668), .A2(n667), .ZN(n669) );
  NOR2_X1 U558 ( .A1(n627), .A2(n762), .ZN(n622) );
  NAND2_X1 U559 ( .A1(n625), .A2(n624), .ZN(n517) );
  NOR2_X1 U560 ( .A1(n955), .A2(n609), .ZN(n611) );
  INV_X1 U561 ( .A(KEYINPUT29), .ZN(n646) );
  AND2_X1 U562 ( .A1(G8), .A2(n677), .ZN(n679) );
  AND2_X1 U563 ( .A1(n596), .A2(n595), .ZN(n648) );
  INV_X1 U564 ( .A(KEYINPUT101), .ZN(n695) );
  INV_X1 U565 ( .A(KEYINPUT90), .ZN(n592) );
  XNOR2_X1 U566 ( .A(n696), .B(n695), .ZN(n703) );
  XNOR2_X1 U567 ( .A(n593), .B(n592), .ZN(n595) );
  NOR2_X1 U568 ( .A1(n571), .A2(G651), .ZN(n794) );
  XOR2_X1 U569 ( .A(KEYINPUT0), .B(G543), .Z(n571) );
  INV_X1 U570 ( .A(G651), .ZN(n521) );
  NOR2_X1 U571 ( .A1(n571), .A2(n521), .ZN(n790) );
  NAND2_X1 U572 ( .A1(n790), .A2(G72), .ZN(n520) );
  NOR2_X1 U573 ( .A1(G651), .A2(G543), .ZN(n518) );
  XNOR2_X1 U574 ( .A(n518), .B(KEYINPUT64), .ZN(n791) );
  NAND2_X1 U575 ( .A1(G85), .A2(n791), .ZN(n519) );
  NAND2_X1 U576 ( .A1(n520), .A2(n519), .ZN(n528) );
  NAND2_X1 U577 ( .A1(n794), .A2(G47), .ZN(n526) );
  XNOR2_X1 U578 ( .A(KEYINPUT68), .B(KEYINPUT1), .ZN(n523) );
  NOR2_X1 U579 ( .A1(G543), .A2(n521), .ZN(n522) );
  XNOR2_X1 U580 ( .A(n523), .B(n522), .ZN(n524) );
  XNOR2_X1 U581 ( .A(KEYINPUT67), .B(n524), .ZN(n795) );
  NAND2_X1 U582 ( .A1(G60), .A2(n795), .ZN(n525) );
  NAND2_X1 U583 ( .A1(n526), .A2(n525), .ZN(n527) );
  OR2_X1 U584 ( .A1(n528), .A2(n527), .ZN(G290) );
  NAND2_X1 U585 ( .A1(G102), .A2(n583), .ZN(n532) );
  XOR2_X1 U586 ( .A(KEYINPUT66), .B(n529), .Z(n530) );
  XNOR2_X1 U587 ( .A(KEYINPUT17), .B(n530), .ZN(n709) );
  NAND2_X1 U588 ( .A1(G138), .A2(n709), .ZN(n531) );
  NAND2_X1 U589 ( .A1(n532), .A2(n531), .ZN(n538) );
  NAND2_X1 U590 ( .A1(G114), .A2(n878), .ZN(n536) );
  NOR2_X1 U591 ( .A1(G2104), .A2(n534), .ZN(n881) );
  NAND2_X1 U592 ( .A1(G126), .A2(n881), .ZN(n535) );
  NAND2_X1 U593 ( .A1(n536), .A2(n535), .ZN(n537) );
  NOR2_X1 U594 ( .A1(n538), .A2(n537), .ZN(G164) );
  NAND2_X1 U595 ( .A1(n794), .A2(G52), .ZN(n540) );
  NAND2_X1 U596 ( .A1(G64), .A2(n795), .ZN(n539) );
  NAND2_X1 U597 ( .A1(n540), .A2(n539), .ZN(n545) );
  NAND2_X1 U598 ( .A1(n790), .A2(G77), .ZN(n542) );
  NAND2_X1 U599 ( .A1(G90), .A2(n791), .ZN(n541) );
  NAND2_X1 U600 ( .A1(n542), .A2(n541), .ZN(n543) );
  XOR2_X1 U601 ( .A(KEYINPUT9), .B(n543), .Z(n544) );
  NOR2_X1 U602 ( .A1(n545), .A2(n544), .ZN(G171) );
  NAND2_X1 U603 ( .A1(n794), .A2(G51), .ZN(n547) );
  NAND2_X1 U604 ( .A1(G63), .A2(n795), .ZN(n546) );
  NAND2_X1 U605 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U606 ( .A(KEYINPUT6), .B(n548), .ZN(n557) );
  NAND2_X1 U607 ( .A1(n790), .A2(G76), .ZN(n549) );
  XNOR2_X1 U608 ( .A(KEYINPUT73), .B(n549), .ZN(n552) );
  NAND2_X1 U609 ( .A1(G89), .A2(n791), .ZN(n550) );
  XOR2_X1 U610 ( .A(n550), .B(KEYINPUT4), .Z(n551) );
  NOR2_X1 U611 ( .A1(n552), .A2(n551), .ZN(n553) );
  XOR2_X1 U612 ( .A(KEYINPUT5), .B(n553), .Z(n555) );
  XNOR2_X1 U613 ( .A(KEYINPUT74), .B(KEYINPUT75), .ZN(n554) );
  XNOR2_X1 U614 ( .A(n555), .B(n554), .ZN(n556) );
  NOR2_X1 U615 ( .A1(n557), .A2(n556), .ZN(n558) );
  XOR2_X1 U616 ( .A(KEYINPUT7), .B(n558), .Z(G168) );
  NAND2_X1 U617 ( .A1(n795), .A2(G62), .ZN(n559) );
  XNOR2_X1 U618 ( .A(n559), .B(KEYINPUT84), .ZN(n566) );
  NAND2_X1 U619 ( .A1(n790), .A2(G75), .ZN(n561) );
  NAND2_X1 U620 ( .A1(G88), .A2(n791), .ZN(n560) );
  NAND2_X1 U621 ( .A1(n561), .A2(n560), .ZN(n564) );
  NAND2_X1 U622 ( .A1(G50), .A2(n794), .ZN(n562) );
  XNOR2_X1 U623 ( .A(KEYINPUT85), .B(n562), .ZN(n563) );
  NOR2_X1 U624 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U625 ( .A1(n566), .A2(n565), .ZN(G303) );
  XOR2_X1 U626 ( .A(G168), .B(KEYINPUT8), .Z(G286) );
  NAND2_X1 U627 ( .A1(G49), .A2(n794), .ZN(n568) );
  NAND2_X1 U628 ( .A1(G74), .A2(G651), .ZN(n567) );
  NAND2_X1 U629 ( .A1(n568), .A2(n567), .ZN(n569) );
  XOR2_X1 U630 ( .A(KEYINPUT81), .B(n569), .Z(n570) );
  NOR2_X1 U631 ( .A1(n795), .A2(n570), .ZN(n573) );
  NAND2_X1 U632 ( .A1(n571), .A2(G87), .ZN(n572) );
  NAND2_X1 U633 ( .A1(n573), .A2(n572), .ZN(G288) );
  NAND2_X1 U634 ( .A1(G86), .A2(n791), .ZN(n575) );
  NAND2_X1 U635 ( .A1(G61), .A2(n795), .ZN(n574) );
  NAND2_X1 U636 ( .A1(n575), .A2(n574), .ZN(n578) );
  NAND2_X1 U637 ( .A1(n790), .A2(G73), .ZN(n576) );
  XOR2_X1 U638 ( .A(KEYINPUT2), .B(n576), .Z(n577) );
  NOR2_X1 U639 ( .A1(n578), .A2(n577), .ZN(n579) );
  XNOR2_X1 U640 ( .A(n579), .B(KEYINPUT82), .ZN(n581) );
  NAND2_X1 U641 ( .A1(G48), .A2(n794), .ZN(n580) );
  NAND2_X1 U642 ( .A1(n581), .A2(n580), .ZN(n582) );
  XOR2_X1 U643 ( .A(KEYINPUT83), .B(n582), .Z(G305) );
  XNOR2_X1 U644 ( .A(G1986), .B(G290), .ZN(n966) );
  NAND2_X1 U645 ( .A1(G101), .A2(n583), .ZN(n584) );
  XOR2_X1 U646 ( .A(KEYINPUT23), .B(n584), .Z(n587) );
  NAND2_X1 U647 ( .A1(G113), .A2(n878), .ZN(n585) );
  XOR2_X1 U648 ( .A(KEYINPUT65), .B(n585), .Z(n586) );
  NAND2_X1 U649 ( .A1(n587), .A2(n586), .ZN(n591) );
  NAND2_X1 U650 ( .A1(G137), .A2(n709), .ZN(n589) );
  NAND2_X1 U651 ( .A1(n881), .A2(G125), .ZN(n588) );
  NAND2_X1 U652 ( .A1(n589), .A2(n588), .ZN(n590) );
  NAND2_X1 U653 ( .A1(G160), .A2(G40), .ZN(n593) );
  INV_X1 U654 ( .A(n595), .ZN(n594) );
  NOR2_X1 U655 ( .A1(G164), .A2(G1384), .ZN(n596) );
  NOR2_X1 U656 ( .A1(n594), .A2(n596), .ZN(n754) );
  NAND2_X1 U657 ( .A1(n966), .A2(n754), .ZN(n741) );
  INV_X1 U658 ( .A(n648), .ZN(n670) );
  NAND2_X1 U659 ( .A1(G8), .A2(n670), .ZN(n706) );
  NOR2_X1 U660 ( .A1(G1966), .A2(n706), .ZN(n668) );
  NAND2_X1 U661 ( .A1(n795), .A2(G56), .ZN(n597) );
  XNOR2_X1 U662 ( .A(n597), .B(KEYINPUT69), .ZN(n598) );
  XNOR2_X1 U663 ( .A(n598), .B(KEYINPUT14), .ZN(n604) );
  NAND2_X1 U664 ( .A1(G81), .A2(n791), .ZN(n599) );
  XNOR2_X1 U665 ( .A(n599), .B(KEYINPUT12), .ZN(n601) );
  NAND2_X1 U666 ( .A1(G68), .A2(n790), .ZN(n600) );
  NAND2_X1 U667 ( .A1(n601), .A2(n600), .ZN(n602) );
  XOR2_X1 U668 ( .A(KEYINPUT13), .B(n602), .Z(n603) );
  NOR2_X1 U669 ( .A1(n604), .A2(n603), .ZN(n606) );
  NAND2_X1 U670 ( .A1(n794), .A2(G43), .ZN(n605) );
  NAND2_X1 U671 ( .A1(n606), .A2(n605), .ZN(n955) );
  INV_X1 U672 ( .A(KEYINPUT26), .ZN(n608) );
  NAND2_X1 U673 ( .A1(G1996), .A2(n648), .ZN(n607) );
  XNOR2_X1 U674 ( .A(n608), .B(n607), .ZN(n609) );
  NAND2_X1 U675 ( .A1(G1341), .A2(n670), .ZN(n610) );
  NAND2_X1 U676 ( .A1(n611), .A2(n610), .ZN(n627) );
  NAND2_X1 U677 ( .A1(G79), .A2(n790), .ZN(n612) );
  XNOR2_X1 U678 ( .A(n612), .B(KEYINPUT72), .ZN(n619) );
  NAND2_X1 U679 ( .A1(n794), .A2(G54), .ZN(n614) );
  NAND2_X1 U680 ( .A1(G66), .A2(n795), .ZN(n613) );
  NAND2_X1 U681 ( .A1(n614), .A2(n613), .ZN(n617) );
  NAND2_X1 U682 ( .A1(G92), .A2(n791), .ZN(n615) );
  XNOR2_X1 U683 ( .A(KEYINPUT71), .B(n615), .ZN(n616) );
  NOR2_X1 U684 ( .A1(n617), .A2(n616), .ZN(n618) );
  NAND2_X1 U685 ( .A1(n619), .A2(n618), .ZN(n620) );
  XNOR2_X1 U686 ( .A(KEYINPUT15), .B(n620), .ZN(n958) );
  INV_X1 U687 ( .A(n958), .ZN(n762) );
  INV_X1 U688 ( .A(KEYINPUT96), .ZN(n621) );
  XNOR2_X1 U689 ( .A(n622), .B(n621), .ZN(n626) );
  NAND2_X1 U690 ( .A1(G1348), .A2(n670), .ZN(n623) );
  XOR2_X1 U691 ( .A(KEYINPUT97), .B(n623), .Z(n625) );
  XOR2_X1 U692 ( .A(KEYINPUT95), .B(n648), .Z(n650) );
  NAND2_X1 U693 ( .A1(G2067), .A2(n650), .ZN(n624) );
  NAND2_X1 U694 ( .A1(n626), .A2(n517), .ZN(n629) );
  NAND2_X1 U695 ( .A1(n762), .A2(n627), .ZN(n628) );
  NAND2_X1 U696 ( .A1(n629), .A2(n628), .ZN(n630) );
  XNOR2_X1 U697 ( .A(n630), .B(KEYINPUT98), .ZN(n641) );
  NAND2_X1 U698 ( .A1(n650), .A2(G2072), .ZN(n631) );
  XNOR2_X1 U699 ( .A(n631), .B(KEYINPUT27), .ZN(n633) );
  INV_X1 U700 ( .A(G1956), .ZN(n840) );
  NOR2_X1 U701 ( .A1(n840), .A2(n650), .ZN(n632) );
  NOR2_X1 U702 ( .A1(n633), .A2(n632), .ZN(n642) );
  NAND2_X1 U703 ( .A1(n794), .A2(G53), .ZN(n635) );
  NAND2_X1 U704 ( .A1(G65), .A2(n795), .ZN(n634) );
  NAND2_X1 U705 ( .A1(n635), .A2(n634), .ZN(n639) );
  NAND2_X1 U706 ( .A1(n790), .A2(G78), .ZN(n637) );
  NAND2_X1 U707 ( .A1(G91), .A2(n791), .ZN(n636) );
  NAND2_X1 U708 ( .A1(n637), .A2(n636), .ZN(n638) );
  NOR2_X1 U709 ( .A1(n639), .A2(n638), .ZN(n960) );
  NAND2_X1 U710 ( .A1(n642), .A2(n960), .ZN(n640) );
  NAND2_X1 U711 ( .A1(n641), .A2(n640), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n642), .A2(n960), .ZN(n643) );
  XOR2_X1 U713 ( .A(n643), .B(KEYINPUT28), .Z(n644) );
  NAND2_X1 U714 ( .A1(n645), .A2(n644), .ZN(n647) );
  XNOR2_X1 U715 ( .A(n647), .B(n646), .ZN(n654) );
  NOR2_X1 U716 ( .A1(n648), .A2(G1961), .ZN(n649) );
  XOR2_X1 U717 ( .A(KEYINPUT94), .B(n649), .Z(n652) );
  XNOR2_X1 U718 ( .A(G2078), .B(KEYINPUT25), .ZN(n981) );
  NAND2_X1 U719 ( .A1(n650), .A2(n981), .ZN(n651) );
  NAND2_X1 U720 ( .A1(n652), .A2(n651), .ZN(n658) );
  NAND2_X1 U721 ( .A1(n658), .A2(G171), .ZN(n653) );
  NAND2_X1 U722 ( .A1(n654), .A2(n653), .ZN(n664) );
  NOR2_X1 U723 ( .A1(G2084), .A2(n670), .ZN(n665) );
  NOR2_X1 U724 ( .A1(n668), .A2(n665), .ZN(n655) );
  NAND2_X1 U725 ( .A1(G8), .A2(n655), .ZN(n656) );
  XNOR2_X1 U726 ( .A(KEYINPUT30), .B(n656), .ZN(n657) );
  NOR2_X1 U727 ( .A1(G168), .A2(n657), .ZN(n660) );
  NOR2_X1 U728 ( .A1(G171), .A2(n658), .ZN(n659) );
  NOR2_X1 U729 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U730 ( .A(n661), .B(KEYINPUT31), .ZN(n662) );
  XNOR2_X1 U731 ( .A(n662), .B(KEYINPUT99), .ZN(n663) );
  NAND2_X1 U732 ( .A1(n664), .A2(n663), .ZN(n674) );
  NAND2_X1 U733 ( .A1(G8), .A2(n665), .ZN(n666) );
  NAND2_X1 U734 ( .A1(n674), .A2(n666), .ZN(n667) );
  XOR2_X1 U735 ( .A(KEYINPUT100), .B(n669), .Z(n681) );
  NOR2_X1 U736 ( .A1(G1971), .A2(n706), .ZN(n672) );
  NOR2_X1 U737 ( .A1(G2090), .A2(n670), .ZN(n671) );
  NOR2_X1 U738 ( .A1(n672), .A2(n671), .ZN(n673) );
  NAND2_X1 U739 ( .A1(n673), .A2(G303), .ZN(n676) );
  NAND2_X1 U740 ( .A1(G286), .A2(n674), .ZN(n675) );
  NAND2_X1 U741 ( .A1(n676), .A2(n675), .ZN(n677) );
  INV_X1 U742 ( .A(KEYINPUT32), .ZN(n678) );
  XNOR2_X1 U743 ( .A(n679), .B(n678), .ZN(n680) );
  NAND2_X1 U744 ( .A1(n681), .A2(n680), .ZN(n699) );
  NOR2_X1 U745 ( .A1(G1976), .A2(G288), .ZN(n687) );
  NOR2_X1 U746 ( .A1(G1971), .A2(G303), .ZN(n682) );
  NOR2_X1 U747 ( .A1(n687), .A2(n682), .ZN(n950) );
  INV_X1 U748 ( .A(KEYINPUT33), .ZN(n683) );
  AND2_X1 U749 ( .A1(n950), .A2(n683), .ZN(n684) );
  NAND2_X1 U750 ( .A1(n699), .A2(n684), .ZN(n694) );
  INV_X1 U751 ( .A(n706), .ZN(n685) );
  NAND2_X1 U752 ( .A1(G1976), .A2(G288), .ZN(n949) );
  AND2_X1 U753 ( .A1(n685), .A2(n949), .ZN(n686) );
  NOR2_X1 U754 ( .A1(KEYINPUT33), .A2(n686), .ZN(n692) );
  XOR2_X1 U755 ( .A(G1981), .B(G305), .Z(n944) );
  INV_X1 U756 ( .A(n944), .ZN(n690) );
  NAND2_X1 U757 ( .A1(n687), .A2(KEYINPUT33), .ZN(n688) );
  NOR2_X1 U758 ( .A1(n706), .A2(n688), .ZN(n689) );
  OR2_X1 U759 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U760 ( .A1(n692), .A2(n691), .ZN(n693) );
  NAND2_X1 U761 ( .A1(n694), .A2(n693), .ZN(n696) );
  NOR2_X1 U762 ( .A1(G2090), .A2(G303), .ZN(n697) );
  XNOR2_X1 U763 ( .A(KEYINPUT102), .B(n697), .ZN(n698) );
  NAND2_X1 U764 ( .A1(n698), .A2(G8), .ZN(n700) );
  NAND2_X1 U765 ( .A1(n700), .A2(n699), .ZN(n701) );
  NAND2_X1 U766 ( .A1(n701), .A2(n706), .ZN(n702) );
  NAND2_X1 U767 ( .A1(n703), .A2(n702), .ZN(n708) );
  NOR2_X1 U768 ( .A1(G1981), .A2(G305), .ZN(n704) );
  XOR2_X1 U769 ( .A(n704), .B(KEYINPUT24), .Z(n705) );
  NOR2_X1 U770 ( .A1(n706), .A2(n705), .ZN(n707) );
  NOR2_X1 U771 ( .A1(n708), .A2(n707), .ZN(n739) );
  NAND2_X1 U772 ( .A1(G117), .A2(n878), .ZN(n711) );
  BUF_X1 U773 ( .A(n709), .Z(n874) );
  NAND2_X1 U774 ( .A1(G141), .A2(n874), .ZN(n710) );
  NAND2_X1 U775 ( .A1(n711), .A2(n710), .ZN(n714) );
  NAND2_X1 U776 ( .A1(n583), .A2(G105), .ZN(n712) );
  XOR2_X1 U777 ( .A(KEYINPUT38), .B(n712), .Z(n713) );
  NOR2_X1 U778 ( .A1(n714), .A2(n713), .ZN(n716) );
  NAND2_X1 U779 ( .A1(n881), .A2(G129), .ZN(n715) );
  NAND2_X1 U780 ( .A1(n716), .A2(n715), .ZN(n891) );
  AND2_X1 U781 ( .A1(n891), .A2(G1996), .ZN(n725) );
  NAND2_X1 U782 ( .A1(G95), .A2(n583), .ZN(n717) );
  XNOR2_X1 U783 ( .A(n717), .B(KEYINPUT92), .ZN(n719) );
  NAND2_X1 U784 ( .A1(n878), .A2(G107), .ZN(n718) );
  NAND2_X1 U785 ( .A1(n719), .A2(n718), .ZN(n723) );
  NAND2_X1 U786 ( .A1(n881), .A2(G119), .ZN(n721) );
  NAND2_X1 U787 ( .A1(G131), .A2(n874), .ZN(n720) );
  NAND2_X1 U788 ( .A1(n721), .A2(n720), .ZN(n722) );
  OR2_X1 U789 ( .A1(n723), .A2(n722), .ZN(n870) );
  XOR2_X1 U790 ( .A(KEYINPUT93), .B(G1991), .Z(n974) );
  AND2_X1 U791 ( .A1(n870), .A2(n974), .ZN(n724) );
  NOR2_X1 U792 ( .A1(n725), .A2(n724), .ZN(n1004) );
  INV_X1 U793 ( .A(n754), .ZN(n726) );
  NOR2_X1 U794 ( .A1(n1004), .A2(n726), .ZN(n746) );
  INV_X1 U795 ( .A(n746), .ZN(n737) );
  XNOR2_X1 U796 ( .A(KEYINPUT37), .B(G2067), .ZN(n752) );
  NAND2_X1 U797 ( .A1(G104), .A2(n583), .ZN(n728) );
  NAND2_X1 U798 ( .A1(G140), .A2(n874), .ZN(n727) );
  NAND2_X1 U799 ( .A1(n728), .A2(n727), .ZN(n729) );
  XNOR2_X1 U800 ( .A(KEYINPUT34), .B(n729), .ZN(n734) );
  NAND2_X1 U801 ( .A1(G116), .A2(n878), .ZN(n731) );
  NAND2_X1 U802 ( .A1(G128), .A2(n881), .ZN(n730) );
  NAND2_X1 U803 ( .A1(n731), .A2(n730), .ZN(n732) );
  XOR2_X1 U804 ( .A(n732), .B(KEYINPUT35), .Z(n733) );
  NOR2_X1 U805 ( .A1(n734), .A2(n733), .ZN(n735) );
  XOR2_X1 U806 ( .A(KEYINPUT36), .B(n735), .Z(n736) );
  XNOR2_X1 U807 ( .A(KEYINPUT91), .B(n736), .ZN(n892) );
  NOR2_X1 U808 ( .A1(n752), .A2(n892), .ZN(n1006) );
  NAND2_X1 U809 ( .A1(n754), .A2(n1006), .ZN(n750) );
  NAND2_X1 U810 ( .A1(n737), .A2(n750), .ZN(n738) );
  NOR2_X1 U811 ( .A1(n739), .A2(n738), .ZN(n740) );
  NAND2_X1 U812 ( .A1(n741), .A2(n740), .ZN(n757) );
  XOR2_X1 U813 ( .A(KEYINPUT39), .B(KEYINPUT105), .Z(n749) );
  NOR2_X1 U814 ( .A1(G1996), .A2(n891), .ZN(n1000) );
  NOR2_X1 U815 ( .A1(n870), .A2(n974), .ZN(n742) );
  XNOR2_X1 U816 ( .A(n742), .B(KEYINPUT104), .ZN(n1010) );
  NOR2_X1 U817 ( .A1(G1986), .A2(G290), .ZN(n743) );
  XOR2_X1 U818 ( .A(n743), .B(KEYINPUT103), .Z(n744) );
  NOR2_X1 U819 ( .A1(n1010), .A2(n744), .ZN(n745) );
  NOR2_X1 U820 ( .A1(n746), .A2(n745), .ZN(n747) );
  NOR2_X1 U821 ( .A1(n1000), .A2(n747), .ZN(n748) );
  XNOR2_X1 U822 ( .A(n749), .B(n748), .ZN(n751) );
  NAND2_X1 U823 ( .A1(n751), .A2(n750), .ZN(n753) );
  NAND2_X1 U824 ( .A1(n752), .A2(n892), .ZN(n1017) );
  NAND2_X1 U825 ( .A1(n753), .A2(n1017), .ZN(n755) );
  NAND2_X1 U826 ( .A1(n755), .A2(n754), .ZN(n756) );
  NAND2_X1 U827 ( .A1(n757), .A2(n756), .ZN(n758) );
  XNOR2_X1 U828 ( .A(n758), .B(KEYINPUT40), .ZN(G329) );
  AND2_X1 U829 ( .A1(G452), .A2(G94), .ZN(G173) );
  INV_X1 U830 ( .A(G57), .ZN(G237) );
  INV_X1 U831 ( .A(G132), .ZN(G219) );
  INV_X1 U832 ( .A(G82), .ZN(G220) );
  NAND2_X1 U833 ( .A1(G7), .A2(G661), .ZN(n760) );
  XOR2_X1 U834 ( .A(n760), .B(KEYINPUT10), .Z(n821) );
  NAND2_X1 U835 ( .A1(n821), .A2(G567), .ZN(n761) );
  XOR2_X1 U836 ( .A(KEYINPUT11), .B(n761), .Z(G234) );
  INV_X1 U837 ( .A(G860), .ZN(n828) );
  OR2_X1 U838 ( .A1(n955), .A2(n828), .ZN(G153) );
  XOR2_X1 U839 ( .A(G171), .B(KEYINPUT70), .Z(G301) );
  NAND2_X1 U840 ( .A1(G868), .A2(G301), .ZN(n764) );
  INV_X1 U841 ( .A(G868), .ZN(n804) );
  NAND2_X1 U842 ( .A1(n762), .A2(n804), .ZN(n763) );
  NAND2_X1 U843 ( .A1(n764), .A2(n763), .ZN(G284) );
  INV_X1 U844 ( .A(n960), .ZN(G299) );
  NOR2_X1 U845 ( .A1(G286), .A2(n804), .ZN(n765) );
  XNOR2_X1 U846 ( .A(n765), .B(KEYINPUT76), .ZN(n767) );
  NOR2_X1 U847 ( .A1(G299), .A2(G868), .ZN(n766) );
  NOR2_X1 U848 ( .A1(n767), .A2(n766), .ZN(n768) );
  XOR2_X1 U849 ( .A(KEYINPUT77), .B(n768), .Z(G297) );
  NAND2_X1 U850 ( .A1(n828), .A2(G559), .ZN(n769) );
  NAND2_X1 U851 ( .A1(n769), .A2(n958), .ZN(n770) );
  XNOR2_X1 U852 ( .A(n770), .B(KEYINPUT16), .ZN(G148) );
  NOR2_X1 U853 ( .A1(G868), .A2(n955), .ZN(n773) );
  NAND2_X1 U854 ( .A1(G868), .A2(n958), .ZN(n771) );
  NOR2_X1 U855 ( .A1(G559), .A2(n771), .ZN(n772) );
  NOR2_X1 U856 ( .A1(n773), .A2(n772), .ZN(n774) );
  XNOR2_X1 U857 ( .A(KEYINPUT78), .B(n774), .ZN(G282) );
  NAND2_X1 U858 ( .A1(G111), .A2(n878), .ZN(n776) );
  NAND2_X1 U859 ( .A1(G135), .A2(n874), .ZN(n775) );
  NAND2_X1 U860 ( .A1(n776), .A2(n775), .ZN(n779) );
  NAND2_X1 U861 ( .A1(n881), .A2(G123), .ZN(n777) );
  XOR2_X1 U862 ( .A(KEYINPUT18), .B(n777), .Z(n778) );
  NOR2_X1 U863 ( .A1(n779), .A2(n778), .ZN(n781) );
  NAND2_X1 U864 ( .A1(n583), .A2(G99), .ZN(n780) );
  NAND2_X1 U865 ( .A1(n781), .A2(n780), .ZN(n1003) );
  XNOR2_X1 U866 ( .A(n1003), .B(G2096), .ZN(n782) );
  XNOR2_X1 U867 ( .A(n782), .B(KEYINPUT79), .ZN(n783) );
  INV_X1 U868 ( .A(G2100), .ZN(n831) );
  NAND2_X1 U869 ( .A1(n783), .A2(n831), .ZN(G156) );
  NAND2_X1 U870 ( .A1(G559), .A2(n958), .ZN(n784) );
  XOR2_X1 U871 ( .A(n955), .B(n784), .Z(n827) );
  XOR2_X1 U872 ( .A(G290), .B(G305), .Z(n785) );
  XNOR2_X1 U873 ( .A(G288), .B(n785), .ZN(n789) );
  XOR2_X1 U874 ( .A(KEYINPUT87), .B(KEYINPUT86), .Z(n787) );
  XOR2_X1 U875 ( .A(G299), .B(KEYINPUT19), .Z(n786) );
  XNOR2_X1 U876 ( .A(n787), .B(n786), .ZN(n788) );
  XOR2_X1 U877 ( .A(n789), .B(n788), .Z(n802) );
  NAND2_X1 U878 ( .A1(n790), .A2(G80), .ZN(n793) );
  NAND2_X1 U879 ( .A1(G93), .A2(n791), .ZN(n792) );
  NAND2_X1 U880 ( .A1(n793), .A2(n792), .ZN(n799) );
  NAND2_X1 U881 ( .A1(n794), .A2(G55), .ZN(n797) );
  NAND2_X1 U882 ( .A1(G67), .A2(n795), .ZN(n796) );
  NAND2_X1 U883 ( .A1(n797), .A2(n796), .ZN(n798) );
  NOR2_X1 U884 ( .A1(n799), .A2(n798), .ZN(n800) );
  XOR2_X1 U885 ( .A(KEYINPUT80), .B(n800), .Z(n829) );
  XOR2_X1 U886 ( .A(G303), .B(n829), .Z(n801) );
  XNOR2_X1 U887 ( .A(n802), .B(n801), .ZN(n898) );
  XNOR2_X1 U888 ( .A(n827), .B(n898), .ZN(n803) );
  NAND2_X1 U889 ( .A1(n803), .A2(G868), .ZN(n806) );
  NAND2_X1 U890 ( .A1(n829), .A2(n804), .ZN(n805) );
  NAND2_X1 U891 ( .A1(n806), .A2(n805), .ZN(G295) );
  NAND2_X1 U892 ( .A1(G2078), .A2(G2084), .ZN(n808) );
  XOR2_X1 U893 ( .A(KEYINPUT88), .B(KEYINPUT20), .Z(n807) );
  XNOR2_X1 U894 ( .A(n808), .B(n807), .ZN(n809) );
  NAND2_X1 U895 ( .A1(G2090), .A2(n809), .ZN(n810) );
  XNOR2_X1 U896 ( .A(KEYINPUT21), .B(n810), .ZN(n811) );
  NAND2_X1 U897 ( .A1(n811), .A2(G2072), .ZN(G158) );
  XNOR2_X1 U898 ( .A(G44), .B(KEYINPUT3), .ZN(G218) );
  NOR2_X1 U899 ( .A1(G220), .A2(G219), .ZN(n812) );
  XOR2_X1 U900 ( .A(KEYINPUT22), .B(n812), .Z(n813) );
  NOR2_X1 U901 ( .A1(G218), .A2(n813), .ZN(n814) );
  NAND2_X1 U902 ( .A1(G96), .A2(n814), .ZN(n825) );
  NAND2_X1 U903 ( .A1(n825), .A2(G2106), .ZN(n818) );
  NAND2_X1 U904 ( .A1(G69), .A2(G120), .ZN(n815) );
  NOR2_X1 U905 ( .A1(G237), .A2(n815), .ZN(n816) );
  NAND2_X1 U906 ( .A1(G108), .A2(n816), .ZN(n826) );
  NAND2_X1 U907 ( .A1(n826), .A2(G567), .ZN(n817) );
  NAND2_X1 U908 ( .A1(n818), .A2(n817), .ZN(n853) );
  NAND2_X1 U909 ( .A1(G483), .A2(G661), .ZN(n819) );
  NOR2_X1 U910 ( .A1(n853), .A2(n819), .ZN(n824) );
  NAND2_X1 U911 ( .A1(n824), .A2(G36), .ZN(n820) );
  XOR2_X1 U912 ( .A(KEYINPUT89), .B(n820), .Z(G176) );
  NAND2_X1 U913 ( .A1(G2106), .A2(n821), .ZN(G217) );
  INV_X1 U914 ( .A(n821), .ZN(G223) );
  AND2_X1 U915 ( .A1(G15), .A2(G2), .ZN(n822) );
  NAND2_X1 U916 ( .A1(G661), .A2(n822), .ZN(G259) );
  NAND2_X1 U917 ( .A1(G3), .A2(G1), .ZN(n823) );
  NAND2_X1 U918 ( .A1(n824), .A2(n823), .ZN(G188) );
  NOR2_X1 U919 ( .A1(n826), .A2(n825), .ZN(G325) );
  XOR2_X1 U920 ( .A(KEYINPUT106), .B(G325), .Z(G261) );
  NAND2_X1 U922 ( .A1(n828), .A2(n827), .ZN(n830) );
  XNOR2_X1 U923 ( .A(n830), .B(n829), .ZN(G145) );
  INV_X1 U924 ( .A(G120), .ZN(G236) );
  INV_X1 U925 ( .A(G96), .ZN(G221) );
  INV_X1 U926 ( .A(G69), .ZN(G235) );
  XNOR2_X1 U927 ( .A(n831), .B(G2096), .ZN(n833) );
  XNOR2_X1 U928 ( .A(KEYINPUT42), .B(G2678), .ZN(n832) );
  XNOR2_X1 U929 ( .A(n833), .B(n832), .ZN(n837) );
  XOR2_X1 U930 ( .A(KEYINPUT43), .B(G2090), .Z(n835) );
  XNOR2_X1 U931 ( .A(G2067), .B(G2072), .ZN(n834) );
  XNOR2_X1 U932 ( .A(n835), .B(n834), .ZN(n836) );
  XOR2_X1 U933 ( .A(n837), .B(n836), .Z(n839) );
  XNOR2_X1 U934 ( .A(G2078), .B(G2084), .ZN(n838) );
  XNOR2_X1 U935 ( .A(n839), .B(n838), .ZN(G227) );
  XNOR2_X1 U936 ( .A(G1981), .B(n840), .ZN(n842) );
  XNOR2_X1 U937 ( .A(G1996), .B(G1991), .ZN(n841) );
  XNOR2_X1 U938 ( .A(n842), .B(n841), .ZN(n852) );
  XOR2_X1 U939 ( .A(KEYINPUT107), .B(KEYINPUT41), .Z(n844) );
  XNOR2_X1 U940 ( .A(G1986), .B(KEYINPUT108), .ZN(n843) );
  XNOR2_X1 U941 ( .A(n844), .B(n843), .ZN(n848) );
  INV_X1 U942 ( .A(G1971), .ZN(n948) );
  XNOR2_X1 U943 ( .A(G1976), .B(n948), .ZN(n846) );
  XNOR2_X1 U944 ( .A(G1966), .B(G1961), .ZN(n845) );
  XNOR2_X1 U945 ( .A(n846), .B(n845), .ZN(n847) );
  XOR2_X1 U946 ( .A(n848), .B(n847), .Z(n850) );
  XNOR2_X1 U947 ( .A(KEYINPUT109), .B(G2474), .ZN(n849) );
  XNOR2_X1 U948 ( .A(n850), .B(n849), .ZN(n851) );
  XOR2_X1 U949 ( .A(n852), .B(n851), .Z(G229) );
  INV_X1 U950 ( .A(n853), .ZN(G319) );
  NAND2_X1 U951 ( .A1(n881), .A2(G124), .ZN(n854) );
  XNOR2_X1 U952 ( .A(n854), .B(KEYINPUT44), .ZN(n856) );
  NAND2_X1 U953 ( .A1(G136), .A2(n874), .ZN(n855) );
  NAND2_X1 U954 ( .A1(n856), .A2(n855), .ZN(n857) );
  XNOR2_X1 U955 ( .A(KEYINPUT110), .B(n857), .ZN(n861) );
  NAND2_X1 U956 ( .A1(G112), .A2(n878), .ZN(n859) );
  NAND2_X1 U957 ( .A1(G100), .A2(n583), .ZN(n858) );
  NAND2_X1 U958 ( .A1(n859), .A2(n858), .ZN(n860) );
  NOR2_X1 U959 ( .A1(n861), .A2(n860), .ZN(n862) );
  XOR2_X1 U960 ( .A(KEYINPUT111), .B(n862), .Z(G162) );
  NAND2_X1 U961 ( .A1(G103), .A2(n583), .ZN(n864) );
  NAND2_X1 U962 ( .A1(G139), .A2(n874), .ZN(n863) );
  NAND2_X1 U963 ( .A1(n864), .A2(n863), .ZN(n869) );
  NAND2_X1 U964 ( .A1(G115), .A2(n878), .ZN(n866) );
  NAND2_X1 U965 ( .A1(G127), .A2(n881), .ZN(n865) );
  NAND2_X1 U966 ( .A1(n866), .A2(n865), .ZN(n867) );
  XOR2_X1 U967 ( .A(KEYINPUT47), .B(n867), .Z(n868) );
  NOR2_X1 U968 ( .A1(n869), .A2(n868), .ZN(n1013) );
  XNOR2_X1 U969 ( .A(n1013), .B(n870), .ZN(n871) );
  XNOR2_X1 U970 ( .A(n871), .B(n1003), .ZN(n890) );
  XOR2_X1 U971 ( .A(KEYINPUT48), .B(KEYINPUT114), .Z(n873) );
  XNOR2_X1 U972 ( .A(KEYINPUT46), .B(KEYINPUT113), .ZN(n872) );
  XNOR2_X1 U973 ( .A(n873), .B(n872), .ZN(n886) );
  NAND2_X1 U974 ( .A1(G106), .A2(n583), .ZN(n876) );
  NAND2_X1 U975 ( .A1(G142), .A2(n874), .ZN(n875) );
  NAND2_X1 U976 ( .A1(n876), .A2(n875), .ZN(n877) );
  XNOR2_X1 U977 ( .A(n877), .B(KEYINPUT45), .ZN(n880) );
  NAND2_X1 U978 ( .A1(G118), .A2(n878), .ZN(n879) );
  NAND2_X1 U979 ( .A1(n880), .A2(n879), .ZN(n884) );
  NAND2_X1 U980 ( .A1(n881), .A2(G130), .ZN(n882) );
  XOR2_X1 U981 ( .A(KEYINPUT112), .B(n882), .Z(n883) );
  NOR2_X1 U982 ( .A1(n884), .A2(n883), .ZN(n885) );
  XOR2_X1 U983 ( .A(n886), .B(n885), .Z(n888) );
  XNOR2_X1 U984 ( .A(G160), .B(G164), .ZN(n887) );
  XNOR2_X1 U985 ( .A(n888), .B(n887), .ZN(n889) );
  XNOR2_X1 U986 ( .A(n890), .B(n889), .ZN(n894) );
  XOR2_X1 U987 ( .A(n892), .B(n891), .Z(n893) );
  XNOR2_X1 U988 ( .A(n894), .B(n893), .ZN(n895) );
  XOR2_X1 U989 ( .A(G162), .B(n895), .Z(n896) );
  NOR2_X1 U990 ( .A1(G37), .A2(n896), .ZN(n897) );
  XOR2_X1 U991 ( .A(KEYINPUT115), .B(n897), .Z(G395) );
  XOR2_X1 U992 ( .A(G286), .B(n898), .Z(n899) );
  XNOR2_X1 U993 ( .A(n955), .B(n899), .ZN(n901) );
  XOR2_X1 U994 ( .A(n958), .B(G171), .Z(n900) );
  XNOR2_X1 U995 ( .A(n901), .B(n900), .ZN(n902) );
  NOR2_X1 U996 ( .A1(G37), .A2(n902), .ZN(G397) );
  XNOR2_X1 U997 ( .A(KEYINPUT116), .B(KEYINPUT49), .ZN(n904) );
  NOR2_X1 U998 ( .A1(G227), .A2(G229), .ZN(n903) );
  XNOR2_X1 U999 ( .A(n904), .B(n903), .ZN(n915) );
  XOR2_X1 U1000 ( .A(G2451), .B(G2430), .Z(n906) );
  XNOR2_X1 U1001 ( .A(G2438), .B(G2443), .ZN(n905) );
  XNOR2_X1 U1002 ( .A(n906), .B(n905), .ZN(n912) );
  XOR2_X1 U1003 ( .A(G2435), .B(G2454), .Z(n908) );
  XNOR2_X1 U1004 ( .A(G1348), .B(G1341), .ZN(n907) );
  XNOR2_X1 U1005 ( .A(n908), .B(n907), .ZN(n910) );
  XOR2_X1 U1006 ( .A(G2446), .B(G2427), .Z(n909) );
  XNOR2_X1 U1007 ( .A(n910), .B(n909), .ZN(n911) );
  XOR2_X1 U1008 ( .A(n912), .B(n911), .Z(n913) );
  NAND2_X1 U1009 ( .A1(G14), .A2(n913), .ZN(n918) );
  NAND2_X1 U1010 ( .A1(G319), .A2(n918), .ZN(n914) );
  NOR2_X1 U1011 ( .A1(n915), .A2(n914), .ZN(n917) );
  NOR2_X1 U1012 ( .A1(G395), .A2(G397), .ZN(n916) );
  NAND2_X1 U1013 ( .A1(n917), .A2(n916), .ZN(G225) );
  INV_X1 U1014 ( .A(G225), .ZN(G308) );
  INV_X1 U1015 ( .A(G303), .ZN(G166) );
  INV_X1 U1016 ( .A(G108), .ZN(G238) );
  INV_X1 U1017 ( .A(n918), .ZN(G401) );
  XOR2_X1 U1018 ( .A(G1956), .B(G20), .Z(n926) );
  XOR2_X1 U1019 ( .A(G1981), .B(G6), .Z(n921) );
  XOR2_X1 U1020 ( .A(G19), .B(KEYINPUT122), .Z(n919) );
  XNOR2_X1 U1021 ( .A(G1341), .B(n919), .ZN(n920) );
  NAND2_X1 U1022 ( .A1(n921), .A2(n920), .ZN(n924) );
  XOR2_X1 U1023 ( .A(KEYINPUT59), .B(G1348), .Z(n922) );
  XNOR2_X1 U1024 ( .A(G4), .B(n922), .ZN(n923) );
  NOR2_X1 U1025 ( .A1(n924), .A2(n923), .ZN(n925) );
  NAND2_X1 U1026 ( .A1(n926), .A2(n925), .ZN(n927) );
  XNOR2_X1 U1027 ( .A(n927), .B(KEYINPUT60), .ZN(n940) );
  XOR2_X1 U1028 ( .A(G1976), .B(KEYINPUT123), .Z(n928) );
  XNOR2_X1 U1029 ( .A(G23), .B(n928), .ZN(n930) );
  XOR2_X1 U1030 ( .A(G22), .B(n948), .Z(n929) );
  NOR2_X1 U1031 ( .A1(n930), .A2(n929), .ZN(n931) );
  XOR2_X1 U1032 ( .A(KEYINPUT124), .B(n931), .Z(n933) );
  XNOR2_X1 U1033 ( .A(G1986), .B(G24), .ZN(n932) );
  NOR2_X1 U1034 ( .A1(n933), .A2(n932), .ZN(n934) );
  XNOR2_X1 U1035 ( .A(KEYINPUT58), .B(n934), .ZN(n938) );
  XNOR2_X1 U1036 ( .A(G1966), .B(G21), .ZN(n936) );
  XNOR2_X1 U1037 ( .A(G1961), .B(G5), .ZN(n935) );
  NOR2_X1 U1038 ( .A1(n936), .A2(n935), .ZN(n937) );
  NAND2_X1 U1039 ( .A1(n938), .A2(n937), .ZN(n939) );
  NOR2_X1 U1040 ( .A1(n940), .A2(n939), .ZN(n941) );
  XOR2_X1 U1041 ( .A(KEYINPUT61), .B(n941), .Z(n942) );
  NOR2_X1 U1042 ( .A1(G16), .A2(n942), .ZN(n943) );
  XNOR2_X1 U1043 ( .A(n943), .B(KEYINPUT125), .ZN(n972) );
  XNOR2_X1 U1044 ( .A(G16), .B(KEYINPUT56), .ZN(n970) );
  XNOR2_X1 U1045 ( .A(G1966), .B(G168), .ZN(n945) );
  NAND2_X1 U1046 ( .A1(n945), .A2(n944), .ZN(n946) );
  XNOR2_X1 U1047 ( .A(n946), .B(KEYINPUT57), .ZN(n947) );
  XNOR2_X1 U1048 ( .A(KEYINPUT120), .B(n947), .ZN(n954) );
  NOR2_X1 U1049 ( .A1(G166), .A2(n948), .ZN(n952) );
  NAND2_X1 U1050 ( .A1(n950), .A2(n949), .ZN(n951) );
  NOR2_X1 U1051 ( .A1(n952), .A2(n951), .ZN(n953) );
  NAND2_X1 U1052 ( .A1(n954), .A2(n953), .ZN(n957) );
  XNOR2_X1 U1053 ( .A(G1341), .B(n955), .ZN(n956) );
  NOR2_X1 U1054 ( .A1(n957), .A2(n956), .ZN(n968) );
  XOR2_X1 U1055 ( .A(n958), .B(G1348), .Z(n959) );
  XNOR2_X1 U1056 ( .A(n959), .B(KEYINPUT121), .ZN(n964) );
  XOR2_X1 U1057 ( .A(G171), .B(G1961), .Z(n962) );
  XOR2_X1 U1058 ( .A(n960), .B(G1956), .Z(n961) );
  NOR2_X1 U1059 ( .A1(n962), .A2(n961), .ZN(n963) );
  NAND2_X1 U1060 ( .A1(n964), .A2(n963), .ZN(n965) );
  NOR2_X1 U1061 ( .A1(n966), .A2(n965), .ZN(n967) );
  NAND2_X1 U1062 ( .A1(n968), .A2(n967), .ZN(n969) );
  NAND2_X1 U1063 ( .A1(n970), .A2(n969), .ZN(n971) );
  NAND2_X1 U1064 ( .A1(n972), .A2(n971), .ZN(n973) );
  XNOR2_X1 U1065 ( .A(n973), .B(KEYINPUT126), .ZN(n996) );
  INV_X1 U1066 ( .A(KEYINPUT55), .ZN(n1022) );
  XNOR2_X1 U1067 ( .A(G2090), .B(G35), .ZN(n989) );
  XOR2_X1 U1068 ( .A(G25), .B(n974), .Z(n980) );
  XOR2_X1 U1069 ( .A(G2067), .B(G26), .Z(n975) );
  NAND2_X1 U1070 ( .A1(n975), .A2(G28), .ZN(n978) );
  XNOR2_X1 U1071 ( .A(KEYINPUT118), .B(G2072), .ZN(n976) );
  XNOR2_X1 U1072 ( .A(G33), .B(n976), .ZN(n977) );
  NOR2_X1 U1073 ( .A1(n978), .A2(n977), .ZN(n979) );
  NAND2_X1 U1074 ( .A1(n980), .A2(n979), .ZN(n986) );
  XOR2_X1 U1075 ( .A(n981), .B(G27), .Z(n983) );
  XNOR2_X1 U1076 ( .A(G1996), .B(G32), .ZN(n982) );
  NOR2_X1 U1077 ( .A1(n983), .A2(n982), .ZN(n984) );
  XNOR2_X1 U1078 ( .A(n984), .B(KEYINPUT119), .ZN(n985) );
  NOR2_X1 U1079 ( .A1(n986), .A2(n985), .ZN(n987) );
  XNOR2_X1 U1080 ( .A(KEYINPUT53), .B(n987), .ZN(n988) );
  NOR2_X1 U1081 ( .A1(n989), .A2(n988), .ZN(n992) );
  XOR2_X1 U1082 ( .A(G2084), .B(G34), .Z(n990) );
  XNOR2_X1 U1083 ( .A(KEYINPUT54), .B(n990), .ZN(n991) );
  NAND2_X1 U1084 ( .A1(n992), .A2(n991), .ZN(n993) );
  XOR2_X1 U1085 ( .A(n1022), .B(n993), .Z(n994) );
  NOR2_X1 U1086 ( .A1(n994), .A2(G29), .ZN(n995) );
  NOR2_X1 U1087 ( .A1(n996), .A2(n995), .ZN(n997) );
  NAND2_X1 U1088 ( .A1(G11), .A2(n997), .ZN(n998) );
  XNOR2_X1 U1089 ( .A(n998), .B(KEYINPUT127), .ZN(n1026) );
  XOR2_X1 U1090 ( .A(G2090), .B(G162), .Z(n999) );
  NOR2_X1 U1091 ( .A1(n1000), .A2(n999), .ZN(n1001) );
  XNOR2_X1 U1092 ( .A(KEYINPUT51), .B(n1001), .ZN(n1002) );
  XNOR2_X1 U1093 ( .A(n1002), .B(KEYINPUT117), .ZN(n1012) );
  XNOR2_X1 U1094 ( .A(G160), .B(G2084), .ZN(n1008) );
  NAND2_X1 U1095 ( .A1(n1004), .A2(n1003), .ZN(n1005) );
  NOR2_X1 U1096 ( .A1(n1006), .A2(n1005), .ZN(n1007) );
  NAND2_X1 U1097 ( .A1(n1008), .A2(n1007), .ZN(n1009) );
  NOR2_X1 U1098 ( .A1(n1010), .A2(n1009), .ZN(n1011) );
  NAND2_X1 U1099 ( .A1(n1012), .A2(n1011), .ZN(n1020) );
  XOR2_X1 U1100 ( .A(G2072), .B(n1013), .Z(n1015) );
  XOR2_X1 U1101 ( .A(G164), .B(G2078), .Z(n1014) );
  NOR2_X1 U1102 ( .A1(n1015), .A2(n1014), .ZN(n1016) );
  XNOR2_X1 U1103 ( .A(n1016), .B(KEYINPUT50), .ZN(n1018) );
  NAND2_X1 U1104 ( .A1(n1018), .A2(n1017), .ZN(n1019) );
  NOR2_X1 U1105 ( .A1(n1020), .A2(n1019), .ZN(n1021) );
  XNOR2_X1 U1106 ( .A(KEYINPUT52), .B(n1021), .ZN(n1023) );
  NAND2_X1 U1107 ( .A1(n1023), .A2(n1022), .ZN(n1024) );
  NAND2_X1 U1108 ( .A1(n1024), .A2(G29), .ZN(n1025) );
  NAND2_X1 U1109 ( .A1(n1026), .A2(n1025), .ZN(n1027) );
  XNOR2_X1 U1110 ( .A(KEYINPUT62), .B(n1027), .ZN(G150) );
  INV_X1 U1111 ( .A(G150), .ZN(G311) );
endmodule

