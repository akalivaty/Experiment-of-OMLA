//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 1 0 1 0 1 1 1 0 1 1 1 1 0 1 0 0 0 0 0 0 0 1 1 0 0 0 1 1 1 1 1 0 0 1 1 1 1 0 1 1 1 0 0 0 0 1 1 0 1 1 1 0 1 0 1 0 0 1 0 1 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:04 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n721, new_n722, new_n723, new_n724,
    new_n725, new_n726, new_n727, new_n728, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n735, new_n736, new_n737, new_n738,
    new_n739, new_n740, new_n741, new_n742, new_n743, new_n744, new_n745,
    new_n746, new_n747, new_n748, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n798, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n808, new_n809, new_n810,
    new_n811, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n822, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n906, new_n907, new_n908, new_n909, new_n910,
    new_n911, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n943, new_n944, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1007,
    new_n1008, new_n1009, new_n1010, new_n1011, new_n1012, new_n1013,
    new_n1014, new_n1015, new_n1016, new_n1017, new_n1018, new_n1019,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1115, new_n1116, new_n1117,
    new_n1118, new_n1119, new_n1120, new_n1121, new_n1122, new_n1123,
    new_n1124, new_n1125, new_n1126, new_n1127, new_n1128, new_n1129,
    new_n1130, new_n1131, new_n1132, new_n1133, new_n1134, new_n1135,
    new_n1136, new_n1137, new_n1138, new_n1139, new_n1140, new_n1141,
    new_n1142, new_n1143, new_n1144, new_n1145, new_n1146, new_n1147,
    new_n1148, new_n1149, new_n1150, new_n1151, new_n1152, new_n1153,
    new_n1154, new_n1155, new_n1157, new_n1158, new_n1159, new_n1160,
    new_n1161, new_n1162, new_n1163, new_n1164, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1173, new_n1174, new_n1175, new_n1176, new_n1177, new_n1178,
    new_n1179, new_n1180, new_n1181, new_n1182, new_n1183, new_n1184,
    new_n1185, new_n1186, new_n1187, new_n1188, new_n1190, new_n1191,
    new_n1192, new_n1193, new_n1194, new_n1195, new_n1196, new_n1197,
    new_n1198, new_n1199, new_n1200, new_n1201, new_n1202, new_n1203,
    new_n1204, new_n1205, new_n1206, new_n1207, new_n1208, new_n1209,
    new_n1210, new_n1211, new_n1212, new_n1213, new_n1214, new_n1215,
    new_n1216, new_n1217, new_n1218, new_n1219, new_n1220, new_n1221,
    new_n1222, new_n1223, new_n1224, new_n1225, new_n1226, new_n1227,
    new_n1228, new_n1229, new_n1230, new_n1231, new_n1232, new_n1233,
    new_n1234, new_n1235, new_n1236, new_n1237, new_n1238, new_n1239,
    new_n1240, new_n1241, new_n1242, new_n1243, new_n1244, new_n1245,
    new_n1246, new_n1247, new_n1248, new_n1250, new_n1251, new_n1252,
    new_n1253, new_n1254, new_n1255, new_n1256, new_n1257, new_n1258,
    new_n1259, new_n1260, new_n1261, new_n1262, new_n1263, new_n1264,
    new_n1265, new_n1266, new_n1267, new_n1268, new_n1269, new_n1270,
    new_n1271, new_n1272, new_n1273, new_n1274, new_n1275, new_n1276,
    new_n1277, new_n1278, new_n1279, new_n1280, new_n1281, new_n1282,
    new_n1283, new_n1284, new_n1285, new_n1286, new_n1287, new_n1288,
    new_n1289, new_n1290, new_n1291, new_n1292, new_n1293, new_n1294,
    new_n1295, new_n1296, new_n1297, new_n1298, new_n1299, new_n1300,
    new_n1301, new_n1302, new_n1303, new_n1304, new_n1305, new_n1306,
    new_n1307, new_n1308, new_n1309, new_n1310, new_n1312, new_n1313,
    new_n1314, new_n1315, new_n1316, new_n1317, new_n1318, new_n1319,
    new_n1320, new_n1321, new_n1322, new_n1323, new_n1324, new_n1325,
    new_n1326, new_n1327, new_n1328, new_n1330, new_n1331, new_n1332,
    new_n1333, new_n1334, new_n1336, new_n1337, new_n1338, new_n1339,
    new_n1340, new_n1342, new_n1343, new_n1344, new_n1345, new_n1346,
    new_n1347, new_n1348, new_n1349, new_n1350, new_n1351, new_n1352,
    new_n1353, new_n1354, new_n1355, new_n1356, new_n1357, new_n1358,
    new_n1359, new_n1360, new_n1361, new_n1362, new_n1363, new_n1364,
    new_n1365, new_n1366, new_n1367, new_n1368, new_n1369, new_n1370,
    new_n1371, new_n1372, new_n1373, new_n1374, new_n1375, new_n1376,
    new_n1377, new_n1378, new_n1379, new_n1380, new_n1381, new_n1382,
    new_n1383, new_n1384, new_n1385, new_n1386, new_n1387, new_n1388,
    new_n1389, new_n1390, new_n1391, new_n1392, new_n1393, new_n1394,
    new_n1395, new_n1396, new_n1397, new_n1398, new_n1399, new_n1400,
    new_n1401, new_n1402, new_n1403, new_n1404, new_n1405, new_n1406,
    new_n1407, new_n1408, new_n1409, new_n1410, new_n1411, new_n1412,
    new_n1414, new_n1415, new_n1416, new_n1417, new_n1418, new_n1419,
    new_n1420, new_n1421;
  INV_X1    g0000(.A(G58), .ZN(new_n201));
  INV_X1    g0001(.A(G68), .ZN(new_n202));
  NAND3_X1  g0002(.A1(new_n201), .A2(new_n202), .A3(KEYINPUT64), .ZN(new_n203));
  INV_X1    g0003(.A(KEYINPUT64), .ZN(new_n204));
  OAI21_X1  g0004(.A(new_n204), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n203), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  OAI21_X1  g0009(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0010(.A(G1), .ZN(new_n211));
  INV_X1    g0011(.A(G20), .ZN(new_n212));
  NOR2_X1   g0012(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g0013(.A(new_n213), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(G13), .ZN(new_n215));
  OAI211_X1 g0015(.A(new_n215), .B(G250), .C1(G257), .C2(G264), .ZN(new_n216));
  XNOR2_X1  g0016(.A(new_n216), .B(KEYINPUT65), .ZN(new_n217));
  XNOR2_X1  g0017(.A(new_n217), .B(KEYINPUT0), .ZN(new_n218));
  AOI22_X1  g0018(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n219));
  INV_X1    g0019(.A(G238), .ZN(new_n220));
  INV_X1    g0020(.A(G87), .ZN(new_n221));
  INV_X1    g0021(.A(G250), .ZN(new_n222));
  OAI221_X1 g0022(.A(new_n219), .B1(new_n202), .B2(new_n220), .C1(new_n221), .C2(new_n222), .ZN(new_n223));
  AOI22_X1  g0023(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n224));
  AOI22_X1  g0024(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n225));
  NAND2_X1  g0025(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  OAI21_X1  g0026(.A(new_n214), .B1(new_n223), .B2(new_n226), .ZN(new_n227));
  OR2_X1    g0027(.A1(new_n227), .A2(KEYINPUT1), .ZN(new_n228));
  XNOR2_X1  g0028(.A(new_n228), .B(KEYINPUT66), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR2_X1   g0030(.A1(new_n230), .A2(new_n212), .ZN(new_n231));
  NOR2_X1   g0031(.A1(new_n206), .A2(new_n207), .ZN(new_n232));
  AOI22_X1  g0032(.A1(new_n227), .A2(KEYINPUT1), .B1(new_n231), .B2(new_n232), .ZN(new_n233));
  AND3_X1   g0033(.A1(new_n218), .A2(new_n229), .A3(new_n233), .ZN(G361));
  XNOR2_X1  g0034(.A(G238), .B(G244), .ZN(new_n235));
  INV_X1    g0035(.A(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT2), .B(G226), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g0042(.A(new_n239), .B(new_n242), .ZN(G358));
  XOR2_X1   g0043(.A(G87), .B(G97), .Z(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n207), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n202), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n246), .B(new_n251), .ZN(G351));
  NAND2_X1  g0052(.A1(G33), .A2(G41), .ZN(new_n253));
  NAND3_X1  g0053(.A1(new_n253), .A2(G1), .A3(G13), .ZN(new_n254));
  INV_X1    g0054(.A(KEYINPUT67), .ZN(new_n255));
  OR2_X1    g0055(.A1(KEYINPUT3), .A2(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(KEYINPUT3), .A2(G33), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n256), .A2(new_n257), .ZN(new_n258));
  INV_X1    g0058(.A(G1698), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(G222), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n255), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  AOI21_X1  g0062(.A(G1698), .B1(new_n256), .B2(new_n257), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n263), .A2(KEYINPUT67), .A3(G222), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n262), .A2(new_n264), .ZN(new_n265));
  AOI21_X1  g0065(.A(new_n259), .B1(new_n256), .B2(new_n257), .ZN(new_n266));
  AND2_X1   g0066(.A1(KEYINPUT3), .A2(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(KEYINPUT3), .A2(G33), .ZN(new_n268));
  NOR2_X1   g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  AOI22_X1  g0069(.A1(new_n266), .A2(G223), .B1(new_n269), .B2(G77), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n254), .B1(new_n265), .B2(new_n270), .ZN(new_n271));
  INV_X1    g0071(.A(G41), .ZN(new_n272));
  INV_X1    g0072(.A(G45), .ZN(new_n273));
  AOI21_X1  g0073(.A(G1), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  NAND3_X1  g0074(.A1(new_n274), .A2(new_n254), .A3(G274), .ZN(new_n275));
  INV_X1    g0075(.A(G226), .ZN(new_n276));
  OAI21_X1  g0076(.A(new_n211), .B1(G41), .B2(G45), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n254), .A2(new_n277), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OR2_X1    g0079(.A1(new_n271), .A2(new_n279), .ZN(new_n280));
  INV_X1    g0080(.A(G169), .ZN(new_n281));
  NAND2_X1  g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n208), .A2(G20), .ZN(new_n283));
  INV_X1    g0083(.A(G150), .ZN(new_n284));
  NOR2_X1   g0084(.A1(G20), .A2(G33), .ZN(new_n285));
  INV_X1    g0085(.A(new_n285), .ZN(new_n286));
  INV_X1    g0086(.A(KEYINPUT8), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(G58), .ZN(new_n288));
  XNOR2_X1  g0088(.A(new_n288), .B(KEYINPUT70), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n201), .A2(KEYINPUT8), .ZN(new_n290));
  INV_X1    g0090(.A(KEYINPUT69), .ZN(new_n291));
  XNOR2_X1  g0091(.A(new_n290), .B(new_n291), .ZN(new_n292));
  AND2_X1   g0092(.A1(new_n289), .A2(new_n292), .ZN(new_n293));
  NAND2_X1  g0093(.A1(new_n212), .A2(G33), .ZN(new_n294));
  OAI221_X1 g0094(.A(new_n283), .B1(new_n284), .B2(new_n286), .C1(new_n293), .C2(new_n294), .ZN(new_n295));
  NAND3_X1  g0095(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT68), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n296), .A2(new_n297), .A3(new_n230), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n296), .B2(new_n230), .ZN(new_n299));
  OR2_X1    g0099(.A1(new_n298), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n295), .A2(new_n300), .ZN(new_n301));
  NOR2_X1   g0101(.A1(new_n298), .A2(new_n299), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n211), .A2(G13), .A3(G20), .ZN(new_n303));
  NAND2_X1  g0103(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g0104(.A1(new_n212), .A2(G1), .ZN(new_n305));
  NOR2_X1   g0105(.A1(new_n305), .A2(new_n207), .ZN(new_n306));
  INV_X1    g0106(.A(new_n306), .ZN(new_n307));
  OAI22_X1  g0107(.A1(new_n304), .A2(new_n307), .B1(G50), .B2(new_n303), .ZN(new_n308));
  INV_X1    g0108(.A(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n301), .A2(new_n309), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n271), .A2(new_n279), .ZN(new_n311));
  INV_X1    g0111(.A(G179), .ZN(new_n312));
  NAND2_X1  g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AND3_X1   g0113(.A1(new_n282), .A2(new_n310), .A3(new_n313), .ZN(new_n314));
  AOI21_X1  g0114(.A(new_n308), .B1(new_n295), .B2(new_n300), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n315), .A2(KEYINPUT9), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n280), .A2(G200), .ZN(new_n317));
  NAND2_X1  g0117(.A1(new_n311), .A2(G190), .ZN(new_n318));
  AND3_X1   g0118(.A1(new_n316), .A2(new_n317), .A3(new_n318), .ZN(new_n319));
  INV_X1    g0119(.A(KEYINPUT9), .ZN(new_n320));
  NAND3_X1  g0120(.A1(new_n310), .A2(KEYINPUT73), .A3(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(KEYINPUT73), .ZN(new_n322));
  OAI21_X1  g0122(.A(new_n322), .B1(new_n315), .B2(KEYINPUT9), .ZN(new_n323));
  NAND2_X1  g0123(.A1(new_n321), .A2(new_n323), .ZN(new_n324));
  NAND2_X1  g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n325), .A2(KEYINPUT10), .ZN(new_n326));
  INV_X1    g0126(.A(KEYINPUT10), .ZN(new_n327));
  NAND3_X1  g0127(.A1(new_n319), .A2(new_n324), .A3(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n314), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  NOR2_X1   g0129(.A1(new_n212), .A2(G68), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n330), .B1(G50), .B2(new_n285), .ZN(new_n331));
  INV_X1    g0131(.A(G77), .ZN(new_n332));
  OAI21_X1  g0132(.A(new_n331), .B1(new_n332), .B2(new_n294), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n333), .A2(new_n300), .A3(KEYINPUT11), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n211), .A2(G13), .ZN(new_n335));
  INV_X1    g0135(.A(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(KEYINPUT12), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n336), .B(new_n330), .C1(KEYINPUT74), .C2(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n337), .A2(KEYINPUT74), .ZN(new_n339));
  XNOR2_X1  g0139(.A(new_n338), .B(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(new_n303), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n296), .A2(new_n230), .ZN(new_n342));
  NOR2_X1   g0142(.A1(new_n341), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n305), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(G68), .A3(new_n344), .ZN(new_n345));
  NAND3_X1  g0145(.A1(new_n334), .A2(new_n340), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g0146(.A(KEYINPUT11), .B1(new_n333), .B2(new_n300), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(KEYINPUT14), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT13), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n276), .A2(new_n259), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n236), .A2(G1698), .ZN(new_n352));
  OAI211_X1 g0152(.A(new_n351), .B(new_n352), .C1(new_n267), .C2(new_n268), .ZN(new_n353));
  NAND2_X1  g0153(.A1(G33), .A2(G97), .ZN(new_n354));
  NAND2_X1  g0154(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  INV_X1    g0155(.A(new_n254), .ZN(new_n356));
  NAND2_X1  g0156(.A1(new_n355), .A2(new_n356), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n254), .A2(G238), .A3(new_n277), .ZN(new_n358));
  AND2_X1   g0158(.A1(new_n275), .A2(new_n358), .ZN(new_n359));
  AOI21_X1  g0159(.A(new_n350), .B1(new_n357), .B2(new_n359), .ZN(new_n360));
  AOI21_X1  g0160(.A(new_n254), .B1(new_n353), .B2(new_n354), .ZN(new_n361));
  NAND2_X1  g0161(.A1(new_n275), .A2(new_n358), .ZN(new_n362));
  NOR3_X1   g0162(.A1(new_n361), .A2(new_n362), .A3(KEYINPUT13), .ZN(new_n363));
  OAI211_X1 g0163(.A(new_n349), .B(G169), .C1(new_n360), .C2(new_n363), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n357), .A2(new_n359), .A3(new_n350), .ZN(new_n365));
  OAI21_X1  g0165(.A(KEYINPUT13), .B1(new_n361), .B2(new_n362), .ZN(new_n366));
  NAND3_X1  g0166(.A1(new_n365), .A2(G179), .A3(new_n366), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n364), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n365), .A2(new_n366), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n349), .B1(new_n369), .B2(G169), .ZN(new_n370));
  OAI21_X1  g0170(.A(KEYINPUT75), .B1(new_n368), .B2(new_n370), .ZN(new_n371));
  NOR2_X1   g0171(.A1(new_n360), .A2(new_n363), .ZN(new_n372));
  OAI21_X1  g0172(.A(KEYINPUT14), .B1(new_n372), .B2(new_n281), .ZN(new_n373));
  INV_X1    g0173(.A(KEYINPUT75), .ZN(new_n374));
  NAND4_X1  g0174(.A1(new_n373), .A2(new_n374), .A3(new_n367), .A4(new_n364), .ZN(new_n375));
  AOI21_X1  g0175(.A(new_n348), .B1(new_n371), .B2(new_n375), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n372), .A2(G190), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n369), .A2(G200), .ZN(new_n378));
  NAND3_X1  g0178(.A1(new_n348), .A2(new_n377), .A3(new_n378), .ZN(new_n379));
  INV_X1    g0179(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g0180(.A1(new_n376), .A2(new_n380), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n289), .A2(new_n292), .ZN(new_n382));
  NAND2_X1  g0182(.A1(new_n382), .A2(new_n344), .ZN(new_n383));
  OAI22_X1  g0183(.A1(new_n383), .A2(new_n304), .B1(new_n382), .B2(new_n303), .ZN(new_n384));
  INV_X1    g0184(.A(new_n342), .ZN(new_n385));
  NAND4_X1  g0185(.A1(new_n256), .A2(KEYINPUT7), .A3(new_n212), .A4(new_n257), .ZN(new_n386));
  NOR3_X1   g0186(.A1(new_n267), .A2(new_n268), .A3(G20), .ZN(new_n387));
  XNOR2_X1  g0187(.A(KEYINPUT76), .B(KEYINPUT7), .ZN(new_n388));
  OAI21_X1  g0188(.A(new_n386), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n389), .A2(G68), .ZN(new_n390));
  NAND2_X1  g0190(.A1(G58), .A2(G68), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n203), .A2(new_n205), .A3(new_n391), .ZN(new_n392));
  AOI22_X1  g0192(.A1(new_n392), .A2(G20), .B1(G159), .B2(new_n285), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n390), .A2(new_n393), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT16), .ZN(new_n395));
  AOI21_X1  g0195(.A(new_n385), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT7), .ZN(new_n397));
  OAI21_X1  g0197(.A(G68), .B1(new_n387), .B2(new_n397), .ZN(new_n398));
  NOR3_X1   g0198(.A1(new_n258), .A2(new_n388), .A3(G20), .ZN(new_n399));
  OAI211_X1 g0199(.A(new_n393), .B(KEYINPUT16), .C1(new_n398), .C2(new_n399), .ZN(new_n400));
  AOI21_X1  g0200(.A(new_n384), .B1(new_n396), .B2(new_n400), .ZN(new_n401));
  OR2_X1    g0201(.A1(G223), .A2(G1698), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n276), .A2(G1698), .ZN(new_n403));
  OAI211_X1 g0203(.A(new_n402), .B(new_n403), .C1(new_n267), .C2(new_n268), .ZN(new_n404));
  NAND2_X1  g0204(.A1(G33), .A2(G87), .ZN(new_n405));
  NAND2_X1  g0205(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n406), .A2(new_n356), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n254), .A2(G232), .A3(new_n277), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n275), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  AOI21_X1  g0210(.A(new_n281), .B1(new_n407), .B2(new_n410), .ZN(new_n411));
  AOI21_X1  g0211(.A(new_n254), .B1(new_n404), .B2(new_n405), .ZN(new_n412));
  NOR3_X1   g0212(.A1(new_n412), .A2(new_n409), .A3(new_n312), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n411), .A2(new_n413), .ZN(new_n414));
  OAI21_X1  g0214(.A(KEYINPUT18), .B1(new_n401), .B2(new_n414), .ZN(new_n415));
  AND2_X1   g0215(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n416));
  NOR2_X1   g0216(.A1(KEYINPUT76), .A2(KEYINPUT7), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  OAI21_X1  g0218(.A(new_n418), .B1(new_n258), .B2(G20), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n202), .B1(new_n419), .B2(new_n386), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n392), .A2(G20), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n285), .A2(G159), .ZN(new_n422));
  NAND2_X1  g0222(.A1(new_n421), .A2(new_n422), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n395), .B1(new_n420), .B2(new_n423), .ZN(new_n424));
  NAND3_X1  g0224(.A1(new_n424), .A2(new_n342), .A3(new_n400), .ZN(new_n425));
  INV_X1    g0225(.A(new_n304), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n305), .B1(new_n289), .B2(new_n292), .ZN(new_n427));
  AOI22_X1  g0227(.A1(new_n426), .A2(new_n427), .B1(new_n293), .B2(new_n341), .ZN(new_n428));
  AOI21_X1  g0228(.A(new_n414), .B1(new_n425), .B2(new_n428), .ZN(new_n429));
  INV_X1    g0229(.A(KEYINPUT18), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g0231(.A(G200), .ZN(new_n432));
  AOI21_X1  g0232(.A(new_n432), .B1(new_n407), .B2(new_n410), .ZN(new_n433));
  INV_X1    g0233(.A(G190), .ZN(new_n434));
  NOR3_X1   g0234(.A1(new_n412), .A2(new_n409), .A3(new_n434), .ZN(new_n435));
  NOR2_X1   g0235(.A1(new_n433), .A2(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n425), .A2(new_n436), .A3(new_n428), .ZN(new_n437));
  INV_X1    g0237(.A(KEYINPUT17), .ZN(new_n438));
  NAND2_X1  g0238(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  NAND4_X1  g0239(.A1(new_n425), .A2(new_n436), .A3(KEYINPUT17), .A4(new_n428), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n415), .A2(new_n431), .A3(new_n439), .A4(new_n440), .ZN(new_n441));
  OR2_X1    g0241(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n288), .A2(new_n290), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n286), .A2(KEYINPUT72), .ZN(new_n444));
  NAND3_X1  g0244(.A1(new_n442), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  XNOR2_X1  g0245(.A(KEYINPUT15), .B(G87), .ZN(new_n446));
  INV_X1    g0246(.A(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n294), .ZN(new_n448));
  AOI22_X1  g0248(.A1(new_n447), .A2(new_n448), .B1(G20), .B2(G77), .ZN(new_n449));
  AOI21_X1  g0249(.A(new_n385), .B1(new_n445), .B2(new_n449), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n343), .A2(G77), .A3(new_n344), .ZN(new_n451));
  OAI21_X1  g0251(.A(new_n451), .B1(G77), .B2(new_n303), .ZN(new_n452));
  NOR2_X1   g0252(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(new_n266), .A2(G238), .ZN(new_n454));
  INV_X1    g0254(.A(G107), .ZN(new_n455));
  OAI221_X1 g0255(.A(new_n454), .B1(new_n455), .B2(new_n258), .C1(new_n236), .C2(new_n260), .ZN(new_n456));
  NAND2_X1  g0256(.A1(new_n456), .A2(new_n356), .ZN(new_n457));
  INV_X1    g0257(.A(G244), .ZN(new_n458));
  NOR2_X1   g0258(.A1(new_n278), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(G274), .ZN(new_n460));
  AND2_X1   g0260(.A1(G1), .A2(G13), .ZN(new_n461));
  AOI21_X1  g0261(.A(new_n460), .B1(new_n461), .B2(new_n253), .ZN(new_n462));
  AOI21_X1  g0262(.A(new_n459), .B1(new_n274), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n457), .A2(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n453), .B1(new_n464), .B2(new_n281), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n465), .B1(G179), .B2(new_n464), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n464), .A2(G200), .ZN(new_n467));
  AND2_X1   g0267(.A1(new_n457), .A2(new_n463), .ZN(new_n468));
  AOI22_X1  g0268(.A1(new_n467), .A2(KEYINPUT71), .B1(new_n468), .B2(G190), .ZN(new_n469));
  NAND4_X1  g0269(.A1(new_n457), .A2(KEYINPUT71), .A3(G190), .A4(new_n463), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n470), .A2(new_n453), .ZN(new_n471));
  OAI21_X1  g0271(.A(new_n466), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  NOR2_X1   g0272(.A1(new_n441), .A2(new_n472), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n329), .A2(new_n381), .A3(new_n473), .ZN(new_n474));
  NOR2_X1   g0274(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n211), .A2(G45), .ZN(new_n476));
  OAI21_X1  g0276(.A(KEYINPUT79), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n273), .A2(G1), .ZN(new_n478));
  INV_X1    g0278(.A(KEYINPUT79), .ZN(new_n479));
  INV_X1    g0279(.A(KEYINPUT5), .ZN(new_n480));
  NAND2_X1  g0280(.A1(new_n480), .A2(G41), .ZN(new_n481));
  NAND3_X1  g0281(.A1(new_n478), .A2(new_n479), .A3(new_n481), .ZN(new_n482));
  NAND2_X1  g0282(.A1(new_n272), .A2(KEYINPUT5), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n477), .A2(new_n482), .A3(new_n462), .A4(new_n483), .ZN(new_n484));
  NAND3_X1  g0284(.A1(new_n478), .A2(new_n481), .A3(new_n483), .ZN(new_n485));
  NAND3_X1  g0285(.A1(new_n485), .A2(G270), .A3(new_n254), .ZN(new_n486));
  AND2_X1   g0286(.A1(new_n484), .A2(new_n486), .ZN(new_n487));
  OAI211_X1 g0287(.A(G264), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n488));
  NAND3_X1  g0288(.A1(new_n256), .A2(G303), .A3(new_n257), .ZN(new_n489));
  NAND2_X1  g0289(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  OAI211_X1 g0290(.A(G257), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n491));
  INV_X1    g0291(.A(KEYINPUT83), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n258), .A2(KEYINPUT83), .A3(G257), .A4(new_n259), .ZN(new_n494));
  AOI21_X1  g0294(.A(new_n490), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  OAI211_X1 g0295(.A(new_n487), .B(G190), .C1(new_n254), .C2(new_n495), .ZN(new_n496));
  INV_X1    g0296(.A(G116), .ZN(new_n497));
  AOI22_X1  g0297(.A1(new_n296), .A2(new_n230), .B1(G20), .B2(new_n497), .ZN(new_n498));
  NAND2_X1  g0298(.A1(G33), .A2(G283), .ZN(new_n499));
  INV_X1    g0299(.A(G97), .ZN(new_n500));
  OAI211_X1 g0300(.A(new_n499), .B(new_n212), .C1(G33), .C2(new_n500), .ZN(new_n501));
  NAND2_X1  g0301(.A1(new_n498), .A2(new_n501), .ZN(new_n502));
  INV_X1    g0302(.A(KEYINPUT20), .ZN(new_n503));
  NAND2_X1  g0303(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  NAND3_X1  g0304(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n501), .ZN(new_n505));
  NAND2_X1  g0305(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND2_X1  g0306(.A1(new_n211), .A2(G33), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(G116), .ZN(new_n508));
  INV_X1    g0308(.A(new_n508), .ZN(new_n509));
  NOR2_X1   g0309(.A1(new_n212), .A2(G116), .ZN(new_n510));
  AOI22_X1  g0310(.A1(new_n343), .A2(new_n509), .B1(new_n336), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g0312(.A(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n484), .A2(new_n486), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n493), .A2(new_n494), .ZN(new_n515));
  INV_X1    g0315(.A(new_n490), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n515), .A2(new_n516), .ZN(new_n517));
  AOI21_X1  g0317(.A(new_n514), .B1(new_n517), .B2(new_n356), .ZN(new_n518));
  OAI211_X1 g0318(.A(new_n496), .B(new_n513), .C1(new_n518), .C2(new_n432), .ZN(new_n519));
  INV_X1    g0319(.A(KEYINPUT84), .ZN(new_n520));
  NAND2_X1  g0320(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n487), .B1(new_n495), .B2(new_n254), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(G200), .ZN(new_n523));
  NAND4_X1  g0323(.A1(new_n523), .A2(KEYINPUT84), .A3(new_n513), .A4(new_n496), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n521), .A2(new_n524), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT85), .ZN(new_n526));
  INV_X1    g0326(.A(KEYINPUT21), .ZN(new_n527));
  AND3_X1   g0327(.A1(new_n498), .A2(KEYINPUT20), .A3(new_n501), .ZN(new_n528));
  AOI21_X1  g0328(.A(KEYINPUT20), .B1(new_n498), .B2(new_n501), .ZN(new_n529));
  NOR2_X1   g0329(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n343), .A2(new_n509), .ZN(new_n531));
  NAND2_X1  g0331(.A1(new_n336), .A2(new_n510), .ZN(new_n532));
  NAND2_X1  g0332(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n530), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n527), .B1(new_n518), .B2(new_n534), .ZN(new_n535));
  AOI21_X1  g0335(.A(new_n281), .B1(new_n506), .B2(new_n511), .ZN(new_n536));
  NAND3_X1  g0336(.A1(new_n522), .A2(KEYINPUT21), .A3(new_n536), .ZN(new_n537));
  NAND2_X1  g0337(.A1(new_n517), .A2(new_n356), .ZN(new_n538));
  NAND4_X1  g0338(.A1(new_n538), .A2(G179), .A3(new_n487), .A4(new_n512), .ZN(new_n539));
  NAND3_X1  g0339(.A1(new_n535), .A2(new_n537), .A3(new_n539), .ZN(new_n540));
  INV_X1    g0340(.A(new_n540), .ZN(new_n541));
  AND3_X1   g0341(.A1(new_n525), .A2(new_n526), .A3(new_n541), .ZN(new_n542));
  AOI21_X1  g0342(.A(new_n526), .B1(new_n525), .B2(new_n541), .ZN(new_n543));
  NOR2_X1   g0343(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  INV_X1    g0344(.A(KEYINPUT6), .ZN(new_n545));
  NOR3_X1   g0345(.A1(new_n545), .A2(G97), .A3(G107), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n500), .A2(KEYINPUT6), .ZN(new_n547));
  AND2_X1   g0347(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n548));
  NOR2_X1   g0348(.A1(new_n455), .A2(KEYINPUT77), .ZN(new_n549));
  OAI22_X1  g0349(.A1(new_n546), .A2(new_n547), .B1(new_n548), .B2(new_n549), .ZN(new_n550));
  XNOR2_X1  g0350(.A(KEYINPUT77), .B(G107), .ZN(new_n551));
  NAND3_X1  g0351(.A1(new_n500), .A2(new_n455), .A3(KEYINPUT6), .ZN(new_n552));
  NAND2_X1  g0352(.A1(new_n545), .A2(G97), .ZN(new_n553));
  NAND3_X1  g0353(.A1(new_n551), .A2(new_n552), .A3(new_n553), .ZN(new_n554));
  NAND3_X1  g0354(.A1(new_n550), .A2(new_n554), .A3(G20), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n285), .A2(G77), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n555), .A2(new_n556), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n455), .B1(new_n419), .B2(new_n386), .ZN(new_n558));
  OAI21_X1  g0358(.A(new_n342), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NOR2_X1   g0359(.A1(new_n303), .A2(G97), .ZN(new_n560));
  AND3_X1   g0360(.A1(new_n302), .A2(new_n303), .A3(new_n507), .ZN(new_n561));
  AOI21_X1  g0361(.A(new_n560), .B1(new_n561), .B2(G97), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n559), .A2(new_n562), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT78), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n499), .B1(new_n564), .B2(KEYINPUT4), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(KEYINPUT4), .ZN(new_n566));
  NAND2_X1  g0366(.A1(new_n259), .A2(G244), .ZN(new_n567));
  OAI22_X1  g0367(.A1(new_n566), .A2(new_n567), .B1(new_n222), .B2(new_n259), .ZN(new_n568));
  AOI21_X1  g0368(.A(new_n565), .B1(new_n568), .B2(new_n258), .ZN(new_n569));
  OAI211_X1 g0369(.A(G244), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n570), .A2(new_n566), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n254), .B1(new_n569), .B2(new_n571), .ZN(new_n572));
  NAND3_X1  g0372(.A1(new_n485), .A2(G257), .A3(new_n254), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n484), .A2(new_n573), .ZN(new_n574));
  OAI21_X1  g0374(.A(new_n281), .B1(new_n572), .B2(new_n574), .ZN(new_n575));
  INV_X1    g0375(.A(new_n565), .ZN(new_n576));
  INV_X1    g0376(.A(KEYINPUT4), .ZN(new_n577));
  NOR2_X1   g0377(.A1(new_n577), .A2(KEYINPUT78), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n458), .A2(G1698), .ZN(new_n579));
  AOI22_X1  g0379(.A1(new_n578), .A2(new_n579), .B1(G250), .B2(G1698), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n576), .B1(new_n580), .B2(new_n269), .ZN(new_n581));
  AOI21_X1  g0381(.A(new_n578), .B1(new_n263), .B2(G244), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n356), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  AND2_X1   g0383(.A1(new_n484), .A2(new_n573), .ZN(new_n584));
  NAND3_X1  g0384(.A1(new_n583), .A2(new_n312), .A3(new_n584), .ZN(new_n585));
  NAND3_X1  g0385(.A1(new_n563), .A2(new_n575), .A3(new_n585), .ZN(new_n586));
  INV_X1    g0386(.A(new_n560), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n302), .A2(new_n303), .A3(new_n507), .ZN(new_n588));
  OAI21_X1  g0388(.A(new_n587), .B1(new_n588), .B2(new_n500), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n389), .A2(G107), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n590), .A2(new_n556), .A3(new_n555), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n589), .B1(new_n342), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n572), .A2(new_n574), .ZN(new_n593));
  AOI21_X1  g0393(.A(KEYINPUT81), .B1(new_n593), .B2(G190), .ZN(new_n594));
  NAND3_X1  g0394(.A1(new_n583), .A2(G190), .A3(new_n584), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT81), .ZN(new_n596));
  NOR2_X1   g0396(.A1(new_n595), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g0397(.A(new_n592), .B1(new_n594), .B2(new_n597), .ZN(new_n598));
  OAI21_X1  g0398(.A(G200), .B1(new_n572), .B2(new_n574), .ZN(new_n599));
  INV_X1    g0399(.A(KEYINPUT80), .ZN(new_n600));
  NAND2_X1  g0400(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n583), .A2(new_n584), .ZN(new_n602));
  NAND3_X1  g0402(.A1(new_n602), .A2(KEYINPUT80), .A3(G200), .ZN(new_n603));
  AND2_X1   g0403(.A1(new_n601), .A2(new_n603), .ZN(new_n604));
  OAI21_X1  g0404(.A(new_n586), .B1(new_n598), .B2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n303), .A2(G107), .ZN(new_n606));
  XNOR2_X1  g0406(.A(KEYINPUT87), .B(KEYINPUT25), .ZN(new_n607));
  XNOR2_X1  g0407(.A(new_n606), .B(new_n607), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n608), .B1(new_n588), .B2(new_n455), .ZN(new_n609));
  INV_X1    g0409(.A(KEYINPUT23), .ZN(new_n610));
  OAI21_X1  g0410(.A(new_n610), .B1(new_n212), .B2(G107), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n455), .A2(KEYINPUT23), .A3(G20), .ZN(new_n612));
  NAND2_X1  g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  INV_X1    g0413(.A(G33), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n614), .A2(new_n497), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n615), .A2(new_n212), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n212), .B(G87), .C1(new_n267), .C2(new_n268), .ZN(new_n617));
  XNOR2_X1  g0417(.A(KEYINPUT86), .B(KEYINPUT22), .ZN(new_n618));
  OAI211_X1 g0418(.A(new_n613), .B(new_n616), .C1(new_n617), .C2(new_n618), .ZN(new_n619));
  NOR2_X1   g0419(.A1(KEYINPUT86), .A2(KEYINPUT22), .ZN(new_n620));
  AND2_X1   g0420(.A1(new_n617), .A2(new_n620), .ZN(new_n621));
  OAI21_X1  g0421(.A(KEYINPUT24), .B1(new_n619), .B2(new_n621), .ZN(new_n622));
  INV_X1    g0422(.A(new_n618), .ZN(new_n623));
  NAND4_X1  g0423(.A1(new_n623), .A2(new_n212), .A3(G87), .A4(new_n258), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n617), .A2(new_n620), .ZN(new_n625));
  INV_X1    g0425(.A(KEYINPUT24), .ZN(new_n626));
  AOI22_X1  g0426(.A1(new_n611), .A2(new_n612), .B1(new_n615), .B2(new_n212), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n624), .A2(new_n625), .A3(new_n626), .A4(new_n627), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n622), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n609), .B1(new_n629), .B2(new_n342), .ZN(new_n630));
  INV_X1    g0430(.A(G294), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n631), .A2(KEYINPUT89), .ZN(new_n632));
  INV_X1    g0432(.A(KEYINPUT89), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n633), .A2(G294), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  AOI22_X1  g0435(.A1(new_n266), .A2(G257), .B1(new_n635), .B2(G33), .ZN(new_n636));
  INV_X1    g0436(.A(KEYINPUT88), .ZN(new_n637));
  AOI21_X1  g0437(.A(new_n637), .B1(new_n263), .B2(G250), .ZN(new_n638));
  OAI211_X1 g0438(.A(G250), .B(new_n259), .C1(new_n267), .C2(new_n268), .ZN(new_n639));
  NOR2_X1   g0439(.A1(new_n639), .A2(KEYINPUT88), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n636), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND3_X1  g0441(.A1(new_n485), .A2(G264), .A3(new_n254), .ZN(new_n642));
  INV_X1    g0442(.A(KEYINPUT90), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND4_X1  g0444(.A1(new_n485), .A2(KEYINPUT90), .A3(G264), .A4(new_n254), .ZN(new_n645));
  AOI22_X1  g0445(.A1(new_n641), .A2(new_n356), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g0446(.A(G200), .B1(new_n646), .B2(new_n484), .ZN(new_n647));
  NAND2_X1  g0447(.A1(new_n639), .A2(KEYINPUT88), .ZN(new_n648));
  NAND4_X1  g0448(.A1(new_n258), .A2(new_n637), .A3(G250), .A4(new_n259), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n648), .A2(new_n649), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n254), .B1(new_n650), .B2(new_n636), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n484), .A2(new_n642), .ZN(new_n652));
  NOR3_X1   g0452(.A1(new_n651), .A2(G190), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g0453(.A(new_n630), .B1(new_n647), .B2(new_n653), .ZN(new_n654));
  OAI21_X1  g0454(.A(G169), .B1(new_n651), .B2(new_n652), .ZN(new_n655));
  NAND2_X1  g0455(.A1(new_n644), .A2(new_n645), .ZN(new_n656));
  OAI211_X1 g0456(.A(G257), .B(G1698), .C1(new_n267), .C2(new_n268), .ZN(new_n657));
  XNOR2_X1  g0457(.A(KEYINPUT89), .B(G294), .ZN(new_n658));
  OAI21_X1  g0458(.A(new_n657), .B1(new_n614), .B2(new_n658), .ZN(new_n659));
  AOI21_X1  g0459(.A(new_n659), .B1(new_n649), .B2(new_n648), .ZN(new_n660));
  OAI211_X1 g0460(.A(new_n484), .B(new_n656), .C1(new_n660), .C2(new_n254), .ZN(new_n661));
  OAI21_X1  g0461(.A(new_n655), .B1(new_n661), .B2(new_n312), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n629), .A2(new_n342), .ZN(new_n663));
  INV_X1    g0463(.A(new_n609), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n663), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n662), .A2(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(KEYINPUT82), .ZN(new_n667));
  NAND2_X1  g0467(.A1(new_n220), .A2(new_n259), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n458), .A2(G1698), .ZN(new_n669));
  OAI211_X1 g0469(.A(new_n668), .B(new_n669), .C1(new_n267), .C2(new_n268), .ZN(new_n670));
  INV_X1    g0470(.A(new_n615), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n254), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  NAND2_X1  g0472(.A1(new_n476), .A2(new_n222), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n211), .A2(new_n460), .A3(G45), .ZN(new_n674));
  NAND3_X1  g0474(.A1(new_n673), .A2(new_n254), .A3(new_n674), .ZN(new_n675));
  INV_X1    g0475(.A(new_n675), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n667), .B1(new_n672), .B2(new_n676), .ZN(new_n677));
  NOR2_X1   g0477(.A1(G238), .A2(G1698), .ZN(new_n678));
  AOI21_X1  g0478(.A(new_n678), .B1(new_n458), .B2(G1698), .ZN(new_n679));
  AOI21_X1  g0479(.A(new_n615), .B1(new_n679), .B2(new_n258), .ZN(new_n680));
  OAI211_X1 g0480(.A(KEYINPUT82), .B(new_n675), .C1(new_n680), .C2(new_n254), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n677), .A2(new_n681), .A3(new_n312), .ZN(new_n682));
  INV_X1    g0482(.A(KEYINPUT19), .ZN(new_n683));
  OAI21_X1  g0483(.A(new_n212), .B1(new_n354), .B2(new_n683), .ZN(new_n684));
  NAND3_X1  g0484(.A1(new_n221), .A2(new_n500), .A3(new_n455), .ZN(new_n685));
  NAND2_X1  g0485(.A1(new_n684), .A2(new_n685), .ZN(new_n686));
  OAI211_X1 g0486(.A(new_n212), .B(G68), .C1(new_n267), .C2(new_n268), .ZN(new_n687));
  OAI21_X1  g0487(.A(new_n683), .B1(new_n294), .B2(new_n500), .ZN(new_n688));
  NAND3_X1  g0488(.A1(new_n686), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n689), .A2(new_n342), .ZN(new_n690));
  NAND2_X1  g0490(.A1(new_n446), .A2(new_n341), .ZN(new_n691));
  OAI211_X1 g0491(.A(new_n690), .B(new_n691), .C1(new_n588), .C2(new_n446), .ZN(new_n692));
  AND2_X1   g0492(.A1(new_n677), .A2(new_n681), .ZN(new_n693));
  OAI211_X1 g0493(.A(new_n682), .B(new_n692), .C1(new_n693), .C2(G169), .ZN(new_n694));
  NAND3_X1  g0494(.A1(new_n677), .A2(new_n681), .A3(G190), .ZN(new_n695));
  NAND4_X1  g0495(.A1(new_n302), .A2(G87), .A3(new_n303), .A4(new_n507), .ZN(new_n696));
  AND3_X1   g0496(.A1(new_n696), .A2(new_n690), .A3(new_n691), .ZN(new_n697));
  OAI211_X1 g0497(.A(new_n695), .B(new_n697), .C1(new_n693), .C2(new_n432), .ZN(new_n698));
  NAND4_X1  g0498(.A1(new_n654), .A2(new_n666), .A3(new_n694), .A4(new_n698), .ZN(new_n699));
  NOR4_X1   g0499(.A1(new_n474), .A2(new_n544), .A3(new_n605), .A4(new_n699), .ZN(G372));
  INV_X1    g0500(.A(new_n474), .ZN(new_n701));
  NAND3_X1  g0501(.A1(new_n646), .A2(G179), .A3(new_n484), .ZN(new_n702));
  AOI21_X1  g0502(.A(new_n630), .B1(new_n655), .B2(new_n702), .ZN(new_n703));
  OAI21_X1  g0503(.A(KEYINPUT91), .B1(new_n703), .B2(new_n540), .ZN(new_n704));
  AND2_X1   g0504(.A1(new_n537), .A2(new_n539), .ZN(new_n705));
  INV_X1    g0505(.A(KEYINPUT91), .ZN(new_n706));
  NAND4_X1  g0506(.A1(new_n666), .A2(new_n705), .A3(new_n706), .A4(new_n535), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n575), .A2(new_n585), .ZN(new_n708));
  NOR2_X1   g0508(.A1(new_n708), .A2(new_n592), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n593), .A2(KEYINPUT81), .A3(G190), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n595), .A2(new_n596), .ZN(new_n711));
  AOI21_X1  g0511(.A(new_n563), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  NAND2_X1  g0512(.A1(new_n601), .A2(new_n603), .ZN(new_n713));
  AOI21_X1  g0513(.A(new_n709), .B1(new_n712), .B2(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n675), .B1(new_n680), .B2(new_n254), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n715), .A2(G200), .ZN(new_n716));
  NAND3_X1  g0516(.A1(new_n695), .A2(new_n697), .A3(new_n716), .ZN(new_n717));
  NAND2_X1  g0517(.A1(new_n715), .A2(new_n281), .ZN(new_n718));
  NAND3_X1  g0518(.A1(new_n682), .A2(new_n718), .A3(new_n692), .ZN(new_n719));
  NAND2_X1  g0519(.A1(new_n717), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n661), .A2(new_n432), .ZN(new_n721));
  OR3_X1    g0521(.A1(new_n651), .A2(G190), .A3(new_n652), .ZN(new_n722));
  NAND2_X1  g0522(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n720), .B1(new_n723), .B2(new_n630), .ZN(new_n724));
  NAND4_X1  g0524(.A1(new_n704), .A2(new_n707), .A3(new_n714), .A4(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n719), .ZN(new_n726));
  INV_X1    g0526(.A(KEYINPUT26), .ZN(new_n727));
  OAI21_X1  g0527(.A(new_n727), .B1(new_n586), .B2(new_n720), .ZN(new_n728));
  XOR2_X1   g0528(.A(KEYINPUT92), .B(KEYINPUT26), .Z(new_n729));
  INV_X1    g0529(.A(new_n729), .ZN(new_n730));
  NAND4_X1  g0530(.A1(new_n709), .A2(new_n694), .A3(new_n698), .A4(new_n730), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n726), .B1(new_n728), .B2(new_n731), .ZN(new_n732));
  NAND2_X1  g0532(.A1(new_n725), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n701), .A2(new_n733), .ZN(new_n734));
  NAND2_X1  g0534(.A1(new_n326), .A2(new_n328), .ZN(new_n735));
  AND2_X1   g0535(.A1(new_n439), .A2(new_n440), .ZN(new_n736));
  NOR2_X1   g0536(.A1(new_n466), .A2(new_n380), .ZN(new_n737));
  OAI21_X1  g0537(.A(new_n736), .B1(new_n376), .B2(new_n737), .ZN(new_n738));
  INV_X1    g0538(.A(KEYINPUT93), .ZN(new_n739));
  AOI211_X1 g0539(.A(KEYINPUT18), .B(new_n414), .C1(new_n428), .C2(new_n425), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n425), .A2(new_n428), .ZN(new_n741));
  INV_X1    g0541(.A(new_n414), .ZN(new_n742));
  AOI21_X1  g0542(.A(new_n430), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  OAI21_X1  g0543(.A(new_n739), .B1(new_n740), .B2(new_n743), .ZN(new_n744));
  NAND3_X1  g0544(.A1(new_n415), .A2(KEYINPUT93), .A3(new_n431), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n738), .A2(new_n746), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n314), .B1(new_n735), .B2(new_n747), .ZN(new_n748));
  NAND2_X1  g0548(.A1(new_n734), .A2(new_n748), .ZN(G369));
  OR3_X1    g0549(.A1(new_n335), .A2(KEYINPUT27), .A3(G20), .ZN(new_n750));
  OAI21_X1  g0550(.A(KEYINPUT27), .B1(new_n335), .B2(G20), .ZN(new_n751));
  NAND3_X1  g0551(.A1(new_n750), .A2(G213), .A3(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(new_n752), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G343), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n513), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g0555(.A1(new_n540), .A2(new_n755), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  OAI21_X1  g0557(.A(new_n757), .B1(new_n544), .B2(new_n755), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n758), .A2(G330), .ZN(new_n759));
  OAI211_X1 g0559(.A(new_n654), .B(new_n666), .C1(new_n630), .C2(new_n754), .ZN(new_n760));
  INV_X1    g0560(.A(new_n754), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n703), .A2(new_n761), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n760), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n759), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(new_n765), .ZN(new_n766));
  NAND4_X1  g0566(.A1(new_n654), .A2(new_n666), .A3(new_n540), .A4(new_n754), .ZN(new_n767));
  NAND2_X1  g0567(.A1(new_n703), .A2(new_n754), .ZN(new_n768));
  AOI21_X1  g0568(.A(KEYINPUT94), .B1(new_n767), .B2(new_n768), .ZN(new_n769));
  NAND3_X1  g0569(.A1(new_n767), .A2(KEYINPUT94), .A3(new_n768), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n766), .B1(new_n769), .B2(new_n771), .ZN(G399));
  NOR2_X1   g0572(.A1(new_n685), .A2(G116), .ZN(new_n773));
  XOR2_X1   g0573(.A(new_n773), .B(KEYINPUT95), .Z(new_n774));
  INV_X1    g0574(.A(new_n215), .ZN(new_n775));
  NOR2_X1   g0575(.A1(new_n775), .A2(G41), .ZN(new_n776));
  NOR3_X1   g0576(.A1(new_n774), .A2(new_n776), .A3(new_n211), .ZN(new_n777));
  AOI21_X1  g0577(.A(new_n777), .B1(new_n232), .B2(new_n776), .ZN(new_n778));
  XOR2_X1   g0578(.A(new_n778), .B(KEYINPUT28), .Z(new_n779));
  INV_X1    g0579(.A(G330), .ZN(new_n780));
  INV_X1    g0580(.A(KEYINPUT30), .ZN(new_n781));
  NAND3_X1  g0581(.A1(new_n693), .A2(new_n646), .A3(new_n593), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n518), .A2(G179), .ZN(new_n783));
  OAI21_X1  g0583(.A(new_n781), .B1(new_n782), .B2(new_n783), .ZN(new_n784));
  NOR2_X1   g0584(.A1(new_n522), .A2(new_n312), .ZN(new_n785));
  AND4_X1   g0585(.A1(new_n583), .A2(new_n584), .A3(new_n677), .A4(new_n681), .ZN(new_n786));
  NAND4_X1  g0586(.A1(new_n785), .A2(new_n786), .A3(KEYINPUT30), .A4(new_n646), .ZN(new_n787));
  NAND3_X1  g0587(.A1(new_n661), .A2(KEYINPUT97), .A3(new_n602), .ZN(new_n788));
  NAND2_X1  g0588(.A1(new_n715), .A2(new_n312), .ZN(new_n789));
  OAI21_X1  g0589(.A(KEYINPUT96), .B1(new_n518), .B2(new_n789), .ZN(new_n790));
  INV_X1    g0590(.A(KEYINPUT96), .ZN(new_n791));
  NAND4_X1  g0591(.A1(new_n522), .A2(new_n791), .A3(new_n312), .A4(new_n715), .ZN(new_n792));
  NAND3_X1  g0592(.A1(new_n788), .A2(new_n790), .A3(new_n792), .ZN(new_n793));
  AOI21_X1  g0593(.A(KEYINPUT97), .B1(new_n661), .B2(new_n602), .ZN(new_n794));
  OAI211_X1 g0594(.A(new_n784), .B(new_n787), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  AND3_X1   g0595(.A1(new_n795), .A2(KEYINPUT31), .A3(new_n761), .ZN(new_n796));
  AOI21_X1  g0596(.A(KEYINPUT31), .B1(new_n795), .B2(new_n761), .ZN(new_n797));
  NOR2_X1   g0597(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n699), .A2(new_n605), .ZN(new_n799));
  OAI211_X1 g0599(.A(new_n799), .B(new_n754), .C1(new_n542), .C2(new_n543), .ZN(new_n800));
  AOI21_X1  g0600(.A(new_n780), .B1(new_n798), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g0601(.A1(new_n666), .A2(new_n705), .A3(new_n535), .ZN(new_n802));
  NAND3_X1  g0602(.A1(new_n714), .A2(new_n802), .A3(new_n724), .ZN(new_n803));
  INV_X1    g0603(.A(KEYINPUT98), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n695), .A2(new_n697), .ZN(new_n805));
  AOI21_X1  g0605(.A(new_n432), .B1(new_n677), .B2(new_n681), .ZN(new_n806));
  NAND2_X1  g0606(.A1(new_n682), .A2(new_n692), .ZN(new_n807));
  AOI21_X1  g0607(.A(G169), .B1(new_n677), .B2(new_n681), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n805), .A2(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI211_X1 g0609(.A(new_n804), .B(new_n729), .C1(new_n809), .C2(new_n586), .ZN(new_n810));
  NAND4_X1  g0610(.A1(new_n709), .A2(KEYINPUT26), .A3(new_n719), .A4(new_n717), .ZN(new_n811));
  NAND2_X1  g0611(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n709), .A2(new_n694), .A3(new_n698), .ZN(new_n813));
  AOI21_X1  g0613(.A(new_n804), .B1(new_n813), .B2(new_n729), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n719), .B(new_n803), .C1(new_n812), .C2(new_n814), .ZN(new_n815));
  AND3_X1   g0615(.A1(new_n815), .A2(KEYINPUT99), .A3(new_n754), .ZN(new_n816));
  AOI21_X1  g0616(.A(KEYINPUT99), .B1(new_n815), .B2(new_n754), .ZN(new_n817));
  OAI21_X1  g0617(.A(KEYINPUT29), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n733), .A2(new_n754), .ZN(new_n819));
  INV_X1    g0619(.A(KEYINPUT29), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  AOI21_X1  g0621(.A(new_n801), .B1(new_n818), .B2(new_n821), .ZN(new_n822));
  OAI21_X1  g0622(.A(new_n779), .B1(new_n822), .B2(G1), .ZN(G364));
  AND2_X1   g0623(.A1(new_n212), .A2(G13), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n824), .A2(G45), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(G1), .ZN(new_n826));
  OR3_X1    g0626(.A1(new_n776), .A2(KEYINPUT100), .A3(new_n826), .ZN(new_n827));
  OAI21_X1  g0627(.A(KEYINPUT100), .B1(new_n776), .B2(new_n826), .ZN(new_n828));
  NAND2_X1  g0628(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  INV_X1    g0629(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n830), .B1(new_n758), .B2(G330), .ZN(new_n831));
  OAI21_X1  g0631(.A(new_n831), .B1(G330), .B2(new_n758), .ZN(new_n832));
  AOI21_X1  g0632(.A(new_n230), .B1(G20), .B2(new_n281), .ZN(new_n833));
  INV_X1    g0633(.A(new_n833), .ZN(new_n834));
  NOR2_X1   g0634(.A1(new_n212), .A2(G190), .ZN(new_n835));
  NOR2_X1   g0635(.A1(new_n312), .A2(G200), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  AND2_X1   g0637(.A1(new_n837), .A2(KEYINPUT103), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n837), .A2(KEYINPUT103), .ZN(new_n839));
  NOR2_X1   g0639(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n840), .A2(new_n332), .ZN(new_n841));
  NAND2_X1  g0641(.A1(new_n312), .A2(new_n432), .ZN(new_n842));
  XNOR2_X1  g0642(.A(new_n842), .B(KEYINPUT104), .ZN(new_n843));
  INV_X1    g0643(.A(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n844), .A2(new_n835), .ZN(new_n845));
  INV_X1    g0645(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n846), .A2(G159), .ZN(new_n847));
  XNOR2_X1  g0647(.A(new_n847), .B(KEYINPUT32), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n212), .A2(G179), .ZN(new_n849));
  NAND3_X1  g0649(.A1(new_n849), .A2(G190), .A3(G200), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n836), .A2(G20), .A3(G190), .ZN(new_n851));
  INV_X1    g0651(.A(KEYINPUT102), .ZN(new_n852));
  NAND2_X1  g0652(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  INV_X1    g0653(.A(new_n853), .ZN(new_n854));
  NOR2_X1   g0654(.A1(new_n851), .A2(new_n852), .ZN(new_n855));
  NOR2_X1   g0655(.A1(new_n854), .A2(new_n855), .ZN(new_n856));
  OAI221_X1 g0656(.A(new_n258), .B1(new_n221), .B2(new_n850), .C1(new_n856), .C2(new_n201), .ZN(new_n857));
  AOI21_X1  g0657(.A(new_n212), .B1(new_n844), .B2(G190), .ZN(new_n858));
  INV_X1    g0658(.A(new_n858), .ZN(new_n859));
  NAND2_X1  g0659(.A1(new_n859), .A2(G97), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n849), .A2(new_n434), .A3(G200), .ZN(new_n861));
  INV_X1    g0661(.A(new_n861), .ZN(new_n862));
  NAND3_X1  g0662(.A1(G20), .A2(G179), .A3(G200), .ZN(new_n863));
  NOR2_X1   g0663(.A1(new_n863), .A2(new_n434), .ZN(new_n864));
  AOI22_X1  g0664(.A1(new_n862), .A2(G107), .B1(G50), .B2(new_n864), .ZN(new_n865));
  NOR2_X1   g0665(.A1(new_n863), .A2(G190), .ZN(new_n866));
  INV_X1    g0666(.A(new_n866), .ZN(new_n867));
  OAI211_X1 g0667(.A(new_n860), .B(new_n865), .C1(new_n202), .C2(new_n867), .ZN(new_n868));
  OR4_X1    g0668(.A1(new_n841), .A2(new_n848), .A3(new_n857), .A4(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(G311), .ZN(new_n870));
  INV_X1    g0670(.A(G283), .ZN(new_n871));
  OAI221_X1 g0671(.A(new_n269), .B1(new_n837), .B2(new_n870), .C1(new_n871), .C2(new_n861), .ZN(new_n872));
  INV_X1    g0672(.A(new_n856), .ZN(new_n873));
  AOI21_X1  g0673(.A(new_n872), .B1(new_n873), .B2(G322), .ZN(new_n874));
  NAND2_X1  g0674(.A1(new_n859), .A2(new_n635), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n846), .A2(G329), .ZN(new_n876));
  INV_X1    g0676(.A(G303), .ZN(new_n877));
  NOR2_X1   g0677(.A1(new_n850), .A2(new_n877), .ZN(new_n878));
  INV_X1    g0678(.A(KEYINPUT33), .ZN(new_n879));
  NOR2_X1   g0679(.A1(new_n879), .A2(G317), .ZN(new_n880));
  AND2_X1   g0680(.A1(new_n879), .A2(G317), .ZN(new_n881));
  NOR3_X1   g0681(.A1(new_n867), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  AOI211_X1 g0682(.A(new_n878), .B(new_n882), .C1(G326), .C2(new_n864), .ZN(new_n883));
  NAND4_X1  g0683(.A1(new_n874), .A2(new_n875), .A3(new_n876), .A4(new_n883), .ZN(new_n884));
  AOI21_X1  g0684(.A(new_n834), .B1(new_n869), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g0685(.A1(G13), .A2(G33), .ZN(new_n886));
  INV_X1    g0686(.A(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n887), .A2(G20), .ZN(new_n888));
  NOR2_X1   g0688(.A1(new_n888), .A2(new_n833), .ZN(new_n889));
  INV_X1    g0689(.A(new_n889), .ZN(new_n890));
  NOR2_X1   g0690(.A1(new_n251), .A2(new_n273), .ZN(new_n891));
  NOR2_X1   g0691(.A1(new_n775), .A2(new_n258), .ZN(new_n892));
  INV_X1    g0692(.A(new_n892), .ZN(new_n893));
  AOI21_X1  g0693(.A(new_n893), .B1(new_n232), .B2(new_n273), .ZN(new_n894));
  INV_X1    g0694(.A(KEYINPUT101), .ZN(new_n895));
  AOI21_X1  g0695(.A(new_n891), .B1(new_n894), .B2(new_n895), .ZN(new_n896));
  OAI21_X1  g0696(.A(new_n896), .B1(new_n895), .B2(new_n894), .ZN(new_n897));
  NOR2_X1   g0697(.A1(new_n775), .A2(new_n269), .ZN(new_n898));
  AOI22_X1  g0698(.A1(new_n898), .A2(G355), .B1(new_n497), .B2(new_n775), .ZN(new_n899));
  AOI21_X1  g0699(.A(new_n890), .B1(new_n897), .B2(new_n899), .ZN(new_n900));
  NOR3_X1   g0700(.A1(new_n885), .A2(new_n900), .A3(new_n829), .ZN(new_n901));
  INV_X1    g0701(.A(new_n888), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n901), .B1(new_n758), .B2(new_n902), .ZN(new_n903));
  AND2_X1   g0703(.A1(new_n832), .A2(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(new_n904), .ZN(G396));
  NOR2_X1   g0705(.A1(new_n833), .A2(new_n886), .ZN(new_n906));
  AOI21_X1  g0706(.A(new_n829), .B1(new_n332), .B2(new_n906), .ZN(new_n907));
  NOR2_X1   g0707(.A1(new_n861), .A2(new_n202), .ZN(new_n908));
  INV_X1    g0708(.A(new_n850), .ZN(new_n909));
  AOI211_X1 g0709(.A(new_n269), .B(new_n908), .C1(G50), .C2(new_n909), .ZN(new_n910));
  INV_X1    g0710(.A(G132), .ZN(new_n911));
  OAI221_X1 g0711(.A(new_n910), .B1(new_n911), .B2(new_n845), .C1(new_n201), .C2(new_n858), .ZN(new_n912));
  AOI22_X1  g0712(.A1(new_n866), .A2(G150), .B1(new_n864), .B2(G137), .ZN(new_n913));
  INV_X1    g0713(.A(G159), .ZN(new_n914));
  INV_X1    g0714(.A(G143), .ZN(new_n915));
  OAI221_X1 g0715(.A(new_n913), .B1(new_n840), .B2(new_n914), .C1(new_n856), .C2(new_n915), .ZN(new_n916));
  INV_X1    g0716(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g0717(.A(new_n912), .B1(new_n917), .B2(KEYINPUT34), .ZN(new_n918));
  OR2_X1    g0718(.A1(new_n917), .A2(KEYINPUT34), .ZN(new_n919));
  OAI22_X1  g0719(.A1(new_n845), .A2(new_n870), .B1(new_n221), .B2(new_n861), .ZN(new_n920));
  XOR2_X1   g0720(.A(new_n920), .B(KEYINPUT105), .Z(new_n921));
  INV_X1    g0721(.A(new_n864), .ZN(new_n922));
  OAI22_X1  g0722(.A1(new_n922), .A2(new_n877), .B1(new_n850), .B2(new_n455), .ZN(new_n923));
  AOI211_X1 g0723(.A(new_n258), .B(new_n923), .C1(G283), .C2(new_n866), .ZN(new_n924));
  INV_X1    g0724(.A(new_n840), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n925), .A2(G116), .ZN(new_n926));
  NAND2_X1  g0726(.A1(new_n873), .A2(G294), .ZN(new_n927));
  AND4_X1   g0727(.A1(new_n860), .A2(new_n924), .A3(new_n926), .A4(new_n927), .ZN(new_n928));
  AOI22_X1  g0728(.A1(new_n918), .A2(new_n919), .B1(new_n921), .B2(new_n928), .ZN(new_n929));
  NOR2_X1   g0729(.A1(new_n466), .A2(new_n761), .ZN(new_n930));
  OAI22_X1  g0730(.A1(new_n469), .A2(new_n471), .B1(new_n453), .B2(new_n754), .ZN(new_n931));
  AOI21_X1  g0731(.A(new_n930), .B1(new_n931), .B2(new_n466), .ZN(new_n932));
  OAI221_X1 g0732(.A(new_n907), .B1(new_n834), .B2(new_n929), .C1(new_n932), .C2(new_n887), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n931), .A2(new_n466), .ZN(new_n934));
  INV_X1    g0734(.A(new_n930), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n934), .A2(new_n935), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n819), .A2(new_n936), .ZN(new_n937));
  NAND3_X1  g0737(.A1(new_n733), .A2(new_n754), .A3(new_n932), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n798), .A2(new_n800), .ZN(new_n940));
  NAND2_X1  g0740(.A1(new_n940), .A2(G330), .ZN(new_n941));
  AOI21_X1  g0741(.A(new_n830), .B1(new_n939), .B2(new_n941), .ZN(new_n942));
  INV_X1    g0742(.A(new_n942), .ZN(new_n943));
  NOR2_X1   g0743(.A1(new_n939), .A2(new_n941), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n933), .B1(new_n943), .B2(new_n944), .ZN(G384));
  NAND2_X1  g0745(.A1(new_n550), .A2(new_n554), .ZN(new_n946));
  INV_X1    g0746(.A(KEYINPUT35), .ZN(new_n947));
  OAI211_X1 g0747(.A(G116), .B(new_n231), .C1(new_n946), .C2(new_n947), .ZN(new_n948));
  AOI21_X1  g0748(.A(new_n948), .B1(new_n947), .B2(new_n946), .ZN(new_n949));
  XNOR2_X1  g0749(.A(new_n949), .B(KEYINPUT36), .ZN(new_n950));
  NAND3_X1  g0750(.A1(new_n232), .A2(G77), .A3(new_n391), .ZN(new_n951));
  AOI211_X1 g0751(.A(new_n211), .B(G13), .C1(new_n951), .C2(new_n247), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n950), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g0753(.A1(new_n348), .A2(new_n754), .ZN(new_n954));
  INV_X1    g0754(.A(new_n954), .ZN(new_n955));
  NAND2_X1  g0755(.A1(new_n381), .A2(new_n955), .ZN(new_n956));
  OAI21_X1  g0756(.A(new_n954), .B1(new_n376), .B2(new_n380), .ZN(new_n957));
  AOI21_X1  g0757(.A(new_n936), .B1(new_n956), .B2(new_n957), .ZN(new_n958));
  AND2_X1   g0758(.A1(new_n940), .A2(new_n958), .ZN(new_n959));
  INV_X1    g0759(.A(KEYINPUT40), .ZN(new_n960));
  INV_X1    g0760(.A(new_n429), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n741), .A2(new_n753), .ZN(new_n962));
  NAND3_X1  g0762(.A1(new_n961), .A2(new_n962), .A3(new_n437), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n963), .A2(KEYINPUT37), .ZN(new_n964));
  INV_X1    g0764(.A(KEYINPUT37), .ZN(new_n965));
  OAI21_X1  g0765(.A(new_n965), .B1(new_n429), .B2(KEYINPUT106), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n741), .A2(KEYINPUT106), .A3(new_n742), .ZN(new_n967));
  NAND3_X1  g0767(.A1(new_n967), .A2(new_n437), .A3(new_n962), .ZN(new_n968));
  OAI21_X1  g0768(.A(new_n964), .B1(new_n966), .B2(new_n968), .ZN(new_n969));
  NAND2_X1  g0769(.A1(new_n439), .A2(new_n440), .ZN(new_n970));
  AOI21_X1  g0770(.A(new_n970), .B1(new_n744), .B2(new_n745), .ZN(new_n971));
  OAI21_X1  g0771(.A(new_n969), .B1(new_n971), .B2(new_n962), .ZN(new_n972));
  INV_X1    g0772(.A(KEYINPUT38), .ZN(new_n973));
  NAND2_X1  g0773(.A1(new_n972), .A2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n400), .A2(new_n300), .ZN(new_n975));
  NAND2_X1  g0775(.A1(new_n387), .A2(new_n418), .ZN(new_n976));
  OAI211_X1 g0776(.A(new_n976), .B(G68), .C1(new_n397), .C2(new_n387), .ZN(new_n977));
  AOI21_X1  g0777(.A(KEYINPUT16), .B1(new_n977), .B2(new_n393), .ZN(new_n978));
  OAI21_X1  g0778(.A(new_n428), .B1(new_n975), .B2(new_n978), .ZN(new_n979));
  NAND2_X1  g0779(.A1(new_n979), .A2(new_n753), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n979), .A2(new_n742), .ZN(new_n981));
  NAND3_X1  g0781(.A1(new_n980), .A2(new_n981), .A3(new_n437), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n982), .A2(KEYINPUT37), .ZN(new_n983));
  OAI21_X1  g0783(.A(new_n983), .B1(new_n966), .B2(new_n968), .ZN(new_n984));
  INV_X1    g0784(.A(new_n980), .ZN(new_n985));
  NAND2_X1  g0785(.A1(new_n441), .A2(new_n985), .ZN(new_n986));
  NAND3_X1  g0786(.A1(new_n984), .A2(new_n986), .A3(KEYINPUT38), .ZN(new_n987));
  AOI21_X1  g0787(.A(new_n960), .B1(new_n974), .B2(new_n987), .ZN(new_n988));
  AND3_X1   g0788(.A1(new_n967), .A2(new_n437), .A3(new_n962), .ZN(new_n989));
  INV_X1    g0789(.A(new_n966), .ZN(new_n990));
  AOI22_X1  g0790(.A1(new_n989), .A2(new_n990), .B1(KEYINPUT37), .B2(new_n982), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n740), .A2(new_n743), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n980), .B1(new_n992), .B2(new_n736), .ZN(new_n993));
  OAI21_X1  g0793(.A(new_n973), .B1(new_n991), .B2(new_n993), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n994), .A2(new_n987), .ZN(new_n995));
  NAND3_X1  g0795(.A1(new_n995), .A2(new_n940), .A3(new_n958), .ZN(new_n996));
  AOI22_X1  g0796(.A1(new_n959), .A2(new_n988), .B1(new_n996), .B2(new_n960), .ZN(new_n997));
  INV_X1    g0797(.A(new_n997), .ZN(new_n998));
  NAND2_X1  g0798(.A1(new_n701), .A2(new_n940), .ZN(new_n999));
  OAI21_X1  g0799(.A(G330), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n1000), .B1(new_n999), .B2(new_n998), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n818), .A2(new_n701), .A3(new_n821), .ZN(new_n1002));
  NAND2_X1  g0802(.A1(new_n1002), .A2(new_n748), .ZN(new_n1003));
  INV_X1    g0803(.A(new_n348), .ZN(new_n1004));
  AOI21_X1  g0804(.A(new_n281), .B1(new_n365), .B2(new_n366), .ZN(new_n1005));
  AOI22_X1  g0805(.A1(new_n349), .A2(new_n1005), .B1(new_n372), .B2(G179), .ZN(new_n1006));
  AOI21_X1  g0806(.A(new_n374), .B1(new_n1006), .B2(new_n373), .ZN(new_n1007));
  NOR3_X1   g0807(.A1(new_n368), .A2(KEYINPUT75), .A3(new_n370), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1004), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g0809(.A1(new_n1009), .A2(new_n761), .ZN(new_n1010));
  NAND3_X1  g0810(.A1(new_n994), .A2(KEYINPUT39), .A3(new_n987), .ZN(new_n1011));
  AND3_X1   g0811(.A1(new_n984), .A2(new_n986), .A3(KEYINPUT38), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n973), .B2(new_n972), .ZN(new_n1013));
  OAI211_X1 g0813(.A(new_n1010), .B(new_n1011), .C1(new_n1013), .C2(KEYINPUT39), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n746), .A2(new_n753), .ZN(new_n1015));
  AOI21_X1  g0815(.A(new_n955), .B1(new_n1009), .B2(new_n379), .ZN(new_n1016));
  NOR3_X1   g0816(.A1(new_n376), .A2(new_n380), .A3(new_n954), .ZN(new_n1017));
  NOR2_X1   g0817(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n1018), .B1(new_n938), .B2(new_n935), .ZN(new_n1019));
  AOI21_X1  g0819(.A(new_n1015), .B1(new_n1019), .B2(new_n995), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1014), .A2(new_n1020), .ZN(new_n1021));
  XOR2_X1   g0821(.A(new_n1003), .B(new_n1021), .Z(new_n1022));
  OAI22_X1  g0822(.A1(new_n1001), .A2(new_n1022), .B1(new_n211), .B2(new_n824), .ZN(new_n1023));
  AND2_X1   g0823(.A1(new_n1001), .A2(new_n1022), .ZN(new_n1024));
  OAI21_X1  g0824(.A(new_n953), .B1(new_n1023), .B2(new_n1024), .ZN(G367));
  NAND2_X1  g0825(.A1(new_n563), .A2(new_n761), .ZN(new_n1026));
  OAI211_X1 g0826(.A(new_n586), .B(new_n1026), .C1(new_n598), .C2(new_n604), .ZN(new_n1027));
  NAND2_X1  g0827(.A1(new_n709), .A2(new_n761), .ZN(new_n1028));
  AND3_X1   g0828(.A1(new_n1027), .A2(KEYINPUT107), .A3(new_n1028), .ZN(new_n1029));
  AOI21_X1  g0829(.A(KEYINPUT107), .B1(new_n1027), .B2(new_n1028), .ZN(new_n1030));
  OAI21_X1  g0830(.A(new_n703), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(new_n586), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1032), .A2(new_n754), .ZN(new_n1033));
  NAND2_X1  g0833(.A1(new_n1027), .A2(new_n1028), .ZN(new_n1034));
  INV_X1    g0834(.A(new_n1034), .ZN(new_n1035));
  NOR2_X1   g0835(.A1(new_n1035), .A2(new_n767), .ZN(new_n1036));
  INV_X1    g0836(.A(KEYINPUT42), .ZN(new_n1037));
  NOR2_X1   g0837(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1038));
  INV_X1    g0838(.A(new_n1038), .ZN(new_n1039));
  NAND3_X1  g0839(.A1(new_n1033), .A2(KEYINPUT108), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g0840(.A(KEYINPUT108), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n761), .B1(new_n1031), .B2(new_n586), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n1041), .B1(new_n1042), .B2(new_n1038), .ZN(new_n1043));
  NAND2_X1  g0843(.A1(new_n1036), .A2(new_n1037), .ZN(new_n1044));
  NAND3_X1  g0844(.A1(new_n1040), .A2(new_n1043), .A3(new_n1044), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n697), .A2(new_n754), .ZN(new_n1046));
  OR2_X1    g0846(.A1(new_n720), .A2(new_n1046), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n726), .A2(new_n1046), .ZN(new_n1048));
  NAND2_X1  g0848(.A1(new_n1047), .A2(new_n1048), .ZN(new_n1049));
  INV_X1    g0849(.A(new_n1049), .ZN(new_n1050));
  INV_X1    g0850(.A(KEYINPUT43), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1050), .A2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n1049), .A2(KEYINPUT43), .ZN(new_n1053));
  NAND3_X1  g0853(.A1(new_n1045), .A2(new_n1052), .A3(new_n1053), .ZN(new_n1054));
  AOI21_X1  g0854(.A(new_n1038), .B1(new_n1032), .B2(new_n754), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1055), .A2(KEYINPUT108), .B1(new_n1037), .B2(new_n1036), .ZN(new_n1056));
  NAND4_X1  g0856(.A1(new_n1056), .A2(new_n1051), .A3(new_n1050), .A4(new_n1043), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  OR2_X1    g0858(.A1(new_n1029), .A2(new_n1030), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n765), .A2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1061));
  NAND4_X1  g0861(.A1(new_n1054), .A2(new_n1057), .A3(new_n765), .A4(new_n1059), .ZN(new_n1062));
  XOR2_X1   g0862(.A(new_n776), .B(KEYINPUT41), .Z(new_n1063));
  OAI21_X1  g0863(.A(new_n1034), .B1(new_n771), .B2(new_n769), .ZN(new_n1064));
  INV_X1    g0864(.A(KEYINPUT45), .ZN(new_n1065));
  XNOR2_X1  g0865(.A(new_n1064), .B(new_n1065), .ZN(new_n1066));
  INV_X1    g0866(.A(new_n769), .ZN(new_n1067));
  NAND3_X1  g0867(.A1(new_n1067), .A2(new_n770), .A3(new_n1035), .ZN(new_n1068));
  INV_X1    g0868(.A(KEYINPUT44), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n1068), .A2(new_n1069), .ZN(new_n1070));
  NAND4_X1  g0870(.A1(new_n1067), .A2(KEYINPUT44), .A3(new_n1035), .A4(new_n770), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n766), .A2(new_n1066), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g0873(.A1(new_n1066), .A2(new_n1072), .ZN(new_n1074));
  NAND2_X1  g0874(.A1(new_n1074), .A2(new_n765), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n540), .A2(new_n754), .ZN(new_n1076));
  INV_X1    g0876(.A(new_n1076), .ZN(new_n1077));
  OAI21_X1  g0877(.A(new_n767), .B1(new_n763), .B2(new_n1077), .ZN(new_n1078));
  NAND3_X1  g0878(.A1(new_n758), .A2(G330), .A3(new_n1078), .ZN(new_n1079));
  INV_X1    g0879(.A(new_n1079), .ZN(new_n1080));
  AOI21_X1  g0880(.A(new_n1078), .B1(new_n758), .B2(G330), .ZN(new_n1081));
  NOR2_X1   g0881(.A1(new_n1080), .A2(new_n1081), .ZN(new_n1082));
  INV_X1    g0882(.A(new_n1082), .ZN(new_n1083));
  NAND4_X1  g0883(.A1(new_n1073), .A2(new_n1075), .A3(new_n1083), .A4(new_n822), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n1063), .B1(new_n1084), .B2(new_n822), .ZN(new_n1085));
  XOR2_X1   g0885(.A(new_n826), .B(KEYINPUT109), .Z(new_n1086));
  OAI211_X1 g0886(.A(new_n1061), .B(new_n1062), .C1(new_n1085), .C2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n892), .A2(new_n242), .ZN(new_n1088));
  AOI21_X1  g0888(.A(new_n890), .B1(new_n775), .B2(new_n447), .ZN(new_n1089));
  AOI21_X1  g0889(.A(new_n829), .B1(new_n1088), .B2(new_n1089), .ZN(new_n1090));
  OAI221_X1 g0890(.A(new_n258), .B1(new_n915), .B2(new_n922), .C1(new_n856), .C2(new_n284), .ZN(new_n1091));
  NOR2_X1   g0891(.A1(new_n858), .A2(new_n202), .ZN(new_n1092));
  INV_X1    g0892(.A(G137), .ZN(new_n1093));
  OAI22_X1  g0893(.A1(new_n845), .A2(new_n1093), .B1(new_n840), .B2(new_n207), .ZN(new_n1094));
  NOR2_X1   g0894(.A1(new_n861), .A2(new_n332), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n850), .A2(new_n201), .ZN(new_n1096));
  NOR2_X1   g0896(.A1(new_n1095), .A2(new_n1096), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1097), .B1(new_n914), .B2(new_n867), .ZN(new_n1098));
  OR4_X1    g0898(.A1(new_n1091), .A2(new_n1092), .A3(new_n1094), .A4(new_n1098), .ZN(new_n1099));
  OAI21_X1  g0899(.A(new_n269), .B1(new_n861), .B2(new_n500), .ZN(new_n1100));
  XOR2_X1   g0900(.A(KEYINPUT110), .B(G317), .Z(new_n1101));
  AOI21_X1  g0901(.A(new_n1100), .B1(new_n846), .B2(new_n1101), .ZN(new_n1102));
  XOR2_X1   g0902(.A(new_n1102), .B(KEYINPUT111), .Z(new_n1103));
  INV_X1    g0903(.A(KEYINPUT46), .ZN(new_n1104));
  OAI21_X1  g0904(.A(new_n1104), .B1(new_n850), .B2(new_n497), .ZN(new_n1105));
  OAI221_X1 g0905(.A(new_n1105), .B1(new_n922), .B2(new_n870), .C1(new_n658), .C2(new_n867), .ZN(new_n1106));
  AOI21_X1  g0906(.A(new_n1106), .B1(new_n859), .B2(G107), .ZN(new_n1107));
  AOI22_X1  g0907(.A1(new_n873), .A2(G303), .B1(new_n925), .B2(G283), .ZN(new_n1108));
  NAND2_X1  g0908(.A1(new_n909), .A2(G116), .ZN(new_n1109));
  OAI211_X1 g0909(.A(new_n1107), .B(new_n1108), .C1(new_n1104), .C2(new_n1109), .ZN(new_n1110));
  OAI21_X1  g0910(.A(new_n1099), .B1(new_n1103), .B2(new_n1110), .ZN(new_n1111));
  XOR2_X1   g0911(.A(new_n1111), .B(KEYINPUT47), .Z(new_n1112));
  OAI221_X1 g0912(.A(new_n1090), .B1(new_n902), .B2(new_n1049), .C1(new_n1112), .C2(new_n834), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1087), .A2(new_n1113), .ZN(G387));
  INV_X1    g0914(.A(KEYINPUT114), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n1115), .B1(new_n1083), .B2(new_n822), .ZN(new_n1116));
  AND2_X1   g0916(.A1(new_n818), .A2(new_n821), .ZN(new_n1117));
  OAI211_X1 g0917(.A(new_n1082), .B(KEYINPUT114), .C1(new_n1117), .C2(new_n801), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1083), .A2(new_n822), .ZN(new_n1119));
  NAND4_X1  g0919(.A1(new_n1116), .A2(new_n1118), .A3(new_n776), .A4(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n764), .A2(new_n888), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n774), .A2(new_n898), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1122), .B1(G107), .B2(new_n215), .ZN(new_n1123));
  OR2_X1    g0923(.A1(new_n774), .A2(KEYINPUT112), .ZN(new_n1124));
  NAND2_X1  g0924(.A1(new_n774), .A2(KEYINPUT112), .ZN(new_n1125));
  NAND2_X1  g0925(.A1(new_n443), .A2(new_n207), .ZN(new_n1126));
  OR2_X1    g0926(.A1(new_n1126), .A2(KEYINPUT50), .ZN(new_n1127));
  OAI21_X1  g0927(.A(new_n273), .B1(new_n202), .B2(new_n332), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1128), .B1(new_n1126), .B2(KEYINPUT50), .ZN(new_n1129));
  NAND4_X1  g0929(.A1(new_n1124), .A2(new_n1125), .A3(new_n1127), .A4(new_n1129), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n893), .B1(new_n239), .B2(G45), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1123), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n830), .B1(new_n1132), .B2(new_n890), .ZN(new_n1133));
  OAI22_X1  g0933(.A1(new_n845), .A2(new_n284), .B1(new_n332), .B2(new_n850), .ZN(new_n1134));
  XNOR2_X1  g0934(.A(new_n1134), .B(KEYINPUT113), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n859), .A2(new_n447), .ZN(new_n1136));
  OAI221_X1 g0936(.A(new_n258), .B1(new_n837), .B2(new_n202), .C1(new_n500), .C2(new_n861), .ZN(new_n1137));
  AOI21_X1  g0937(.A(new_n1137), .B1(G159), .B2(new_n864), .ZN(new_n1138));
  AOI22_X1  g0938(.A1(new_n873), .A2(G50), .B1(new_n382), .B2(new_n866), .ZN(new_n1139));
  NAND4_X1  g0939(.A1(new_n1135), .A2(new_n1136), .A3(new_n1138), .A4(new_n1139), .ZN(new_n1140));
  NAND2_X1  g0940(.A1(new_n846), .A2(G326), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n258), .B1(new_n862), .B2(G116), .ZN(new_n1142));
  OAI22_X1  g0942(.A1(new_n858), .A2(new_n871), .B1(new_n658), .B2(new_n850), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n873), .A2(new_n1101), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n866), .A2(G311), .B1(new_n864), .B2(G322), .ZN(new_n1145));
  OAI211_X1 g0945(.A(new_n1144), .B(new_n1145), .C1(new_n877), .C2(new_n840), .ZN(new_n1146));
  INV_X1    g0946(.A(KEYINPUT48), .ZN(new_n1147));
  AOI21_X1  g0947(.A(new_n1143), .B1(new_n1146), .B2(new_n1147), .ZN(new_n1148));
  OAI21_X1  g0948(.A(new_n1148), .B1(new_n1147), .B2(new_n1146), .ZN(new_n1149));
  INV_X1    g0949(.A(KEYINPUT49), .ZN(new_n1150));
  OAI211_X1 g0950(.A(new_n1141), .B(new_n1142), .C1(new_n1149), .C2(new_n1150), .ZN(new_n1151));
  AND2_X1   g0951(.A1(new_n1149), .A2(new_n1150), .ZN(new_n1152));
  OAI21_X1  g0952(.A(new_n1140), .B1(new_n1151), .B2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1133), .B1(new_n1153), .B2(new_n833), .ZN(new_n1154));
  AOI22_X1  g0954(.A1(new_n1083), .A2(new_n1086), .B1(new_n1121), .B2(new_n1154), .ZN(new_n1155));
  NAND2_X1  g0955(.A1(new_n1120), .A2(new_n1155), .ZN(G393));
  INV_X1    g0956(.A(new_n1086), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1073), .A2(new_n1075), .A3(KEYINPUT115), .ZN(new_n1158));
  OR3_X1    g0958(.A1(new_n1074), .A2(KEYINPUT115), .A3(new_n765), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1158), .A2(new_n1159), .ZN(new_n1160));
  INV_X1    g0960(.A(KEYINPUT116), .ZN(new_n1161));
  AOI21_X1  g0961(.A(new_n1157), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  OAI21_X1  g0962(.A(new_n1162), .B1(new_n1161), .B2(new_n1160), .ZN(new_n1163));
  NOR2_X1   g0963(.A1(new_n1059), .A2(new_n902), .ZN(new_n1164));
  AOI22_X1  g0964(.A1(new_n873), .A2(G311), .B1(G317), .B2(new_n864), .ZN(new_n1165));
  XOR2_X1   g0965(.A(new_n1165), .B(KEYINPUT52), .Z(new_n1166));
  OAI221_X1 g0966(.A(new_n269), .B1(new_n861), .B2(new_n455), .C1(new_n871), .C2(new_n850), .ZN(new_n1167));
  AOI21_X1  g0967(.A(new_n1167), .B1(new_n846), .B2(G322), .ZN(new_n1168));
  XOR2_X1   g0968(.A(new_n1168), .B(KEYINPUT119), .Z(new_n1169));
  OAI22_X1  g0969(.A1(new_n867), .A2(new_n877), .B1(new_n837), .B2(new_n631), .ZN(new_n1170));
  AOI21_X1  g0970(.A(new_n1170), .B1(new_n859), .B2(G116), .ZN(new_n1171));
  NAND3_X1  g0971(.A1(new_n1166), .A2(new_n1169), .A3(new_n1171), .ZN(new_n1172));
  AOI22_X1  g0972(.A1(new_n925), .A2(new_n443), .B1(G50), .B2(new_n866), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT118), .ZN(new_n1174));
  OAI22_X1  g0974(.A1(new_n856), .A2(new_n914), .B1(new_n284), .B2(new_n922), .ZN(new_n1175));
  XNOR2_X1  g0975(.A(new_n1175), .B(KEYINPUT51), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n269), .B1(new_n862), .B2(G87), .ZN(new_n1177));
  OAI221_X1 g0977(.A(new_n1177), .B1(new_n202), .B2(new_n850), .C1(new_n845), .C2(new_n915), .ZN(new_n1178));
  AOI21_X1  g0978(.A(new_n1178), .B1(G77), .B2(new_n859), .ZN(new_n1179));
  NAND3_X1  g0979(.A1(new_n1174), .A2(new_n1176), .A3(new_n1179), .ZN(new_n1180));
  AOI21_X1  g0980(.A(new_n834), .B1(new_n1172), .B2(new_n1180), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n889), .B1(new_n500), .B2(new_n215), .C1(new_n893), .C2(new_n246), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n830), .A2(new_n1182), .ZN(new_n1183));
  XOR2_X1   g0983(.A(new_n1183), .B(KEYINPUT117), .Z(new_n1184));
  NOR3_X1   g0984(.A1(new_n1164), .A2(new_n1181), .A3(new_n1184), .ZN(new_n1185));
  AND2_X1   g0985(.A1(new_n1084), .A2(new_n776), .ZN(new_n1186));
  NAND3_X1  g0986(.A1(new_n1158), .A2(new_n1159), .A3(new_n1119), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n1185), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g0988(.A1(new_n1163), .A2(new_n1188), .ZN(G390));
  OAI21_X1  g0989(.A(new_n1018), .B1(new_n941), .B2(new_n936), .ZN(new_n1190));
  OAI211_X1 g0990(.A(new_n801), .B(new_n932), .C1(new_n1017), .C2(new_n1016), .ZN(new_n1191));
  NAND2_X1  g0991(.A1(new_n1190), .A2(new_n1191), .ZN(new_n1192));
  NAND2_X1  g0992(.A1(new_n938), .A2(new_n935), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n1192), .A2(new_n1193), .ZN(new_n1194));
  NAND2_X1  g0994(.A1(new_n815), .A2(new_n754), .ZN(new_n1195));
  INV_X1    g0995(.A(KEYINPUT99), .ZN(new_n1196));
  NAND2_X1  g0996(.A1(new_n1195), .A2(new_n1196), .ZN(new_n1197));
  NAND3_X1  g0997(.A1(new_n815), .A2(KEYINPUT99), .A3(new_n754), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1197), .A2(new_n1198), .A3(new_n935), .ZN(new_n1199));
  NAND2_X1  g0999(.A1(new_n1199), .A2(new_n934), .ZN(new_n1200));
  NAND3_X1  g1000(.A1(new_n1200), .A2(new_n1191), .A3(new_n1190), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1194), .A2(new_n1201), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n701), .A2(new_n801), .ZN(new_n1203));
  NAND3_X1  g1003(.A1(new_n1002), .A2(new_n748), .A3(new_n1203), .ZN(new_n1204));
  INV_X1    g1004(.A(new_n1204), .ZN(new_n1205));
  NAND2_X1  g1005(.A1(new_n1202), .A2(new_n1205), .ZN(new_n1206));
  NOR2_X1   g1006(.A1(new_n1013), .A2(new_n1010), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1200), .B2(new_n1018), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1011), .B1(new_n1013), .B2(KEYINPUT39), .ZN(new_n1209));
  OAI21_X1  g1009(.A(new_n1209), .B1(new_n1010), .B2(new_n1019), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1208), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(KEYINPUT120), .ZN(new_n1212));
  NOR2_X1   g1012(.A1(new_n1191), .A2(new_n1212), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1211), .A2(new_n1214), .ZN(new_n1215));
  NAND3_X1  g1015(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1216));
  NAND3_X1  g1016(.A1(new_n1206), .A2(new_n1215), .A3(new_n1216), .ZN(new_n1217));
  AOI21_X1  g1017(.A(new_n1204), .B1(new_n1194), .B2(new_n1201), .ZN(new_n1218));
  AND3_X1   g1018(.A1(new_n1208), .A2(new_n1210), .A3(new_n1213), .ZN(new_n1219));
  AOI21_X1  g1019(.A(new_n1213), .B1(new_n1208), .B2(new_n1210), .ZN(new_n1220));
  OAI21_X1  g1020(.A(new_n1218), .B1(new_n1219), .B2(new_n1220), .ZN(new_n1221));
  NAND3_X1  g1021(.A1(new_n1217), .A2(new_n1221), .A3(new_n776), .ZN(new_n1222));
  NAND2_X1  g1022(.A1(new_n1215), .A2(new_n1216), .ZN(new_n1223));
  NAND2_X1  g1023(.A1(new_n1223), .A2(new_n1086), .ZN(new_n1224));
  INV_X1    g1024(.A(new_n906), .ZN(new_n1225));
  OAI21_X1  g1025(.A(new_n830), .B1(new_n382), .B2(new_n1225), .ZN(new_n1226));
  OAI22_X1  g1026(.A1(new_n858), .A2(new_n332), .B1(new_n856), .B2(new_n497), .ZN(new_n1227));
  XOR2_X1   g1027(.A(new_n1227), .B(KEYINPUT121), .Z(new_n1228));
  OAI21_X1  g1028(.A(new_n269), .B1(new_n850), .B2(new_n221), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1229), .B1(new_n925), .B2(G97), .ZN(new_n1230));
  NOR2_X1   g1030(.A1(new_n922), .A2(new_n871), .ZN(new_n1231));
  AOI211_X1 g1031(.A(new_n908), .B(new_n1231), .C1(G107), .C2(new_n866), .ZN(new_n1232));
  OAI211_X1 g1032(.A(new_n1230), .B(new_n1232), .C1(new_n631), .C2(new_n845), .ZN(new_n1233));
  OR3_X1    g1033(.A1(new_n850), .A2(KEYINPUT53), .A3(new_n284), .ZN(new_n1234));
  OAI21_X1  g1034(.A(KEYINPUT53), .B1(new_n850), .B2(new_n284), .ZN(new_n1235));
  INV_X1    g1035(.A(G125), .ZN(new_n1236));
  OAI211_X1 g1036(.A(new_n1234), .B(new_n1235), .C1(new_n845), .C2(new_n1236), .ZN(new_n1237));
  XNOR2_X1  g1037(.A(KEYINPUT54), .B(G143), .ZN(new_n1238));
  INV_X1    g1038(.A(new_n1238), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n873), .A2(G132), .B1(new_n925), .B2(new_n1239), .ZN(new_n1240));
  INV_X1    g1040(.A(G128), .ZN(new_n1241));
  OAI22_X1  g1041(.A1(new_n922), .A2(new_n1241), .B1(new_n861), .B2(new_n207), .ZN(new_n1242));
  AOI211_X1 g1042(.A(new_n269), .B(new_n1242), .C1(G137), .C2(new_n866), .ZN(new_n1243));
  OAI211_X1 g1043(.A(new_n1240), .B(new_n1243), .C1(new_n914), .C2(new_n858), .ZN(new_n1244));
  OAI22_X1  g1044(.A1(new_n1228), .A2(new_n1233), .B1(new_n1237), .B2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(new_n1226), .B1(new_n1245), .B2(new_n833), .ZN(new_n1246));
  INV_X1    g1046(.A(new_n1209), .ZN(new_n1247));
  OAI21_X1  g1047(.A(new_n1246), .B1(new_n1247), .B2(new_n887), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1222), .A2(new_n1224), .A3(new_n1248), .ZN(G378));
  AOI21_X1  g1049(.A(new_n1204), .B1(new_n1223), .B2(new_n1202), .ZN(new_n1250));
  AOI22_X1  g1050(.A1(new_n989), .A2(new_n990), .B1(new_n963), .B2(KEYINPUT37), .ZN(new_n1251));
  NOR3_X1   g1051(.A1(new_n740), .A2(new_n743), .A3(new_n739), .ZN(new_n1252));
  AOI21_X1  g1052(.A(KEYINPUT93), .B1(new_n415), .B2(new_n431), .ZN(new_n1253));
  OAI21_X1  g1053(.A(new_n736), .B1(new_n1252), .B2(new_n1253), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n962), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1251), .B1(new_n1254), .B2(new_n1255), .ZN(new_n1256));
  OAI21_X1  g1056(.A(new_n987), .B1(new_n1256), .B2(KEYINPUT38), .ZN(new_n1257));
  NAND4_X1  g1057(.A1(new_n1257), .A2(KEYINPUT40), .A3(new_n940), .A4(new_n958), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n996), .A2(new_n960), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1258), .A2(new_n1259), .A3(G330), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1260), .A2(new_n1014), .A3(new_n1020), .ZN(new_n1261));
  NAND3_X1  g1061(.A1(new_n1021), .A2(G330), .A3(new_n997), .ZN(new_n1262));
  INV_X1    g1062(.A(new_n314), .ZN(new_n1263));
  NAND2_X1  g1063(.A1(new_n735), .A2(new_n1263), .ZN(new_n1264));
  NOR2_X1   g1064(.A1(new_n315), .A2(new_n752), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  OAI21_X1  g1066(.A(new_n329), .B1(new_n315), .B2(new_n752), .ZN(new_n1267));
  XNOR2_X1  g1067(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1268));
  AND3_X1   g1068(.A1(new_n1266), .A2(new_n1267), .A3(new_n1268), .ZN(new_n1269));
  AOI21_X1  g1069(.A(new_n1268), .B1(new_n1266), .B2(new_n1267), .ZN(new_n1270));
  NOR2_X1   g1070(.A1(new_n1269), .A2(new_n1270), .ZN(new_n1271));
  NAND3_X1  g1071(.A1(new_n1261), .A2(new_n1262), .A3(new_n1271), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  AOI21_X1  g1073(.A(new_n1271), .B1(new_n1261), .B2(new_n1262), .ZN(new_n1274));
  OAI21_X1  g1074(.A(KEYINPUT57), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1275));
  OAI21_X1  g1075(.A(new_n776), .B1(new_n1250), .B2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1221), .A2(new_n1205), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1271), .ZN(new_n1279));
  NAND2_X1  g1079(.A1(new_n1278), .A2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1272), .ZN(new_n1281));
  AOI21_X1  g1081(.A(KEYINPUT57), .B1(new_n1277), .B2(new_n1281), .ZN(new_n1282));
  OR2_X1    g1082(.A1(new_n1276), .A2(new_n1282), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1157), .B1(new_n1280), .B2(new_n1272), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1279), .A2(new_n887), .ZN(new_n1285));
  OAI22_X1  g1085(.A1(new_n922), .A2(new_n1236), .B1(new_n837), .B2(new_n1093), .ZN(new_n1286));
  OAI22_X1  g1086(.A1(new_n867), .A2(new_n911), .B1(new_n850), .B2(new_n1238), .ZN(new_n1287));
  AOI211_X1 g1087(.A(new_n1286), .B(new_n1287), .C1(new_n873), .C2(G128), .ZN(new_n1288));
  OAI21_X1  g1088(.A(new_n1288), .B1(new_n284), .B2(new_n858), .ZN(new_n1289));
  OR2_X1    g1089(.A1(new_n1289), .A2(KEYINPUT59), .ZN(new_n1290));
  NAND2_X1  g1090(.A1(new_n1289), .A2(KEYINPUT59), .ZN(new_n1291));
  OAI211_X1 g1091(.A(new_n614), .B(new_n272), .C1(new_n861), .C2(new_n914), .ZN(new_n1292));
  AOI21_X1  g1092(.A(new_n1292), .B1(new_n846), .B2(G124), .ZN(new_n1293));
  NAND3_X1  g1093(.A1(new_n1290), .A2(new_n1291), .A3(new_n1293), .ZN(new_n1294));
  NOR2_X1   g1094(.A1(new_n258), .A2(G41), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1295), .B1(new_n446), .B2(new_n837), .ZN(new_n1296));
  AOI21_X1  g1096(.A(new_n1296), .B1(G77), .B2(new_n909), .ZN(new_n1297));
  OAI221_X1 g1097(.A(new_n1297), .B1(new_n455), .B2(new_n856), .C1(new_n871), .C2(new_n845), .ZN(new_n1298));
  NOR2_X1   g1098(.A1(new_n861), .A2(new_n201), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1299), .B1(G116), .B2(new_n864), .ZN(new_n1300));
  OAI21_X1  g1100(.A(new_n1300), .B1(new_n500), .B2(new_n867), .ZN(new_n1301));
  NOR3_X1   g1101(.A1(new_n1298), .A2(new_n1092), .A3(new_n1301), .ZN(new_n1302));
  NAND2_X1  g1102(.A1(new_n1302), .A2(KEYINPUT58), .ZN(new_n1303));
  OR2_X1    g1103(.A1(new_n1302), .A2(KEYINPUT58), .ZN(new_n1304));
  INV_X1    g1104(.A(new_n1295), .ZN(new_n1305));
  OAI211_X1 g1105(.A(new_n1305), .B(new_n207), .C1(G33), .C2(G41), .ZN(new_n1306));
  AND4_X1   g1106(.A1(new_n1294), .A2(new_n1303), .A3(new_n1304), .A4(new_n1306), .ZN(new_n1307));
  OAI221_X1 g1107(.A(new_n830), .B1(G50), .B2(new_n1225), .C1(new_n1307), .C2(new_n834), .ZN(new_n1308));
  NOR2_X1   g1108(.A1(new_n1285), .A2(new_n1308), .ZN(new_n1309));
  NOR2_X1   g1109(.A1(new_n1284), .A2(new_n1309), .ZN(new_n1310));
  NAND2_X1  g1110(.A1(new_n1283), .A2(new_n1310), .ZN(G375));
  INV_X1    g1111(.A(new_n1063), .ZN(new_n1312));
  NAND3_X1  g1112(.A1(new_n1194), .A2(new_n1204), .A3(new_n1201), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1206), .A2(new_n1312), .A3(new_n1313), .ZN(new_n1314));
  NAND2_X1  g1114(.A1(new_n1018), .A2(new_n886), .ZN(new_n1315));
  OAI21_X1  g1115(.A(new_n830), .B1(G68), .B2(new_n1225), .ZN(new_n1316));
  AOI211_X1 g1116(.A(new_n258), .B(new_n1095), .C1(new_n925), .C2(G107), .ZN(new_n1317));
  OAI221_X1 g1117(.A(new_n1317), .B1(new_n871), .B2(new_n856), .C1(new_n877), .C2(new_n845), .ZN(new_n1318));
  AOI22_X1  g1118(.A1(new_n866), .A2(G116), .B1(new_n864), .B2(G294), .ZN(new_n1319));
  OAI211_X1 g1119(.A(new_n1136), .B(new_n1319), .C1(new_n500), .C2(new_n850), .ZN(new_n1320));
  OAI21_X1  g1120(.A(new_n258), .B1(new_n837), .B2(new_n284), .ZN(new_n1321));
  AOI211_X1 g1121(.A(new_n1299), .B(new_n1321), .C1(new_n846), .C2(G128), .ZN(new_n1322));
  OAI21_X1  g1122(.A(new_n1322), .B1(new_n1093), .B2(new_n856), .ZN(new_n1323));
  AOI22_X1  g1123(.A1(new_n909), .A2(G159), .B1(new_n1239), .B2(new_n866), .ZN(new_n1324));
  OAI221_X1 g1124(.A(new_n1324), .B1(new_n911), .B2(new_n922), .C1(new_n858), .C2(new_n207), .ZN(new_n1325));
  OAI22_X1  g1125(.A1(new_n1318), .A2(new_n1320), .B1(new_n1323), .B2(new_n1325), .ZN(new_n1326));
  AOI21_X1  g1126(.A(new_n1316), .B1(new_n1326), .B2(new_n833), .ZN(new_n1327));
  AOI22_X1  g1127(.A1(new_n1202), .A2(new_n1086), .B1(new_n1315), .B2(new_n1327), .ZN(new_n1328));
  NAND2_X1  g1128(.A1(new_n1314), .A2(new_n1328), .ZN(G381));
  INV_X1    g1129(.A(G375), .ZN(new_n1330));
  INV_X1    g1130(.A(G378), .ZN(new_n1331));
  AND3_X1   g1131(.A1(new_n1120), .A2(new_n904), .A3(new_n1155), .ZN(new_n1332));
  NAND3_X1  g1132(.A1(new_n1332), .A2(new_n1328), .A3(new_n1314), .ZN(new_n1333));
  NOR4_X1   g1133(.A1(G390), .A2(new_n1333), .A3(G387), .A4(G384), .ZN(new_n1334));
  NAND3_X1  g1134(.A1(new_n1330), .A2(new_n1331), .A3(new_n1334), .ZN(G407));
  INV_X1    g1135(.A(G343), .ZN(new_n1336));
  NAND2_X1  g1136(.A1(new_n1336), .A2(G213), .ZN(new_n1337));
  INV_X1    g1137(.A(new_n1337), .ZN(new_n1338));
  NAND3_X1  g1138(.A1(new_n1330), .A2(new_n1331), .A3(new_n1338), .ZN(new_n1339));
  NAND3_X1  g1139(.A1(G407), .A2(new_n1339), .A3(G213), .ZN(new_n1340));
  XOR2_X1   g1140(.A(new_n1340), .B(KEYINPUT122), .Z(G409));
  AOI21_X1  g1141(.A(new_n904), .B1(new_n1120), .B2(new_n1155), .ZN(new_n1342));
  NOR2_X1   g1142(.A1(new_n1332), .A2(new_n1342), .ZN(new_n1343));
  NAND2_X1  g1143(.A1(G387), .A2(new_n1343), .ZN(new_n1344));
  OAI211_X1 g1144(.A(new_n1087), .B(new_n1113), .C1(new_n1332), .C2(new_n1342), .ZN(new_n1345));
  NAND2_X1  g1145(.A1(new_n1344), .A2(new_n1345), .ZN(new_n1346));
  NAND2_X1  g1146(.A1(new_n1346), .A2(G390), .ZN(new_n1347));
  NAND4_X1  g1147(.A1(new_n1344), .A2(new_n1163), .A3(new_n1188), .A4(new_n1345), .ZN(new_n1348));
  NAND2_X1  g1148(.A1(new_n1347), .A2(new_n1348), .ZN(new_n1349));
  OAI21_X1  g1149(.A(KEYINPUT123), .B1(new_n1284), .B2(new_n1309), .ZN(new_n1350));
  OAI21_X1  g1150(.A(new_n1086), .B1(new_n1273), .B2(new_n1274), .ZN(new_n1351));
  INV_X1    g1151(.A(new_n1309), .ZN(new_n1352));
  INV_X1    g1152(.A(KEYINPUT123), .ZN(new_n1353));
  NAND3_X1  g1153(.A1(new_n1351), .A2(new_n1352), .A3(new_n1353), .ZN(new_n1354));
  NAND3_X1  g1154(.A1(new_n1277), .A2(new_n1312), .A3(new_n1281), .ZN(new_n1355));
  NAND3_X1  g1155(.A1(new_n1350), .A2(new_n1354), .A3(new_n1355), .ZN(new_n1356));
  NAND2_X1  g1156(.A1(new_n1356), .A2(new_n1331), .ZN(new_n1357));
  OAI211_X1 g1157(.A(G378), .B(new_n1310), .C1(new_n1276), .C2(new_n1282), .ZN(new_n1358));
  NAND2_X1  g1158(.A1(new_n1357), .A2(new_n1358), .ZN(new_n1359));
  NAND2_X1  g1159(.A1(new_n1206), .A2(KEYINPUT60), .ZN(new_n1360));
  NAND2_X1  g1160(.A1(new_n1360), .A2(new_n1313), .ZN(new_n1361));
  NAND4_X1  g1161(.A1(new_n1194), .A2(new_n1204), .A3(KEYINPUT60), .A4(new_n1201), .ZN(new_n1362));
  NAND2_X1  g1162(.A1(new_n1362), .A2(new_n776), .ZN(new_n1363));
  INV_X1    g1163(.A(new_n1363), .ZN(new_n1364));
  NAND2_X1  g1164(.A1(new_n1361), .A2(new_n1364), .ZN(new_n1365));
  AOI21_X1  g1165(.A(G384), .B1(new_n1365), .B2(new_n1328), .ZN(new_n1366));
  AOI21_X1  g1166(.A(new_n1363), .B1(new_n1360), .B2(new_n1313), .ZN(new_n1367));
  INV_X1    g1167(.A(G384), .ZN(new_n1368));
  INV_X1    g1168(.A(new_n1328), .ZN(new_n1369));
  NOR3_X1   g1169(.A1(new_n1367), .A2(new_n1368), .A3(new_n1369), .ZN(new_n1370));
  NOR2_X1   g1170(.A1(new_n1366), .A2(new_n1370), .ZN(new_n1371));
  NAND3_X1  g1171(.A1(new_n1359), .A2(new_n1337), .A3(new_n1371), .ZN(new_n1372));
  INV_X1    g1172(.A(KEYINPUT62), .ZN(new_n1373));
  NAND2_X1  g1173(.A1(new_n1372), .A2(new_n1373), .ZN(new_n1374));
  AOI21_X1  g1174(.A(new_n1338), .B1(new_n1357), .B2(new_n1358), .ZN(new_n1375));
  NAND3_X1  g1175(.A1(new_n1375), .A2(KEYINPUT62), .A3(new_n1371), .ZN(new_n1376));
  AND3_X1   g1176(.A1(new_n1374), .A2(KEYINPUT125), .A3(new_n1376), .ZN(new_n1377));
  INV_X1    g1177(.A(KEYINPUT125), .ZN(new_n1378));
  NAND3_X1  g1178(.A1(new_n1372), .A2(new_n1378), .A3(new_n1373), .ZN(new_n1379));
  INV_X1    g1179(.A(KEYINPUT61), .ZN(new_n1380));
  NAND2_X1  g1180(.A1(new_n1359), .A2(new_n1337), .ZN(new_n1381));
  NAND2_X1  g1181(.A1(new_n1338), .A2(G2897), .ZN(new_n1382));
  INV_X1    g1182(.A(new_n1382), .ZN(new_n1383));
  OAI21_X1  g1183(.A(new_n1383), .B1(new_n1366), .B2(new_n1370), .ZN(new_n1384));
  NAND3_X1  g1184(.A1(new_n1365), .A2(G384), .A3(new_n1328), .ZN(new_n1385));
  OAI21_X1  g1185(.A(new_n1368), .B1(new_n1367), .B2(new_n1369), .ZN(new_n1386));
  NAND3_X1  g1186(.A1(new_n1385), .A2(new_n1386), .A3(new_n1382), .ZN(new_n1387));
  NAND2_X1  g1187(.A1(new_n1384), .A2(new_n1387), .ZN(new_n1388));
  INV_X1    g1188(.A(new_n1388), .ZN(new_n1389));
  NAND2_X1  g1189(.A1(new_n1381), .A2(new_n1389), .ZN(new_n1390));
  NAND3_X1  g1190(.A1(new_n1379), .A2(new_n1380), .A3(new_n1390), .ZN(new_n1391));
  OAI21_X1  g1191(.A(new_n1349), .B1(new_n1377), .B2(new_n1391), .ZN(new_n1392));
  NAND2_X1  g1192(.A1(new_n1390), .A2(KEYINPUT63), .ZN(new_n1393));
  NAND2_X1  g1193(.A1(new_n1393), .A2(new_n1372), .ZN(new_n1394));
  NAND3_X1  g1194(.A1(new_n1375), .A2(KEYINPUT63), .A3(new_n1371), .ZN(new_n1395));
  NAND3_X1  g1195(.A1(new_n1347), .A2(new_n1380), .A3(new_n1348), .ZN(new_n1396));
  INV_X1    g1196(.A(KEYINPUT124), .ZN(new_n1397));
  NAND2_X1  g1197(.A1(new_n1396), .A2(new_n1397), .ZN(new_n1398));
  NAND4_X1  g1198(.A1(new_n1347), .A2(KEYINPUT124), .A3(new_n1380), .A4(new_n1348), .ZN(new_n1399));
  AND2_X1   g1199(.A1(new_n1398), .A2(new_n1399), .ZN(new_n1400));
  NAND3_X1  g1200(.A1(new_n1394), .A2(new_n1395), .A3(new_n1400), .ZN(new_n1401));
  NAND3_X1  g1201(.A1(new_n1392), .A2(KEYINPUT126), .A3(new_n1401), .ZN(new_n1402));
  INV_X1    g1202(.A(KEYINPUT126), .ZN(new_n1403));
  INV_X1    g1203(.A(new_n1349), .ZN(new_n1404));
  OAI21_X1  g1204(.A(new_n1380), .B1(new_n1375), .B2(new_n1388), .ZN(new_n1405));
  AOI21_X1  g1205(.A(KEYINPUT62), .B1(new_n1375), .B2(new_n1371), .ZN(new_n1406));
  AOI21_X1  g1206(.A(new_n1405), .B1(new_n1378), .B2(new_n1406), .ZN(new_n1407));
  NAND3_X1  g1207(.A1(new_n1374), .A2(KEYINPUT125), .A3(new_n1376), .ZN(new_n1408));
  AOI21_X1  g1208(.A(new_n1404), .B1(new_n1407), .B2(new_n1408), .ZN(new_n1409));
  NAND3_X1  g1209(.A1(new_n1398), .A2(new_n1395), .A3(new_n1399), .ZN(new_n1410));
  AOI21_X1  g1210(.A(new_n1410), .B1(new_n1372), .B2(new_n1393), .ZN(new_n1411));
  OAI21_X1  g1211(.A(new_n1403), .B1(new_n1409), .B2(new_n1411), .ZN(new_n1412));
  NAND2_X1  g1212(.A1(new_n1402), .A2(new_n1412), .ZN(G405));
  XNOR2_X1  g1213(.A(G375), .B(new_n1331), .ZN(new_n1414));
  INV_X1    g1214(.A(new_n1371), .ZN(new_n1415));
  OR2_X1    g1215(.A1(new_n1414), .A2(new_n1415), .ZN(new_n1416));
  INV_X1    g1216(.A(KEYINPUT127), .ZN(new_n1417));
  NAND2_X1  g1217(.A1(new_n1414), .A2(new_n1415), .ZN(new_n1418));
  NAND4_X1  g1218(.A1(new_n1416), .A2(new_n1417), .A3(new_n1349), .A4(new_n1418), .ZN(new_n1419));
  AND2_X1   g1219(.A1(new_n1416), .A2(new_n1418), .ZN(new_n1420));
  XNOR2_X1  g1220(.A(new_n1349), .B(new_n1417), .ZN(new_n1421));
  OAI21_X1  g1221(.A(new_n1419), .B1(new_n1420), .B2(new_n1421), .ZN(G402));
endmodule


