//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 1 0 0 1 0 1 0 0 0 1 1 0 0 1 0 0 1 1 0 1 0 0 0 0 0 0 1 0 1 1 0 0 0 1 0 1 1 1 1 1 1 1 0 1 1 1 0 0 0 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:48 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n210, new_n211, new_n212, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n233, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n242, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n691, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1059, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1212,
    new_n1213, new_n1214, new_n1215, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1283, new_n1284, new_n1285, new_n1286, new_n1287,
    new_n1288;
  INV_X1    g0000(.A(KEYINPUT64), .ZN(new_n201));
  INV_X1    g0001(.A(G58), .ZN(new_n202));
  INV_X1    g0002(.A(G68), .ZN(new_n203));
  NAND3_X1  g0003(.A1(new_n201), .A2(new_n202), .A3(new_n203), .ZN(new_n204));
  OAI21_X1  g0004(.A(KEYINPUT64), .B1(G58), .B2(G68), .ZN(new_n205));
  NAND2_X1  g0005(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  INV_X1    g0006(.A(G50), .ZN(new_n207));
  NAND2_X1  g0007(.A1(new_n206), .A2(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G77), .ZN(G353));
  INV_X1    g0009(.A(G97), .ZN(new_n210));
  INV_X1    g0010(.A(G107), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n210), .A2(new_n211), .ZN(new_n212));
  NAND2_X1  g0012(.A1(new_n212), .A2(G87), .ZN(G355));
  INV_X1    g0013(.A(G1), .ZN(new_n214));
  INV_X1    g0014(.A(G20), .ZN(new_n215));
  NOR2_X1   g0015(.A1(new_n214), .A2(new_n215), .ZN(new_n216));
  INV_X1    g0016(.A(new_n216), .ZN(new_n217));
  NOR2_X1   g0017(.A1(new_n217), .A2(G13), .ZN(new_n218));
  OAI211_X1 g0018(.A(new_n218), .B(G250), .C1(G257), .C2(G264), .ZN(new_n219));
  XNOR2_X1  g0019(.A(new_n219), .B(KEYINPUT0), .ZN(new_n220));
  NOR2_X1   g0020(.A1(new_n206), .A2(new_n207), .ZN(new_n221));
  NAND2_X1  g0021(.A1(G1), .A2(G13), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n222), .A2(new_n215), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n221), .A2(new_n223), .ZN(new_n224));
  XOR2_X1   g0024(.A(KEYINPUT65), .B(G238), .Z(new_n225));
  NOR2_X1   g0025(.A1(new_n225), .A2(new_n203), .ZN(new_n226));
  AOI22_X1  g0026(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n227));
  AOI22_X1  g0027(.A1(G58), .A2(G232), .B1(G77), .B2(G244), .ZN(new_n228));
  AOI22_X1  g0028(.A1(G50), .A2(G226), .B1(G97), .B2(G257), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G107), .A2(G264), .ZN(new_n230));
  NAND4_X1  g0030(.A1(new_n227), .A2(new_n228), .A3(new_n229), .A4(new_n230), .ZN(new_n231));
  OAI21_X1  g0031(.A(new_n217), .B1(new_n226), .B2(new_n231), .ZN(new_n232));
  OAI211_X1 g0032(.A(new_n220), .B(new_n224), .C1(KEYINPUT1), .C2(new_n232), .ZN(new_n233));
  AOI21_X1  g0033(.A(new_n233), .B1(KEYINPUT1), .B2(new_n232), .ZN(G361));
  XOR2_X1   g0034(.A(G238), .B(G244), .Z(new_n235));
  XNOR2_X1  g0035(.A(G226), .B(G232), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(KEYINPUT66), .B(KEYINPUT2), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(G264), .B(G270), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G358));
  XNOR2_X1  g0043(.A(G87), .B(G97), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G107), .B(G116), .ZN(new_n245));
  XNOR2_X1  g0045(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n207), .A2(G68), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n203), .A2(G50), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  XNOR2_X1  g0049(.A(G58), .B(G77), .ZN(new_n250));
  XNOR2_X1  g0050(.A(new_n249), .B(new_n250), .ZN(new_n251));
  XOR2_X1   g0051(.A(new_n246), .B(new_n251), .Z(G351));
  AND2_X1   g0052(.A1(KEYINPUT67), .A2(G41), .ZN(new_n253));
  NOR2_X1   g0053(.A1(KEYINPUT67), .A2(G41), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n253), .A2(new_n254), .A3(G45), .ZN(new_n255));
  OAI21_X1  g0055(.A(KEYINPUT68), .B1(new_n255), .B2(G1), .ZN(new_n256));
  NAND2_X1  g0056(.A1(G33), .A2(G41), .ZN(new_n257));
  NAND3_X1  g0057(.A1(new_n257), .A2(G1), .A3(G13), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n258), .A2(G274), .ZN(new_n259));
  INV_X1    g0059(.A(new_n259), .ZN(new_n260));
  OR2_X1    g0060(.A1(KEYINPUT67), .A2(G41), .ZN(new_n261));
  INV_X1    g0061(.A(G45), .ZN(new_n262));
  NAND2_X1  g0062(.A1(KEYINPUT67), .A2(G41), .ZN(new_n263));
  NAND3_X1  g0063(.A1(new_n261), .A2(new_n262), .A3(new_n263), .ZN(new_n264));
  INV_X1    g0064(.A(KEYINPUT68), .ZN(new_n265));
  NAND3_X1  g0065(.A1(new_n264), .A2(new_n265), .A3(new_n214), .ZN(new_n266));
  NAND3_X1  g0066(.A1(new_n256), .A2(new_n260), .A3(new_n266), .ZN(new_n267));
  INV_X1    g0067(.A(KEYINPUT3), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n268), .A2(G33), .ZN(new_n269));
  INV_X1    g0069(.A(G33), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT3), .ZN(new_n271));
  NAND2_X1  g0071(.A1(new_n269), .A2(new_n271), .ZN(new_n272));
  INV_X1    g0072(.A(G77), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n258), .B1(new_n272), .B2(new_n273), .ZN(new_n274));
  XNOR2_X1  g0074(.A(KEYINPUT3), .B(G33), .ZN(new_n275));
  NOR2_X1   g0075(.A1(G222), .A2(G1698), .ZN(new_n276));
  INV_X1    g0076(.A(G1698), .ZN(new_n277));
  NOR2_X1   g0077(.A1(new_n277), .A2(G223), .ZN(new_n278));
  OAI21_X1  g0078(.A(new_n275), .B1(new_n276), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g0079(.A(new_n214), .B1(G41), .B2(G45), .ZN(new_n280));
  AND2_X1   g0080(.A1(new_n258), .A2(new_n280), .ZN(new_n281));
  AOI22_X1  g0081(.A1(new_n274), .A2(new_n279), .B1(new_n281), .B2(G226), .ZN(new_n282));
  NAND2_X1  g0082(.A1(new_n267), .A2(new_n282), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n283), .A2(G179), .ZN(new_n284));
  XNOR2_X1  g0084(.A(KEYINPUT8), .B(G58), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n215), .A2(G33), .ZN(new_n286));
  INV_X1    g0086(.A(G150), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n215), .A2(new_n270), .ZN(new_n288));
  OAI22_X1  g0088(.A1(new_n285), .A2(new_n286), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NAND2_X1  g0089(.A1(new_n289), .A2(KEYINPUT69), .ZN(new_n290));
  NAND2_X1  g0090(.A1(new_n208), .A2(G20), .ZN(new_n291));
  INV_X1    g0091(.A(KEYINPUT69), .ZN(new_n292));
  OAI221_X1 g0092(.A(new_n292), .B1(new_n287), .B2(new_n288), .C1(new_n285), .C2(new_n286), .ZN(new_n293));
  NAND3_X1  g0093(.A1(new_n290), .A2(new_n291), .A3(new_n293), .ZN(new_n294));
  NAND3_X1  g0094(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n295));
  NAND2_X1  g0095(.A1(new_n295), .A2(new_n222), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(new_n296), .ZN(new_n297));
  INV_X1    g0097(.A(G13), .ZN(new_n298));
  NOR3_X1   g0098(.A1(new_n298), .A2(new_n215), .A3(G1), .ZN(new_n299));
  NOR2_X1   g0099(.A1(new_n299), .A2(new_n296), .ZN(new_n300));
  INV_X1    g0100(.A(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n214), .A2(G20), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n302), .A2(G50), .ZN(new_n303));
  INV_X1    g0103(.A(new_n299), .ZN(new_n304));
  OAI22_X1  g0104(.A1(new_n301), .A2(new_n303), .B1(G50), .B2(new_n304), .ZN(new_n305));
  INV_X1    g0105(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n297), .A2(new_n306), .ZN(new_n307));
  INV_X1    g0107(.A(new_n307), .ZN(new_n308));
  INV_X1    g0108(.A(G169), .ZN(new_n309));
  AOI211_X1 g0109(.A(new_n284), .B(new_n308), .C1(new_n309), .C2(new_n283), .ZN(new_n310));
  NAND2_X1  g0110(.A1(new_n283), .A2(G200), .ZN(new_n311));
  INV_X1    g0111(.A(KEYINPUT72), .ZN(new_n312));
  NOR2_X1   g0112(.A1(new_n311), .A2(new_n312), .ZN(new_n313));
  AOI21_X1  g0113(.A(KEYINPUT72), .B1(new_n283), .B2(G200), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n313), .A2(KEYINPUT10), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g0115(.A1(new_n307), .A2(KEYINPUT9), .ZN(new_n316));
  INV_X1    g0116(.A(KEYINPUT71), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT9), .ZN(new_n318));
  NAND3_X1  g0118(.A1(new_n297), .A2(new_n318), .A3(new_n306), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n316), .A2(new_n317), .A3(new_n319), .ZN(new_n320));
  AOI211_X1 g0120(.A(KEYINPUT9), .B(new_n305), .C1(new_n294), .C2(new_n296), .ZN(new_n321));
  AOI21_X1  g0121(.A(new_n318), .B1(new_n297), .B2(new_n306), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT71), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND3_X1  g0123(.A1(new_n267), .A2(G190), .A3(new_n282), .ZN(new_n324));
  INV_X1    g0124(.A(KEYINPUT73), .ZN(new_n325));
  XNOR2_X1  g0125(.A(new_n324), .B(new_n325), .ZN(new_n326));
  NAND4_X1  g0126(.A1(new_n315), .A2(new_n320), .A3(new_n323), .A4(new_n326), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n311), .ZN(new_n328));
  NOR2_X1   g0128(.A1(new_n321), .A2(new_n322), .ZN(new_n329));
  OAI21_X1  g0129(.A(KEYINPUT10), .B1(new_n328), .B2(new_n329), .ZN(new_n330));
  AOI21_X1  g0130(.A(new_n310), .B1(new_n327), .B2(new_n330), .ZN(new_n331));
  NAND2_X1  g0131(.A1(new_n202), .A2(KEYINPUT8), .ZN(new_n332));
  INV_X1    g0132(.A(KEYINPUT8), .ZN(new_n333));
  NAND2_X1  g0133(.A1(new_n333), .A2(G58), .ZN(new_n334));
  NAND2_X1  g0134(.A1(new_n332), .A2(new_n334), .ZN(new_n335));
  AND2_X1   g0135(.A1(new_n335), .A2(new_n302), .ZN(new_n336));
  AOI22_X1  g0136(.A1(new_n336), .A2(new_n300), .B1(new_n299), .B2(new_n285), .ZN(new_n337));
  INV_X1    g0137(.A(new_n337), .ZN(new_n338));
  NAND2_X1  g0138(.A1(G58), .A2(G68), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n204), .A2(new_n205), .A3(new_n339), .ZN(new_n340));
  INV_X1    g0140(.A(G159), .ZN(new_n341));
  OAI21_X1  g0141(.A(KEYINPUT77), .B1(new_n288), .B2(new_n341), .ZN(new_n342));
  NOR2_X1   g0142(.A1(G20), .A2(G33), .ZN(new_n343));
  INV_X1    g0143(.A(KEYINPUT77), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n343), .A2(new_n344), .A3(G159), .ZN(new_n345));
  AOI22_X1  g0145(.A1(G20), .A2(new_n340), .B1(new_n342), .B2(new_n345), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT76), .ZN(new_n347));
  AND3_X1   g0147(.A1(new_n269), .A2(new_n271), .A3(new_n347), .ZN(new_n348));
  AOI21_X1  g0148(.A(new_n347), .B1(new_n269), .B2(new_n271), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT7), .ZN(new_n350));
  NAND2_X1  g0150(.A1(new_n350), .A2(new_n215), .ZN(new_n351));
  NOR3_X1   g0151(.A1(new_n348), .A2(new_n349), .A3(new_n351), .ZN(new_n352));
  AOI21_X1  g0152(.A(G20), .B1(new_n269), .B2(new_n271), .ZN(new_n353));
  OAI21_X1  g0153(.A(G68), .B1(new_n353), .B2(new_n350), .ZN(new_n354));
  OAI211_X1 g0154(.A(KEYINPUT16), .B(new_n346), .C1(new_n352), .C2(new_n354), .ZN(new_n355));
  AND2_X1   g0155(.A1(new_n355), .A2(new_n296), .ZN(new_n356));
  INV_X1    g0156(.A(KEYINPUT16), .ZN(new_n357));
  OAI21_X1  g0157(.A(KEYINPUT78), .B1(new_n270), .B2(KEYINPUT3), .ZN(new_n358));
  INV_X1    g0158(.A(KEYINPUT78), .ZN(new_n359));
  NAND3_X1  g0159(.A1(new_n359), .A2(new_n268), .A3(G33), .ZN(new_n360));
  NAND3_X1  g0160(.A1(new_n358), .A2(new_n360), .A3(new_n271), .ZN(new_n361));
  NOR2_X1   g0161(.A1(new_n350), .A2(G20), .ZN(new_n362));
  NAND2_X1  g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  OAI21_X1  g0163(.A(new_n350), .B1(new_n275), .B2(G20), .ZN(new_n364));
  AOI21_X1  g0164(.A(new_n203), .B1(new_n363), .B2(new_n364), .ZN(new_n365));
  NAND2_X1  g0165(.A1(new_n340), .A2(G20), .ZN(new_n366));
  NAND2_X1  g0166(.A1(new_n342), .A2(new_n345), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  OAI21_X1  g0168(.A(new_n357), .B1(new_n365), .B2(new_n368), .ZN(new_n369));
  AOI21_X1  g0169(.A(new_n338), .B1(new_n356), .B2(new_n369), .ZN(new_n370));
  OR2_X1    g0170(.A1(G223), .A2(G1698), .ZN(new_n371));
  OAI21_X1  g0171(.A(new_n371), .B1(G226), .B2(new_n277), .ZN(new_n372));
  INV_X1    g0172(.A(G87), .ZN(new_n373));
  OAI22_X1  g0173(.A1(new_n372), .A2(new_n272), .B1(new_n270), .B2(new_n373), .ZN(new_n374));
  AOI21_X1  g0174(.A(new_n222), .B1(G33), .B2(G41), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n374), .A2(new_n375), .ZN(new_n376));
  INV_X1    g0176(.A(KEYINPUT79), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n258), .A2(new_n280), .ZN(new_n378));
  INV_X1    g0178(.A(G232), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  NAND4_X1  g0180(.A1(new_n258), .A2(new_n280), .A3(KEYINPUT79), .A4(G232), .ZN(new_n381));
  NAND2_X1  g0181(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  NAND3_X1  g0182(.A1(new_n267), .A2(new_n376), .A3(new_n382), .ZN(new_n383));
  NAND2_X1  g0183(.A1(new_n383), .A2(G169), .ZN(new_n384));
  AOI22_X1  g0184(.A1(new_n380), .A2(new_n381), .B1(new_n374), .B2(new_n375), .ZN(new_n385));
  NAND3_X1  g0185(.A1(new_n385), .A2(G179), .A3(new_n267), .ZN(new_n386));
  AND2_X1   g0186(.A1(new_n384), .A2(new_n386), .ZN(new_n387));
  OAI21_X1  g0187(.A(KEYINPUT18), .B1(new_n370), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n383), .A2(G200), .ZN(new_n389));
  NAND3_X1  g0189(.A1(new_n385), .A2(G190), .A3(new_n267), .ZN(new_n390));
  AND2_X1   g0190(.A1(new_n389), .A2(new_n390), .ZN(new_n391));
  NAND3_X1  g0191(.A1(new_n370), .A2(new_n391), .A3(KEYINPUT17), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n369), .A2(new_n296), .A3(new_n355), .ZN(new_n393));
  NAND4_X1  g0193(.A1(new_n393), .A2(new_n337), .A3(new_n389), .A4(new_n390), .ZN(new_n394));
  INV_X1    g0194(.A(KEYINPUT17), .ZN(new_n395));
  NAND2_X1  g0195(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g0196(.A1(new_n355), .A2(new_n296), .ZN(new_n397));
  NAND2_X1  g0197(.A1(new_n363), .A2(new_n364), .ZN(new_n398));
  NAND2_X1  g0198(.A1(new_n398), .A2(G68), .ZN(new_n399));
  AOI21_X1  g0199(.A(KEYINPUT16), .B1(new_n399), .B2(new_n346), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n337), .B1(new_n397), .B2(new_n400), .ZN(new_n401));
  INV_X1    g0201(.A(KEYINPUT18), .ZN(new_n402));
  NAND2_X1  g0202(.A1(new_n384), .A2(new_n386), .ZN(new_n403));
  NAND3_X1  g0203(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  NAND4_X1  g0204(.A1(new_n388), .A2(new_n392), .A3(new_n396), .A4(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(new_n405), .ZN(new_n406));
  NAND3_X1  g0206(.A1(new_n275), .A2(G232), .A3(new_n277), .ZN(new_n407));
  NAND2_X1  g0207(.A1(new_n275), .A2(G1698), .ZN(new_n408));
  OAI221_X1 g0208(.A(new_n407), .B1(new_n211), .B2(new_n275), .C1(new_n408), .C2(new_n225), .ZN(new_n409));
  AOI21_X1  g0209(.A(new_n258), .B1(new_n409), .B2(KEYINPUT70), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(KEYINPUT70), .B2(new_n409), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n264), .A2(new_n214), .ZN(new_n412));
  AOI21_X1  g0212(.A(new_n259), .B1(new_n412), .B2(KEYINPUT68), .ZN(new_n413));
  AOI22_X1  g0213(.A1(new_n413), .A2(new_n266), .B1(G244), .B2(new_n281), .ZN(new_n414));
  AND2_X1   g0214(.A1(new_n411), .A2(new_n414), .ZN(new_n415));
  INV_X1    g0215(.A(G179), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n415), .A2(new_n416), .ZN(new_n417));
  AOI22_X1  g0217(.A1(new_n335), .A2(new_n343), .B1(G20), .B2(G77), .ZN(new_n418));
  XOR2_X1   g0218(.A(KEYINPUT15), .B(G87), .Z(new_n419));
  INV_X1    g0219(.A(new_n419), .ZN(new_n420));
  OAI21_X1  g0220(.A(new_n418), .B1(new_n420), .B2(new_n286), .ZN(new_n421));
  AND2_X1   g0221(.A1(new_n421), .A2(new_n296), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n300), .A2(G77), .A3(new_n302), .ZN(new_n423));
  OAI21_X1  g0223(.A(new_n423), .B1(G77), .B2(new_n304), .ZN(new_n424));
  NOR2_X1   g0224(.A1(new_n422), .A2(new_n424), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n411), .A2(new_n414), .ZN(new_n426));
  AOI21_X1  g0226(.A(new_n425), .B1(new_n426), .B2(new_n309), .ZN(new_n427));
  NAND2_X1  g0227(.A1(new_n417), .A2(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(new_n425), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n415), .B2(G190), .ZN(new_n430));
  NAND2_X1  g0230(.A1(new_n426), .A2(G200), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n430), .A2(new_n431), .ZN(new_n432));
  NAND4_X1  g0232(.A1(new_n331), .A2(new_n406), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  NAND2_X1  g0233(.A1(new_n299), .A2(new_n203), .ZN(new_n434));
  XNOR2_X1  g0234(.A(new_n434), .B(KEYINPUT12), .ZN(new_n435));
  AOI22_X1  g0235(.A1(new_n343), .A2(G50), .B1(G20), .B2(new_n203), .ZN(new_n436));
  OAI21_X1  g0236(.A(new_n436), .B1(new_n273), .B2(new_n286), .ZN(new_n437));
  NAND3_X1  g0237(.A1(new_n437), .A2(KEYINPUT11), .A3(new_n296), .ZN(new_n438));
  NAND3_X1  g0238(.A1(new_n300), .A2(G68), .A3(new_n302), .ZN(new_n439));
  NAND3_X1  g0239(.A1(new_n435), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  AOI21_X1  g0240(.A(KEYINPUT11), .B1(new_n437), .B2(new_n296), .ZN(new_n441));
  NOR2_X1   g0241(.A1(new_n440), .A2(new_n441), .ZN(new_n442));
  INV_X1    g0242(.A(new_n442), .ZN(new_n443));
  INV_X1    g0243(.A(KEYINPUT14), .ZN(new_n444));
  INV_X1    g0244(.A(KEYINPUT13), .ZN(new_n445));
  INV_X1    g0245(.A(KEYINPUT74), .ZN(new_n446));
  NAND2_X1  g0246(.A1(new_n267), .A2(new_n446), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n413), .A2(KEYINPUT74), .A3(new_n266), .ZN(new_n448));
  NAND2_X1  g0248(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n378), .A2(KEYINPUT75), .ZN(new_n450));
  INV_X1    g0250(.A(KEYINPUT75), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n258), .A2(new_n451), .A3(new_n280), .ZN(new_n452));
  NAND3_X1  g0252(.A1(new_n450), .A2(G238), .A3(new_n452), .ZN(new_n453));
  NAND2_X1  g0253(.A1(G33), .A2(G97), .ZN(new_n454));
  NAND2_X1  g0254(.A1(new_n379), .A2(G1698), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n455), .B1(G226), .B2(G1698), .ZN(new_n456));
  OAI21_X1  g0256(.A(new_n454), .B1(new_n456), .B2(new_n272), .ZN(new_n457));
  NAND2_X1  g0257(.A1(new_n457), .A2(new_n375), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n453), .A2(new_n458), .ZN(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  AOI21_X1  g0260(.A(new_n445), .B1(new_n449), .B2(new_n460), .ZN(new_n461));
  AOI211_X1 g0261(.A(KEYINPUT13), .B(new_n459), .C1(new_n447), .C2(new_n448), .ZN(new_n462));
  OAI211_X1 g0262(.A(new_n444), .B(G169), .C1(new_n461), .C2(new_n462), .ZN(new_n463));
  NOR2_X1   g0263(.A1(new_n267), .A2(new_n446), .ZN(new_n464));
  AOI21_X1  g0264(.A(KEYINPUT74), .B1(new_n413), .B2(new_n266), .ZN(new_n465));
  OAI21_X1  g0265(.A(new_n460), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g0266(.A1(new_n466), .A2(KEYINPUT13), .ZN(new_n467));
  NAND3_X1  g0267(.A1(new_n449), .A2(new_n445), .A3(new_n460), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n467), .A2(G179), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n463), .A2(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n467), .A2(new_n468), .ZN(new_n471));
  AOI21_X1  g0271(.A(new_n444), .B1(new_n471), .B2(G169), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n443), .B1(new_n470), .B2(new_n472), .ZN(new_n473));
  OAI21_X1  g0273(.A(G200), .B1(new_n461), .B2(new_n462), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n467), .A2(G190), .A3(new_n468), .ZN(new_n475));
  NAND3_X1  g0275(.A1(new_n474), .A2(new_n442), .A3(new_n475), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n473), .A2(new_n476), .ZN(new_n477));
  NOR2_X1   g0277(.A1(new_n433), .A2(new_n477), .ZN(new_n478));
  NAND4_X1  g0278(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(G1698), .ZN(new_n479));
  NAND2_X1  g0279(.A1(G33), .A2(G283), .ZN(new_n480));
  NAND4_X1  g0280(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(new_n277), .ZN(new_n481));
  INV_X1    g0281(.A(KEYINPUT4), .ZN(new_n482));
  OAI211_X1 g0282(.A(new_n479), .B(new_n480), .C1(new_n481), .C2(new_n482), .ZN(new_n483));
  XNOR2_X1  g0283(.A(KEYINPUT80), .B(KEYINPUT4), .ZN(new_n484));
  AND2_X1   g0284(.A1(new_n481), .A2(new_n484), .ZN(new_n485));
  OAI21_X1  g0285(.A(new_n375), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  INV_X1    g0286(.A(KEYINPUT81), .ZN(new_n487));
  INV_X1    g0287(.A(KEYINPUT5), .ZN(new_n488));
  OAI211_X1 g0288(.A(new_n214), .B(G45), .C1(new_n488), .C2(G41), .ZN(new_n489));
  INV_X1    g0289(.A(new_n489), .ZN(new_n490));
  OAI21_X1  g0290(.A(new_n488), .B1(new_n253), .B2(new_n254), .ZN(new_n491));
  AOI21_X1  g0291(.A(new_n375), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  NAND2_X1  g0292(.A1(new_n261), .A2(new_n263), .ZN(new_n493));
  AOI21_X1  g0293(.A(new_n489), .B1(new_n493), .B2(new_n488), .ZN(new_n494));
  AOI22_X1  g0294(.A1(new_n492), .A2(G257), .B1(new_n494), .B2(new_n260), .ZN(new_n495));
  AND3_X1   g0295(.A1(new_n486), .A2(new_n487), .A3(new_n495), .ZN(new_n496));
  AOI21_X1  g0296(.A(new_n487), .B1(new_n486), .B2(new_n495), .ZN(new_n497));
  OAI21_X1  g0297(.A(new_n309), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  NAND3_X1  g0298(.A1(new_n486), .A2(new_n416), .A3(new_n495), .ZN(new_n499));
  NAND2_X1  g0299(.A1(new_n499), .A2(KEYINPUT82), .ZN(new_n500));
  INV_X1    g0300(.A(KEYINPUT82), .ZN(new_n501));
  NAND4_X1  g0301(.A1(new_n486), .A2(new_n495), .A3(new_n501), .A4(new_n416), .ZN(new_n502));
  NAND2_X1  g0302(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(KEYINPUT6), .ZN(new_n504));
  NOR3_X1   g0304(.A1(new_n504), .A2(new_n210), .A3(G107), .ZN(new_n505));
  XNOR2_X1  g0305(.A(G97), .B(G107), .ZN(new_n506));
  AOI21_X1  g0306(.A(new_n505), .B1(new_n504), .B2(new_n506), .ZN(new_n507));
  OAI22_X1  g0307(.A1(new_n507), .A2(new_n215), .B1(new_n273), .B2(new_n288), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n211), .B1(new_n363), .B2(new_n364), .ZN(new_n509));
  OAI21_X1  g0309(.A(new_n296), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NOR2_X1   g0310(.A1(new_n304), .A2(G97), .ZN(new_n511));
  NAND2_X1  g0311(.A1(new_n214), .A2(G33), .ZN(new_n512));
  NAND2_X1  g0312(.A1(new_n300), .A2(new_n512), .ZN(new_n513));
  INV_X1    g0313(.A(new_n513), .ZN(new_n514));
  AOI21_X1  g0314(.A(new_n511), .B1(new_n514), .B2(G97), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n510), .A2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n498), .A2(new_n503), .A3(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n486), .A2(new_n495), .ZN(new_n518));
  NAND2_X1  g0318(.A1(new_n518), .A2(KEYINPUT81), .ZN(new_n519));
  NAND3_X1  g0319(.A1(new_n486), .A2(new_n487), .A3(new_n495), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n519), .A2(G190), .A3(new_n520), .ZN(new_n521));
  INV_X1    g0321(.A(new_n516), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n518), .A2(G200), .ZN(new_n523));
  NAND3_X1  g0323(.A1(new_n521), .A2(new_n522), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g0324(.A1(new_n275), .A2(new_n215), .A3(G68), .ZN(new_n525));
  INV_X1    g0325(.A(KEYINPUT19), .ZN(new_n526));
  OAI21_X1  g0326(.A(new_n215), .B1(new_n454), .B2(new_n526), .ZN(new_n527));
  OAI21_X1  g0327(.A(new_n527), .B1(G87), .B2(new_n212), .ZN(new_n528));
  OAI21_X1  g0328(.A(new_n526), .B1(new_n286), .B2(new_n210), .ZN(new_n529));
  NAND3_X1  g0329(.A1(new_n525), .A2(new_n528), .A3(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT83), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT83), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n525), .A2(new_n528), .A3(new_n532), .A4(new_n529), .ZN(new_n533));
  NAND3_X1  g0333(.A1(new_n531), .A2(new_n296), .A3(new_n533), .ZN(new_n534));
  NOR2_X1   g0334(.A1(new_n304), .A2(new_n419), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n514), .A2(G87), .ZN(new_n537));
  AND3_X1   g0337(.A1(new_n534), .A2(new_n536), .A3(new_n537), .ZN(new_n538));
  INV_X1    g0338(.A(G250), .ZN(new_n539));
  OAI21_X1  g0339(.A(new_n539), .B1(new_n262), .B2(G1), .ZN(new_n540));
  INV_X1    g0340(.A(G274), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n214), .A2(new_n541), .A3(G45), .ZN(new_n542));
  AND3_X1   g0342(.A1(new_n258), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND4_X1  g0343(.A1(new_n269), .A2(new_n271), .A3(G244), .A4(G1698), .ZN(new_n544));
  NAND4_X1  g0344(.A1(new_n269), .A2(new_n271), .A3(G238), .A4(new_n277), .ZN(new_n545));
  NAND2_X1  g0345(.A1(G33), .A2(G116), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n544), .A2(new_n545), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n543), .B1(new_n547), .B2(new_n375), .ZN(new_n548));
  INV_X1    g0348(.A(G200), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  AOI21_X1  g0350(.A(new_n550), .B1(G190), .B2(new_n548), .ZN(new_n551));
  AND2_X1   g0351(.A1(new_n548), .A2(new_n416), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n548), .A2(G169), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n514), .A2(new_n419), .ZN(new_n555));
  NAND3_X1  g0355(.A1(new_n534), .A2(new_n555), .A3(new_n536), .ZN(new_n556));
  AOI22_X1  g0356(.A1(new_n538), .A2(new_n551), .B1(new_n554), .B2(new_n556), .ZN(new_n557));
  AND3_X1   g0357(.A1(new_n517), .A2(new_n524), .A3(new_n557), .ZN(new_n558));
  AND3_X1   g0358(.A1(new_n211), .A2(KEYINPUT23), .A3(G20), .ZN(new_n559));
  AOI21_X1  g0359(.A(KEYINPUT23), .B1(new_n211), .B2(G20), .ZN(new_n560));
  OAI22_X1  g0360(.A1(new_n559), .A2(new_n560), .B1(G20), .B2(new_n546), .ZN(new_n561));
  NAND4_X1  g0361(.A1(new_n269), .A2(new_n271), .A3(new_n215), .A4(G87), .ZN(new_n562));
  NAND2_X1  g0362(.A1(new_n562), .A2(KEYINPUT22), .ZN(new_n563));
  INV_X1    g0363(.A(KEYINPUT22), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n275), .A2(new_n564), .A3(new_n215), .A4(G87), .ZN(new_n565));
  AOI211_X1 g0365(.A(KEYINPUT24), .B(new_n561), .C1(new_n563), .C2(new_n565), .ZN(new_n566));
  INV_X1    g0366(.A(KEYINPUT24), .ZN(new_n567));
  NAND2_X1  g0367(.A1(new_n563), .A2(new_n565), .ZN(new_n568));
  INV_X1    g0368(.A(new_n561), .ZN(new_n569));
  AOI21_X1  g0369(.A(new_n567), .B1(new_n568), .B2(new_n569), .ZN(new_n570));
  OAI21_X1  g0370(.A(new_n296), .B1(new_n566), .B2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(KEYINPUT25), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n304), .B2(G107), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n299), .A2(KEYINPUT25), .A3(new_n211), .ZN(new_n574));
  AOI22_X1  g0374(.A1(new_n514), .A2(G107), .B1(new_n573), .B2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n571), .A2(new_n575), .ZN(new_n576));
  NAND4_X1  g0376(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(G1698), .ZN(new_n577));
  NAND4_X1  g0377(.A1(new_n269), .A2(new_n271), .A3(G250), .A4(new_n277), .ZN(new_n578));
  NAND2_X1  g0378(.A1(G33), .A2(G294), .ZN(new_n579));
  NAND3_X1  g0379(.A1(new_n577), .A2(new_n578), .A3(new_n579), .ZN(new_n580));
  AOI21_X1  g0380(.A(new_n258), .B1(new_n580), .B2(KEYINPUT84), .ZN(new_n581));
  INV_X1    g0381(.A(KEYINPUT84), .ZN(new_n582));
  NAND4_X1  g0382(.A1(new_n577), .A2(new_n578), .A3(new_n582), .A4(new_n579), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n581), .A2(new_n583), .ZN(new_n584));
  NAND2_X1  g0384(.A1(new_n494), .A2(new_n260), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n492), .A2(G264), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g0387(.A1(new_n587), .A2(new_n309), .ZN(new_n588));
  AOI22_X1  g0388(.A1(new_n581), .A2(new_n583), .B1(G264), .B2(new_n492), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n589), .A2(new_n416), .A3(new_n585), .ZN(new_n590));
  NAND3_X1  g0390(.A1(new_n576), .A2(new_n588), .A3(new_n590), .ZN(new_n591));
  INV_X1    g0391(.A(new_n591), .ZN(new_n592));
  INV_X1    g0392(.A(G190), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n589), .A2(new_n593), .A3(new_n585), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n587), .A2(new_n549), .ZN(new_n595));
  AOI21_X1  g0395(.A(new_n576), .B1(new_n594), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n492), .A2(G270), .B1(new_n494), .B2(new_n260), .ZN(new_n597));
  NAND4_X1  g0397(.A1(new_n269), .A2(new_n271), .A3(G264), .A4(G1698), .ZN(new_n598));
  NAND4_X1  g0398(.A1(new_n269), .A2(new_n271), .A3(G257), .A4(new_n277), .ZN(new_n599));
  INV_X1    g0399(.A(G303), .ZN(new_n600));
  OAI211_X1 g0400(.A(new_n598), .B(new_n599), .C1(new_n600), .C2(new_n275), .ZN(new_n601));
  NAND2_X1  g0401(.A1(new_n601), .A2(new_n375), .ZN(new_n602));
  NAND2_X1  g0402(.A1(new_n597), .A2(new_n602), .ZN(new_n603));
  NAND3_X1  g0403(.A1(new_n300), .A2(G116), .A3(new_n512), .ZN(new_n604));
  INV_X1    g0404(.A(G116), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n299), .A2(new_n605), .ZN(new_n606));
  AOI22_X1  g0406(.A1(new_n295), .A2(new_n222), .B1(G20), .B2(new_n605), .ZN(new_n607));
  OAI211_X1 g0407(.A(new_n480), .B(new_n215), .C1(G33), .C2(new_n210), .ZN(new_n608));
  AND3_X1   g0408(.A1(new_n607), .A2(KEYINPUT20), .A3(new_n608), .ZN(new_n609));
  AOI21_X1  g0409(.A(KEYINPUT20), .B1(new_n607), .B2(new_n608), .ZN(new_n610));
  OAI211_X1 g0410(.A(new_n604), .B(new_n606), .C1(new_n609), .C2(new_n610), .ZN(new_n611));
  NAND3_X1  g0411(.A1(new_n603), .A2(G169), .A3(new_n611), .ZN(new_n612));
  INV_X1    g0412(.A(KEYINPUT21), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  AND2_X1   g0414(.A1(new_n601), .A2(new_n375), .ZN(new_n615));
  AOI21_X1  g0415(.A(KEYINPUT5), .B1(new_n261), .B2(new_n263), .ZN(new_n616));
  OAI211_X1 g0416(.A(G270), .B(new_n258), .C1(new_n616), .C2(new_n489), .ZN(new_n617));
  NAND2_X1  g0417(.A1(new_n585), .A2(new_n617), .ZN(new_n618));
  OAI21_X1  g0418(.A(G200), .B1(new_n615), .B2(new_n618), .ZN(new_n619));
  INV_X1    g0419(.A(new_n611), .ZN(new_n620));
  NAND3_X1  g0420(.A1(new_n597), .A2(G190), .A3(new_n602), .ZN(new_n621));
  NAND3_X1  g0421(.A1(new_n619), .A2(new_n620), .A3(new_n621), .ZN(new_n622));
  NAND4_X1  g0422(.A1(new_n603), .A2(KEYINPUT21), .A3(G169), .A4(new_n611), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n416), .B1(new_n601), .B2(new_n375), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n611), .A2(new_n597), .A3(new_n624), .ZN(new_n625));
  NAND4_X1  g0425(.A1(new_n614), .A2(new_n622), .A3(new_n623), .A4(new_n625), .ZN(new_n626));
  NOR3_X1   g0426(.A1(new_n592), .A2(new_n596), .A3(new_n626), .ZN(new_n627));
  AND3_X1   g0427(.A1(new_n478), .A2(new_n558), .A3(new_n627), .ZN(G372));
  INV_X1    g0428(.A(KEYINPUT86), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n629), .B1(new_n370), .B2(new_n387), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n401), .A2(KEYINPUT86), .A3(new_n403), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  XNOR2_X1  g0432(.A(KEYINPUT87), .B(KEYINPUT18), .ZN(new_n633));
  INV_X1    g0433(.A(new_n633), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n632), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n630), .A2(new_n631), .A3(new_n633), .ZN(new_n636));
  AND2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(new_n428), .ZN(new_n638));
  OAI21_X1  g0438(.A(G169), .B1(new_n461), .B2(new_n462), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n639), .A2(KEYINPUT14), .ZN(new_n640));
  NAND3_X1  g0440(.A1(new_n640), .A2(new_n469), .A3(new_n463), .ZN(new_n641));
  AOI21_X1  g0441(.A(new_n638), .B1(new_n641), .B2(new_n443), .ZN(new_n642));
  AND2_X1   g0442(.A1(new_n392), .A2(new_n396), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n643), .A2(new_n476), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n637), .B1(new_n642), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n327), .A2(new_n330), .ZN(new_n646));
  AOI21_X1  g0446(.A(new_n310), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  NAND3_X1  g0447(.A1(new_n614), .A2(new_n623), .A3(new_n625), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n592), .A2(new_n648), .ZN(new_n649));
  NAND2_X1  g0449(.A1(new_n595), .A2(new_n594), .ZN(new_n650));
  INV_X1    g0450(.A(new_n576), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n650), .A2(new_n651), .ZN(new_n652));
  NAND4_X1  g0452(.A1(new_n652), .A2(new_n517), .A3(new_n524), .A4(new_n557), .ZN(new_n653));
  AOI21_X1  g0453(.A(new_n649), .B1(new_n653), .B2(KEYINPUT85), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n654), .B1(KEYINPUT85), .B2(new_n653), .ZN(new_n655));
  INV_X1    g0455(.A(new_n554), .ZN(new_n656));
  INV_X1    g0456(.A(new_n556), .ZN(new_n657));
  NOR2_X1   g0457(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  INV_X1    g0458(.A(KEYINPUT26), .ZN(new_n659));
  INV_X1    g0459(.A(new_n557), .ZN(new_n660));
  OAI21_X1  g0460(.A(new_n659), .B1(new_n660), .B2(new_n517), .ZN(new_n661));
  INV_X1    g0461(.A(new_n517), .ZN(new_n662));
  NAND3_X1  g0462(.A1(new_n662), .A2(KEYINPUT26), .A3(new_n557), .ZN(new_n663));
  AOI21_X1  g0463(.A(new_n658), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  NAND2_X1  g0464(.A1(new_n655), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n665), .A2(new_n478), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n647), .A2(new_n666), .ZN(G369));
  NOR2_X1   g0467(.A1(new_n592), .A2(new_n596), .ZN(new_n668));
  NAND3_X1  g0468(.A1(new_n214), .A2(new_n215), .A3(G13), .ZN(new_n669));
  OR2_X1    g0469(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n670));
  NAND2_X1  g0470(.A1(new_n669), .A2(KEYINPUT27), .ZN(new_n671));
  NAND3_X1  g0471(.A1(new_n670), .A2(G213), .A3(new_n671), .ZN(new_n672));
  INV_X1    g0472(.A(G343), .ZN(new_n673));
  NOR2_X1   g0473(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  INV_X1    g0474(.A(new_n674), .ZN(new_n675));
  AND2_X1   g0475(.A1(new_n648), .A2(new_n675), .ZN(new_n676));
  AOI22_X1  g0476(.A1(new_n668), .A2(new_n676), .B1(new_n592), .B2(new_n675), .ZN(new_n677));
  NOR2_X1   g0477(.A1(new_n620), .A2(new_n675), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n648), .A2(new_n678), .ZN(new_n679));
  OAI21_X1  g0479(.A(new_n679), .B1(new_n626), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g0480(.A(new_n680), .B(KEYINPUT88), .ZN(new_n681));
  AOI21_X1  g0481(.A(KEYINPUT89), .B1(new_n681), .B2(G330), .ZN(new_n682));
  INV_X1    g0482(.A(new_n682), .ZN(new_n683));
  NAND3_X1  g0483(.A1(new_n681), .A2(KEYINPUT89), .A3(G330), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  INV_X1    g0485(.A(new_n685), .ZN(new_n686));
  OAI21_X1  g0486(.A(new_n668), .B1(new_n651), .B2(new_n675), .ZN(new_n687));
  NAND2_X1  g0487(.A1(new_n592), .A2(new_n674), .ZN(new_n688));
  NAND2_X1  g0488(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  INV_X1    g0489(.A(new_n689), .ZN(new_n690));
  OAI21_X1  g0490(.A(new_n677), .B1(new_n686), .B2(new_n690), .ZN(new_n691));
  XOR2_X1   g0491(.A(new_n691), .B(KEYINPUT90), .Z(G399));
  INV_X1    g0492(.A(new_n218), .ZN(new_n693));
  NOR2_X1   g0493(.A1(new_n693), .A2(new_n493), .ZN(new_n694));
  NAND2_X1  g0494(.A1(new_n694), .A2(new_n221), .ZN(new_n695));
  INV_X1    g0495(.A(new_n694), .ZN(new_n696));
  NAND2_X1  g0496(.A1(new_n696), .A2(G1), .ZN(new_n697));
  NOR3_X1   g0497(.A1(new_n212), .A2(G87), .A3(G116), .ZN(new_n698));
  XOR2_X1   g0498(.A(new_n698), .B(KEYINPUT91), .Z(new_n699));
  OAI21_X1  g0499(.A(new_n695), .B1(new_n697), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g0500(.A(new_n700), .B(KEYINPUT28), .ZN(new_n701));
  INV_X1    g0501(.A(new_n664), .ZN(new_n702));
  NOR2_X1   g0502(.A1(new_n653), .A2(new_n649), .ZN(new_n703));
  OAI211_X1 g0503(.A(KEYINPUT29), .B(new_n675), .C1(new_n702), .C2(new_n703), .ZN(new_n704));
  AOI21_X1  g0504(.A(new_n674), .B1(new_n655), .B2(new_n664), .ZN(new_n705));
  OAI21_X1  g0505(.A(new_n704), .B1(new_n705), .B2(KEYINPUT29), .ZN(new_n706));
  NAND3_X1  g0506(.A1(new_n627), .A2(new_n558), .A3(new_n675), .ZN(new_n707));
  AND3_X1   g0507(.A1(new_n624), .A2(new_n597), .A3(new_n548), .ZN(new_n708));
  NAND4_X1  g0508(.A1(new_n519), .A2(new_n520), .A3(new_n708), .A4(new_n589), .ZN(new_n709));
  INV_X1    g0509(.A(KEYINPUT30), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  NAND2_X1  g0511(.A1(new_n584), .A2(new_n586), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n624), .A2(new_n597), .A3(new_n548), .ZN(new_n713));
  NOR2_X1   g0513(.A1(new_n712), .A2(new_n713), .ZN(new_n714));
  NAND4_X1  g0514(.A1(new_n714), .A2(KEYINPUT30), .A3(new_n519), .A4(new_n520), .ZN(new_n715));
  NOR2_X1   g0515(.A1(new_n548), .A2(G179), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n587), .A2(new_n518), .A3(new_n603), .A4(new_n716), .ZN(new_n717));
  NAND3_X1  g0517(.A1(new_n711), .A2(new_n715), .A3(new_n717), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(new_n674), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT31), .ZN(new_n720));
  NAND2_X1  g0520(.A1(new_n719), .A2(new_n720), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n718), .A2(KEYINPUT31), .A3(new_n674), .ZN(new_n722));
  NAND3_X1  g0522(.A1(new_n707), .A2(new_n721), .A3(new_n722), .ZN(new_n723));
  NAND2_X1  g0523(.A1(new_n723), .A2(G330), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n706), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n701), .B1(new_n726), .B2(G1), .ZN(G364));
  NOR2_X1   g0527(.A1(new_n298), .A2(G20), .ZN(new_n728));
  AOI21_X1  g0528(.A(new_n214), .B1(new_n728), .B2(G45), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n696), .A2(KEYINPUT92), .A3(new_n729), .ZN(new_n730));
  INV_X1    g0530(.A(KEYINPUT92), .ZN(new_n731));
  INV_X1    g0531(.A(new_n729), .ZN(new_n732));
  OAI21_X1  g0532(.A(new_n731), .B1(new_n694), .B2(new_n732), .ZN(new_n733));
  NAND2_X1  g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  OAI211_X1 g0534(.A(new_n686), .B(new_n734), .C1(G330), .C2(new_n681), .ZN(new_n735));
  NOR2_X1   g0535(.A1(G13), .A2(G33), .ZN(new_n736));
  INV_X1    g0536(.A(new_n736), .ZN(new_n737));
  NOR2_X1   g0537(.A1(new_n737), .A2(G20), .ZN(new_n738));
  AOI21_X1  g0538(.A(new_n222), .B1(G20), .B2(new_n309), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  NOR2_X1   g0541(.A1(new_n348), .A2(new_n349), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(new_n218), .ZN(new_n743));
  XNOR2_X1  g0543(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  NAND2_X1  g0544(.A1(new_n221), .A2(new_n262), .ZN(new_n745));
  OAI211_X1 g0545(.A(new_n744), .B(new_n745), .C1(new_n262), .C2(new_n251), .ZN(new_n746));
  NAND2_X1  g0546(.A1(new_n218), .A2(new_n275), .ZN(new_n747));
  XNOR2_X1  g0547(.A(new_n747), .B(KEYINPUT93), .ZN(new_n748));
  XOR2_X1   g0548(.A(G355), .B(KEYINPUT94), .Z(new_n749));
  AOI22_X1  g0549(.A1(new_n748), .A2(new_n749), .B1(new_n605), .B2(new_n693), .ZN(new_n750));
  AOI21_X1  g0550(.A(new_n741), .B1(new_n746), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(new_n739), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n215), .A2(new_n416), .ZN(new_n753));
  NAND2_X1  g0553(.A1(new_n753), .A2(G200), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n754), .A2(G190), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n215), .A2(G179), .ZN(new_n757));
  NAND3_X1  g0557(.A1(new_n757), .A2(G190), .A3(G200), .ZN(new_n758));
  OAI22_X1  g0558(.A1(new_n756), .A2(new_n203), .B1(new_n373), .B2(new_n758), .ZN(new_n759));
  NOR2_X1   g0559(.A1(new_n754), .A2(new_n593), .ZN(new_n760));
  INV_X1    g0560(.A(new_n760), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND2_X1  g0562(.A1(new_n757), .A2(new_n762), .ZN(new_n763));
  INV_X1    g0563(.A(new_n763), .ZN(new_n764));
  NAND2_X1  g0564(.A1(new_n764), .A2(G159), .ZN(new_n765));
  OAI22_X1  g0565(.A1(new_n761), .A2(new_n207), .B1(new_n765), .B2(KEYINPUT32), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n759), .A2(new_n766), .ZN(new_n767));
  NAND3_X1  g0567(.A1(new_n757), .A2(new_n593), .A3(G200), .ZN(new_n768));
  XNOR2_X1  g0568(.A(new_n768), .B(KEYINPUT96), .ZN(new_n769));
  NAND2_X1  g0569(.A1(new_n769), .A2(G107), .ZN(new_n770));
  NAND3_X1  g0570(.A1(new_n753), .A2(G190), .A3(new_n549), .ZN(new_n771));
  OAI21_X1  g0571(.A(new_n275), .B1(new_n771), .B2(new_n202), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n753), .A2(new_n762), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n772), .B1(G77), .B2(new_n774), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n593), .A2(G179), .A3(G200), .ZN(new_n776));
  NOR2_X1   g0576(.A1(new_n776), .A2(new_n215), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n765), .A2(KEYINPUT32), .B1(new_n778), .B2(G97), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n767), .A2(new_n770), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  INV_X1    g0580(.A(new_n771), .ZN(new_n781));
  AOI22_X1  g0581(.A1(new_n781), .A2(G322), .B1(new_n764), .B2(G329), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n275), .B1(new_n774), .B2(G311), .ZN(new_n783));
  AND2_X1   g0583(.A1(new_n782), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n769), .A2(G283), .ZN(new_n785));
  XNOR2_X1  g0585(.A(KEYINPUT33), .B(G317), .ZN(new_n786));
  AOI22_X1  g0586(.A1(G294), .A2(new_n778), .B1(new_n755), .B2(new_n786), .ZN(new_n787));
  INV_X1    g0587(.A(new_n758), .ZN(new_n788));
  AOI22_X1  g0588(.A1(new_n760), .A2(G326), .B1(new_n788), .B2(G303), .ZN(new_n789));
  NAND4_X1  g0589(.A1(new_n784), .A2(new_n785), .A3(new_n787), .A4(new_n789), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n752), .B1(new_n780), .B2(new_n790), .ZN(new_n791));
  NOR3_X1   g0591(.A1(new_n751), .A2(new_n791), .A3(new_n734), .ZN(new_n792));
  INV_X1    g0592(.A(new_n738), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n792), .B1(new_n680), .B2(new_n793), .ZN(new_n794));
  AND2_X1   g0594(.A1(new_n735), .A2(new_n794), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(G396));
  NAND3_X1  g0596(.A1(new_n417), .A2(new_n427), .A3(new_n675), .ZN(new_n797));
  AOI22_X1  g0597(.A1(new_n430), .A2(new_n431), .B1(new_n429), .B2(new_n674), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n797), .B1(new_n798), .B2(new_n638), .ZN(new_n799));
  INV_X1    g0599(.A(new_n799), .ZN(new_n800));
  XNOR2_X1  g0600(.A(new_n705), .B(new_n800), .ZN(new_n801));
  NOR2_X1   g0601(.A1(new_n801), .A2(new_n724), .ZN(new_n802));
  XNOR2_X1  g0602(.A(new_n802), .B(KEYINPUT97), .ZN(new_n803));
  INV_X1    g0603(.A(new_n734), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n804), .B1(new_n801), .B2(new_n724), .ZN(new_n805));
  NAND2_X1  g0605(.A1(new_n803), .A2(new_n805), .ZN(new_n806));
  INV_X1    g0606(.A(G294), .ZN(new_n807));
  INV_X1    g0607(.A(G311), .ZN(new_n808));
  OAI22_X1  g0608(.A1(new_n771), .A2(new_n807), .B1(new_n763), .B2(new_n808), .ZN(new_n809));
  AOI211_X1 g0609(.A(new_n275), .B(new_n809), .C1(G116), .C2(new_n774), .ZN(new_n810));
  NAND2_X1  g0610(.A1(new_n769), .A2(G87), .ZN(new_n811));
  AOI22_X1  g0611(.A1(new_n778), .A2(G97), .B1(new_n788), .B2(G107), .ZN(new_n812));
  AOI22_X1  g0612(.A1(G283), .A2(new_n755), .B1(new_n760), .B2(G303), .ZN(new_n813));
  NAND4_X1  g0613(.A1(new_n810), .A2(new_n811), .A3(new_n812), .A4(new_n813), .ZN(new_n814));
  AOI22_X1  g0614(.A1(new_n781), .A2(G143), .B1(new_n774), .B2(G159), .ZN(new_n815));
  INV_X1    g0615(.A(G137), .ZN(new_n816));
  OAI221_X1 g0616(.A(new_n815), .B1(new_n756), .B2(new_n287), .C1(new_n816), .C2(new_n761), .ZN(new_n817));
  INV_X1    g0617(.A(KEYINPUT34), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n769), .A2(G68), .ZN(new_n820));
  AOI21_X1  g0620(.A(new_n742), .B1(G132), .B2(new_n764), .ZN(new_n821));
  AOI22_X1  g0621(.A1(new_n778), .A2(G58), .B1(new_n788), .B2(G50), .ZN(new_n822));
  NAND4_X1  g0622(.A1(new_n819), .A2(new_n820), .A3(new_n821), .A4(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n817), .A2(new_n818), .ZN(new_n824));
  OAI21_X1  g0624(.A(new_n814), .B1(new_n823), .B2(new_n824), .ZN(new_n825));
  NAND2_X1  g0625(.A1(new_n825), .A2(new_n739), .ZN(new_n826));
  NOR2_X1   g0626(.A1(new_n739), .A2(new_n736), .ZN(new_n827));
  AOI21_X1  g0627(.A(new_n734), .B1(new_n273), .B2(new_n827), .ZN(new_n828));
  OAI211_X1 g0628(.A(new_n826), .B(new_n828), .C1(new_n800), .C2(new_n737), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n806), .A2(new_n829), .ZN(G384));
  INV_X1    g0630(.A(new_n507), .ZN(new_n831));
  OR2_X1    g0631(.A1(new_n831), .A2(KEYINPUT35), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(KEYINPUT35), .ZN(new_n833));
  NAND4_X1  g0633(.A1(new_n832), .A2(G116), .A3(new_n223), .A4(new_n833), .ZN(new_n834));
  XOR2_X1   g0634(.A(new_n834), .B(KEYINPUT36), .Z(new_n835));
  NAND3_X1  g0635(.A1(new_n221), .A2(G77), .A3(new_n339), .ZN(new_n836));
  XNOR2_X1  g0636(.A(new_n247), .B(KEYINPUT98), .ZN(new_n837));
  AOI211_X1 g0637(.A(new_n214), .B(G13), .C1(new_n836), .C2(new_n837), .ZN(new_n838));
  NOR2_X1   g0638(.A1(new_n835), .A2(new_n838), .ZN(new_n839));
  NAND2_X1  g0639(.A1(new_n272), .A2(KEYINPUT76), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n275), .A2(new_n347), .ZN(new_n841));
  NAND4_X1  g0641(.A1(new_n840), .A2(new_n841), .A3(new_n350), .A4(new_n215), .ZN(new_n842));
  NAND2_X1  g0642(.A1(new_n272), .A2(new_n215), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n203), .B1(new_n843), .B2(KEYINPUT7), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n842), .A2(new_n844), .ZN(new_n845));
  AOI21_X1  g0645(.A(KEYINPUT16), .B1(new_n845), .B2(new_n346), .ZN(new_n846));
  OAI21_X1  g0646(.A(new_n337), .B1(new_n397), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n672), .ZN(new_n848));
  AND2_X1   g0648(.A1(new_n847), .A2(new_n848), .ZN(new_n849));
  NAND2_X1  g0649(.A1(new_n405), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g0650(.A1(new_n384), .A2(new_n386), .A3(new_n672), .ZN(new_n851));
  AND2_X1   g0651(.A1(new_n851), .A2(new_n847), .ZN(new_n852));
  INV_X1    g0652(.A(new_n394), .ZN(new_n853));
  OAI21_X1  g0653(.A(KEYINPUT37), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g0654(.A1(new_n401), .A2(new_n851), .ZN(new_n855));
  INV_X1    g0655(.A(KEYINPUT37), .ZN(new_n856));
  NAND3_X1  g0656(.A1(new_n855), .A2(new_n856), .A3(new_n394), .ZN(new_n857));
  NAND2_X1  g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  AND4_X1   g0658(.A1(KEYINPUT101), .A2(new_n850), .A3(KEYINPUT38), .A4(new_n858), .ZN(new_n859));
  AOI22_X1  g0659(.A1(new_n405), .A2(new_n849), .B1(new_n854), .B2(new_n857), .ZN(new_n860));
  AOI21_X1  g0660(.A(KEYINPUT101), .B1(new_n860), .B2(KEYINPUT38), .ZN(new_n861));
  NOR2_X1   g0661(.A1(new_n859), .A2(new_n861), .ZN(new_n862));
  INV_X1    g0662(.A(KEYINPUT100), .ZN(new_n863));
  AND3_X1   g0663(.A1(new_n401), .A2(KEYINPUT86), .A3(new_n403), .ZN(new_n864));
  AOI21_X1  g0664(.A(KEYINPUT86), .B1(new_n401), .B2(new_n403), .ZN(new_n865));
  OAI211_X1 g0665(.A(new_n863), .B(new_n394), .C1(new_n864), .C2(new_n865), .ZN(new_n866));
  NOR2_X1   g0666(.A1(new_n370), .A2(new_n672), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  NAND2_X1  g0668(.A1(new_n866), .A2(new_n868), .ZN(new_n869));
  AOI21_X1  g0669(.A(new_n863), .B1(new_n632), .B2(new_n394), .ZN(new_n870));
  OAI21_X1  g0670(.A(KEYINPUT37), .B1(new_n869), .B2(new_n870), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n635), .A2(new_n643), .A3(new_n636), .ZN(new_n872));
  AOI22_X1  g0672(.A1(new_n871), .A2(new_n857), .B1(new_n867), .B2(new_n872), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n862), .B1(new_n873), .B2(KEYINPUT38), .ZN(new_n874));
  INV_X1    g0674(.A(KEYINPUT39), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n641), .A2(new_n443), .A3(new_n675), .ZN(new_n877));
  INV_X1    g0677(.A(new_n877), .ZN(new_n878));
  OR2_X1    g0678(.A1(new_n860), .A2(KEYINPUT38), .ZN(new_n879));
  NAND2_X1  g0679(.A1(new_n860), .A2(KEYINPUT38), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n879), .A2(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(new_n875), .ZN(new_n882));
  INV_X1    g0682(.A(new_n882), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n876), .A2(new_n878), .A3(new_n883), .ZN(new_n884));
  XNOR2_X1  g0684(.A(new_n797), .B(KEYINPUT99), .ZN(new_n885));
  INV_X1    g0685(.A(new_n885), .ZN(new_n886));
  INV_X1    g0686(.A(new_n705), .ZN(new_n887));
  OAI21_X1  g0687(.A(new_n886), .B1(new_n887), .B2(new_n799), .ZN(new_n888));
  NAND2_X1  g0688(.A1(new_n443), .A2(new_n674), .ZN(new_n889));
  NAND3_X1  g0689(.A1(new_n473), .A2(new_n476), .A3(new_n889), .ZN(new_n890));
  INV_X1    g0690(.A(new_n476), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n443), .B(new_n674), .C1(new_n641), .C2(new_n891), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n890), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g0693(.A1(new_n888), .A2(new_n881), .A3(new_n893), .ZN(new_n894));
  OR2_X1    g0694(.A1(new_n637), .A2(new_n848), .ZN(new_n895));
  NAND3_X1  g0695(.A1(new_n884), .A2(new_n894), .A3(new_n895), .ZN(new_n896));
  OAI211_X1 g0696(.A(new_n478), .B(new_n704), .C1(new_n705), .C2(KEYINPUT29), .ZN(new_n897));
  AND2_X1   g0697(.A1(new_n897), .A2(new_n647), .ZN(new_n898));
  XOR2_X1   g0698(.A(new_n896), .B(new_n898), .Z(new_n899));
  AOI21_X1  g0699(.A(new_n799), .B1(new_n890), .B2(new_n892), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n723), .A2(KEYINPUT102), .ZN(new_n901));
  INV_X1    g0701(.A(KEYINPUT102), .ZN(new_n902));
  NAND4_X1  g0702(.A1(new_n707), .A2(new_n721), .A3(new_n902), .A4(new_n722), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n900), .A2(new_n901), .A3(new_n903), .ZN(new_n904));
  INV_X1    g0704(.A(KEYINPUT103), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NAND4_X1  g0706(.A1(new_n900), .A2(new_n901), .A3(KEYINPUT103), .A4(new_n903), .ZN(new_n907));
  NAND4_X1  g0707(.A1(new_n906), .A2(new_n874), .A3(KEYINPUT40), .A4(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n881), .A2(new_n900), .A3(new_n901), .A4(new_n903), .ZN(new_n909));
  INV_X1    g0709(.A(KEYINPUT40), .ZN(new_n910));
  NAND2_X1  g0710(.A1(new_n909), .A2(new_n910), .ZN(new_n911));
  NAND2_X1  g0711(.A1(new_n908), .A2(new_n911), .ZN(new_n912));
  AND2_X1   g0712(.A1(new_n901), .A2(new_n903), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n913), .A2(new_n478), .ZN(new_n914));
  OR2_X1    g0714(.A1(new_n912), .A2(new_n914), .ZN(new_n915));
  NAND2_X1  g0715(.A1(new_n912), .A2(new_n914), .ZN(new_n916));
  NAND3_X1  g0716(.A1(new_n915), .A2(G330), .A3(new_n916), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n899), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n214), .B2(new_n728), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n899), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n839), .B1(new_n919), .B2(new_n920), .ZN(G367));
  NOR2_X1   g0721(.A1(new_n686), .A2(new_n690), .ZN(new_n922));
  OAI211_X1 g0722(.A(new_n517), .B(new_n524), .C1(new_n522), .C2(new_n675), .ZN(new_n923));
  OAI21_X1  g0723(.A(new_n923), .B1(new_n517), .B2(new_n675), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n677), .A2(new_n924), .ZN(new_n925));
  XOR2_X1   g0725(.A(new_n925), .B(KEYINPUT45), .Z(new_n926));
  OR3_X1    g0726(.A1(new_n677), .A2(new_n924), .A3(KEYINPUT104), .ZN(new_n927));
  OAI21_X1  g0727(.A(KEYINPUT104), .B1(new_n677), .B2(new_n924), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n927), .A2(KEYINPUT44), .A3(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  AOI21_X1  g0730(.A(KEYINPUT44), .B1(new_n927), .B2(new_n928), .ZN(new_n931));
  OR3_X1    g0731(.A1(new_n922), .A2(new_n930), .A3(new_n931), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n922), .B1(new_n930), .B2(new_n931), .ZN(new_n933));
  NAND2_X1  g0733(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  AND2_X1   g0734(.A1(new_n668), .A2(new_n676), .ZN(new_n935));
  INV_X1    g0735(.A(new_n676), .ZN(new_n936));
  AOI21_X1  g0736(.A(new_n935), .B1(new_n690), .B2(new_n936), .ZN(new_n937));
  OR2_X1    g0737(.A1(new_n685), .A2(new_n937), .ZN(new_n938));
  NAND2_X1  g0738(.A1(new_n685), .A2(new_n937), .ZN(new_n939));
  NAND2_X1  g0739(.A1(new_n938), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n726), .B1(new_n934), .B2(new_n940), .ZN(new_n941));
  XNOR2_X1  g0741(.A(new_n694), .B(KEYINPUT41), .ZN(new_n942));
  NAND2_X1  g0742(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n943), .A2(new_n729), .ZN(new_n944));
  NAND2_X1  g0744(.A1(new_n922), .A2(new_n924), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n935), .A2(new_n924), .ZN(new_n946));
  OR2_X1    g0746(.A1(new_n946), .A2(KEYINPUT42), .ZN(new_n947));
  INV_X1    g0747(.A(new_n524), .ZN(new_n948));
  OAI21_X1  g0748(.A(new_n517), .B1(new_n948), .B2(new_n591), .ZN(new_n949));
  AOI22_X1  g0749(.A1(new_n946), .A2(KEYINPUT42), .B1(new_n675), .B2(new_n949), .ZN(new_n950));
  OR2_X1    g0750(.A1(new_n538), .A2(new_n675), .ZN(new_n951));
  OR3_X1    g0751(.A1(new_n951), .A2(new_n657), .A3(new_n656), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n951), .A2(new_n557), .ZN(new_n953));
  NAND2_X1  g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  AOI22_X1  g0754(.A1(new_n947), .A2(new_n950), .B1(KEYINPUT43), .B2(new_n954), .ZN(new_n955));
  NOR2_X1   g0755(.A1(new_n954), .A2(KEYINPUT43), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  XNOR2_X1  g0757(.A(new_n945), .B(new_n957), .ZN(new_n958));
  NAND3_X1  g0758(.A1(new_n952), .A2(new_n738), .A3(new_n953), .ZN(new_n959));
  OAI22_X1  g0759(.A1(new_n773), .A2(new_n207), .B1(new_n763), .B2(new_n816), .ZN(new_n960));
  AOI211_X1 g0760(.A(new_n272), .B(new_n960), .C1(G150), .C2(new_n781), .ZN(new_n961));
  INV_X1    g0761(.A(new_n768), .ZN(new_n962));
  NAND2_X1  g0762(.A1(new_n962), .A2(G77), .ZN(new_n963));
  AOI22_X1  g0763(.A1(G68), .A2(new_n778), .B1(new_n760), .B2(G143), .ZN(new_n964));
  AOI22_X1  g0764(.A1(new_n755), .A2(G159), .B1(new_n788), .B2(G58), .ZN(new_n965));
  NAND4_X1  g0765(.A1(new_n961), .A2(new_n963), .A3(new_n964), .A4(new_n965), .ZN(new_n966));
  OAI22_X1  g0766(.A1(new_n761), .A2(new_n808), .B1(new_n211), .B2(new_n777), .ZN(new_n967));
  AOI21_X1  g0767(.A(new_n967), .B1(G97), .B2(new_n962), .ZN(new_n968));
  NAND2_X1  g0768(.A1(new_n774), .A2(G283), .ZN(new_n969));
  AOI22_X1  g0769(.A1(new_n781), .A2(G303), .B1(new_n764), .B2(G317), .ZN(new_n970));
  INV_X1    g0770(.A(new_n742), .ZN(new_n971));
  AOI21_X1  g0771(.A(new_n971), .B1(G294), .B2(new_n755), .ZN(new_n972));
  NAND4_X1  g0772(.A1(new_n968), .A2(new_n969), .A3(new_n970), .A4(new_n972), .ZN(new_n973));
  NOR2_X1   g0773(.A1(new_n758), .A2(new_n605), .ZN(new_n974));
  XNOR2_X1  g0774(.A(new_n974), .B(KEYINPUT46), .ZN(new_n975));
  OAI21_X1  g0775(.A(new_n966), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g0776(.A(KEYINPUT47), .ZN(new_n977));
  AND2_X1   g0777(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  NOR2_X1   g0778(.A1(new_n976), .A2(new_n977), .ZN(new_n979));
  NOR3_X1   g0779(.A1(new_n978), .A2(new_n979), .A3(new_n752), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n744), .A2(new_n242), .ZN(new_n981));
  AOI21_X1  g0781(.A(new_n741), .B1(new_n693), .B2(new_n419), .ZN(new_n982));
  AOI21_X1  g0782(.A(new_n734), .B1(new_n981), .B2(new_n982), .ZN(new_n983));
  XOR2_X1   g0783(.A(new_n983), .B(KEYINPUT105), .Z(new_n984));
  NOR2_X1   g0784(.A1(new_n980), .A2(new_n984), .ZN(new_n985));
  XOR2_X1   g0785(.A(new_n985), .B(KEYINPUT106), .Z(new_n986));
  AOI22_X1  g0786(.A1(new_n944), .A2(new_n958), .B1(new_n959), .B2(new_n986), .ZN(new_n987));
  INV_X1    g0787(.A(new_n987), .ZN(G387));
  INV_X1    g0788(.A(new_n940), .ZN(new_n989));
  NAND2_X1  g0789(.A1(new_n989), .A2(new_n726), .ZN(new_n990));
  NAND2_X1  g0790(.A1(new_n940), .A2(new_n725), .ZN(new_n991));
  NAND3_X1  g0791(.A1(new_n990), .A2(new_n694), .A3(new_n991), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n761), .A2(new_n341), .B1(new_n420), .B2(new_n777), .ZN(new_n993));
  NOR2_X1   g0793(.A1(new_n758), .A2(new_n273), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n993), .A2(new_n994), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n769), .A2(G97), .ZN(new_n996));
  OAI22_X1  g0796(.A1(new_n773), .A2(new_n203), .B1(new_n763), .B2(new_n287), .ZN(new_n997));
  AOI21_X1  g0797(.A(new_n997), .B1(G50), .B2(new_n781), .ZN(new_n998));
  AOI21_X1  g0798(.A(new_n742), .B1(new_n335), .B2(new_n755), .ZN(new_n999));
  NAND4_X1  g0799(.A1(new_n995), .A2(new_n996), .A3(new_n998), .A4(new_n999), .ZN(new_n1000));
  AOI21_X1  g0800(.A(new_n971), .B1(G326), .B2(new_n764), .ZN(new_n1001));
  INV_X1    g0801(.A(G283), .ZN(new_n1002));
  OAI22_X1  g0802(.A1(new_n777), .A2(new_n1002), .B1(new_n758), .B2(new_n807), .ZN(new_n1003));
  AOI22_X1  g0803(.A1(new_n781), .A2(G317), .B1(new_n774), .B2(G303), .ZN(new_n1004));
  XOR2_X1   g0804(.A(KEYINPUT108), .B(G322), .Z(new_n1005));
  OAI221_X1 g0805(.A(new_n1004), .B1(new_n756), .B2(new_n808), .C1(new_n761), .C2(new_n1005), .ZN(new_n1006));
  INV_X1    g0806(.A(KEYINPUT48), .ZN(new_n1007));
  AOI21_X1  g0807(.A(new_n1003), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  OAI21_X1  g0808(.A(new_n1008), .B1(new_n1007), .B2(new_n1006), .ZN(new_n1009));
  INV_X1    g0809(.A(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n1001), .B1(new_n605), .B2(new_n768), .C1(new_n1009), .C2(new_n1010), .ZN(new_n1011));
  AND2_X1   g0811(.A1(new_n1009), .A2(new_n1010), .ZN(new_n1012));
  OAI21_X1  g0812(.A(new_n1000), .B1(new_n1011), .B2(new_n1012), .ZN(new_n1013));
  INV_X1    g0813(.A(KEYINPUT109), .ZN(new_n1014));
  AOI21_X1  g0814(.A(new_n752), .B1(new_n1013), .B2(new_n1014), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n1015), .B1(new_n1014), .B2(new_n1013), .ZN(new_n1016));
  AOI22_X1  g0816(.A1(new_n748), .A2(new_n699), .B1(new_n211), .B2(new_n693), .ZN(new_n1017));
  AOI211_X1 g0817(.A(G45), .B(new_n699), .C1(G68), .C2(G77), .ZN(new_n1018));
  NOR2_X1   g0818(.A1(new_n285), .A2(G50), .ZN(new_n1019));
  XNOR2_X1  g0819(.A(new_n1019), .B(KEYINPUT50), .ZN(new_n1020));
  NAND2_X1  g0820(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n1021), .A2(new_n744), .ZN(new_n1022));
  NOR2_X1   g0822(.A1(new_n239), .A2(new_n262), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1017), .B1(new_n1022), .B2(new_n1023), .ZN(new_n1024));
  INV_X1    g0824(.A(KEYINPUT107), .ZN(new_n1025));
  AND2_X1   g0825(.A1(new_n1024), .A2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n740), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1027));
  OAI211_X1 g0827(.A(new_n1016), .B(new_n804), .C1(new_n1026), .C2(new_n1027), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n690), .B2(new_n738), .ZN(new_n1029));
  AOI21_X1  g0829(.A(new_n1029), .B1(new_n989), .B2(new_n732), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n992), .A2(new_n1030), .ZN(G393));
  OR2_X1    g0831(.A1(new_n934), .A2(new_n990), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n934), .A2(new_n990), .ZN(new_n1033));
  NAND3_X1  g0833(.A1(new_n1032), .A2(new_n694), .A3(new_n1033), .ZN(new_n1034));
  NOR2_X1   g0834(.A1(new_n934), .A2(new_n729), .ZN(new_n1035));
  OR2_X1    g0835(.A1(new_n924), .A2(new_n793), .ZN(new_n1036));
  NAND2_X1  g0836(.A1(new_n744), .A2(new_n246), .ZN(new_n1037));
  OAI211_X1 g0837(.A(new_n1037), .B(new_n740), .C1(new_n210), .C2(new_n218), .ZN(new_n1038));
  AOI22_X1  g0838(.A1(G116), .A2(new_n778), .B1(new_n755), .B2(G303), .ZN(new_n1039));
  INV_X1    g0839(.A(KEYINPUT111), .ZN(new_n1040));
  OAI22_X1  g0840(.A1(new_n1039), .A2(new_n1040), .B1(new_n807), .B2(new_n773), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(G317), .A2(new_n760), .B1(new_n781), .B2(G311), .ZN(new_n1042));
  XNOR2_X1  g0842(.A(new_n1042), .B(KEYINPUT52), .ZN(new_n1043));
  AOI211_X1 g0843(.A(new_n1041), .B(new_n1043), .C1(new_n1040), .C2(new_n1039), .ZN(new_n1044));
  INV_X1    g0844(.A(new_n1005), .ZN(new_n1045));
  AOI21_X1  g0845(.A(new_n275), .B1(new_n1045), .B2(new_n764), .ZN(new_n1046));
  OAI211_X1 g0846(.A(new_n770), .B(new_n1046), .C1(new_n1002), .C2(new_n758), .ZN(new_n1047));
  XOR2_X1   g0847(.A(new_n1047), .B(KEYINPUT110), .Z(new_n1048));
  OAI22_X1  g0848(.A1(new_n761), .A2(new_n287), .B1(new_n341), .B2(new_n771), .ZN(new_n1049));
  XNOR2_X1  g0849(.A(new_n1049), .B(KEYINPUT51), .ZN(new_n1050));
  AOI22_X1  g0850(.A1(new_n335), .A2(new_n774), .B1(new_n764), .B2(G143), .ZN(new_n1051));
  NAND2_X1  g0851(.A1(new_n1051), .A2(new_n971), .ZN(new_n1052));
  NAND2_X1  g0852(.A1(new_n778), .A2(G77), .ZN(new_n1053));
  OAI221_X1 g0853(.A(new_n1053), .B1(new_n203), .B2(new_n758), .C1(new_n756), .C2(new_n207), .ZN(new_n1054));
  AOI211_X1 g0854(.A(new_n1052), .B(new_n1054), .C1(G87), .C2(new_n769), .ZN(new_n1055));
  AOI22_X1  g0855(.A1(new_n1044), .A2(new_n1048), .B1(new_n1050), .B2(new_n1055), .ZN(new_n1056));
  OAI211_X1 g0856(.A(new_n804), .B(new_n1038), .C1(new_n1056), .C2(new_n752), .ZN(new_n1057));
  XOR2_X1   g0857(.A(new_n1057), .B(KEYINPUT112), .Z(new_n1058));
  AOI21_X1  g0858(.A(new_n1035), .B1(new_n1036), .B2(new_n1058), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1034), .A2(new_n1059), .ZN(G390));
  NOR2_X1   g0860(.A1(new_n702), .A2(new_n703), .ZN(new_n1061));
  NOR2_X1   g0861(.A1(new_n1061), .A2(new_n674), .ZN(new_n1062));
  AOI21_X1  g0862(.A(new_n885), .B1(new_n1062), .B2(new_n800), .ZN(new_n1063));
  INV_X1    g0863(.A(new_n893), .ZN(new_n1064));
  OAI211_X1 g0864(.A(new_n877), .B(new_n874), .C1(new_n1063), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n878), .B1(new_n888), .B2(new_n893), .ZN(new_n1066));
  AOI21_X1  g0866(.A(new_n882), .B1(new_n874), .B2(new_n875), .ZN(new_n1067));
  OAI21_X1  g0867(.A(new_n1065), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g0868(.A(G330), .ZN(new_n1069));
  NOR2_X1   g0869(.A1(new_n799), .A2(new_n1069), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n913), .A2(new_n1070), .ZN(new_n1071));
  NOR2_X1   g0871(.A1(new_n1071), .A2(new_n1064), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1068), .A2(new_n1072), .ZN(new_n1073));
  NAND3_X1  g0873(.A1(new_n893), .A2(new_n1070), .A3(new_n723), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1065), .B(new_n1074), .C1(new_n1066), .C2(new_n1067), .ZN(new_n1075));
  NAND2_X1  g0875(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  OR3_X1    g0876(.A1(new_n1076), .A2(KEYINPUT116), .A3(new_n729), .ZN(new_n1077));
  OAI21_X1  g0877(.A(KEYINPUT116), .B1(new_n1076), .B2(new_n729), .ZN(new_n1078));
  NAND2_X1  g0878(.A1(new_n1077), .A2(new_n1078), .ZN(new_n1079));
  NAND4_X1  g0879(.A1(new_n901), .A2(new_n478), .A3(G330), .A4(new_n903), .ZN(new_n1080));
  XNOR2_X1  g0880(.A(new_n1080), .B(KEYINPUT113), .ZN(new_n1081));
  AND3_X1   g0881(.A1(new_n1081), .A2(KEYINPUT114), .A3(new_n898), .ZN(new_n1082));
  AOI21_X1  g0882(.A(KEYINPUT114), .B1(new_n1081), .B2(new_n898), .ZN(new_n1083));
  NOR2_X1   g0883(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1084));
  AOI21_X1  g0884(.A(new_n893), .B1(new_n723), .B2(new_n1070), .ZN(new_n1085));
  OR2_X1    g0885(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1086));
  NAND2_X1  g0886(.A1(new_n1085), .A2(KEYINPUT115), .ZN(new_n1087));
  NAND2_X1  g0887(.A1(new_n1086), .A2(new_n1087), .ZN(new_n1088));
  OAI21_X1  g0888(.A(new_n888), .B1(new_n1088), .B2(new_n1072), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1071), .A2(new_n1064), .ZN(new_n1090));
  NAND3_X1  g0890(.A1(new_n1090), .A2(new_n1074), .A3(new_n1063), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1089), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g0893(.A1(new_n1093), .A2(new_n1076), .ZN(new_n1094));
  NAND4_X1  g0894(.A1(new_n1084), .A2(new_n1075), .A3(new_n1073), .A4(new_n1092), .ZN(new_n1095));
  NAND3_X1  g0895(.A1(new_n1094), .A2(new_n694), .A3(new_n1095), .ZN(new_n1096));
  OAI221_X1 g0896(.A(new_n272), .B1(new_n763), .B2(new_n807), .C1(new_n771), .C2(new_n605), .ZN(new_n1097));
  OAI21_X1  g0897(.A(new_n1053), .B1(new_n373), .B2(new_n758), .ZN(new_n1098));
  AOI211_X1 g0898(.A(new_n1097), .B(new_n1098), .C1(G283), .C2(new_n760), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n756), .A2(new_n211), .B1(new_n773), .B2(new_n210), .ZN(new_n1100));
  NAND2_X1  g0900(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1101));
  OR2_X1    g0901(.A1(new_n1100), .A2(KEYINPUT117), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1099), .A2(new_n820), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  OR2_X1    g0903(.A1(new_n1103), .A2(KEYINPUT118), .ZN(new_n1104));
  AOI22_X1  g0904(.A1(new_n781), .A2(G132), .B1(new_n764), .B2(G125), .ZN(new_n1105));
  OAI21_X1  g0905(.A(KEYINPUT53), .B1(new_n758), .B2(new_n287), .ZN(new_n1106));
  XNOR2_X1  g0906(.A(KEYINPUT54), .B(G143), .ZN(new_n1107));
  INV_X1    g0907(.A(new_n1107), .ZN(new_n1108));
  AOI21_X1  g0908(.A(new_n272), .B1(new_n774), .B2(new_n1108), .ZN(new_n1109));
  NAND3_X1  g0909(.A1(new_n1105), .A2(new_n1106), .A3(new_n1109), .ZN(new_n1110));
  OAI22_X1  g0910(.A1(new_n756), .A2(new_n816), .B1(new_n207), .B2(new_n768), .ZN(new_n1111));
  INV_X1    g0911(.A(G128), .ZN(new_n1112));
  OAI22_X1  g0912(.A1(new_n761), .A2(new_n1112), .B1(new_n341), .B2(new_n777), .ZN(new_n1113));
  NOR3_X1   g0913(.A1(new_n758), .A2(KEYINPUT53), .A3(new_n287), .ZN(new_n1114));
  NOR4_X1   g0914(.A1(new_n1110), .A2(new_n1111), .A3(new_n1113), .A4(new_n1114), .ZN(new_n1115));
  AOI21_X1  g0915(.A(new_n1115), .B1(new_n1103), .B2(KEYINPUT118), .ZN(new_n1116));
  AOI21_X1  g0916(.A(new_n752), .B1(new_n1104), .B2(new_n1116), .ZN(new_n1117));
  AOI211_X1 g0917(.A(new_n734), .B(new_n1117), .C1(new_n285), .C2(new_n827), .ZN(new_n1118));
  XOR2_X1   g0918(.A(new_n1118), .B(KEYINPUT119), .Z(new_n1119));
  OAI21_X1  g0919(.A(new_n1119), .B1(new_n1067), .B2(new_n737), .ZN(new_n1120));
  NAND3_X1  g0920(.A1(new_n1079), .A2(new_n1096), .A3(new_n1120), .ZN(G378));
  NOR2_X1   g0921(.A1(new_n308), .A2(new_n672), .ZN(new_n1122));
  INV_X1    g0922(.A(new_n1122), .ZN(new_n1123));
  XNOR2_X1  g0923(.A(new_n331), .B(new_n1123), .ZN(new_n1124));
  XNOR2_X1  g0924(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1125));
  XNOR2_X1  g0925(.A(new_n1124), .B(new_n1125), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1126), .A2(new_n736), .ZN(new_n1127));
  AOI21_X1  g0927(.A(new_n734), .B1(new_n207), .B2(new_n827), .ZN(new_n1128));
  XOR2_X1   g0928(.A(new_n1128), .B(KEYINPUT121), .Z(new_n1129));
  NOR2_X1   g0929(.A1(new_n971), .A2(new_n493), .ZN(new_n1130));
  NOR2_X1   g0930(.A1(G33), .A2(G41), .ZN(new_n1131));
  XNOR2_X1  g0931(.A(new_n1131), .B(KEYINPUT120), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1132), .ZN(new_n1133));
  NOR3_X1   g0933(.A1(new_n1130), .A2(G50), .A3(new_n1133), .ZN(new_n1134));
  AOI22_X1  g0934(.A1(new_n781), .A2(G107), .B1(new_n764), .B2(G283), .ZN(new_n1135));
  OAI21_X1  g0935(.A(new_n1135), .B1(new_n420), .B2(new_n773), .ZN(new_n1136));
  AOI211_X1 g0936(.A(new_n994), .B(new_n1136), .C1(G68), .C2(new_n778), .ZN(new_n1137));
  OAI22_X1  g0937(.A1(new_n761), .A2(new_n605), .B1(new_n202), .B2(new_n768), .ZN(new_n1138));
  AOI21_X1  g0938(.A(new_n1138), .B1(G97), .B2(new_n755), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1137), .A2(new_n1139), .A3(new_n1130), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT58), .ZN(new_n1141));
  AOI21_X1  g0941(.A(new_n1134), .B1(new_n1140), .B2(new_n1141), .ZN(new_n1142));
  AOI21_X1  g0942(.A(new_n1132), .B1(G124), .B2(new_n764), .ZN(new_n1143));
  OAI22_X1  g0943(.A1(new_n771), .A2(new_n1112), .B1(new_n773), .B2(new_n816), .ZN(new_n1144));
  AOI22_X1  g0944(.A1(new_n755), .A2(G132), .B1(new_n788), .B2(new_n1108), .ZN(new_n1145));
  INV_X1    g0945(.A(G125), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n1145), .B1(new_n1146), .B2(new_n761), .ZN(new_n1147));
  AOI211_X1 g0947(.A(new_n1144), .B(new_n1147), .C1(G150), .C2(new_n778), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT59), .ZN(new_n1149));
  OAI221_X1 g0949(.A(new_n1143), .B1(new_n341), .B2(new_n768), .C1(new_n1148), .C2(new_n1149), .ZN(new_n1150));
  INV_X1    g0950(.A(new_n1148), .ZN(new_n1151));
  NOR2_X1   g0951(.A1(new_n1151), .A2(KEYINPUT59), .ZN(new_n1152));
  OAI221_X1 g0952(.A(new_n1142), .B1(new_n1141), .B2(new_n1140), .C1(new_n1150), .C2(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1129), .B1(new_n1153), .B2(new_n739), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1127), .A2(new_n1154), .ZN(new_n1155));
  INV_X1    g0955(.A(new_n896), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1069), .B1(new_n909), .B2(new_n910), .ZN(new_n1157));
  INV_X1    g0957(.A(new_n1126), .ZN(new_n1158));
  NAND3_X1  g0958(.A1(new_n908), .A2(new_n1157), .A3(new_n1158), .ZN(new_n1159));
  INV_X1    g0959(.A(KEYINPUT122), .ZN(new_n1160));
  NAND2_X1  g0960(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  NAND4_X1  g0961(.A1(new_n908), .A2(new_n1157), .A3(KEYINPUT122), .A4(new_n1158), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n1161), .A2(new_n1162), .ZN(new_n1163));
  AOI21_X1  g0963(.A(new_n1158), .B1(new_n908), .B2(new_n1157), .ZN(new_n1164));
  INV_X1    g0964(.A(new_n1164), .ZN(new_n1165));
  AOI21_X1  g0965(.A(new_n1156), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1166));
  NOR2_X1   g0966(.A1(new_n896), .A2(new_n1164), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1163), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT123), .ZN(new_n1169));
  INV_X1    g0969(.A(KEYINPUT123), .ZN(new_n1170));
  NAND3_X1  g0970(.A1(new_n1163), .A2(new_n1167), .A3(new_n1170), .ZN(new_n1171));
  AOI21_X1  g0971(.A(new_n1166), .B1(new_n1169), .B2(new_n1171), .ZN(new_n1172));
  OAI21_X1  g0972(.A(new_n1155), .B1(new_n1172), .B2(new_n729), .ZN(new_n1173));
  NAND2_X1  g0973(.A1(new_n1173), .A2(KEYINPUT124), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1175), .A2(new_n896), .ZN(new_n1176));
  AND3_X1   g0976(.A1(new_n1163), .A2(new_n1170), .A3(new_n1167), .ZN(new_n1177));
  AOI21_X1  g0977(.A(new_n1170), .B1(new_n1163), .B2(new_n1167), .ZN(new_n1178));
  OAI21_X1  g0978(.A(new_n1176), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1179), .A2(new_n732), .ZN(new_n1180));
  INV_X1    g0980(.A(KEYINPUT124), .ZN(new_n1181));
  NAND3_X1  g0981(.A1(new_n1180), .A2(new_n1181), .A3(new_n1155), .ZN(new_n1182));
  INV_X1    g0982(.A(KEYINPUT57), .ZN(new_n1183));
  AND2_X1   g0983(.A1(new_n1095), .A2(new_n1084), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1183), .B1(new_n1172), .B2(new_n1184), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1183), .B1(new_n1095), .B2(new_n1084), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1176), .A2(new_n1168), .ZN(new_n1187));
  AOI21_X1  g0987(.A(new_n696), .B1(new_n1186), .B2(new_n1187), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n1174), .A2(new_n1182), .B1(new_n1185), .B2(new_n1188), .ZN(new_n1189));
  INV_X1    g0989(.A(new_n1189), .ZN(G375));
  NAND2_X1  g0990(.A1(new_n1064), .A2(new_n736), .ZN(new_n1191));
  OAI22_X1  g0991(.A1(new_n771), .A2(new_n1002), .B1(new_n773), .B2(new_n211), .ZN(new_n1192));
  AOI211_X1 g0992(.A(new_n275), .B(new_n1192), .C1(G303), .C2(new_n764), .ZN(new_n1193));
  NAND2_X1  g0993(.A1(new_n769), .A2(G77), .ZN(new_n1194));
  AOI22_X1  g0994(.A1(new_n419), .A2(new_n778), .B1(new_n755), .B2(G116), .ZN(new_n1195));
  AOI22_X1  g0995(.A1(new_n760), .A2(G294), .B1(new_n788), .B2(G97), .ZN(new_n1196));
  NAND4_X1  g0996(.A1(new_n1193), .A2(new_n1194), .A3(new_n1195), .A4(new_n1196), .ZN(new_n1197));
  OAI22_X1  g0997(.A1(new_n771), .A2(new_n816), .B1(new_n763), .B2(new_n1112), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n1198), .B1(G150), .B2(new_n774), .ZN(new_n1199));
  AOI21_X1  g0999(.A(new_n742), .B1(G58), .B2(new_n962), .ZN(new_n1200));
  AOI22_X1  g1000(.A1(new_n755), .A2(new_n1108), .B1(new_n788), .B2(G159), .ZN(new_n1201));
  AOI22_X1  g1001(.A1(G50), .A2(new_n778), .B1(new_n760), .B2(G132), .ZN(new_n1202));
  NAND4_X1  g1002(.A1(new_n1199), .A2(new_n1200), .A3(new_n1201), .A4(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n752), .B1(new_n1197), .B2(new_n1203), .ZN(new_n1204));
  AOI211_X1 g1004(.A(new_n734), .B(new_n1204), .C1(new_n203), .C2(new_n827), .ZN(new_n1205));
  AOI22_X1  g1005(.A1(new_n1092), .A2(new_n732), .B1(new_n1191), .B2(new_n1205), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1093), .A2(new_n942), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1084), .A2(new_n1092), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1206), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  INV_X1    g1009(.A(G378), .ZN(new_n1210));
  NAND2_X1  g1010(.A1(new_n1189), .A2(new_n1210), .ZN(new_n1211));
  INV_X1    g1011(.A(G384), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n992), .A2(new_n795), .A3(new_n1030), .ZN(new_n1213));
  INV_X1    g1013(.A(new_n1213), .ZN(new_n1214));
  NAND4_X1  g1014(.A1(new_n1034), .A2(new_n1059), .A3(new_n1212), .A4(new_n1214), .ZN(new_n1215));
  OR4_X1    g1015(.A1(G387), .A2(new_n1211), .A3(G381), .A4(new_n1215), .ZN(G407));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G343), .C2(new_n1211), .ZN(G409));
  NAND2_X1  g1017(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n1181), .B1(new_n1180), .B2(new_n1155), .ZN(new_n1219));
  INV_X1    g1019(.A(new_n1155), .ZN(new_n1220));
  AOI211_X1 g1020(.A(KEYINPUT124), .B(new_n1220), .C1(new_n1179), .C2(new_n732), .ZN(new_n1221));
  OAI211_X1 g1021(.A(G378), .B(new_n1218), .C1(new_n1219), .C2(new_n1221), .ZN(new_n1222));
  INV_X1    g1022(.A(new_n1184), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1223), .A2(new_n942), .A3(new_n1179), .ZN(new_n1224));
  AOI21_X1  g1024(.A(new_n1220), .B1(new_n1187), .B2(new_n732), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1224), .A2(new_n1225), .ZN(new_n1226));
  NAND2_X1  g1026(.A1(new_n1226), .A2(new_n1210), .ZN(new_n1227));
  NAND2_X1  g1027(.A1(new_n1222), .A2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n673), .A2(G213), .ZN(new_n1229));
  AOI21_X1  g1029(.A(new_n1208), .B1(KEYINPUT60), .B2(new_n1093), .ZN(new_n1230));
  OR2_X1    g1030(.A1(new_n1082), .A2(new_n1083), .ZN(new_n1231));
  INV_X1    g1031(.A(new_n1092), .ZN(new_n1232));
  NAND3_X1  g1032(.A1(new_n1231), .A2(KEYINPUT60), .A3(new_n1232), .ZN(new_n1233));
  NAND2_X1  g1033(.A1(new_n1233), .A2(new_n694), .ZN(new_n1234));
  OAI21_X1  g1034(.A(new_n1206), .B1(new_n1230), .B2(new_n1234), .ZN(new_n1235));
  OR2_X1    g1035(.A1(new_n1212), .A2(KEYINPUT125), .ZN(new_n1236));
  NAND2_X1  g1036(.A1(new_n1212), .A2(KEYINPUT125), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1235), .A2(new_n1236), .A3(new_n1237), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1093), .A2(KEYINPUT60), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1231), .A2(new_n1232), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1239), .A2(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(new_n694), .A3(new_n1233), .ZN(new_n1242));
  NAND4_X1  g1042(.A1(new_n1242), .A2(KEYINPUT125), .A3(new_n1212), .A4(new_n1206), .ZN(new_n1243));
  NAND2_X1  g1043(.A1(new_n1238), .A2(new_n1243), .ZN(new_n1244));
  NAND3_X1  g1044(.A1(new_n1228), .A2(new_n1229), .A3(new_n1244), .ZN(new_n1245));
  NAND2_X1  g1045(.A1(new_n1245), .A2(KEYINPUT62), .ZN(new_n1246));
  INV_X1    g1046(.A(KEYINPUT61), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1229), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1248), .A2(KEYINPUT126), .A3(G2897), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(KEYINPUT126), .B1(new_n1248), .B2(G2897), .ZN(new_n1251));
  NOR2_X1   g1051(.A1(new_n1250), .A2(new_n1251), .ZN(new_n1252));
  NAND3_X1  g1052(.A1(new_n1238), .A2(new_n1243), .A3(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1244), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1254), .B2(new_n1249), .ZN(new_n1255));
  AOI21_X1  g1055(.A(G378), .B1(new_n1224), .B2(new_n1225), .ZN(new_n1256));
  AOI21_X1  g1056(.A(new_n1256), .B1(new_n1189), .B2(G378), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1255), .B1(new_n1257), .B2(new_n1248), .ZN(new_n1258));
  AOI21_X1  g1058(.A(new_n1248), .B1(new_n1222), .B2(new_n1227), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT62), .ZN(new_n1260));
  NAND3_X1  g1060(.A1(new_n1259), .A2(new_n1260), .A3(new_n1244), .ZN(new_n1261));
  NAND4_X1  g1061(.A1(new_n1246), .A2(new_n1247), .A3(new_n1258), .A4(new_n1261), .ZN(new_n1262));
  XNOR2_X1  g1062(.A(G393), .B(new_n795), .ZN(new_n1263));
  OR2_X1    g1063(.A1(new_n1263), .A2(G390), .ZN(new_n1264));
  NAND2_X1  g1064(.A1(new_n1263), .A2(G390), .ZN(new_n1265));
  AND3_X1   g1065(.A1(new_n1264), .A2(new_n987), .A3(new_n1265), .ZN(new_n1266));
  AOI21_X1  g1066(.A(new_n987), .B1(new_n1264), .B2(new_n1265), .ZN(new_n1267));
  NOR2_X1   g1067(.A1(new_n1266), .A2(new_n1267), .ZN(new_n1268));
  INV_X1    g1068(.A(new_n1268), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1262), .A2(new_n1269), .ZN(new_n1270));
  AND3_X1   g1070(.A1(new_n1238), .A2(new_n1243), .A3(new_n1252), .ZN(new_n1271));
  AOI21_X1  g1071(.A(new_n1249), .B1(new_n1238), .B2(new_n1243), .ZN(new_n1272));
  NOR2_X1   g1072(.A1(new_n1271), .A2(new_n1272), .ZN(new_n1273));
  OAI211_X1 g1073(.A(new_n1247), .B(new_n1268), .C1(new_n1259), .C2(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  INV_X1    g1075(.A(KEYINPUT63), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1245), .A2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(KEYINPUT127), .ZN(new_n1278));
  OAI21_X1  g1078(.A(new_n1278), .B1(new_n1245), .B2(new_n1276), .ZN(new_n1279));
  NAND4_X1  g1079(.A1(new_n1259), .A2(KEYINPUT127), .A3(KEYINPUT63), .A4(new_n1244), .ZN(new_n1280));
  NAND4_X1  g1080(.A1(new_n1275), .A2(new_n1277), .A3(new_n1279), .A4(new_n1280), .ZN(new_n1281));
  NAND2_X1  g1081(.A1(new_n1270), .A2(new_n1281), .ZN(G405));
  NAND2_X1  g1082(.A1(G375), .A2(new_n1210), .ZN(new_n1283));
  NAND3_X1  g1083(.A1(new_n1283), .A2(new_n1222), .A3(new_n1244), .ZN(new_n1284));
  NOR2_X1   g1084(.A1(new_n1189), .A2(G378), .ZN(new_n1285));
  INV_X1    g1085(.A(new_n1222), .ZN(new_n1286));
  OAI21_X1  g1086(.A(new_n1254), .B1(new_n1285), .B2(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1284), .A2(new_n1287), .ZN(new_n1288));
  XNOR2_X1  g1088(.A(new_n1288), .B(new_n1268), .ZN(G402));
endmodule


