

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
         n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600,
         n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611,
         n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
         n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633,
         n634, n635, n636, n637, n638, n639, n640, n641, n642, n643, n644,
         n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655,
         n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, n666,
         n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677,
         n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
         n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699,
         n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710,
         n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
         n722, n723, n724, n725, n726;

  INV_X1 U370 ( .A(G953), .ZN(n717) );
  AND2_X1 U371 ( .A1(n545), .A2(n512), .ZN(n513) );
  INV_X1 U372 ( .A(n554), .ZN(n447) );
  XNOR2_X2 U373 ( .A(n513), .B(KEYINPUT108), .ZN(n726) );
  XNOR2_X2 U374 ( .A(n423), .B(KEYINPUT4), .ZN(n708) );
  XNOR2_X2 U375 ( .A(KEYINPUT64), .B(KEYINPUT68), .ZN(n423) );
  NOR2_X1 U376 ( .A1(n581), .A2(n654), .ZN(n561) );
  XNOR2_X1 U377 ( .A(n527), .B(n526), .ZN(n606) );
  NOR2_X1 U378 ( .A1(n649), .A2(n654), .ZN(n556) );
  NOR2_X1 U379 ( .A1(n641), .A2(n640), .ZN(n535) );
  INV_X1 U380 ( .A(n519), .ZN(n640) );
  NAND2_X1 U381 ( .A1(n409), .A2(n357), .ZN(n408) );
  OR2_X1 U382 ( .A1(n715), .A2(n693), .ZN(n409) );
  XNOR2_X1 U383 ( .A(n715), .B(n593), .ZN(n358) );
  NOR2_X2 U384 ( .A1(n348), .A2(n362), .ZN(n548) );
  XNOR2_X1 U385 ( .A(n394), .B(KEYINPUT22), .ZN(n517) );
  XNOR2_X1 U386 ( .A(n542), .B(KEYINPUT105), .ZN(n626) );
  XNOR2_X1 U387 ( .A(G478), .B(n480), .ZN(n541) );
  NOR2_X1 U388 ( .A1(n517), .A2(n519), .ZN(n545) );
  NOR2_X1 U389 ( .A1(n549), .A2(G900), .ZN(n550) );
  NOR2_X1 U390 ( .A1(n723), .A2(n725), .ZN(n563) );
  XNOR2_X1 U391 ( .A(KEYINPUT67), .B(G101), .ZN(n424) );
  XNOR2_X1 U392 ( .A(n474), .B(n465), .ZN(n709) );
  XNOR2_X1 U393 ( .A(n709), .B(G146), .ZN(n491) );
  NOR2_X1 U394 ( .A1(n379), .A2(n559), .ZN(n572) );
  NAND2_X1 U395 ( .A1(n380), .A2(n635), .ZN(n379) );
  XNOR2_X1 U396 ( .A(n360), .B(n359), .ZN(n653) );
  INV_X1 U397 ( .A(KEYINPUT107), .ZN(n359) );
  NOR2_X1 U398 ( .A1(n541), .A2(n539), .ZN(n360) );
  INV_X1 U399 ( .A(n724), .ZN(n398) );
  XNOR2_X1 U400 ( .A(n377), .B(KEYINPUT81), .ZN(n559) );
  NAND2_X1 U401 ( .A1(n349), .A2(n378), .ZN(n377) );
  INV_X1 U402 ( .A(n551), .ZN(n378) );
  XNOR2_X1 U403 ( .A(n632), .B(KEYINPUT85), .ZN(n367) );
  AND2_X1 U404 ( .A1(n570), .A2(n361), .ZN(n368) );
  XNOR2_X1 U405 ( .A(n433), .B(n402), .ZN(n474) );
  INV_X1 U406 ( .A(G134), .ZN(n402) );
  NOR2_X1 U407 ( .A1(G953), .A2(G237), .ZN(n483) );
  XOR2_X1 U408 ( .A(KEYINPUT101), .B(KEYINPUT12), .Z(n417) );
  XNOR2_X1 U409 ( .A(n420), .B(n419), .ZN(n421) );
  INV_X1 U410 ( .A(KEYINPUT79), .ZN(n419) );
  XOR2_X1 U411 ( .A(G137), .B(G140), .Z(n493) );
  XNOR2_X1 U412 ( .A(n489), .B(n426), .ZN(n440) );
  XNOR2_X1 U413 ( .A(n403), .B(G128), .ZN(n433) );
  INV_X1 U414 ( .A(G143), .ZN(n403) );
  NAND2_X1 U415 ( .A1(n387), .A2(n385), .ZN(n564) );
  AND2_X1 U416 ( .A1(n390), .A2(n388), .ZN(n387) );
  NAND2_X1 U417 ( .A1(n447), .A2(n386), .ZN(n385) );
  XNOR2_X1 U418 ( .A(n370), .B(n491), .ZN(n608) );
  XNOR2_X1 U419 ( .A(n381), .B(KEYINPUT112), .ZN(n565) );
  NAND2_X1 U420 ( .A1(n383), .A2(n382), .ZN(n381) );
  XNOR2_X1 U421 ( .A(n552), .B(KEYINPUT28), .ZN(n383) );
  XNOR2_X1 U422 ( .A(n468), .B(n467), .ZN(n682) );
  XNOR2_X1 U423 ( .A(n415), .B(n466), .ZN(n467) );
  AND2_X1 U424 ( .A1(n350), .A2(n569), .ZN(n361) );
  INV_X1 U425 ( .A(n594), .ZN(n410) );
  NAND2_X1 U426 ( .A1(n374), .A2(G953), .ZN(n549) );
  XNOR2_X1 U427 ( .A(n376), .B(n375), .ZN(n374) );
  INV_X1 U428 ( .A(KEYINPUT92), .ZN(n375) );
  XNOR2_X1 U429 ( .A(KEYINPUT15), .B(G902), .ZN(n594) );
  INV_X1 U430 ( .A(n651), .ZN(n389) );
  NOR2_X1 U431 ( .A1(n449), .A2(n389), .ZN(n386) );
  NAND2_X1 U432 ( .A1(KEYINPUT65), .A2(KEYINPUT44), .ZN(n396) );
  XNOR2_X1 U433 ( .A(n384), .B(n431), .ZN(n487) );
  XOR2_X1 U434 ( .A(KEYINPUT71), .B(G119), .Z(n431) );
  XNOR2_X1 U435 ( .A(n365), .B(G116), .ZN(n384) );
  XNOR2_X1 U436 ( .A(G113), .B(KEYINPUT3), .ZN(n365) );
  XOR2_X1 U437 ( .A(KEYINPUT10), .B(n457), .Z(n494) );
  NOR2_X1 U438 ( .A1(n693), .A2(n405), .ZN(n404) );
  NAND2_X1 U439 ( .A1(n410), .A2(n406), .ZN(n405) );
  INV_X1 U440 ( .A(KEYINPUT2), .ZN(n406) );
  XNOR2_X1 U441 ( .A(G146), .B(G125), .ZN(n456) );
  INV_X1 U442 ( .A(G237), .ZN(n442) );
  INV_X1 U443 ( .A(G902), .ZN(n443) );
  INV_X1 U444 ( .A(n559), .ZN(n414) );
  INV_X1 U445 ( .A(KEYINPUT1), .ZN(n430) );
  NAND2_X1 U446 ( .A1(n400), .A2(n592), .ZN(n715) );
  XNOR2_X1 U447 ( .A(n366), .B(n401), .ZN(n400) );
  INV_X1 U448 ( .A(KEYINPUT48), .ZN(n401) );
  XNOR2_X1 U449 ( .A(n487), .B(n432), .ZN(n702) );
  XNOR2_X1 U450 ( .A(KEYINPUT16), .B(G122), .ZN(n432) );
  XNOR2_X1 U451 ( .A(G116), .B(G107), .ZN(n471) );
  XOR2_X1 U452 ( .A(KEYINPUT7), .B(G122), .Z(n472) );
  XOR2_X1 U453 ( .A(KEYINPUT69), .B(G131), .Z(n465) );
  XNOR2_X1 U454 ( .A(G122), .B(KEYINPUT102), .ZN(n458) );
  XNOR2_X1 U455 ( .A(G143), .B(G113), .ZN(n463) );
  XOR2_X1 U456 ( .A(G140), .B(G104), .Z(n464) );
  XNOR2_X1 U457 ( .A(n363), .B(n491), .ZN(n674) );
  XNOR2_X1 U458 ( .A(n440), .B(n427), .ZN(n363) );
  XNOR2_X1 U459 ( .A(n373), .B(n574), .ZN(n586) );
  NOR2_X1 U460 ( .A1(n573), .A2(n626), .ZN(n373) );
  NOR2_X2 U461 ( .A1(n564), .A2(n453), .ZN(n455) );
  OR2_X1 U462 ( .A1(n608), .A2(G902), .ZN(n369) );
  OR2_X1 U463 ( .A1(n686), .A2(G902), .ZN(n480) );
  XNOR2_X1 U464 ( .A(n509), .B(n508), .ZN(n510) );
  NOR2_X1 U465 ( .A1(n689), .A2(G902), .ZN(n511) );
  XNOR2_X1 U466 ( .A(n557), .B(KEYINPUT42), .ZN(n723) );
  NOR2_X1 U467 ( .A1(n576), .A2(n640), .ZN(n632) );
  XNOR2_X1 U468 ( .A(n372), .B(n371), .ZN(n576) );
  INV_X1 U469 ( .A(KEYINPUT36), .ZN(n371) );
  NOR2_X1 U470 ( .A1(n586), .A2(n575), .ZN(n372) );
  NOR2_X1 U471 ( .A1(n685), .A2(n692), .ZN(n364) );
  NOR2_X1 U472 ( .A1(n600), .A2(n692), .ZN(n602) );
  AND2_X1 U473 ( .A1(n530), .A2(n529), .ZN(n348) );
  XNOR2_X1 U474 ( .A(KEYINPUT109), .B(n550), .ZN(n349) );
  XOR2_X1 U475 ( .A(n584), .B(KEYINPUT82), .Z(n350) );
  XOR2_X1 U476 ( .A(n536), .B(KEYINPUT93), .Z(n351) );
  AND2_X1 U477 ( .A1(n653), .A2(n635), .ZN(n352) );
  NOR2_X1 U478 ( .A1(n655), .A2(n654), .ZN(n353) );
  AND2_X1 U479 ( .A1(n547), .A2(n615), .ZN(n354) );
  AND2_X1 U480 ( .A1(n395), .A2(n398), .ZN(n355) );
  XNOR2_X1 U481 ( .A(KEYINPUT30), .B(KEYINPUT111), .ZN(n356) );
  AND2_X1 U482 ( .A1(n410), .A2(KEYINPUT2), .ZN(n357) );
  NAND2_X1 U483 ( .A1(n404), .A2(n358), .ZN(n407) );
  NAND2_X1 U484 ( .A1(n391), .A2(n354), .ZN(n362) );
  XNOR2_X1 U485 ( .A(n364), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U486 ( .A1(n368), .A2(n367), .ZN(n366) );
  XNOR2_X2 U487 ( .A(n369), .B(n492), .ZN(n558) );
  XNOR2_X1 U488 ( .A(n490), .B(n489), .ZN(n370) );
  NAND2_X1 U489 ( .A1(n451), .A2(G902), .ZN(n376) );
  INV_X1 U490 ( .A(n636), .ZN(n380) );
  NOR2_X1 U491 ( .A1(n664), .A2(n565), .ZN(n557) );
  INV_X1 U492 ( .A(n553), .ZN(n382) );
  NAND2_X1 U493 ( .A1(n447), .A2(n651), .ZN(n575) );
  NAND2_X1 U494 ( .A1(n449), .A2(n389), .ZN(n388) );
  NAND2_X1 U495 ( .A1(n554), .A2(n449), .ZN(n390) );
  NAND2_X1 U496 ( .A1(n355), .A2(n392), .ZN(n391) );
  NAND2_X1 U497 ( .A1(n393), .A2(n532), .ZN(n392) );
  NAND2_X1 U498 ( .A1(n606), .A2(n531), .ZN(n393) );
  NAND2_X2 U499 ( .A1(n408), .A2(n407), .ZN(n680) );
  NOR2_X2 U500 ( .A1(G902), .A2(n674), .ZN(n429) );
  XNOR2_X2 U501 ( .A(n521), .B(n520), .ZN(n665) );
  NAND2_X1 U502 ( .A1(n536), .A2(n352), .ZN(n394) );
  INV_X1 U503 ( .A(n726), .ZN(n395) );
  NAND2_X1 U504 ( .A1(n397), .A2(n396), .ZN(n528) );
  NAND2_X1 U505 ( .A1(n399), .A2(n398), .ZN(n397) );
  NOR2_X1 U506 ( .A1(n726), .A2(n531), .ZN(n399) );
  INV_X1 U507 ( .A(n409), .ZN(n634) );
  NAND2_X1 U508 ( .A1(n413), .A2(n411), .ZN(n581) );
  XNOR2_X1 U509 ( .A(n412), .B(n356), .ZN(n411) );
  NAND2_X1 U510 ( .A1(n558), .A2(n651), .ZN(n412) );
  AND2_X1 U511 ( .A1(n560), .A2(n414), .ZN(n413) );
  XNOR2_X2 U512 ( .A(n548), .B(KEYINPUT45), .ZN(n693) );
  XOR2_X1 U513 ( .A(n464), .B(n463), .Z(n415) );
  XOR2_X1 U514 ( .A(n454), .B(KEYINPUT0), .Z(n416) );
  XNOR2_X1 U515 ( .A(n421), .B(n493), .ZN(n422) );
  XNOR2_X1 U516 ( .A(n682), .B(n681), .ZN(n683) );
  NOR2_X1 U517 ( .A1(n558), .A2(n636), .ZN(n512) );
  INV_X1 U518 ( .A(G952), .ZN(n418) );
  AND2_X1 U519 ( .A1(n418), .A2(G953), .ZN(n692) );
  NAND2_X1 U520 ( .A1(n717), .A2(G227), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n422), .B(KEYINPUT94), .ZN(n427) );
  XNOR2_X1 U522 ( .A(n708), .B(n424), .ZN(n489) );
  XNOR2_X1 U523 ( .A(G110), .B(G107), .ZN(n425) );
  XNOR2_X1 U524 ( .A(n425), .B(G104), .ZN(n701) );
  XNOR2_X1 U525 ( .A(n701), .B(KEYINPUT73), .ZN(n426) );
  XNOR2_X1 U526 ( .A(KEYINPUT70), .B(G469), .ZN(n428) );
  XNOR2_X2 U527 ( .A(n429), .B(n428), .ZN(n553) );
  XNOR2_X2 U528 ( .A(n553), .B(n430), .ZN(n519) );
  XNOR2_X1 U529 ( .A(n456), .B(n433), .ZN(n438) );
  XOR2_X1 U530 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n435) );
  NAND2_X1 U531 ( .A1(G224), .A2(n717), .ZN(n434) );
  XNOR2_X1 U532 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U533 ( .A(n436), .B(KEYINPUT91), .ZN(n437) );
  XNOR2_X1 U534 ( .A(n438), .B(n437), .ZN(n439) );
  XNOR2_X1 U535 ( .A(n702), .B(n439), .ZN(n441) );
  XNOR2_X1 U536 ( .A(n441), .B(n440), .ZN(n595) );
  NAND2_X1 U537 ( .A1(n595), .A2(n594), .ZN(n445) );
  NAND2_X1 U538 ( .A1(n443), .A2(n442), .ZN(n446) );
  NAND2_X1 U539 ( .A1(n446), .A2(G210), .ZN(n444) );
  XNOR2_X2 U540 ( .A(n445), .B(n444), .ZN(n554) );
  NAND2_X1 U541 ( .A1(n446), .A2(G214), .ZN(n651) );
  XNOR2_X1 U542 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n448) );
  XNOR2_X1 U543 ( .A(n448), .B(KEYINPUT66), .ZN(n449) );
  NAND2_X1 U544 ( .A1(G234), .A2(G237), .ZN(n450) );
  XNOR2_X1 U545 ( .A(n450), .B(KEYINPUT14), .ZN(n451) );
  NOR2_X1 U546 ( .A1(n549), .A2(G898), .ZN(n452) );
  NAND2_X1 U547 ( .A1(G952), .A2(n451), .ZN(n663) );
  NOR2_X1 U548 ( .A1(n663), .A2(G953), .ZN(n551) );
  NOR2_X1 U549 ( .A1(n452), .A2(n551), .ZN(n453) );
  INV_X1 U550 ( .A(KEYINPUT88), .ZN(n454) );
  XNOR2_X2 U551 ( .A(n455), .B(n416), .ZN(n536) );
  INV_X1 U552 ( .A(n456), .ZN(n457) );
  INV_X1 U553 ( .A(n494), .ZN(n462) );
  XNOR2_X1 U554 ( .A(n417), .B(n458), .ZN(n460) );
  NAND2_X1 U555 ( .A1(G214), .A2(n483), .ZN(n459) );
  XNOR2_X1 U556 ( .A(n460), .B(n459), .ZN(n461) );
  XNOR2_X1 U557 ( .A(n462), .B(n461), .ZN(n468) );
  XNOR2_X1 U558 ( .A(n465), .B(KEYINPUT11), .ZN(n466) );
  NOR2_X1 U559 ( .A1(G902), .A2(n682), .ZN(n470) );
  XNOR2_X1 U560 ( .A(KEYINPUT13), .B(G475), .ZN(n469) );
  XNOR2_X1 U561 ( .A(n470), .B(n469), .ZN(n539) );
  XNOR2_X1 U562 ( .A(KEYINPUT9), .B(KEYINPUT104), .ZN(n479) );
  XNOR2_X1 U563 ( .A(n472), .B(n471), .ZN(n473) );
  XOR2_X1 U564 ( .A(n474), .B(n473), .Z(n477) );
  NAND2_X1 U565 ( .A1(G234), .A2(n717), .ZN(n475) );
  XOR2_X1 U566 ( .A(KEYINPUT8), .B(n475), .Z(n501) );
  NAND2_X1 U567 ( .A1(G217), .A2(n501), .ZN(n476) );
  XNOR2_X1 U568 ( .A(n477), .B(n476), .ZN(n478) );
  XNOR2_X1 U569 ( .A(n479), .B(n478), .ZN(n686) );
  NAND2_X1 U570 ( .A1(G234), .A2(n594), .ZN(n481) );
  XNOR2_X1 U571 ( .A(KEYINPUT20), .B(n481), .ZN(n505) );
  NAND2_X1 U572 ( .A1(n505), .A2(G221), .ZN(n482) );
  XOR2_X1 U573 ( .A(n482), .B(KEYINPUT21), .Z(n635) );
  XOR2_X1 U574 ( .A(KEYINPUT100), .B(KEYINPUT5), .Z(n485) );
  NAND2_X1 U575 ( .A1(n483), .A2(G210), .ZN(n484) );
  XNOR2_X1 U576 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X1 U577 ( .A(n486), .B(G137), .ZN(n488) );
  XNOR2_X1 U578 ( .A(n488), .B(n487), .ZN(n490) );
  XNOR2_X1 U579 ( .A(G472), .B(KEYINPUT74), .ZN(n492) );
  INV_X1 U580 ( .A(n558), .ZN(n639) );
  XOR2_X1 U581 ( .A(n494), .B(n493), .Z(n711) );
  XNOR2_X1 U582 ( .A(KEYINPUT96), .B(G110), .ZN(n496) );
  XNOR2_X1 U583 ( .A(G128), .B(G119), .ZN(n495) );
  XNOR2_X1 U584 ( .A(n496), .B(n495), .ZN(n500) );
  XOR2_X1 U585 ( .A(KEYINPUT24), .B(KEYINPUT95), .Z(n498) );
  XNOR2_X1 U586 ( .A(KEYINPUT23), .B(KEYINPUT72), .ZN(n497) );
  XNOR2_X1 U587 ( .A(n498), .B(n497), .ZN(n499) );
  XNOR2_X1 U588 ( .A(n500), .B(n499), .ZN(n503) );
  NAND2_X1 U589 ( .A1(G221), .A2(n501), .ZN(n502) );
  XNOR2_X1 U590 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U591 ( .A(n711), .B(n504), .ZN(n689) );
  NAND2_X1 U592 ( .A1(n505), .A2(G217), .ZN(n509) );
  XOR2_X1 U593 ( .A(KEYINPUT97), .B(KEYINPUT98), .Z(n507) );
  XNOR2_X1 U594 ( .A(KEYINPUT78), .B(KEYINPUT25), .ZN(n506) );
  XNOR2_X1 U595 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X2 U596 ( .A(n511), .B(n510), .ZN(n636) );
  XOR2_X1 U597 ( .A(n558), .B(KEYINPUT6), .Z(n571) );
  INV_X1 U598 ( .A(n571), .ZN(n544) );
  NAND2_X1 U599 ( .A1(n519), .A2(n544), .ZN(n514) );
  NOR2_X1 U600 ( .A1(n636), .A2(n514), .ZN(n515) );
  XOR2_X1 U601 ( .A(KEYINPUT80), .B(n515), .Z(n516) );
  NOR2_X1 U602 ( .A1(n517), .A2(n516), .ZN(n518) );
  XNOR2_X1 U603 ( .A(n518), .B(KEYINPUT32), .ZN(n724) );
  INV_X1 U604 ( .A(KEYINPUT65), .ZN(n532) );
  NAND2_X1 U605 ( .A1(n635), .A2(n636), .ZN(n641) );
  NAND2_X1 U606 ( .A1(n535), .A2(n571), .ZN(n521) );
  XNOR2_X1 U607 ( .A(KEYINPUT89), .B(KEYINPUT33), .ZN(n520) );
  INV_X1 U608 ( .A(n665), .ZN(n522) );
  NAND2_X1 U609 ( .A1(n522), .A2(n351), .ZN(n524) );
  INV_X1 U610 ( .A(KEYINPUT34), .ZN(n523) );
  XNOR2_X1 U611 ( .A(n524), .B(n523), .ZN(n525) );
  AND2_X1 U612 ( .A1(n539), .A2(n541), .ZN(n579) );
  NAND2_X1 U613 ( .A1(n525), .A2(n579), .ZN(n527) );
  XNOR2_X1 U614 ( .A(KEYINPUT83), .B(KEYINPUT35), .ZN(n526) );
  NAND2_X1 U615 ( .A1(n528), .A2(n606), .ZN(n530) );
  INV_X1 U616 ( .A(KEYINPUT44), .ZN(n531) );
  NAND2_X1 U617 ( .A1(n532), .A2(n531), .ZN(n529) );
  NOR2_X1 U618 ( .A1(n553), .A2(n641), .ZN(n560) );
  NAND2_X1 U619 ( .A1(n351), .A2(n560), .ZN(n533) );
  XNOR2_X1 U620 ( .A(n533), .B(KEYINPUT99), .ZN(n534) );
  NAND2_X1 U621 ( .A1(n534), .A2(n639), .ZN(n617) );
  AND2_X1 U622 ( .A1(n558), .A2(n535), .ZN(n646) );
  NAND2_X1 U623 ( .A1(n536), .A2(n646), .ZN(n538) );
  INV_X1 U624 ( .A(KEYINPUT31), .ZN(n537) );
  XNOR2_X1 U625 ( .A(n538), .B(n537), .ZN(n629) );
  NAND2_X1 U626 ( .A1(n617), .A2(n629), .ZN(n543) );
  XNOR2_X1 U627 ( .A(n539), .B(KEYINPUT103), .ZN(n540) );
  NAND2_X1 U628 ( .A1(n540), .A2(n541), .ZN(n630) );
  XNOR2_X1 U629 ( .A(KEYINPUT106), .B(n630), .ZN(n590) );
  NOR2_X1 U630 ( .A1(n541), .A2(n540), .ZN(n542) );
  NAND2_X1 U631 ( .A1(n590), .A2(n626), .ZN(n650) );
  NAND2_X1 U632 ( .A1(n543), .A2(n650), .ZN(n547) );
  AND2_X1 U633 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U634 ( .A1(n546), .A2(n636), .ZN(n615) );
  AND2_X1 U635 ( .A1(n558), .A2(n572), .ZN(n552) );
  NAND2_X1 U636 ( .A1(n653), .A2(n651), .ZN(n649) );
  INV_X1 U637 ( .A(KEYINPUT38), .ZN(n555) );
  XNOR2_X1 U638 ( .A(n554), .B(n555), .ZN(n654) );
  XNOR2_X1 U639 ( .A(n556), .B(KEYINPUT41), .ZN(n664) );
  XNOR2_X1 U640 ( .A(n561), .B(KEYINPUT39), .ZN(n589) );
  NOR2_X1 U641 ( .A1(n589), .A2(n626), .ZN(n562) );
  XNOR2_X1 U642 ( .A(n562), .B(KEYINPUT40), .ZN(n725) );
  XNOR2_X1 U643 ( .A(n563), .B(KEYINPUT46), .ZN(n570) );
  NOR2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n577) );
  INV_X1 U645 ( .A(n577), .ZN(n624) );
  INV_X1 U646 ( .A(n650), .ZN(n566) );
  NOR2_X1 U647 ( .A1(n566), .A2(KEYINPUT47), .ZN(n567) );
  XNOR2_X1 U648 ( .A(n567), .B(KEYINPUT75), .ZN(n568) );
  OR2_X1 U649 ( .A1(n624), .A2(n568), .ZN(n569) );
  NAND2_X1 U650 ( .A1(n572), .A2(n571), .ZN(n573) );
  INV_X1 U651 ( .A(KEYINPUT110), .ZN(n574) );
  NAND2_X1 U652 ( .A1(n577), .A2(n650), .ZN(n578) );
  NAND2_X1 U653 ( .A1(n578), .A2(KEYINPUT47), .ZN(n583) );
  INV_X1 U654 ( .A(n579), .ZN(n580) );
  NOR2_X1 U655 ( .A1(n581), .A2(n580), .ZN(n582) );
  NAND2_X1 U656 ( .A1(n582), .A2(n447), .ZN(n603) );
  NAND2_X1 U657 ( .A1(n583), .A2(n603), .ZN(n584) );
  NAND2_X1 U658 ( .A1(n651), .A2(n640), .ZN(n585) );
  NOR2_X1 U659 ( .A1(n586), .A2(n585), .ZN(n587) );
  XNOR2_X1 U660 ( .A(n587), .B(KEYINPUT43), .ZN(n588) );
  OR2_X1 U661 ( .A1(n588), .A2(n447), .ZN(n604) );
  NOR2_X1 U662 ( .A1(n590), .A2(n589), .ZN(n591) );
  XNOR2_X1 U663 ( .A(n591), .B(KEYINPUT113), .ZN(n721) );
  AND2_X1 U664 ( .A1(n604), .A2(n721), .ZN(n592) );
  INV_X1 U665 ( .A(KEYINPUT76), .ZN(n593) );
  NAND2_X1 U666 ( .A1(n680), .A2(G210), .ZN(n599) );
  XNOR2_X1 U667 ( .A(KEYINPUT55), .B(KEYINPUT54), .ZN(n596) );
  XOR2_X1 U668 ( .A(n596), .B(KEYINPUT87), .Z(n597) );
  XNOR2_X1 U669 ( .A(n595), .B(n597), .ZN(n598) );
  XNOR2_X1 U670 ( .A(n599), .B(n598), .ZN(n600) );
  XNOR2_X1 U671 ( .A(KEYINPUT84), .B(KEYINPUT56), .ZN(n601) );
  XNOR2_X1 U672 ( .A(n602), .B(n601), .ZN(G51) );
  XNOR2_X1 U673 ( .A(n603), .B(G143), .ZN(G45) );
  XNOR2_X1 U674 ( .A(n604), .B(G140), .ZN(G42) );
  XOR2_X1 U675 ( .A(G122), .B(KEYINPUT125), .Z(n605) );
  XNOR2_X1 U676 ( .A(n606), .B(n605), .ZN(G24) );
  NAND2_X1 U677 ( .A1(n680), .A2(G472), .ZN(n610) );
  XNOR2_X1 U678 ( .A(KEYINPUT114), .B(KEYINPUT62), .ZN(n607) );
  XNOR2_X1 U679 ( .A(n608), .B(n607), .ZN(n609) );
  XNOR2_X1 U680 ( .A(n610), .B(n609), .ZN(n611) );
  NOR2_X1 U681 ( .A1(n611), .A2(n692), .ZN(n614) );
  XNOR2_X1 U682 ( .A(KEYINPUT90), .B(KEYINPUT63), .ZN(n612) );
  XOR2_X1 U683 ( .A(n612), .B(KEYINPUT86), .Z(n613) );
  XNOR2_X1 U684 ( .A(n614), .B(n613), .ZN(G57) );
  XNOR2_X1 U685 ( .A(G101), .B(n615), .ZN(G3) );
  NOR2_X1 U686 ( .A1(n626), .A2(n617), .ZN(n616) );
  XOR2_X1 U687 ( .A(G104), .B(n616), .Z(G6) );
  NOR2_X1 U688 ( .A1(n630), .A2(n617), .ZN(n619) );
  XNOR2_X1 U689 ( .A(KEYINPUT27), .B(KEYINPUT26), .ZN(n618) );
  XNOR2_X1 U690 ( .A(n619), .B(n618), .ZN(n620) );
  XNOR2_X1 U691 ( .A(G107), .B(n620), .ZN(G9) );
  NOR2_X1 U692 ( .A1(n624), .A2(n630), .ZN(n622) );
  XNOR2_X1 U693 ( .A(KEYINPUT115), .B(KEYINPUT29), .ZN(n621) );
  XNOR2_X1 U694 ( .A(n622), .B(n621), .ZN(n623) );
  XOR2_X1 U695 ( .A(G128), .B(n623), .Z(G30) );
  NOR2_X1 U696 ( .A1(n624), .A2(n626), .ZN(n625) );
  XOR2_X1 U697 ( .A(G146), .B(n625), .Z(G48) );
  NOR2_X1 U698 ( .A1(n626), .A2(n629), .ZN(n627) );
  XOR2_X1 U699 ( .A(KEYINPUT116), .B(n627), .Z(n628) );
  XNOR2_X1 U700 ( .A(G113), .B(n628), .ZN(G15) );
  NOR2_X1 U701 ( .A1(n630), .A2(n629), .ZN(n631) );
  XOR2_X1 U702 ( .A(G116), .B(n631), .Z(G18) );
  XNOR2_X1 U703 ( .A(G125), .B(n632), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n633), .B(KEYINPUT37), .ZN(G27) );
  XNOR2_X1 U705 ( .A(n634), .B(KEYINPUT2), .ZN(n669) );
  NOR2_X1 U706 ( .A1(n636), .A2(n635), .ZN(n637) );
  XNOR2_X1 U707 ( .A(n637), .B(KEYINPUT49), .ZN(n638) );
  NAND2_X1 U708 ( .A1(n639), .A2(n638), .ZN(n644) );
  AND2_X1 U709 ( .A1(n641), .A2(n640), .ZN(n642) );
  XNOR2_X1 U710 ( .A(n642), .B(KEYINPUT50), .ZN(n643) );
  NOR2_X1 U711 ( .A1(n644), .A2(n643), .ZN(n645) );
  NOR2_X1 U712 ( .A1(n646), .A2(n645), .ZN(n647) );
  XOR2_X1 U713 ( .A(KEYINPUT51), .B(n647), .Z(n648) );
  NOR2_X1 U714 ( .A1(n664), .A2(n648), .ZN(n660) );
  INV_X1 U715 ( .A(n649), .ZN(n656) );
  AND2_X1 U716 ( .A1(n651), .A2(n650), .ZN(n652) );
  NOR2_X1 U717 ( .A1(n653), .A2(n652), .ZN(n655) );
  NOR2_X1 U718 ( .A1(n656), .A2(n353), .ZN(n657) );
  NOR2_X1 U719 ( .A1(n665), .A2(n657), .ZN(n658) );
  XOR2_X1 U720 ( .A(KEYINPUT117), .B(n658), .Z(n659) );
  NOR2_X1 U721 ( .A1(n660), .A2(n659), .ZN(n661) );
  XNOR2_X1 U722 ( .A(n661), .B(KEYINPUT52), .ZN(n662) );
  NOR2_X1 U723 ( .A1(n663), .A2(n662), .ZN(n667) );
  NOR2_X1 U724 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U725 ( .A1(n667), .A2(n666), .ZN(n668) );
  NAND2_X1 U726 ( .A1(n669), .A2(n668), .ZN(n670) );
  NOR2_X1 U727 ( .A1(G953), .A2(n670), .ZN(n672) );
  XNOR2_X1 U728 ( .A(KEYINPUT53), .B(KEYINPUT118), .ZN(n671) );
  XNOR2_X1 U729 ( .A(n672), .B(n671), .ZN(G75) );
  BUF_X1 U730 ( .A(n680), .Z(n673) );
  NAND2_X1 U731 ( .A1(n673), .A2(G469), .ZN(n678) );
  XNOR2_X1 U732 ( .A(KEYINPUT58), .B(KEYINPUT119), .ZN(n676) );
  XNOR2_X1 U733 ( .A(n674), .B(KEYINPUT57), .ZN(n675) );
  XNOR2_X1 U734 ( .A(n676), .B(n675), .ZN(n677) );
  XNOR2_X1 U735 ( .A(n678), .B(n677), .ZN(n679) );
  NOR2_X1 U736 ( .A1(n692), .A2(n679), .ZN(G54) );
  NAND2_X1 U737 ( .A1(n680), .A2(G475), .ZN(n684) );
  XOR2_X1 U738 ( .A(KEYINPUT59), .B(KEYINPUT120), .Z(n681) );
  XNOR2_X1 U739 ( .A(n684), .B(n683), .ZN(n685) );
  NAND2_X1 U740 ( .A1(n673), .A2(G478), .ZN(n687) );
  XNOR2_X1 U741 ( .A(n687), .B(n686), .ZN(n688) );
  NOR2_X1 U742 ( .A1(n692), .A2(n688), .ZN(G63) );
  NAND2_X1 U743 ( .A1(n673), .A2(G217), .ZN(n690) );
  XNOR2_X1 U744 ( .A(n690), .B(n689), .ZN(n691) );
  NOR2_X1 U745 ( .A1(n692), .A2(n691), .ZN(G66) );
  NOR2_X1 U746 ( .A1(n693), .A2(G953), .ZN(n694) );
  XNOR2_X1 U747 ( .A(n694), .B(KEYINPUT123), .ZN(n700) );
  XOR2_X1 U748 ( .A(KEYINPUT121), .B(KEYINPUT61), .Z(n696) );
  NAND2_X1 U749 ( .A1(G224), .A2(G953), .ZN(n695) );
  XNOR2_X1 U750 ( .A(n696), .B(n695), .ZN(n697) );
  NAND2_X1 U751 ( .A1(G898), .A2(n697), .ZN(n698) );
  XNOR2_X1 U752 ( .A(KEYINPUT122), .B(n698), .ZN(n699) );
  NAND2_X1 U753 ( .A1(n700), .A2(n699), .ZN(n707) );
  XNOR2_X1 U754 ( .A(G101), .B(n701), .ZN(n703) );
  XNOR2_X1 U755 ( .A(n703), .B(n702), .ZN(n705) );
  NOR2_X1 U756 ( .A1(G898), .A2(n717), .ZN(n704) );
  NOR2_X1 U757 ( .A1(n705), .A2(n704), .ZN(n706) );
  XNOR2_X1 U758 ( .A(n707), .B(n706), .ZN(G69) );
  XNOR2_X1 U759 ( .A(n708), .B(n709), .ZN(n710) );
  XOR2_X1 U760 ( .A(n711), .B(n710), .Z(n716) );
  XNOR2_X1 U761 ( .A(n716), .B(KEYINPUT124), .ZN(n712) );
  XNOR2_X1 U762 ( .A(G227), .B(n712), .ZN(n713) );
  NAND2_X1 U763 ( .A1(G900), .A2(n713), .ZN(n714) );
  NAND2_X1 U764 ( .A1(n714), .A2(G953), .ZN(n720) );
  XNOR2_X1 U765 ( .A(n716), .B(n715), .ZN(n718) );
  NAND2_X1 U766 ( .A1(n718), .A2(n717), .ZN(n719) );
  NAND2_X1 U767 ( .A1(n720), .A2(n719), .ZN(G72) );
  XNOR2_X1 U768 ( .A(G134), .B(n721), .ZN(G36) );
  XOR2_X1 U769 ( .A(G137), .B(KEYINPUT126), .Z(n722) );
  XNOR2_X1 U770 ( .A(n723), .B(n722), .ZN(G39) );
  XOR2_X1 U771 ( .A(G119), .B(n724), .Z(G21) );
  XOR2_X1 U772 ( .A(n725), .B(G131), .Z(G33) );
  XOR2_X1 U773 ( .A(G110), .B(n726), .Z(G12) );
endmodule

