//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 1 0 0 0 0 0 0 1 1 0 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 1 0 1 1 1 0 0 1 0 1 0 1 1 1 0 0 0 0 1 0 1 1 0 1 0 0 1 1 0 0 1 0 0 1 0 0 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:16:34 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n624,
    new_n625, new_n626, new_n628, new_n629, new_n630, new_n631, new_n632,
    new_n633, new_n634, new_n635, new_n636, new_n637, new_n638, new_n639,
    new_n640, new_n641, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n655, new_n656, new_n657, new_n658, new_n659, new_n660, new_n661,
    new_n662, new_n663, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n700, new_n701,
    new_n702, new_n704, new_n706, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n747, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n773, new_n774, new_n776, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n798, new_n799, new_n800, new_n801, new_n802,
    new_n803, new_n804, new_n805, new_n806, new_n807, new_n808, new_n809,
    new_n810, new_n812, new_n813, new_n814, new_n815, new_n816, new_n817,
    new_n818, new_n819, new_n820, new_n821, new_n823, new_n824, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n853, new_n854, new_n855, new_n856, new_n857,
    new_n858, new_n860, new_n861, new_n862, new_n863, new_n864, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n895, new_n896, new_n897;
  NAND2_X1  g000(.A1(G229gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G43gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G50gat), .ZN(new_n204));
  INV_X1    g003(.A(G50gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G43gat), .ZN(new_n206));
  AND3_X1   g005(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT15), .ZN(new_n207));
  AOI21_X1  g006(.A(new_n207), .B1(G29gat), .B2(G36gat), .ZN(new_n208));
  INV_X1    g007(.A(KEYINPUT15), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT78), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n206), .B1(new_n204), .B2(new_n210), .ZN(new_n211));
  NOR2_X1   g010(.A1(new_n205), .A2(G43gat), .ZN(new_n212));
  NOR2_X1   g011(.A1(new_n212), .A2(KEYINPUT78), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n209), .B1(new_n211), .B2(new_n213), .ZN(new_n214));
  OAI21_X1  g013(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  INV_X1    g015(.A(KEYINPUT14), .ZN(new_n217));
  INV_X1    g016(.A(G29gat), .ZN(new_n218));
  INV_X1    g017(.A(G36gat), .ZN(new_n219));
  NAND3_X1  g018(.A1(new_n217), .A2(new_n218), .A3(new_n219), .ZN(new_n220));
  XNOR2_X1  g019(.A(new_n220), .B(KEYINPUT79), .ZN(new_n221));
  OAI211_X1 g020(.A(new_n208), .B(new_n214), .C1(new_n216), .C2(new_n221), .ZN(new_n222));
  AOI22_X1  g021(.A1(new_n220), .A2(new_n215), .B1(G29gat), .B2(G36gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n204), .A2(new_n206), .A3(KEYINPUT15), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT77), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n225), .A2(new_n226), .ZN(new_n227));
  OAI21_X1  g026(.A(KEYINPUT77), .B1(new_n223), .B2(new_n224), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n222), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(KEYINPUT80), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n230), .A2(new_n231), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n222), .A2(new_n229), .A3(KEYINPUT80), .ZN(new_n233));
  XNOR2_X1  g032(.A(G15gat), .B(G22gat), .ZN(new_n234));
  INV_X1    g033(.A(G1gat), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT16), .A3(new_n235), .ZN(new_n236));
  OAI221_X1 g035(.A(new_n236), .B1(KEYINPUT81), .B2(G8gat), .C1(new_n235), .C2(new_n234), .ZN(new_n237));
  NAND2_X1  g036(.A1(KEYINPUT81), .A2(G8gat), .ZN(new_n238));
  XNOR2_X1  g037(.A(new_n237), .B(new_n238), .ZN(new_n239));
  NAND3_X1  g038(.A1(new_n232), .A2(new_n233), .A3(new_n239), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT17), .ZN(new_n241));
  AND3_X1   g040(.A1(new_n232), .A2(new_n241), .A3(new_n233), .ZN(new_n242));
  INV_X1    g041(.A(new_n239), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n222), .A2(new_n229), .A3(KEYINPUT17), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n202), .B(new_n240), .C1(new_n242), .C2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(KEYINPUT18), .ZN(new_n247));
  NAND2_X1  g046(.A1(new_n246), .A2(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n232), .A2(new_n233), .ZN(new_n249));
  OAI211_X1 g048(.A(new_n243), .B(new_n244), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n250), .A2(KEYINPUT18), .A3(new_n202), .A4(new_n240), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n243), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n252), .A2(new_n240), .ZN(new_n253));
  XOR2_X1   g052(.A(new_n202), .B(KEYINPUT13), .Z(new_n254));
  NAND2_X1  g053(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND3_X1  g054(.A1(new_n248), .A2(new_n251), .A3(new_n255), .ZN(new_n256));
  XNOR2_X1  g055(.A(G113gat), .B(G141gat), .ZN(new_n257));
  XNOR2_X1  g056(.A(new_n257), .B(G197gat), .ZN(new_n258));
  XOR2_X1   g057(.A(KEYINPUT11), .B(G169gat), .Z(new_n259));
  XNOR2_X1  g058(.A(new_n258), .B(new_n259), .ZN(new_n260));
  XNOR2_X1  g059(.A(new_n260), .B(KEYINPUT12), .ZN(new_n261));
  INV_X1    g060(.A(new_n261), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n256), .A2(new_n262), .ZN(new_n263));
  NAND4_X1  g062(.A1(new_n248), .A2(new_n251), .A3(new_n261), .A4(new_n255), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(new_n265), .ZN(new_n266));
  XNOR2_X1  g065(.A(G1gat), .B(G29gat), .ZN(new_n267));
  XNOR2_X1  g066(.A(G57gat), .B(G85gat), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(new_n268), .ZN(new_n269));
  XNOR2_X1  g068(.A(KEYINPUT71), .B(KEYINPUT0), .ZN(new_n270));
  XNOR2_X1  g069(.A(new_n269), .B(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G141gat), .B(G148gat), .ZN(new_n272));
  INV_X1    g071(.A(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G155gat), .ZN(new_n274));
  INV_X1    g073(.A(G162gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND2_X1  g075(.A1(G155gat), .A2(G162gat), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n276), .A2(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n277), .A2(KEYINPUT2), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n273), .A2(new_n278), .A3(new_n279), .ZN(new_n280));
  OAI211_X1 g079(.A(new_n277), .B(new_n276), .C1(new_n272), .C2(KEYINPUT2), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT70), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  AOI21_X1  g082(.A(KEYINPUT70), .B1(new_n280), .B2(new_n281), .ZN(new_n284));
  OAI21_X1  g083(.A(KEYINPUT3), .B1(new_n283), .B2(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n280), .A2(new_n281), .ZN(new_n286));
  NOR2_X1   g085(.A1(new_n286), .A2(KEYINPUT3), .ZN(new_n287));
  XNOR2_X1  g086(.A(G113gat), .B(G120gat), .ZN(new_n288));
  NOR2_X1   g087(.A1(new_n288), .A2(KEYINPUT1), .ZN(new_n289));
  OR2_X1    g088(.A1(G127gat), .A2(G134gat), .ZN(new_n290));
  NAND2_X1  g089(.A1(G127gat), .A2(G134gat), .ZN(new_n291));
  NAND2_X1  g090(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT1), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n293), .A2(KEYINPUT64), .ZN(new_n294));
  NAND2_X1  g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(new_n289), .A2(new_n295), .ZN(new_n296));
  OAI211_X1 g095(.A(new_n292), .B(new_n294), .C1(new_n288), .C2(KEYINPUT1), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NOR2_X1   g097(.A1(new_n287), .A2(new_n298), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n285), .A2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(G225gat), .A2(G233gat), .ZN(new_n301));
  AND2_X1   g100(.A1(new_n280), .A2(new_n281), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n302), .A2(new_n298), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT4), .ZN(new_n304));
  NAND2_X1  g103(.A1(new_n303), .A2(new_n304), .ZN(new_n305));
  NAND3_X1  g104(.A1(new_n302), .A2(new_n298), .A3(KEYINPUT4), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n300), .A2(new_n301), .A3(new_n305), .A4(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(KEYINPUT5), .ZN(new_n308));
  AND2_X1   g107(.A1(new_n296), .A2(new_n297), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n309), .B1(new_n283), .B2(new_n284), .ZN(new_n310));
  NAND2_X1  g109(.A1(new_n310), .A2(new_n303), .ZN(new_n311));
  INV_X1    g110(.A(new_n301), .ZN(new_n312));
  AOI21_X1  g111(.A(new_n308), .B1(new_n311), .B2(new_n312), .ZN(new_n313));
  NAND2_X1  g112(.A1(new_n307), .A2(new_n313), .ZN(new_n314));
  AND2_X1   g113(.A1(new_n305), .A2(new_n306), .ZN(new_n315));
  NAND4_X1  g114(.A1(new_n315), .A2(new_n308), .A3(new_n300), .A4(new_n301), .ZN(new_n316));
  AOI21_X1  g115(.A(new_n271), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(KEYINPUT75), .ZN(new_n318));
  OAI21_X1  g117(.A(new_n309), .B1(KEYINPUT3), .B2(new_n286), .ZN(new_n319));
  INV_X1    g118(.A(new_n284), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n320), .A2(new_n282), .ZN(new_n321));
  AOI21_X1  g120(.A(new_n319), .B1(new_n321), .B2(KEYINPUT3), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n305), .A2(new_n306), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n318), .B1(new_n324), .B2(new_n301), .ZN(new_n325));
  OAI211_X1 g124(.A(KEYINPUT75), .B(new_n312), .C1(new_n322), .C2(new_n323), .ZN(new_n326));
  NOR2_X1   g125(.A1(new_n311), .A2(new_n312), .ZN(new_n327));
  INV_X1    g126(.A(KEYINPUT39), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n325), .A2(new_n326), .A3(new_n329), .ZN(new_n330));
  AND2_X1   g129(.A1(new_n325), .A2(new_n326), .ZN(new_n331));
  OAI211_X1 g130(.A(new_n271), .B(new_n330), .C1(new_n331), .C2(KEYINPUT39), .ZN(new_n332));
  INV_X1    g131(.A(KEYINPUT40), .ZN(new_n333));
  AOI21_X1  g132(.A(new_n317), .B1(new_n332), .B2(new_n333), .ZN(new_n334));
  XNOR2_X1  g133(.A(G197gat), .B(G204gat), .ZN(new_n335));
  AND2_X1   g134(.A1(G211gat), .A2(G218gat), .ZN(new_n336));
  OAI21_X1  g135(.A(new_n335), .B1(KEYINPUT22), .B2(new_n336), .ZN(new_n337));
  XNOR2_X1  g136(.A(G211gat), .B(G218gat), .ZN(new_n338));
  XNOR2_X1  g137(.A(new_n337), .B(new_n338), .ZN(new_n339));
  NAND2_X1  g138(.A1(G226gat), .A2(G233gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(new_n340), .B(KEYINPUT67), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT68), .ZN(new_n342));
  INV_X1    g141(.A(G169gat), .ZN(new_n343));
  INV_X1    g142(.A(G176gat), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n343), .A2(new_n344), .ZN(new_n345));
  NOR2_X1   g144(.A1(G169gat), .A2(G176gat), .ZN(new_n346));
  OR3_X1    g145(.A1(new_n345), .A2(KEYINPUT26), .A3(new_n346), .ZN(new_n347));
  AOI22_X1  g146(.A1(new_n346), .A2(KEYINPUT26), .B1(G183gat), .B2(G190gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(KEYINPUT27), .B(G183gat), .ZN(new_n349));
  INV_X1    g148(.A(G190gat), .ZN(new_n350));
  AND3_X1   g149(.A1(new_n349), .A2(KEYINPUT28), .A3(new_n350), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT28), .B1(new_n349), .B2(new_n350), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n347), .B(new_n348), .C1(new_n351), .C2(new_n352), .ZN(new_n353));
  NAND2_X1  g152(.A1(G183gat), .A2(G190gat), .ZN(new_n354));
  OAI22_X1  g153(.A1(new_n354), .A2(KEYINPUT24), .B1(new_n343), .B2(new_n344), .ZN(new_n355));
  OAI21_X1  g154(.A(KEYINPUT23), .B1(G169gat), .B2(G176gat), .ZN(new_n356));
  INV_X1    g155(.A(KEYINPUT23), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n346), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g157(.A(new_n355), .B1(new_n356), .B2(new_n358), .ZN(new_n359));
  OR2_X1    g158(.A1(G183gat), .A2(G190gat), .ZN(new_n360));
  NAND3_X1  g159(.A1(new_n360), .A2(KEYINPUT24), .A3(new_n354), .ZN(new_n361));
  AOI21_X1  g160(.A(KEYINPUT25), .B1(new_n359), .B2(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(new_n355), .ZN(new_n363));
  NAND2_X1  g162(.A1(new_n358), .A2(new_n356), .ZN(new_n364));
  NAND3_X1  g163(.A1(new_n363), .A2(new_n361), .A3(new_n364), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT25), .ZN(new_n366));
  NOR2_X1   g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  OAI211_X1 g166(.A(new_n342), .B(new_n353), .C1(new_n362), .C2(new_n367), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  NAND3_X1  g168(.A1(new_n359), .A2(KEYINPUT25), .A3(new_n361), .ZN(new_n370));
  NAND2_X1  g169(.A1(new_n365), .A2(new_n366), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n370), .A2(new_n371), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n342), .B1(new_n372), .B2(new_n353), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n341), .B1(new_n369), .B2(new_n373), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n353), .B1(new_n362), .B2(new_n367), .ZN(new_n375));
  INV_X1    g174(.A(KEYINPUT29), .ZN(new_n376));
  INV_X1    g175(.A(new_n341), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n375), .A2(new_n376), .A3(new_n377), .ZN(new_n378));
  AOI21_X1  g177(.A(new_n339), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  NAND2_X1  g178(.A1(new_n375), .A2(KEYINPUT68), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n380), .A2(new_n376), .A3(new_n368), .ZN(new_n381));
  NAND2_X1  g180(.A1(new_n381), .A2(new_n377), .ZN(new_n382));
  NAND2_X1  g181(.A1(new_n375), .A2(new_n341), .ZN(new_n383));
  NAND2_X1  g182(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  AOI21_X1  g183(.A(new_n379), .B1(new_n384), .B2(new_n339), .ZN(new_n385));
  XNOR2_X1  g184(.A(G8gat), .B(G36gat), .ZN(new_n386));
  XNOR2_X1  g185(.A(G64gat), .B(G92gat), .ZN(new_n387));
  XOR2_X1   g186(.A(new_n386), .B(new_n387), .Z(new_n388));
  NAND4_X1  g187(.A1(new_n385), .A2(KEYINPUT69), .A3(KEYINPUT30), .A4(new_n388), .ZN(new_n389));
  INV_X1    g188(.A(KEYINPUT69), .ZN(new_n390));
  INV_X1    g189(.A(new_n339), .ZN(new_n391));
  AOI21_X1  g190(.A(new_n377), .B1(new_n380), .B2(new_n368), .ZN(new_n392));
  INV_X1    g191(.A(new_n378), .ZN(new_n393));
  OAI21_X1  g192(.A(new_n391), .B1(new_n392), .B2(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n383), .ZN(new_n395));
  AOI21_X1  g194(.A(new_n395), .B1(new_n381), .B2(new_n377), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n394), .B(new_n388), .C1(new_n396), .C2(new_n391), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  OAI21_X1  g197(.A(new_n390), .B1(new_n397), .B2(new_n398), .ZN(new_n399));
  NAND2_X1  g198(.A1(new_n389), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n397), .A2(new_n398), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n394), .B1(new_n396), .B2(new_n391), .ZN(new_n402));
  INV_X1    g201(.A(new_n388), .ZN(new_n403));
  NAND2_X1  g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g203(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n400), .A2(new_n405), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n334), .B(new_n406), .C1(new_n333), .C2(new_n332), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT37), .ZN(new_n408));
  AOI21_X1  g207(.A(new_n388), .B1(new_n385), .B2(new_n408), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n409), .B1(new_n408), .B2(new_n385), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n410), .A2(KEYINPUT38), .ZN(new_n411));
  INV_X1    g210(.A(KEYINPUT76), .ZN(new_n412));
  AOI21_X1  g211(.A(new_n412), .B1(new_n317), .B2(KEYINPUT6), .ZN(new_n413));
  NAND2_X1  g212(.A1(new_n314), .A2(new_n316), .ZN(new_n414));
  INV_X1    g213(.A(new_n271), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n414), .A2(KEYINPUT6), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n314), .A2(new_n316), .A3(new_n271), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT6), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  OAI21_X1  g218(.A(new_n416), .B1(new_n419), .B2(new_n317), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n413), .B1(new_n420), .B2(new_n412), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n384), .A2(new_n391), .ZN(new_n422));
  NAND2_X1  g221(.A1(new_n374), .A2(new_n378), .ZN(new_n423));
  AOI21_X1  g222(.A(new_n408), .B1(new_n423), .B2(new_n339), .ZN(new_n424));
  AOI21_X1  g223(.A(KEYINPUT38), .B1(new_n422), .B2(new_n424), .ZN(new_n425));
  AOI22_X1  g224(.A1(new_n409), .A2(new_n425), .B1(new_n385), .B2(new_n388), .ZN(new_n426));
  NAND3_X1  g225(.A1(new_n411), .A2(new_n421), .A3(new_n426), .ZN(new_n427));
  INV_X1    g226(.A(KEYINPUT3), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n428), .B1(new_n339), .B2(KEYINPUT29), .ZN(new_n429));
  NAND2_X1  g228(.A1(new_n429), .A2(new_n286), .ZN(new_n430));
  NAND2_X1  g229(.A1(G228gat), .A2(G233gat), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n339), .B1(new_n287), .B2(KEYINPUT29), .ZN(new_n432));
  AND3_X1   g231(.A1(new_n430), .A2(new_n431), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n321), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n431), .B1(new_n434), .B2(new_n432), .ZN(new_n435));
  INV_X1    g234(.A(G22gat), .ZN(new_n436));
  OR3_X1    g235(.A1(new_n433), .A2(new_n435), .A3(new_n436), .ZN(new_n437));
  XNOR2_X1  g236(.A(G78gat), .B(G106gat), .ZN(new_n438));
  XNOR2_X1  g237(.A(new_n438), .B(KEYINPUT73), .ZN(new_n439));
  XNOR2_X1  g238(.A(KEYINPUT31), .B(G50gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(new_n439), .B(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT74), .ZN(new_n442));
  XNOR2_X1  g241(.A(new_n441), .B(new_n442), .ZN(new_n443));
  OAI21_X1  g242(.A(new_n436), .B1(new_n433), .B2(new_n435), .ZN(new_n444));
  AND3_X1   g243(.A1(new_n437), .A2(new_n443), .A3(new_n444), .ZN(new_n445));
  AOI22_X1  g244(.A1(new_n437), .A2(new_n444), .B1(new_n442), .B2(new_n441), .ZN(new_n446));
  NOR2_X1   g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  INV_X1    g246(.A(new_n447), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n407), .A2(new_n427), .A3(new_n448), .ZN(new_n449));
  INV_X1    g248(.A(new_n449), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n420), .A2(new_n404), .A3(new_n401), .ZN(new_n451));
  AND2_X1   g250(.A1(new_n389), .A2(new_n399), .ZN(new_n452));
  OAI21_X1  g251(.A(KEYINPUT72), .B1(new_n451), .B2(new_n452), .ZN(new_n453));
  INV_X1    g252(.A(KEYINPUT72), .ZN(new_n454));
  NAND4_X1  g253(.A1(new_n400), .A2(new_n405), .A3(new_n454), .A4(new_n420), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n448), .B1(new_n453), .B2(new_n455), .ZN(new_n456));
  INV_X1    g255(.A(KEYINPUT34), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n375), .A2(new_n298), .ZN(new_n458));
  NAND3_X1  g257(.A1(new_n372), .A2(new_n309), .A3(new_n353), .ZN(new_n459));
  AOI22_X1  g258(.A1(new_n458), .A2(new_n459), .B1(G227gat), .B2(G233gat), .ZN(new_n460));
  OAI21_X1  g259(.A(new_n457), .B1(new_n460), .B2(KEYINPUT65), .ZN(new_n461));
  NAND4_X1  g260(.A1(new_n458), .A2(G227gat), .A3(G233gat), .A4(new_n459), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n462), .A2(KEYINPUT32), .ZN(new_n463));
  INV_X1    g262(.A(KEYINPUT33), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n462), .A2(new_n464), .ZN(new_n465));
  XOR2_X1   g264(.A(G15gat), .B(G43gat), .Z(new_n466));
  XNOR2_X1  g265(.A(G71gat), .B(G99gat), .ZN(new_n467));
  XNOR2_X1  g266(.A(new_n466), .B(new_n467), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n463), .A2(new_n465), .A3(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n468), .ZN(new_n470));
  OAI211_X1 g269(.A(new_n462), .B(KEYINPUT32), .C1(new_n464), .C2(new_n470), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n461), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  INV_X1    g271(.A(new_n472), .ZN(new_n473));
  NAND3_X1  g272(.A1(new_n469), .A2(new_n471), .A3(new_n461), .ZN(new_n474));
  NAND4_X1  g273(.A1(new_n473), .A2(KEYINPUT65), .A3(new_n460), .A4(new_n474), .ZN(new_n475));
  NAND2_X1  g274(.A1(new_n460), .A2(KEYINPUT65), .ZN(new_n476));
  INV_X1    g275(.A(new_n474), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n476), .B1(new_n477), .B2(new_n472), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n475), .A2(new_n478), .ZN(new_n479));
  INV_X1    g278(.A(KEYINPUT66), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n480), .A2(KEYINPUT36), .ZN(new_n482));
  NAND3_X1  g281(.A1(new_n479), .A2(new_n481), .A3(new_n482), .ZN(new_n483));
  NAND4_X1  g282(.A1(new_n475), .A2(new_n478), .A3(new_n480), .A4(KEYINPUT36), .ZN(new_n484));
  NAND2_X1  g283(.A1(new_n483), .A2(new_n484), .ZN(new_n485));
  NOR2_X1   g284(.A1(new_n456), .A2(new_n485), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n450), .A2(new_n486), .ZN(new_n487));
  AOI21_X1  g286(.A(new_n447), .B1(new_n475), .B2(new_n478), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n453), .A2(new_n455), .A3(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(KEYINPUT35), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n421), .A2(KEYINPUT35), .ZN(new_n491));
  INV_X1    g290(.A(new_n406), .ZN(new_n492));
  NAND3_X1  g291(.A1(new_n491), .A2(new_n488), .A3(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n490), .A2(new_n493), .ZN(new_n494));
  AOI21_X1  g293(.A(new_n266), .B1(new_n487), .B2(new_n494), .ZN(new_n495));
  NOR2_X1   g294(.A1(G71gat), .A2(G78gat), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT9), .ZN(new_n497));
  NAND2_X1  g296(.A1(G71gat), .A2(G78gat), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT83), .ZN(new_n500));
  INV_X1    g299(.A(G57gat), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  NAND2_X1  g301(.A1(KEYINPUT83), .A2(G57gat), .ZN(new_n503));
  NAND3_X1  g302(.A1(new_n502), .A2(G64gat), .A3(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(G64gat), .ZN(new_n505));
  AOI21_X1  g304(.A(KEYINPUT84), .B1(new_n505), .B2(G57gat), .ZN(new_n506));
  NAND2_X1  g305(.A1(new_n504), .A2(new_n506), .ZN(new_n507));
  NAND4_X1  g306(.A1(new_n502), .A2(KEYINPUT84), .A3(G64gat), .A4(new_n503), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n507), .A2(KEYINPUT85), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT85), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n499), .B1(new_n509), .B2(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n496), .B1(KEYINPUT82), .B2(new_n498), .ZN(new_n512));
  XNOR2_X1  g311(.A(G57gat), .B(G64gat), .ZN(new_n513));
  NOR2_X1   g312(.A1(KEYINPUT82), .A2(KEYINPUT9), .ZN(new_n514));
  OAI221_X1 g313(.A(new_n512), .B1(KEYINPUT82), .B2(new_n498), .C1(new_n513), .C2(new_n514), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n511), .A2(new_n515), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT21), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NAND2_X1  g317(.A1(G231gat), .A2(G233gat), .ZN(new_n519));
  XNOR2_X1  g318(.A(new_n518), .B(new_n519), .ZN(new_n520));
  XNOR2_X1  g319(.A(new_n520), .B(G127gat), .ZN(new_n521));
  OAI21_X1  g320(.A(new_n243), .B1(new_n517), .B2(new_n516), .ZN(new_n522));
  XNOR2_X1  g321(.A(new_n522), .B(KEYINPUT87), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  INV_X1    g323(.A(new_n524), .ZN(new_n525));
  NOR2_X1   g324(.A1(new_n521), .A2(new_n523), .ZN(new_n526));
  XNOR2_X1  g325(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n527));
  XNOR2_X1  g326(.A(new_n527), .B(KEYINPUT86), .ZN(new_n528));
  XNOR2_X1  g327(.A(new_n528), .B(G155gat), .ZN(new_n529));
  XOR2_X1   g328(.A(G183gat), .B(G211gat), .Z(new_n530));
  XNOR2_X1  g329(.A(new_n530), .B(KEYINPUT88), .ZN(new_n531));
  XNOR2_X1  g330(.A(new_n529), .B(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(new_n532), .ZN(new_n533));
  OR3_X1    g332(.A1(new_n525), .A2(new_n526), .A3(new_n533), .ZN(new_n534));
  OAI21_X1  g333(.A(new_n533), .B1(new_n525), .B2(new_n526), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n534), .A2(new_n535), .ZN(new_n536));
  INV_X1    g335(.A(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n538));
  INV_X1    g337(.A(G85gat), .ZN(new_n539));
  NAND2_X1  g338(.A1(KEYINPUT90), .A2(G92gat), .ZN(new_n540));
  NAND3_X1  g339(.A1(new_n538), .A2(new_n539), .A3(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G99gat), .ZN(new_n542));
  INV_X1    g341(.A(G106gat), .ZN(new_n543));
  OAI21_X1  g342(.A(KEYINPUT8), .B1(new_n542), .B2(new_n543), .ZN(new_n544));
  AND2_X1   g343(.A1(new_n541), .A2(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(G99gat), .B(G106gat), .ZN(new_n546));
  NAND3_X1  g345(.A1(KEYINPUT89), .A2(G85gat), .A3(G92gat), .ZN(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(KEYINPUT7), .ZN(new_n548));
  AND3_X1   g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  AOI21_X1  g348(.A(new_n546), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g349(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  NAND2_X1  g350(.A1(new_n551), .A2(KEYINPUT91), .ZN(new_n552));
  INV_X1    g351(.A(KEYINPUT91), .ZN(new_n553));
  OAI21_X1  g352(.A(new_n553), .B1(new_n549), .B2(new_n550), .ZN(new_n554));
  NAND2_X1  g353(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NOR2_X1   g354(.A1(new_n249), .A2(new_n555), .ZN(new_n556));
  AND2_X1   g355(.A1(G232gat), .A2(G233gat), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(KEYINPUT41), .B2(new_n557), .ZN(new_n558));
  OAI211_X1 g357(.A(new_n244), .B(new_n555), .C1(new_n249), .C2(KEYINPUT17), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  XOR2_X1   g359(.A(G190gat), .B(G218gat), .Z(new_n561));
  NAND2_X1  g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NOR2_X1   g361(.A1(new_n557), .A2(KEYINPUT41), .ZN(new_n563));
  XNOR2_X1  g362(.A(G134gat), .B(G162gat), .ZN(new_n564));
  XNOR2_X1  g363(.A(new_n563), .B(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n561), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n558), .A2(new_n566), .A3(new_n559), .ZN(new_n567));
  AND3_X1   g366(.A1(new_n562), .A2(new_n565), .A3(new_n567), .ZN(new_n568));
  AOI21_X1  g367(.A(new_n565), .B1(new_n562), .B2(new_n567), .ZN(new_n569));
  NOR2_X1   g368(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n537), .A2(new_n571), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n511), .A2(new_n515), .A3(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n551), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT10), .ZN(new_n577));
  NAND4_X1  g376(.A1(new_n551), .A2(new_n511), .A3(new_n515), .A4(new_n573), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n576), .A2(new_n577), .A3(new_n578), .ZN(new_n579));
  INV_X1    g378(.A(new_n516), .ZN(new_n580));
  NAND4_X1  g379(.A1(new_n580), .A2(new_n552), .A3(KEYINPUT10), .A4(new_n554), .ZN(new_n581));
  NAND2_X1  g380(.A1(new_n579), .A2(new_n581), .ZN(new_n582));
  NAND2_X1  g381(.A1(G230gat), .A2(G233gat), .ZN(new_n583));
  XOR2_X1   g382(.A(new_n583), .B(KEYINPUT93), .Z(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  NAND2_X1  g384(.A1(new_n582), .A2(new_n585), .ZN(new_n586));
  AOI21_X1  g385(.A(new_n585), .B1(new_n576), .B2(new_n578), .ZN(new_n587));
  INV_X1    g386(.A(new_n587), .ZN(new_n588));
  XNOR2_X1  g387(.A(G120gat), .B(G148gat), .ZN(new_n589));
  XNOR2_X1  g388(.A(G176gat), .B(G204gat), .ZN(new_n590));
  XOR2_X1   g389(.A(new_n589), .B(new_n590), .Z(new_n591));
  NAND3_X1  g390(.A1(new_n586), .A2(new_n588), .A3(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n592), .A2(KEYINPUT94), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT94), .ZN(new_n594));
  NAND4_X1  g393(.A1(new_n586), .A2(new_n594), .A3(new_n588), .A4(new_n591), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n593), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n591), .ZN(new_n597));
  AOI21_X1  g396(.A(new_n584), .B1(new_n579), .B2(new_n581), .ZN(new_n598));
  OAI21_X1  g397(.A(new_n597), .B1(new_n598), .B2(new_n587), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT95), .ZN(new_n600));
  NAND2_X1  g399(.A1(new_n599), .A2(new_n600), .ZN(new_n601));
  OAI211_X1 g400(.A(KEYINPUT95), .B(new_n597), .C1(new_n598), .C2(new_n587), .ZN(new_n602));
  NAND2_X1  g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(KEYINPUT96), .B1(new_n596), .B2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(new_n604), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n596), .A2(KEYINPUT96), .A3(new_n603), .ZN(new_n606));
  NAND2_X1  g405(.A1(new_n605), .A2(new_n606), .ZN(new_n607));
  NOR2_X1   g406(.A1(new_n572), .A2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n495), .A2(new_n608), .ZN(new_n609));
  NOR2_X1   g408(.A1(new_n609), .A2(new_n420), .ZN(new_n610));
  XOR2_X1   g409(.A(KEYINPUT97), .B(G1gat), .Z(new_n611));
  XNOR2_X1  g410(.A(new_n610), .B(new_n611), .ZN(G1324gat));
  NAND3_X1  g411(.A1(new_n495), .A2(new_n406), .A3(new_n608), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n613), .A2(G8gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(KEYINPUT16), .B(G8gat), .ZN(new_n615));
  NOR2_X1   g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(KEYINPUT42), .B1(new_n614), .B2(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(new_n617), .B1(KEYINPUT42), .B2(new_n616), .ZN(G1325gat));
  INV_X1    g417(.A(new_n485), .ZN(new_n619));
  OAI21_X1  g418(.A(G15gat), .B1(new_n609), .B2(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n479), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n621), .A2(G15gat), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n609), .B2(new_n622), .ZN(G1326gat));
  NOR2_X1   g422(.A1(new_n609), .A2(new_n448), .ZN(new_n624));
  XNOR2_X1  g423(.A(new_n624), .B(KEYINPUT98), .ZN(new_n625));
  XNOR2_X1  g424(.A(KEYINPUT43), .B(G22gat), .ZN(new_n626));
  XNOR2_X1  g425(.A(new_n625), .B(new_n626), .ZN(G1327gat));
  AND3_X1   g426(.A1(new_n596), .A2(KEYINPUT96), .A3(new_n603), .ZN(new_n628));
  NOR2_X1   g427(.A1(new_n628), .A2(new_n604), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n536), .A2(new_n629), .A3(new_n570), .ZN(new_n630));
  XOR2_X1   g429(.A(new_n630), .B(KEYINPUT99), .Z(new_n631));
  INV_X1    g430(.A(new_n420), .ZN(new_n632));
  NAND4_X1  g431(.A1(new_n495), .A2(new_n631), .A3(new_n218), .A4(new_n632), .ZN(new_n633));
  XNOR2_X1  g432(.A(new_n633), .B(KEYINPUT45), .ZN(new_n634));
  NOR3_X1   g433(.A1(new_n449), .A2(new_n485), .A3(new_n456), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n494), .A2(KEYINPUT101), .ZN(new_n636));
  INV_X1    g435(.A(KEYINPUT101), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n490), .A2(new_n637), .A3(new_n493), .ZN(new_n638));
  AOI21_X1  g437(.A(new_n635), .B1(new_n636), .B2(new_n638), .ZN(new_n639));
  NOR2_X1   g438(.A1(new_n571), .A2(KEYINPUT44), .ZN(new_n640));
  INV_X1    g439(.A(new_n640), .ZN(new_n641));
  OAI21_X1  g440(.A(KEYINPUT102), .B1(new_n639), .B2(new_n641), .ZN(new_n642));
  INV_X1    g441(.A(new_n638), .ZN(new_n643));
  AOI21_X1  g442(.A(new_n637), .B1(new_n490), .B2(new_n493), .ZN(new_n644));
  OAI21_X1  g443(.A(new_n487), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(KEYINPUT102), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n645), .A2(new_n646), .A3(new_n640), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n487), .A2(new_n494), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n570), .ZN(new_n649));
  AOI22_X1  g448(.A1(new_n642), .A2(new_n647), .B1(KEYINPUT44), .B2(new_n649), .ZN(new_n650));
  XNOR2_X1  g449(.A(new_n607), .B(KEYINPUT100), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n651), .A2(new_n265), .A3(new_n536), .ZN(new_n652));
  NOR3_X1   g451(.A1(new_n650), .A2(new_n420), .A3(new_n652), .ZN(new_n653));
  OAI21_X1  g452(.A(new_n634), .B1(new_n653), .B2(new_n218), .ZN(G1328gat));
  INV_X1    g453(.A(KEYINPUT104), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n642), .A2(new_n647), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n649), .A2(KEYINPUT44), .ZN(new_n657));
  AOI21_X1  g456(.A(new_n652), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AOI21_X1  g457(.A(new_n219), .B1(new_n658), .B2(new_n406), .ZN(new_n659));
  NAND4_X1  g458(.A1(new_n631), .A2(new_n495), .A3(new_n219), .A4(new_n406), .ZN(new_n660));
  NAND2_X1  g459(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n661));
  INV_X1    g460(.A(new_n661), .ZN(new_n662));
  OR2_X1    g461(.A1(new_n660), .A2(new_n662), .ZN(new_n663));
  NOR2_X1   g462(.A1(KEYINPUT103), .A2(KEYINPUT46), .ZN(new_n664));
  OAI21_X1  g463(.A(new_n660), .B1(new_n662), .B2(new_n664), .ZN(new_n665));
  NAND2_X1  g464(.A1(new_n663), .A2(new_n665), .ZN(new_n666));
  OAI21_X1  g465(.A(new_n655), .B1(new_n659), .B2(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n666), .ZN(new_n668));
  NOR3_X1   g467(.A1(new_n650), .A2(new_n492), .A3(new_n652), .ZN(new_n669));
  OAI211_X1 g468(.A(new_n668), .B(KEYINPUT104), .C1(new_n669), .C2(new_n219), .ZN(new_n670));
  NAND2_X1  g469(.A1(new_n667), .A2(new_n670), .ZN(G1329gat));
  NAND2_X1  g470(.A1(new_n656), .A2(new_n657), .ZN(new_n672));
  INV_X1    g471(.A(new_n652), .ZN(new_n673));
  NAND4_X1  g472(.A1(new_n672), .A2(G43gat), .A3(new_n485), .A4(new_n673), .ZN(new_n674));
  NAND3_X1  g473(.A1(new_n495), .A2(new_n631), .A3(new_n479), .ZN(new_n675));
  AOI22_X1  g474(.A1(new_n675), .A2(new_n203), .B1(KEYINPUT105), .B2(KEYINPUT47), .ZN(new_n676));
  NOR2_X1   g475(.A1(KEYINPUT105), .A2(KEYINPUT47), .ZN(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT106), .ZN(new_n678));
  AND3_X1   g477(.A1(new_n674), .A2(new_n676), .A3(new_n678), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n678), .B1(new_n674), .B2(new_n676), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n679), .A2(new_n680), .ZN(G1330gat));
  NAND4_X1  g480(.A1(new_n631), .A2(new_n495), .A3(new_n205), .A4(new_n447), .ZN(new_n682));
  XOR2_X1   g481(.A(new_n682), .B(KEYINPUT108), .Z(new_n683));
  NAND3_X1  g482(.A1(new_n672), .A2(new_n447), .A3(new_n673), .ZN(new_n684));
  AOI21_X1  g483(.A(new_n683), .B1(new_n684), .B2(G50gat), .ZN(new_n685));
  XOR2_X1   g484(.A(KEYINPUT107), .B(KEYINPUT48), .Z(new_n686));
  AOI21_X1  g485(.A(new_n205), .B1(new_n658), .B2(new_n447), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n682), .A2(KEYINPUT48), .ZN(new_n688));
  OAI22_X1  g487(.A1(new_n685), .A2(new_n686), .B1(new_n687), .B2(new_n688), .ZN(G1331gat));
  NOR4_X1   g488(.A1(new_n639), .A2(new_n265), .A3(new_n572), .A4(new_n651), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n690), .A2(new_n632), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n502), .A2(new_n503), .ZN(new_n692));
  XNOR2_X1  g491(.A(new_n691), .B(new_n692), .ZN(G1332gat));
  XNOR2_X1  g492(.A(new_n406), .B(KEYINPUT109), .ZN(new_n694));
  INV_X1    g493(.A(new_n694), .ZN(new_n695));
  NAND2_X1  g494(.A1(new_n690), .A2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n697));
  XOR2_X1   g496(.A(KEYINPUT49), .B(G64gat), .Z(new_n698));
  OAI21_X1  g497(.A(new_n697), .B1(new_n696), .B2(new_n698), .ZN(G1333gat));
  NAND2_X1  g498(.A1(new_n690), .A2(new_n485), .ZN(new_n700));
  NOR2_X1   g499(.A1(new_n621), .A2(G71gat), .ZN(new_n701));
  AOI22_X1  g500(.A1(new_n700), .A2(G71gat), .B1(new_n690), .B2(new_n701), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n702), .B(KEYINPUT50), .ZN(G1334gat));
  NAND2_X1  g502(.A1(new_n690), .A2(new_n447), .ZN(new_n704));
  XNOR2_X1  g503(.A(new_n704), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g504(.A1(new_n537), .A2(new_n265), .ZN(new_n706));
  NAND2_X1  g505(.A1(new_n706), .A2(new_n607), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n707), .B1(new_n656), .B2(new_n657), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(G85gat), .B1(new_n709), .B2(new_n420), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT110), .ZN(new_n711));
  INV_X1    g510(.A(KEYINPUT51), .ZN(new_n712));
  NOR2_X1   g511(.A1(new_n711), .A2(new_n712), .ZN(new_n713));
  AOI21_X1  g512(.A(new_n571), .B1(new_n711), .B2(new_n712), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n706), .A2(new_n714), .ZN(new_n715));
  OR3_X1    g514(.A1(new_n639), .A2(new_n713), .A3(new_n715), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n713), .B1(new_n639), .B2(new_n715), .ZN(new_n717));
  AND2_X1   g516(.A1(new_n716), .A2(new_n717), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n718), .A2(new_n607), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n632), .A2(new_n539), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n710), .B1(new_n719), .B2(new_n720), .ZN(G1336gat));
  INV_X1    g520(.A(new_n651), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n694), .A2(G92gat), .ZN(new_n723));
  NAND4_X1  g522(.A1(new_n716), .A2(new_n722), .A3(new_n717), .A4(new_n723), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n707), .ZN(new_n726));
  NAND3_X1  g525(.A1(new_n672), .A2(new_n406), .A3(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n538), .A2(new_n540), .ZN(new_n728));
  AOI21_X1  g527(.A(new_n725), .B1(new_n727), .B2(new_n728), .ZN(new_n729));
  INV_X1    g528(.A(KEYINPUT52), .ZN(new_n730));
  AOI22_X1  g529(.A1(new_n708), .A2(new_n695), .B1(new_n538), .B2(new_n540), .ZN(new_n731));
  XOR2_X1   g530(.A(KEYINPUT111), .B(KEYINPUT52), .Z(new_n732));
  NAND2_X1  g531(.A1(new_n724), .A2(new_n732), .ZN(new_n733));
  OAI22_X1  g532(.A1(new_n729), .A2(new_n730), .B1(new_n731), .B2(new_n733), .ZN(G1337gat));
  OAI21_X1  g533(.A(G99gat), .B1(new_n709), .B2(new_n619), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n479), .A2(new_n542), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n735), .B1(new_n719), .B2(new_n736), .ZN(G1338gat));
  AOI21_X1  g536(.A(new_n543), .B1(new_n708), .B2(new_n447), .ZN(new_n738));
  NOR2_X1   g537(.A1(new_n448), .A2(G106gat), .ZN(new_n739));
  AND4_X1   g538(.A1(new_n722), .A2(new_n716), .A3(new_n717), .A4(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(KEYINPUT53), .B1(new_n738), .B2(new_n740), .ZN(new_n741));
  INV_X1    g540(.A(new_n740), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT53), .ZN(new_n743));
  NOR3_X1   g542(.A1(new_n650), .A2(new_n448), .A3(new_n707), .ZN(new_n744));
  OAI211_X1 g543(.A(new_n742), .B(new_n743), .C1(new_n744), .C2(new_n543), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n741), .A2(new_n745), .ZN(G1339gat));
  AOI21_X1  g545(.A(new_n202), .B1(new_n250), .B2(new_n240), .ZN(new_n747));
  NOR2_X1   g546(.A1(new_n253), .A2(new_n254), .ZN(new_n748));
  OAI21_X1  g547(.A(new_n260), .B1(new_n747), .B2(new_n748), .ZN(new_n749));
  AND2_X1   g548(.A1(new_n264), .A2(new_n749), .ZN(new_n750));
  OAI21_X1  g549(.A(new_n750), .B1(new_n628), .B2(new_n604), .ZN(new_n751));
  NAND3_X1  g550(.A1(new_n579), .A2(new_n584), .A3(new_n581), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n586), .A2(KEYINPUT54), .A3(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(KEYINPUT54), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n591), .B1(new_n598), .B2(new_n754), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(KEYINPUT55), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n753), .A2(new_n755), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT55), .ZN(new_n758));
  NAND2_X1  g557(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND4_X1  g558(.A1(new_n265), .A2(new_n596), .A3(new_n756), .A4(new_n759), .ZN(new_n760));
  AOI21_X1  g559(.A(new_n570), .B1(new_n751), .B2(new_n760), .ZN(new_n761));
  AND2_X1   g560(.A1(new_n596), .A2(new_n756), .ZN(new_n762));
  AND4_X1   g561(.A1(new_n570), .A2(new_n750), .A3(new_n762), .A4(new_n759), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n536), .B1(new_n761), .B2(new_n763), .ZN(new_n764));
  NAND4_X1  g563(.A1(new_n537), .A2(new_n266), .A3(new_n571), .A4(new_n629), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  AND2_X1   g565(.A1(new_n766), .A2(new_n488), .ZN(new_n767));
  NOR2_X1   g566(.A1(new_n695), .A2(new_n420), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(new_n769), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n770), .A2(new_n265), .ZN(new_n771));
  XNOR2_X1  g570(.A(new_n771), .B(G113gat), .ZN(G1340gat));
  AND3_X1   g571(.A1(new_n770), .A2(G120gat), .A3(new_n722), .ZN(new_n773));
  AOI21_X1  g572(.A(G120gat), .B1(new_n770), .B2(new_n607), .ZN(new_n774));
  NOR2_X1   g573(.A1(new_n773), .A2(new_n774), .ZN(G1341gat));
  NAND2_X1  g574(.A1(new_n770), .A2(new_n537), .ZN(new_n776));
  XNOR2_X1  g575(.A(new_n776), .B(G127gat), .ZN(G1342gat));
  NAND3_X1  g576(.A1(new_n570), .A2(new_n632), .A3(new_n492), .ZN(new_n778));
  NOR2_X1   g577(.A1(new_n778), .A2(G134gat), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n767), .A2(new_n779), .ZN(new_n780));
  XOR2_X1   g579(.A(new_n780), .B(KEYINPUT56), .Z(new_n781));
  OAI21_X1  g580(.A(G134gat), .B1(new_n769), .B2(new_n571), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(G1343gat));
  AOI21_X1  g582(.A(new_n448), .B1(new_n764), .B2(new_n765), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n768), .A2(new_n619), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n784), .A2(new_n786), .ZN(new_n787));
  OR2_X1    g586(.A1(new_n266), .A2(G141gat), .ZN(new_n788));
  NOR2_X1   g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  INV_X1    g588(.A(new_n789), .ZN(new_n790));
  OR2_X1    g589(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT57), .ZN(new_n792));
  AOI21_X1  g591(.A(new_n785), .B1(new_n784), .B2(new_n792), .ZN(new_n793));
  AND4_X1   g592(.A1(new_n265), .A2(new_n596), .A3(new_n756), .A4(new_n759), .ZN(new_n794));
  AOI21_X1  g593(.A(new_n794), .B1(new_n751), .B2(KEYINPUT112), .ZN(new_n795));
  INV_X1    g594(.A(KEYINPUT112), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n607), .A2(new_n796), .A3(new_n750), .ZN(new_n797));
  AOI21_X1  g596(.A(new_n570), .B1(new_n795), .B2(new_n797), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n536), .B1(new_n798), .B2(new_n763), .ZN(new_n799));
  AOI21_X1  g598(.A(new_n448), .B1(new_n799), .B2(new_n765), .ZN(new_n800));
  OAI211_X1 g599(.A(new_n265), .B(new_n793), .C1(new_n800), .C2(new_n792), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(G141gat), .ZN(new_n802));
  INV_X1    g601(.A(KEYINPUT58), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n790), .A2(KEYINPUT114), .ZN(new_n804));
  NAND4_X1  g603(.A1(new_n791), .A2(new_n802), .A3(new_n803), .A4(new_n804), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT113), .ZN(new_n806));
  NAND2_X1  g605(.A1(new_n802), .A2(new_n790), .ZN(new_n807));
  AOI21_X1  g606(.A(new_n806), .B1(new_n807), .B2(KEYINPUT58), .ZN(new_n808));
  AOI21_X1  g607(.A(new_n789), .B1(new_n801), .B2(G141gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n809), .A2(KEYINPUT113), .A3(new_n803), .ZN(new_n810));
  OAI21_X1  g609(.A(new_n805), .B1(new_n808), .B2(new_n810), .ZN(G1344gat));
  NAND2_X1  g610(.A1(new_n784), .A2(KEYINPUT57), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n812), .B1(new_n800), .B2(KEYINPUT57), .ZN(new_n813));
  NAND3_X1  g612(.A1(new_n813), .A2(new_n607), .A3(new_n786), .ZN(new_n814));
  NAND3_X1  g613(.A1(new_n814), .A2(KEYINPUT59), .A3(G148gat), .ZN(new_n815));
  INV_X1    g614(.A(G148gat), .ZN(new_n816));
  NAND2_X1  g615(.A1(new_n607), .A2(new_n816), .ZN(new_n817));
  INV_X1    g616(.A(new_n793), .ZN(new_n818));
  INV_X1    g617(.A(new_n800), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n818), .B1(new_n819), .B2(KEYINPUT57), .ZN(new_n820));
  AOI21_X1  g619(.A(new_n816), .B1(new_n820), .B2(new_n607), .ZN(new_n821));
  OAI221_X1 g620(.A(new_n815), .B1(new_n787), .B2(new_n817), .C1(new_n821), .C2(KEYINPUT59), .ZN(G1345gat));
  AOI21_X1  g621(.A(new_n274), .B1(new_n820), .B2(new_n537), .ZN(new_n823));
  NOR3_X1   g622(.A1(new_n787), .A2(G155gat), .A3(new_n536), .ZN(new_n824));
  OR2_X1    g623(.A1(new_n823), .A2(new_n824), .ZN(G1346gat));
  OAI211_X1 g624(.A(new_n570), .B(new_n793), .C1(new_n800), .C2(new_n792), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n275), .B1(new_n826), .B2(KEYINPUT115), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n827), .B1(KEYINPUT115), .B2(new_n826), .ZN(new_n828));
  INV_X1    g627(.A(new_n784), .ZN(new_n829));
  OR3_X1    g628(.A1(new_n485), .A2(new_n778), .A3(G162gat), .ZN(new_n830));
  OAI21_X1  g629(.A(new_n828), .B1(new_n829), .B2(new_n830), .ZN(G1347gat));
  NOR2_X1   g630(.A1(new_n492), .A2(new_n632), .ZN(new_n832));
  AND3_X1   g631(.A1(new_n832), .A2(KEYINPUT118), .A3(new_n479), .ZN(new_n833));
  AOI21_X1  g632(.A(KEYINPUT118), .B1(new_n832), .B2(new_n479), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n833), .A2(new_n834), .A3(new_n447), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n766), .A2(new_n835), .ZN(new_n836));
  NOR3_X1   g635(.A1(new_n836), .A2(new_n343), .A3(new_n266), .ZN(new_n837));
  NOR3_X1   g636(.A1(new_n694), .A2(new_n447), .A3(new_n621), .ZN(new_n838));
  XNOR2_X1  g637(.A(new_n838), .B(KEYINPUT116), .ZN(new_n839));
  AOI21_X1  g638(.A(new_n632), .B1(new_n764), .B2(new_n765), .ZN(new_n840));
  NAND2_X1  g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g640(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n841), .A2(KEYINPUT117), .ZN(new_n843));
  NAND3_X1  g642(.A1(new_n842), .A2(new_n265), .A3(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n837), .B1(new_n844), .B2(new_n343), .ZN(G1348gat));
  NOR3_X1   g644(.A1(new_n836), .A2(new_n344), .A3(new_n651), .ZN(new_n846));
  NAND3_X1  g645(.A1(new_n842), .A2(new_n607), .A3(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(new_n344), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT119), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND3_X1  g649(.A1(new_n847), .A2(KEYINPUT119), .A3(new_n344), .ZN(new_n851));
  AOI21_X1  g650(.A(new_n846), .B1(new_n850), .B2(new_n851), .ZN(G1349gat));
  OAI21_X1  g651(.A(G183gat), .B1(new_n836), .B2(new_n536), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT120), .ZN(new_n854));
  NAND2_X1  g653(.A1(new_n854), .A2(KEYINPUT60), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n537), .A2(new_n349), .ZN(new_n856));
  OAI211_X1 g655(.A(new_n853), .B(new_n855), .C1(new_n841), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g656(.A1(new_n854), .A2(KEYINPUT60), .ZN(new_n858));
  XOR2_X1   g657(.A(new_n857), .B(new_n858), .Z(G1350gat));
  NAND4_X1  g658(.A1(new_n842), .A2(new_n350), .A3(new_n570), .A4(new_n843), .ZN(new_n860));
  INV_X1    g659(.A(KEYINPUT121), .ZN(new_n861));
  XNOR2_X1  g660(.A(new_n860), .B(new_n861), .ZN(new_n862));
  OAI21_X1  g661(.A(G190gat), .B1(new_n836), .B2(new_n571), .ZN(new_n863));
  XNOR2_X1  g662(.A(new_n863), .B(KEYINPUT61), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n862), .A2(new_n864), .ZN(G1351gat));
  INV_X1    g664(.A(G197gat), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n619), .A2(new_n832), .ZN(new_n867));
  XNOR2_X1  g666(.A(new_n867), .B(KEYINPUT124), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n813), .A2(new_n265), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n866), .B1(new_n869), .B2(KEYINPUT125), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n870), .B1(KEYINPUT125), .B2(new_n869), .ZN(new_n871));
  NAND3_X1  g670(.A1(new_n695), .A2(new_n619), .A3(new_n447), .ZN(new_n872));
  XNOR2_X1  g671(.A(new_n872), .B(KEYINPUT122), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n873), .A2(new_n840), .ZN(new_n874));
  INV_X1    g673(.A(new_n874), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n875), .A2(new_n866), .A3(new_n265), .ZN(new_n876));
  XNOR2_X1  g675(.A(new_n876), .B(KEYINPUT123), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n871), .A2(new_n877), .ZN(G1352gat));
  NAND3_X1  g677(.A1(new_n813), .A2(new_n722), .A3(new_n868), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n879), .A2(G204gat), .ZN(new_n880));
  OR3_X1    g679(.A1(new_n874), .A2(G204gat), .A3(new_n629), .ZN(new_n881));
  AND2_X1   g680(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n882));
  NOR2_X1   g681(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n883));
  OAI21_X1  g682(.A(new_n881), .B1(new_n882), .B2(new_n883), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n880), .B(new_n884), .C1(new_n881), .C2(new_n882), .ZN(G1353gat));
  INV_X1    g684(.A(new_n813), .ZN(new_n886));
  NAND3_X1  g685(.A1(new_n619), .A2(new_n537), .A3(new_n832), .ZN(new_n887));
  OAI21_X1  g686(.A(G211gat), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(KEYINPUT63), .ZN(new_n889));
  NOR3_X1   g688(.A1(new_n874), .A2(G211gat), .A3(new_n536), .ZN(new_n890));
  XNOR2_X1  g689(.A(new_n890), .B(KEYINPUT127), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT63), .ZN(new_n892));
  OAI211_X1 g691(.A(new_n892), .B(G211gat), .C1(new_n886), .C2(new_n887), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n889), .A2(new_n891), .A3(new_n893), .ZN(G1354gat));
  INV_X1    g693(.A(G218gat), .ZN(new_n895));
  NAND3_X1  g694(.A1(new_n875), .A2(new_n895), .A3(new_n570), .ZN(new_n896));
  AND3_X1   g695(.A1(new_n813), .A2(new_n570), .A3(new_n868), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n896), .B1(new_n897), .B2(new_n895), .ZN(G1355gat));
endmodule


