//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 0 0 0 0 0 0 0 1 1 0 0 1 0 1 1 1 1 0 0 0 0 1 1 1 1 0 0 0 0 0 0 1 0 1 0 0 1 0 0 1 1 0 0 0 1 1 1 0 0 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:42:29 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n203, new_n204, new_n205, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n232, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n241, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n248, new_n249, new_n250, new_n251, new_n252, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n630, new_n631, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n650, new_n651, new_n652, new_n653, new_n654, new_n655,
    new_n656, new_n657, new_n658, new_n659, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1021,
    new_n1022, new_n1023, new_n1024, new_n1025, new_n1026, new_n1027,
    new_n1028, new_n1029, new_n1030, new_n1031, new_n1032, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1050, new_n1051, new_n1052,
    new_n1053, new_n1054, new_n1055, new_n1056, new_n1057, new_n1058,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1201, new_n1202, new_n1203, new_n1204, new_n1205,
    new_n1206, new_n1207, new_n1208, new_n1210, new_n1211, new_n1213,
    new_n1214, new_n1215, new_n1216, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1259, new_n1260, new_n1261, new_n1262, new_n1263;
  XOR2_X1   g0000(.A(KEYINPUT64), .B(G50), .Z(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  INV_X1    g0002(.A(G58), .ZN(new_n203));
  INV_X1    g0003(.A(G68), .ZN(new_n204));
  NAND2_X1  g0004(.A1(new_n203), .A2(new_n204), .ZN(new_n205));
  NOR3_X1   g0005(.A1(new_n202), .A2(G77), .A3(new_n205), .ZN(G353));
  OAI21_X1  g0006(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0007(.A(G1), .ZN(new_n208));
  INV_X1    g0008(.A(G20), .ZN(new_n209));
  NOR2_X1   g0009(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  INV_X1    g0010(.A(new_n210), .ZN(new_n211));
  AOI22_X1  g0011(.A1(G50), .A2(G226), .B1(G116), .B2(G270), .ZN(new_n212));
  INV_X1    g0012(.A(G238), .ZN(new_n213));
  INV_X1    g0013(.A(G87), .ZN(new_n214));
  INV_X1    g0014(.A(G250), .ZN(new_n215));
  OAI221_X1 g0015(.A(new_n212), .B1(new_n204), .B2(new_n213), .C1(new_n214), .C2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  OAI21_X1  g0019(.A(new_n211), .B1(new_n216), .B2(new_n219), .ZN(new_n220));
  XNOR2_X1  g0020(.A(new_n220), .B(KEYINPUT65), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n221), .A2(KEYINPUT1), .ZN(new_n222));
  XNOR2_X1  g0022(.A(new_n222), .B(KEYINPUT66), .ZN(new_n223));
  NAND2_X1  g0023(.A1(new_n205), .A2(G50), .ZN(new_n224));
  INV_X1    g0024(.A(new_n224), .ZN(new_n225));
  NAND2_X1  g0025(.A1(G1), .A2(G13), .ZN(new_n226));
  NOR2_X1   g0026(.A1(new_n226), .A2(new_n209), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g0028(.A1(new_n211), .A2(G13), .ZN(new_n229));
  OAI211_X1 g0029(.A(new_n229), .B(G250), .C1(G257), .C2(G264), .ZN(new_n230));
  XNOR2_X1  g0030(.A(new_n230), .B(KEYINPUT0), .ZN(new_n231));
  OAI211_X1 g0031(.A(new_n228), .B(new_n231), .C1(new_n221), .C2(KEYINPUT1), .ZN(new_n232));
  NOR2_X1   g0032(.A1(new_n223), .A2(new_n232), .ZN(G361));
  XNOR2_X1  g0033(.A(G238), .B(G244), .ZN(new_n234));
  INV_X1    g0034(.A(G232), .ZN(new_n235));
  XNOR2_X1  g0035(.A(new_n234), .B(new_n235), .ZN(new_n236));
  XNOR2_X1  g0036(.A(KEYINPUT2), .B(G226), .ZN(new_n237));
  XNOR2_X1  g0037(.A(new_n236), .B(new_n237), .ZN(new_n238));
  XOR2_X1   g0038(.A(G264), .B(G270), .Z(new_n239));
  XNOR2_X1  g0039(.A(G250), .B(G257), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n239), .B(new_n240), .ZN(new_n241));
  XOR2_X1   g0041(.A(new_n238), .B(new_n241), .Z(G358));
  XOR2_X1   g0042(.A(G68), .B(G77), .Z(new_n243));
  XOR2_X1   g0043(.A(G50), .B(G58), .Z(new_n244));
  XNOR2_X1  g0044(.A(new_n243), .B(new_n244), .ZN(new_n245));
  INV_X1    g0045(.A(G107), .ZN(new_n246));
  NAND2_X1  g0046(.A1(new_n246), .A2(G97), .ZN(new_n247));
  INV_X1    g0047(.A(G97), .ZN(new_n248));
  NAND2_X1  g0048(.A1(new_n248), .A2(G107), .ZN(new_n249));
  NAND2_X1  g0049(.A1(new_n247), .A2(new_n249), .ZN(new_n250));
  XNOR2_X1  g0050(.A(G87), .B(G116), .ZN(new_n251));
  XNOR2_X1  g0051(.A(new_n250), .B(new_n251), .ZN(new_n252));
  XOR2_X1   g0052(.A(new_n245), .B(new_n252), .Z(G351));
  INV_X1    g0053(.A(G13), .ZN(new_n254));
  NOR3_X1   g0054(.A1(new_n254), .A2(new_n209), .A3(G1), .ZN(new_n255));
  NAND3_X1  g0055(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n256));
  NAND2_X1  g0056(.A1(new_n256), .A2(new_n226), .ZN(new_n257));
  NOR2_X1   g0057(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g0058(.A1(new_n208), .A2(G20), .ZN(new_n259));
  NAND3_X1  g0059(.A1(new_n258), .A2(G50), .A3(new_n259), .ZN(new_n260));
  INV_X1    g0060(.A(new_n255), .ZN(new_n261));
  OAI21_X1  g0061(.A(new_n260), .B1(G50), .B2(new_n261), .ZN(new_n262));
  XNOR2_X1  g0062(.A(new_n262), .B(KEYINPUT69), .ZN(new_n263));
  INV_X1    g0063(.A(new_n205), .ZN(new_n264));
  AOI21_X1  g0064(.A(new_n209), .B1(new_n201), .B2(new_n264), .ZN(new_n265));
  XNOR2_X1  g0065(.A(KEYINPUT8), .B(G58), .ZN(new_n266));
  INV_X1    g0066(.A(G33), .ZN(new_n267));
  NOR2_X1   g0067(.A1(new_n267), .A2(G20), .ZN(new_n268));
  INV_X1    g0068(.A(new_n268), .ZN(new_n269));
  INV_X1    g0069(.A(G150), .ZN(new_n270));
  NOR2_X1   g0070(.A1(G20), .A2(G33), .ZN(new_n271));
  INV_X1    g0071(.A(new_n271), .ZN(new_n272));
  OAI22_X1  g0072(.A1(new_n266), .A2(new_n269), .B1(new_n270), .B2(new_n272), .ZN(new_n273));
  OAI21_X1  g0073(.A(new_n257), .B1(new_n265), .B2(new_n273), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n263), .A2(new_n274), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n275), .B(KEYINPUT9), .ZN(new_n276));
  INV_X1    g0076(.A(new_n226), .ZN(new_n277));
  NAND2_X1  g0077(.A1(G33), .A2(G41), .ZN(new_n278));
  NAND2_X1  g0078(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g0079(.A1(KEYINPUT3), .A2(G33), .ZN(new_n280));
  NOR2_X1   g0080(.A1(KEYINPUT3), .A2(G33), .ZN(new_n281));
  NOR2_X1   g0081(.A1(new_n280), .A2(new_n281), .ZN(new_n282));
  INV_X1    g0082(.A(G1698), .ZN(new_n283));
  NOR2_X1   g0083(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n284), .A2(G223), .B1(G77), .B2(new_n282), .ZN(new_n285));
  INV_X1    g0085(.A(G222), .ZN(new_n286));
  NOR2_X1   g0086(.A1(new_n282), .A2(G1698), .ZN(new_n287));
  INV_X1    g0087(.A(new_n287), .ZN(new_n288));
  OAI21_X1  g0088(.A(new_n285), .B1(new_n286), .B2(new_n288), .ZN(new_n289));
  INV_X1    g0089(.A(KEYINPUT68), .ZN(new_n290));
  AOI21_X1  g0090(.A(new_n279), .B1(new_n289), .B2(new_n290), .ZN(new_n291));
  OAI21_X1  g0091(.A(new_n291), .B1(new_n290), .B2(new_n289), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n279), .A2(G274), .ZN(new_n293));
  OAI21_X1  g0093(.A(new_n208), .B1(G41), .B2(G45), .ZN(new_n294));
  NOR2_X1   g0094(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  OR2_X1    g0095(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n296));
  NAND2_X1  g0096(.A1(new_n294), .A2(KEYINPUT67), .ZN(new_n297));
  NAND3_X1  g0097(.A1(new_n296), .A2(new_n279), .A3(new_n297), .ZN(new_n298));
  INV_X1    g0098(.A(new_n298), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n295), .B1(new_n299), .B2(G226), .ZN(new_n300));
  AND2_X1   g0100(.A1(new_n292), .A2(new_n300), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(G190), .ZN(new_n302));
  INV_X1    g0102(.A(G200), .ZN(new_n303));
  OAI211_X1 g0103(.A(new_n276), .B(new_n302), .C1(new_n303), .C2(new_n301), .ZN(new_n304));
  XNOR2_X1  g0104(.A(new_n304), .B(KEYINPUT10), .ZN(new_n305));
  INV_X1    g0105(.A(G179), .ZN(new_n306));
  NAND2_X1  g0106(.A1(new_n301), .A2(new_n306), .ZN(new_n307));
  OAI211_X1 g0107(.A(new_n307), .B(new_n275), .C1(G169), .C2(new_n301), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n305), .A2(new_n308), .ZN(new_n309));
  INV_X1    g0109(.A(new_n309), .ZN(new_n310));
  OAI21_X1  g0110(.A(KEYINPUT75), .B1(new_n261), .B2(G68), .ZN(new_n311));
  XOR2_X1   g0111(.A(new_n311), .B(KEYINPUT12), .Z(new_n312));
  INV_X1    g0112(.A(G77), .ZN(new_n313));
  OAI22_X1  g0113(.A1(new_n269), .A2(new_n313), .B1(new_n209), .B2(G68), .ZN(new_n314));
  INV_X1    g0114(.A(G50), .ZN(new_n315));
  NOR2_X1   g0115(.A1(new_n272), .A2(new_n315), .ZN(new_n316));
  OAI21_X1  g0116(.A(new_n257), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(KEYINPUT11), .ZN(new_n318));
  OR2_X1    g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND3_X1  g0119(.A1(new_n258), .A2(G68), .A3(new_n259), .ZN(new_n320));
  NAND2_X1  g0120(.A1(new_n317), .A2(new_n318), .ZN(new_n321));
  NAND4_X1  g0121(.A1(new_n312), .A2(new_n319), .A3(new_n320), .A4(new_n321), .ZN(new_n322));
  OAI21_X1  g0122(.A(KEYINPUT73), .B1(new_n267), .B2(new_n248), .ZN(new_n323));
  INV_X1    g0123(.A(KEYINPUT73), .ZN(new_n324));
  NAND3_X1  g0124(.A1(new_n324), .A2(G33), .A3(G97), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n323), .A2(new_n325), .ZN(new_n326));
  AOI21_X1  g0126(.A(new_n326), .B1(new_n284), .B2(G232), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n287), .A2(G226), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n279), .B1(new_n327), .B2(new_n328), .ZN(new_n329));
  OR2_X1    g0129(.A1(new_n293), .A2(new_n294), .ZN(new_n330));
  OAI21_X1  g0130(.A(new_n330), .B1(new_n298), .B2(new_n213), .ZN(new_n331));
  OAI21_X1  g0131(.A(KEYINPUT13), .B1(new_n329), .B2(new_n331), .ZN(new_n332));
  AND2_X1   g0132(.A1(new_n332), .A2(G190), .ZN(new_n333));
  INV_X1    g0133(.A(new_n329), .ZN(new_n334));
  INV_X1    g0134(.A(KEYINPUT13), .ZN(new_n335));
  AOI21_X1  g0135(.A(new_n295), .B1(new_n299), .B2(G238), .ZN(new_n336));
  NAND3_X1  g0136(.A1(new_n334), .A2(new_n335), .A3(new_n336), .ZN(new_n337));
  AOI21_X1  g0137(.A(new_n322), .B1(new_n333), .B2(new_n337), .ZN(new_n338));
  INV_X1    g0138(.A(KEYINPUT74), .ZN(new_n339));
  NAND3_X1  g0139(.A1(new_n337), .A2(new_n339), .A3(new_n332), .ZN(new_n340));
  NAND4_X1  g0140(.A1(new_n334), .A2(KEYINPUT74), .A3(new_n335), .A4(new_n336), .ZN(new_n341));
  NAND3_X1  g0141(.A1(new_n340), .A2(G200), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n338), .A2(new_n342), .ZN(new_n343));
  INV_X1    g0143(.A(new_n343), .ZN(new_n344));
  NAND3_X1  g0144(.A1(new_n340), .A2(G169), .A3(new_n341), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n345), .A2(KEYINPUT14), .ZN(new_n346));
  INV_X1    g0146(.A(KEYINPUT14), .ZN(new_n347));
  NAND4_X1  g0147(.A1(new_n340), .A2(new_n347), .A3(G169), .A4(new_n341), .ZN(new_n348));
  NAND3_X1  g0148(.A1(new_n337), .A2(G179), .A3(new_n332), .ZN(new_n349));
  NAND3_X1  g0149(.A1(new_n346), .A2(new_n348), .A3(new_n349), .ZN(new_n350));
  AOI21_X1  g0150(.A(new_n344), .B1(new_n350), .B2(new_n322), .ZN(new_n351));
  INV_X1    g0151(.A(new_n281), .ZN(new_n352));
  XNOR2_X1  g0152(.A(KEYINPUT76), .B(G33), .ZN(new_n353));
  INV_X1    g0153(.A(KEYINPUT3), .ZN(new_n354));
  OAI21_X1  g0154(.A(new_n352), .B1(new_n353), .B2(new_n354), .ZN(new_n355));
  MUX2_X1   g0155(.A(G223), .B(G226), .S(G1698), .Z(new_n356));
  AOI22_X1  g0156(.A1(new_n355), .A2(new_n356), .B1(G33), .B2(G87), .ZN(new_n357));
  NOR2_X1   g0157(.A1(new_n357), .A2(new_n279), .ZN(new_n358));
  OAI21_X1  g0158(.A(new_n330), .B1(new_n298), .B2(new_n235), .ZN(new_n359));
  NOR2_X1   g0159(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n360), .A2(G179), .ZN(new_n361));
  INV_X1    g0161(.A(G169), .ZN(new_n362));
  OAI21_X1  g0162(.A(new_n361), .B1(new_n362), .B2(new_n360), .ZN(new_n363));
  AOI21_X1  g0163(.A(new_n266), .B1(new_n208), .B2(G20), .ZN(new_n364));
  AOI22_X1  g0164(.A1(new_n364), .A2(new_n258), .B1(new_n255), .B2(new_n266), .ZN(new_n365));
  XNOR2_X1  g0165(.A(G58), .B(G68), .ZN(new_n366));
  AOI22_X1  g0166(.A1(new_n366), .A2(G20), .B1(G159), .B2(new_n271), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n209), .B(new_n352), .C1(new_n353), .C2(new_n354), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n368), .A2(KEYINPUT7), .ZN(new_n369));
  INV_X1    g0169(.A(new_n369), .ZN(new_n370));
  OAI21_X1  g0170(.A(G68), .B1(new_n368), .B2(KEYINPUT7), .ZN(new_n371));
  OAI211_X1 g0171(.A(KEYINPUT16), .B(new_n367), .C1(new_n370), .C2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n372), .A2(new_n257), .ZN(new_n373));
  AOI21_X1  g0173(.A(G20), .B1(KEYINPUT3), .B2(G33), .ZN(new_n374));
  NAND2_X1  g0174(.A1(new_n267), .A2(KEYINPUT76), .ZN(new_n375));
  INV_X1    g0175(.A(KEYINPUT76), .ZN(new_n376));
  NAND2_X1  g0176(.A1(new_n376), .A2(G33), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  OAI211_X1 g0178(.A(KEYINPUT7), .B(new_n374), .C1(new_n378), .C2(KEYINPUT3), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n352), .A2(new_n374), .ZN(new_n380));
  INV_X1    g0180(.A(KEYINPUT7), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n380), .A2(KEYINPUT77), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g0182(.A(KEYINPUT77), .B1(new_n380), .B2(new_n381), .ZN(new_n383));
  OAI21_X1  g0183(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  NAND2_X1  g0184(.A1(new_n384), .A2(G68), .ZN(new_n385));
  AOI21_X1  g0185(.A(KEYINPUT16), .B1(new_n385), .B2(new_n367), .ZN(new_n386));
  OAI21_X1  g0186(.A(new_n365), .B1(new_n373), .B2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n363), .A2(new_n387), .ZN(new_n388));
  NAND2_X1  g0188(.A1(new_n388), .A2(KEYINPUT18), .ZN(new_n389));
  AND2_X1   g0189(.A1(new_n385), .A2(new_n367), .ZN(new_n390));
  OAI211_X1 g0190(.A(new_n257), .B(new_n372), .C1(new_n390), .C2(KEYINPUT16), .ZN(new_n391));
  AOI21_X1  g0191(.A(new_n295), .B1(new_n299), .B2(G232), .ZN(new_n392));
  OAI211_X1 g0192(.A(new_n392), .B(G190), .C1(new_n279), .C2(new_n357), .ZN(new_n393));
  OAI21_X1  g0193(.A(G200), .B1(new_n358), .B2(new_n359), .ZN(new_n394));
  AND2_X1   g0194(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  NAND4_X1  g0195(.A1(new_n391), .A2(new_n395), .A3(KEYINPUT17), .A4(new_n365), .ZN(new_n396));
  INV_X1    g0196(.A(KEYINPUT18), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n363), .A2(new_n387), .A3(new_n397), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT17), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n393), .A2(new_n394), .ZN(new_n400));
  OAI21_X1  g0200(.A(new_n399), .B1(new_n387), .B2(new_n400), .ZN(new_n401));
  NAND4_X1  g0201(.A1(new_n389), .A2(new_n396), .A3(new_n398), .A4(new_n401), .ZN(new_n402));
  INV_X1    g0202(.A(new_n402), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n284), .A2(G238), .B1(G107), .B2(new_n282), .ZN(new_n404));
  OAI21_X1  g0204(.A(new_n404), .B1(new_n235), .B2(new_n288), .ZN(new_n405));
  INV_X1    g0205(.A(new_n279), .ZN(new_n406));
  NAND2_X1  g0206(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  AOI21_X1  g0207(.A(new_n295), .B1(new_n299), .B2(G244), .ZN(new_n408));
  AOI21_X1  g0208(.A(G169), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND3_X1  g0209(.A1(new_n258), .A2(G77), .A3(new_n259), .ZN(new_n410));
  OAI21_X1  g0210(.A(new_n410), .B1(G77), .B2(new_n261), .ZN(new_n411));
  INV_X1    g0211(.A(KEYINPUT70), .ZN(new_n412));
  XNOR2_X1  g0212(.A(new_n266), .B(new_n412), .ZN(new_n413));
  NAND2_X1  g0213(.A1(new_n413), .A2(new_n271), .ZN(new_n414));
  XOR2_X1   g0214(.A(KEYINPUT15), .B(G87), .Z(new_n415));
  AOI22_X1  g0215(.A1(new_n415), .A2(new_n268), .B1(G20), .B2(G77), .ZN(new_n416));
  NAND2_X1  g0216(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g0217(.A(new_n411), .B1(new_n417), .B2(new_n257), .ZN(new_n418));
  OR3_X1    g0218(.A1(new_n409), .A2(KEYINPUT71), .A3(new_n418), .ZN(new_n419));
  AND2_X1   g0219(.A1(new_n407), .A2(new_n408), .ZN(new_n420));
  NAND2_X1  g0220(.A1(new_n420), .A2(new_n306), .ZN(new_n421));
  OAI21_X1  g0221(.A(KEYINPUT71), .B1(new_n409), .B2(new_n418), .ZN(new_n422));
  NAND3_X1  g0222(.A1(new_n419), .A2(new_n421), .A3(new_n422), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n420), .A2(G190), .ZN(new_n424));
  OAI211_X1 g0224(.A(new_n424), .B(new_n418), .C1(new_n303), .C2(new_n420), .ZN(new_n425));
  NAND2_X1  g0225(.A1(new_n423), .A2(new_n425), .ZN(new_n426));
  XOR2_X1   g0226(.A(new_n426), .B(KEYINPUT72), .Z(new_n427));
  NAND4_X1  g0227(.A1(new_n310), .A2(new_n351), .A3(new_n403), .A4(new_n427), .ZN(new_n428));
  INV_X1    g0228(.A(G45), .ZN(new_n429));
  NOR2_X1   g0229(.A1(new_n429), .A2(G1), .ZN(new_n430));
  NOR2_X1   g0230(.A1(new_n430), .A2(new_n215), .ZN(new_n431));
  NAND2_X1  g0231(.A1(new_n431), .A2(new_n279), .ZN(new_n432));
  INV_X1    g0232(.A(new_n430), .ZN(new_n433));
  OAI21_X1  g0233(.A(new_n432), .B1(new_n293), .B2(new_n433), .ZN(new_n434));
  NAND3_X1  g0234(.A1(new_n355), .A2(G238), .A3(new_n283), .ZN(new_n435));
  INV_X1    g0235(.A(G116), .ZN(new_n436));
  AOI21_X1  g0236(.A(new_n436), .B1(new_n375), .B2(new_n377), .ZN(new_n437));
  INV_X1    g0237(.A(new_n437), .ZN(new_n438));
  AOI21_X1  g0238(.A(new_n354), .B1(new_n375), .B2(new_n377), .ZN(new_n439));
  OAI211_X1 g0239(.A(G244), .B(G1698), .C1(new_n439), .C2(new_n281), .ZN(new_n440));
  NAND3_X1  g0240(.A1(new_n435), .A2(new_n438), .A3(new_n440), .ZN(new_n441));
  AOI21_X1  g0241(.A(new_n434), .B1(new_n441), .B2(new_n406), .ZN(new_n442));
  NAND2_X1  g0242(.A1(new_n442), .A2(G190), .ZN(new_n443));
  NOR2_X1   g0243(.A1(new_n261), .A2(new_n415), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n208), .A2(G33), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n258), .A2(new_n445), .ZN(new_n446));
  NOR2_X1   g0246(.A1(new_n446), .A2(new_n214), .ZN(new_n447));
  NAND3_X1  g0247(.A1(new_n355), .A2(new_n209), .A3(G68), .ZN(new_n448));
  OR2_X1    g0248(.A1(new_n214), .A2(KEYINPUT81), .ZN(new_n449));
  NOR2_X1   g0249(.A1(G97), .A2(G107), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n214), .A2(KEYINPUT81), .ZN(new_n451));
  NAND3_X1  g0251(.A1(new_n449), .A2(new_n450), .A3(new_n451), .ZN(new_n452));
  INV_X1    g0252(.A(KEYINPUT19), .ZN(new_n453));
  AOI21_X1  g0253(.A(new_n453), .B1(new_n323), .B2(new_n325), .ZN(new_n454));
  OAI21_X1  g0254(.A(new_n452), .B1(new_n454), .B2(G20), .ZN(new_n455));
  OAI21_X1  g0255(.A(new_n453), .B1(new_n269), .B2(new_n248), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n448), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  AOI211_X1 g0257(.A(new_n444), .B(new_n447), .C1(new_n457), .C2(new_n257), .ZN(new_n458));
  OAI211_X1 g0258(.A(new_n443), .B(new_n458), .C1(new_n303), .C2(new_n442), .ZN(new_n459));
  NAND2_X1  g0259(.A1(new_n442), .A2(new_n306), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n457), .A2(new_n257), .ZN(new_n461));
  INV_X1    g0261(.A(new_n444), .ZN(new_n462));
  INV_X1    g0262(.A(new_n446), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n463), .A2(new_n415), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n461), .A2(new_n462), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g0265(.A(new_n460), .B(new_n465), .C1(G169), .C2(new_n442), .ZN(new_n466));
  INV_X1    g0266(.A(KEYINPUT24), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n437), .A2(new_n209), .ZN(new_n468));
  INV_X1    g0268(.A(KEYINPUT22), .ZN(new_n469));
  NAND2_X1  g0269(.A1(new_n209), .A2(G87), .ZN(new_n470));
  OAI21_X1  g0270(.A(new_n469), .B1(new_n282), .B2(new_n470), .ZN(new_n471));
  INV_X1    g0271(.A(KEYINPUT23), .ZN(new_n472));
  OAI21_X1  g0272(.A(new_n472), .B1(new_n209), .B2(G107), .ZN(new_n473));
  NAND3_X1  g0273(.A1(new_n246), .A2(KEYINPUT23), .A3(G20), .ZN(new_n474));
  NAND2_X1  g0274(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  AND3_X1   g0275(.A1(new_n468), .A2(new_n471), .A3(new_n475), .ZN(new_n476));
  NOR2_X1   g0276(.A1(new_n469), .A2(new_n214), .ZN(new_n477));
  OAI211_X1 g0277(.A(new_n209), .B(new_n477), .C1(new_n439), .C2(new_n281), .ZN(new_n478));
  AOI21_X1  g0278(.A(new_n467), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  AOI22_X1  g0279(.A1(new_n437), .A2(new_n209), .B1(new_n473), .B2(new_n474), .ZN(new_n480));
  NAND3_X1  g0280(.A1(new_n478), .A2(new_n480), .A3(new_n471), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n481), .A2(KEYINPUT24), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n257), .B1(new_n479), .B2(new_n482), .ZN(new_n483));
  OAI211_X1 g0283(.A(G257), .B(G1698), .C1(new_n439), .C2(new_n281), .ZN(new_n484));
  OAI211_X1 g0284(.A(G250), .B(new_n283), .C1(new_n439), .C2(new_n281), .ZN(new_n485));
  NAND2_X1  g0285(.A1(new_n378), .A2(G294), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n484), .A2(new_n485), .A3(new_n486), .ZN(new_n487));
  NAND2_X1  g0287(.A1(new_n487), .A2(new_n406), .ZN(new_n488));
  XNOR2_X1  g0288(.A(KEYINPUT5), .B(G41), .ZN(new_n489));
  NAND4_X1  g0289(.A1(new_n279), .A2(new_n489), .A3(G274), .A4(new_n430), .ZN(new_n490));
  AOI22_X1  g0290(.A1(new_n489), .A2(new_n430), .B1(new_n277), .B2(new_n278), .ZN(new_n491));
  AND2_X1   g0291(.A1(new_n491), .A2(G264), .ZN(new_n492));
  INV_X1    g0292(.A(new_n492), .ZN(new_n493));
  NAND4_X1  g0293(.A1(new_n488), .A2(G190), .A3(new_n490), .A4(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n255), .A2(new_n246), .ZN(new_n495));
  XOR2_X1   g0295(.A(KEYINPUT87), .B(KEYINPUT25), .Z(new_n496));
  XNOR2_X1  g0296(.A(new_n495), .B(new_n496), .ZN(new_n497));
  NOR2_X1   g0297(.A1(new_n446), .A2(new_n246), .ZN(new_n498));
  NOR2_X1   g0298(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND3_X1  g0299(.A1(new_n483), .A2(new_n494), .A3(new_n499), .ZN(new_n500));
  INV_X1    g0300(.A(new_n490), .ZN(new_n501));
  AOI211_X1 g0301(.A(new_n501), .B(new_n492), .C1(new_n487), .C2(new_n406), .ZN(new_n502));
  NOR2_X1   g0302(.A1(new_n502), .A2(new_n303), .ZN(new_n503));
  OAI211_X1 g0303(.A(new_n459), .B(new_n466), .C1(new_n500), .C2(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(new_n504), .ZN(new_n505));
  INV_X1    g0305(.A(KEYINPUT80), .ZN(new_n506));
  OAI211_X1 g0306(.A(G244), .B(new_n283), .C1(new_n439), .C2(new_n281), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(KEYINPUT78), .ZN(new_n508));
  INV_X1    g0308(.A(KEYINPUT4), .ZN(new_n509));
  INV_X1    g0309(.A(KEYINPUT78), .ZN(new_n510));
  NAND4_X1  g0310(.A1(new_n355), .A2(new_n510), .A3(G244), .A4(new_n283), .ZN(new_n511));
  NAND3_X1  g0311(.A1(new_n508), .A2(new_n509), .A3(new_n511), .ZN(new_n512));
  NAND3_X1  g0312(.A1(new_n287), .A2(KEYINPUT4), .A3(G244), .ZN(new_n513));
  NAND2_X1  g0313(.A1(G33), .A2(G283), .ZN(new_n514));
  NAND2_X1  g0314(.A1(new_n284), .A2(G250), .ZN(new_n515));
  AND3_X1   g0315(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND2_X1  g0316(.A1(new_n512), .A2(new_n516), .ZN(new_n517));
  NAND2_X1  g0317(.A1(new_n517), .A2(new_n406), .ZN(new_n518));
  AND2_X1   g0318(.A1(KEYINPUT5), .A2(G41), .ZN(new_n519));
  NOR2_X1   g0319(.A1(KEYINPUT5), .A2(G41), .ZN(new_n520));
  OAI21_X1  g0320(.A(new_n430), .B1(new_n519), .B2(new_n520), .ZN(new_n521));
  NAND3_X1  g0321(.A1(new_n521), .A2(G257), .A3(new_n279), .ZN(new_n522));
  NAND2_X1  g0322(.A1(new_n522), .A2(new_n490), .ZN(new_n523));
  INV_X1    g0323(.A(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n506), .B1(new_n518), .B2(new_n524), .ZN(new_n525));
  AOI21_X1  g0325(.A(new_n279), .B1(new_n512), .B2(new_n516), .ZN(new_n526));
  NOR3_X1   g0326(.A1(new_n526), .A2(KEYINPUT80), .A3(new_n523), .ZN(new_n527));
  OAI21_X1  g0327(.A(G190), .B1(new_n525), .B2(new_n527), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n255), .A2(new_n248), .ZN(new_n529));
  OAI21_X1  g0329(.A(new_n529), .B1(new_n446), .B2(new_n248), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n384), .A2(G107), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT6), .ZN(new_n532));
  NOR2_X1   g0332(.A1(new_n248), .A2(new_n246), .ZN(new_n533));
  OAI21_X1  g0333(.A(new_n532), .B1(new_n533), .B2(new_n450), .ZN(new_n534));
  OAI21_X1  g0334(.A(new_n534), .B1(new_n532), .B2(new_n247), .ZN(new_n535));
  AOI22_X1  g0335(.A1(new_n535), .A2(G20), .B1(G77), .B2(new_n271), .ZN(new_n536));
  NAND2_X1  g0336(.A1(new_n531), .A2(new_n536), .ZN(new_n537));
  AOI21_X1  g0337(.A(new_n530), .B1(new_n537), .B2(new_n257), .ZN(new_n538));
  INV_X1    g0338(.A(KEYINPUT79), .ZN(new_n539));
  XNOR2_X1  g0339(.A(new_n523), .B(new_n539), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n540), .B1(new_n517), .B2(new_n406), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n538), .B1(new_n541), .B2(new_n303), .ZN(new_n542));
  INV_X1    g0342(.A(new_n542), .ZN(new_n543));
  NAND2_X1  g0343(.A1(new_n528), .A2(new_n543), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n518), .A2(new_n506), .A3(new_n524), .ZN(new_n545));
  OAI21_X1  g0345(.A(KEYINPUT80), .B1(new_n526), .B2(new_n523), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n545), .A2(new_n362), .A3(new_n546), .ZN(new_n547));
  AOI21_X1  g0347(.A(new_n538), .B1(new_n541), .B2(new_n306), .ZN(new_n548));
  NAND2_X1  g0348(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND3_X1  g0349(.A1(new_n505), .A2(new_n544), .A3(new_n549), .ZN(new_n550));
  INV_X1    g0350(.A(KEYINPUT82), .ZN(new_n551));
  AOI21_X1  g0351(.A(new_n551), .B1(new_n491), .B2(G270), .ZN(new_n552));
  NAND4_X1  g0352(.A1(new_n521), .A2(new_n551), .A3(G270), .A4(new_n279), .ZN(new_n553));
  NAND2_X1  g0353(.A1(new_n553), .A2(new_n490), .ZN(new_n554));
  OAI21_X1  g0354(.A(KEYINPUT83), .B1(new_n552), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n521), .A2(new_n279), .ZN(new_n556));
  INV_X1    g0356(.A(G270), .ZN(new_n557));
  OAI21_X1  g0357(.A(KEYINPUT82), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  INV_X1    g0358(.A(KEYINPUT83), .ZN(new_n559));
  NAND4_X1  g0359(.A1(new_n558), .A2(new_n559), .A3(new_n490), .A4(new_n553), .ZN(new_n560));
  AND2_X1   g0360(.A1(new_n555), .A2(new_n560), .ZN(new_n561));
  OAI211_X1 g0361(.A(G257), .B(new_n283), .C1(new_n439), .C2(new_n281), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT84), .ZN(new_n563));
  NAND2_X1  g0363(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  NAND4_X1  g0364(.A1(new_n355), .A2(KEYINPUT84), .A3(G257), .A4(new_n283), .ZN(new_n565));
  NAND2_X1  g0365(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  OAI211_X1 g0366(.A(G264), .B(G1698), .C1(new_n439), .C2(new_n281), .ZN(new_n567));
  XNOR2_X1  g0367(.A(KEYINPUT85), .B(G303), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n282), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n567), .A2(new_n569), .ZN(new_n570));
  INV_X1    g0370(.A(new_n570), .ZN(new_n571));
  AOI21_X1  g0371(.A(new_n279), .B1(new_n566), .B2(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(new_n561), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g0373(.A1(new_n573), .A2(G190), .ZN(new_n574));
  OAI21_X1  g0374(.A(G200), .B1(new_n561), .B2(new_n572), .ZN(new_n575));
  OAI211_X1 g0375(.A(new_n514), .B(new_n209), .C1(G33), .C2(new_n248), .ZN(new_n576));
  OAI211_X1 g0376(.A(new_n576), .B(new_n257), .C1(new_n209), .C2(G116), .ZN(new_n577));
  XNOR2_X1  g0377(.A(new_n577), .B(KEYINPUT20), .ZN(new_n578));
  NOR2_X1   g0378(.A1(new_n261), .A2(G116), .ZN(new_n579));
  INV_X1    g0379(.A(new_n579), .ZN(new_n580));
  OAI21_X1  g0380(.A(new_n580), .B1(new_n446), .B2(new_n436), .ZN(new_n581));
  NOR2_X1   g0381(.A1(new_n578), .A2(new_n581), .ZN(new_n582));
  AND3_X1   g0382(.A1(new_n574), .A2(new_n575), .A3(new_n582), .ZN(new_n583));
  NAND4_X1  g0383(.A1(new_n488), .A2(G179), .A3(new_n490), .A4(new_n493), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n584), .B1(new_n502), .B2(new_n362), .ZN(new_n585));
  NAND2_X1  g0385(.A1(new_n483), .A2(new_n499), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  OAI21_X1  g0387(.A(G169), .B1(new_n578), .B2(new_n581), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n566), .A2(new_n571), .ZN(new_n589));
  NAND2_X1  g0389(.A1(new_n589), .A2(new_n406), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n555), .A2(new_n560), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n588), .B1(new_n590), .B2(new_n591), .ZN(new_n592));
  NOR2_X1   g0392(.A1(new_n582), .A2(new_n306), .ZN(new_n593));
  AOI22_X1  g0393(.A1(new_n592), .A2(KEYINPUT21), .B1(new_n573), .B2(new_n593), .ZN(new_n594));
  NOR3_X1   g0394(.A1(new_n592), .A2(KEYINPUT86), .A3(KEYINPUT21), .ZN(new_n595));
  INV_X1    g0395(.A(KEYINPUT86), .ZN(new_n596));
  XOR2_X1   g0396(.A(new_n577), .B(KEYINPUT20), .Z(new_n597));
  AOI21_X1  g0397(.A(new_n579), .B1(new_n463), .B2(G116), .ZN(new_n598));
  AOI21_X1  g0398(.A(new_n362), .B1(new_n597), .B2(new_n598), .ZN(new_n599));
  OAI21_X1  g0399(.A(new_n599), .B1(new_n561), .B2(new_n572), .ZN(new_n600));
  INV_X1    g0400(.A(KEYINPUT21), .ZN(new_n601));
  AOI21_X1  g0401(.A(new_n596), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI211_X1 g0402(.A(new_n587), .B(new_n594), .C1(new_n595), .C2(new_n602), .ZN(new_n603));
  NOR4_X1   g0403(.A1(new_n428), .A2(new_n550), .A3(new_n583), .A4(new_n603), .ZN(G372));
  INV_X1    g0404(.A(new_n428), .ZN(new_n605));
  INV_X1    g0405(.A(KEYINPUT89), .ZN(new_n606));
  OAI21_X1  g0406(.A(new_n594), .B1(new_n595), .B2(new_n602), .ZN(new_n607));
  AND3_X1   g0407(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT88), .ZN(new_n608));
  AOI21_X1  g0408(.A(KEYINPUT88), .B1(new_n585), .B2(new_n586), .ZN(new_n609));
  NOR2_X1   g0409(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n607), .A2(new_n610), .ZN(new_n611));
  OAI21_X1  g0411(.A(new_n606), .B1(new_n611), .B2(new_n550), .ZN(new_n612));
  AND2_X1   g0412(.A1(new_n547), .A2(new_n548), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n459), .A2(new_n466), .ZN(new_n614));
  INV_X1    g0414(.A(new_n614), .ZN(new_n615));
  NAND3_X1  g0415(.A1(new_n613), .A2(KEYINPUT26), .A3(new_n615), .ZN(new_n616));
  INV_X1    g0416(.A(KEYINPUT90), .ZN(new_n617));
  INV_X1    g0417(.A(KEYINPUT26), .ZN(new_n618));
  OAI21_X1  g0418(.A(new_n618), .B1(new_n549), .B2(new_n614), .ZN(new_n619));
  NAND3_X1  g0419(.A1(new_n616), .A2(new_n617), .A3(new_n619), .ZN(new_n620));
  OAI211_X1 g0420(.A(KEYINPUT90), .B(new_n618), .C1(new_n549), .C2(new_n614), .ZN(new_n621));
  AND2_X1   g0421(.A1(new_n621), .A2(new_n466), .ZN(new_n622));
  INV_X1    g0422(.A(KEYINPUT88), .ZN(new_n623));
  AOI211_X1 g0423(.A(new_n306), .B(new_n492), .C1(new_n487), .C2(new_n406), .ZN(new_n624));
  NAND3_X1  g0424(.A1(new_n488), .A2(new_n490), .A3(new_n493), .ZN(new_n625));
  AOI22_X1  g0425(.A1(new_n490), .A2(new_n624), .B1(new_n625), .B2(G169), .ZN(new_n626));
  INV_X1    g0426(.A(new_n499), .ZN(new_n627));
  XNOR2_X1  g0427(.A(new_n481), .B(KEYINPUT24), .ZN(new_n628));
  AOI21_X1  g0428(.A(new_n627), .B1(new_n628), .B2(new_n257), .ZN(new_n629));
  OAI21_X1  g0429(.A(new_n623), .B1(new_n626), .B2(new_n629), .ZN(new_n630));
  NAND3_X1  g0430(.A1(new_n585), .A2(new_n586), .A3(KEYINPUT88), .ZN(new_n631));
  NAND2_X1  g0431(.A1(new_n630), .A2(new_n631), .ZN(new_n632));
  OAI21_X1  g0432(.A(KEYINPUT86), .B1(new_n592), .B2(KEYINPUT21), .ZN(new_n633));
  NAND3_X1  g0433(.A1(new_n600), .A2(new_n596), .A3(new_n601), .ZN(new_n634));
  NAND2_X1  g0434(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  NAND3_X1  g0435(.A1(new_n632), .A2(new_n635), .A3(new_n594), .ZN(new_n636));
  AOI22_X1  g0436(.A1(new_n528), .A2(new_n543), .B1(new_n547), .B2(new_n548), .ZN(new_n637));
  NAND4_X1  g0437(.A1(new_n636), .A2(KEYINPUT89), .A3(new_n637), .A4(new_n505), .ZN(new_n638));
  NAND4_X1  g0438(.A1(new_n612), .A2(new_n620), .A3(new_n622), .A4(new_n638), .ZN(new_n639));
  NAND2_X1  g0439(.A1(new_n605), .A2(new_n639), .ZN(new_n640));
  XNOR2_X1  g0440(.A(new_n640), .B(KEYINPUT91), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n396), .A2(new_n401), .ZN(new_n642));
  OR2_X1    g0442(.A1(new_n344), .A2(new_n423), .ZN(new_n643));
  NAND2_X1  g0443(.A1(new_n350), .A2(new_n322), .ZN(new_n644));
  AOI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n389), .A2(new_n398), .ZN(new_n646));
  OAI21_X1  g0446(.A(new_n305), .B1(new_n645), .B2(new_n646), .ZN(new_n647));
  AND2_X1   g0447(.A1(new_n647), .A2(new_n308), .ZN(new_n648));
  NAND2_X1  g0448(.A1(new_n641), .A2(new_n648), .ZN(G369));
  INV_X1    g0449(.A(new_n587), .ZN(new_n650));
  OR2_X1    g0450(.A1(new_n500), .A2(new_n503), .ZN(new_n651));
  NAND3_X1  g0451(.A1(new_n208), .A2(new_n209), .A3(G13), .ZN(new_n652));
  OR2_X1    g0452(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n653));
  NAND2_X1  g0453(.A1(new_n652), .A2(KEYINPUT27), .ZN(new_n654));
  NAND3_X1  g0454(.A1(new_n653), .A2(G213), .A3(new_n654), .ZN(new_n655));
  INV_X1    g0455(.A(G343), .ZN(new_n656));
  NOR2_X1   g0456(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  NAND2_X1  g0457(.A1(new_n586), .A2(new_n657), .ZN(new_n658));
  AOI21_X1  g0458(.A(new_n650), .B1(new_n651), .B2(new_n658), .ZN(new_n659));
  INV_X1    g0459(.A(new_n657), .ZN(new_n660));
  AOI21_X1  g0460(.A(new_n659), .B1(new_n650), .B2(new_n660), .ZN(new_n661));
  XNOR2_X1  g0461(.A(new_n661), .B(KEYINPUT92), .ZN(new_n662));
  NAND2_X1  g0462(.A1(new_n607), .A2(new_n660), .ZN(new_n663));
  XOR2_X1   g0463(.A(new_n663), .B(KEYINPUT93), .Z(new_n664));
  NAND2_X1  g0464(.A1(new_n662), .A2(new_n664), .ZN(new_n665));
  NAND2_X1  g0465(.A1(new_n610), .A2(new_n660), .ZN(new_n666));
  NAND2_X1  g0466(.A1(new_n665), .A2(new_n666), .ZN(new_n667));
  INV_X1    g0467(.A(new_n667), .ZN(new_n668));
  NOR2_X1   g0468(.A1(new_n582), .A2(new_n660), .ZN(new_n669));
  INV_X1    g0469(.A(new_n607), .ZN(new_n670));
  INV_X1    g0470(.A(new_n583), .ZN(new_n671));
  AOI21_X1  g0471(.A(new_n669), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  AOI21_X1  g0472(.A(new_n672), .B1(new_n670), .B2(new_n669), .ZN(new_n673));
  NAND3_X1  g0473(.A1(new_n662), .A2(G330), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g0474(.A1(new_n668), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g0475(.A(new_n675), .B(KEYINPUT94), .ZN(G399));
  INV_X1    g0476(.A(G41), .ZN(new_n677));
  NAND2_X1  g0477(.A1(new_n229), .A2(new_n677), .ZN(new_n678));
  NOR2_X1   g0478(.A1(new_n452), .A2(G116), .ZN(new_n679));
  NAND3_X1  g0479(.A1(new_n678), .A2(new_n679), .A3(G1), .ZN(new_n680));
  OAI21_X1  g0480(.A(new_n680), .B1(new_n224), .B2(new_n678), .ZN(new_n681));
  XNOR2_X1  g0481(.A(new_n681), .B(KEYINPUT28), .ZN(new_n682));
  INV_X1    g0482(.A(G330), .ZN(new_n683));
  NOR2_X1   g0483(.A1(new_n603), .A2(new_n583), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n545), .A2(new_n546), .ZN(new_n685));
  AOI21_X1  g0485(.A(new_n542), .B1(new_n685), .B2(G190), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n613), .A2(new_n686), .A3(new_n504), .ZN(new_n687));
  NAND3_X1  g0487(.A1(new_n684), .A2(new_n687), .A3(new_n660), .ZN(new_n688));
  INV_X1    g0488(.A(KEYINPUT96), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n688), .A2(new_n689), .ZN(new_n690));
  NAND4_X1  g0490(.A1(new_n684), .A2(new_n687), .A3(KEYINPUT96), .A4(new_n660), .ZN(new_n691));
  NAND2_X1  g0491(.A1(new_n690), .A2(new_n691), .ZN(new_n692));
  NOR3_X1   g0492(.A1(new_n573), .A2(G179), .A3(new_n442), .ZN(new_n693));
  INV_X1    g0493(.A(KEYINPUT95), .ZN(new_n694));
  INV_X1    g0494(.A(new_n541), .ZN(new_n695));
  AOI21_X1  g0495(.A(new_n694), .B1(new_n695), .B2(new_n625), .ZN(new_n696));
  OAI211_X1 g0496(.A(new_n694), .B(new_n625), .C1(new_n526), .C2(new_n540), .ZN(new_n697));
  INV_X1    g0497(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g0498(.A(new_n693), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  AND4_X1   g0499(.A1(new_n442), .A2(new_n590), .A3(new_n591), .A4(new_n624), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n685), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT30), .ZN(new_n702));
  NAND2_X1  g0502(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  NAND3_X1  g0503(.A1(new_n685), .A2(new_n700), .A3(KEYINPUT30), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n699), .A2(new_n703), .A3(new_n704), .ZN(new_n705));
  AND3_X1   g0505(.A1(new_n705), .A2(KEYINPUT31), .A3(new_n657), .ZN(new_n706));
  AOI21_X1  g0506(.A(KEYINPUT31), .B1(new_n705), .B2(new_n657), .ZN(new_n707));
  NOR2_X1   g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g0508(.A(new_n683), .B1(new_n692), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g0509(.A1(new_n639), .A2(new_n660), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT97), .ZN(new_n711));
  INV_X1    g0511(.A(KEYINPUT29), .ZN(new_n712));
  NAND3_X1  g0512(.A1(new_n710), .A2(new_n711), .A3(new_n712), .ZN(new_n713));
  INV_X1    g0513(.A(KEYINPUT99), .ZN(new_n714));
  INV_X1    g0514(.A(new_n603), .ZN(new_n715));
  OAI21_X1  g0515(.A(new_n714), .B1(new_n715), .B2(new_n550), .ZN(new_n716));
  INV_X1    g0516(.A(KEYINPUT98), .ZN(new_n717));
  NOR4_X1   g0517(.A1(new_n549), .A2(new_n614), .A3(new_n717), .A4(new_n618), .ZN(new_n718));
  INV_X1    g0518(.A(new_n466), .ZN(new_n719));
  NOR2_X1   g0519(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND4_X1  g0520(.A1(new_n603), .A2(new_n637), .A3(KEYINPUT99), .A4(new_n505), .ZN(new_n721));
  NAND3_X1  g0521(.A1(new_n616), .A2(new_n717), .A3(new_n619), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n716), .A2(new_n720), .A3(new_n721), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n723), .A2(KEYINPUT29), .A3(new_n660), .ZN(new_n724));
  AND2_X1   g0524(.A1(new_n713), .A2(new_n724), .ZN(new_n725));
  NAND2_X1  g0525(.A1(new_n710), .A2(new_n712), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n726), .A2(KEYINPUT97), .ZN(new_n727));
  AOI21_X1  g0527(.A(new_n709), .B1(new_n725), .B2(new_n727), .ZN(new_n728));
  OAI21_X1  g0528(.A(new_n682), .B1(new_n728), .B2(G1), .ZN(G364));
  INV_X1    g0529(.A(new_n678), .ZN(new_n730));
  NOR2_X1   g0530(.A1(new_n254), .A2(G20), .ZN(new_n731));
  AOI21_X1  g0531(.A(new_n208), .B1(new_n731), .B2(G45), .ZN(new_n732));
  INV_X1    g0532(.A(new_n732), .ZN(new_n733));
  NOR2_X1   g0533(.A1(new_n730), .A2(new_n733), .ZN(new_n734));
  XNOR2_X1  g0534(.A(new_n734), .B(KEYINPUT100), .ZN(new_n735));
  INV_X1    g0535(.A(new_n282), .ZN(new_n736));
  NAND2_X1  g0536(.A1(new_n229), .A2(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(G355), .ZN(new_n738));
  OAI22_X1  g0538(.A1(new_n737), .A2(new_n738), .B1(G116), .B2(new_n229), .ZN(new_n739));
  INV_X1    g0539(.A(new_n355), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n740), .A2(new_n229), .ZN(new_n741));
  AOI21_X1  g0541(.A(new_n741), .B1(new_n429), .B2(new_n225), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n245), .A2(G45), .ZN(new_n743));
  AOI21_X1  g0543(.A(new_n739), .B1(new_n742), .B2(new_n743), .ZN(new_n744));
  NOR2_X1   g0544(.A1(G13), .A2(G33), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR2_X1   g0546(.A1(new_n746), .A2(G20), .ZN(new_n747));
  AOI21_X1  g0547(.A(new_n226), .B1(G20), .B2(new_n362), .ZN(new_n748));
  NOR2_X1   g0548(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  INV_X1    g0549(.A(new_n749), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n735), .B1(new_n744), .B2(new_n750), .ZN(new_n751));
  INV_X1    g0551(.A(G303), .ZN(new_n752));
  INV_X1    g0552(.A(G190), .ZN(new_n753));
  NOR2_X1   g0553(.A1(new_n753), .A2(new_n303), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n209), .A2(G179), .ZN(new_n755));
  NAND2_X1  g0555(.A1(new_n754), .A2(new_n755), .ZN(new_n756));
  NOR2_X1   g0556(.A1(new_n209), .A2(new_n306), .ZN(new_n757));
  NOR2_X1   g0557(.A1(G190), .A2(G200), .ZN(new_n758));
  NAND2_X1  g0558(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  INV_X1    g0559(.A(G311), .ZN(new_n760));
  OAI22_X1  g0560(.A1(new_n752), .A2(new_n756), .B1(new_n759), .B2(new_n760), .ZN(new_n761));
  NAND3_X1  g0561(.A1(new_n755), .A2(new_n753), .A3(G200), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  AND2_X1   g0563(.A1(new_n763), .A2(G283), .ZN(new_n764));
  INV_X1    g0564(.A(new_n757), .ZN(new_n765));
  NOR3_X1   g0565(.A1(new_n765), .A2(new_n303), .A3(G190), .ZN(new_n766));
  XNOR2_X1  g0566(.A(KEYINPUT33), .B(G317), .ZN(new_n767));
  AOI211_X1 g0567(.A(new_n761), .B(new_n764), .C1(new_n766), .C2(new_n767), .ZN(new_n768));
  NOR3_X1   g0568(.A1(new_n753), .A2(G179), .A3(G200), .ZN(new_n769));
  NOR2_X1   g0569(.A1(new_n769), .A2(new_n209), .ZN(new_n770));
  INV_X1    g0570(.A(new_n770), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n771), .A2(G294), .ZN(new_n772));
  NAND2_X1  g0572(.A1(new_n757), .A2(new_n754), .ZN(new_n773));
  INV_X1    g0573(.A(new_n773), .ZN(new_n774));
  AOI21_X1  g0574(.A(new_n736), .B1(new_n774), .B2(G326), .ZN(new_n775));
  NOR3_X1   g0575(.A1(new_n765), .A2(new_n753), .A3(G200), .ZN(new_n776));
  NAND2_X1  g0576(.A1(new_n755), .A2(new_n758), .ZN(new_n777));
  INV_X1    g0577(.A(new_n777), .ZN(new_n778));
  AOI22_X1  g0578(.A1(new_n776), .A2(G322), .B1(G329), .B2(new_n778), .ZN(new_n779));
  NAND4_X1  g0579(.A1(new_n768), .A2(new_n772), .A3(new_n775), .A4(new_n779), .ZN(new_n780));
  NOR2_X1   g0580(.A1(new_n770), .A2(new_n248), .ZN(new_n781));
  AOI21_X1  g0581(.A(new_n781), .B1(G68), .B2(new_n766), .ZN(new_n782));
  XOR2_X1   g0582(.A(new_n782), .B(KEYINPUT101), .Z(new_n783));
  NOR2_X1   g0583(.A1(new_n762), .A2(new_n246), .ZN(new_n784));
  OAI22_X1  g0584(.A1(new_n773), .A2(new_n315), .B1(new_n759), .B2(new_n313), .ZN(new_n785));
  AOI211_X1 g0585(.A(new_n784), .B(new_n785), .C1(G58), .C2(new_n776), .ZN(new_n786));
  INV_X1    g0586(.A(KEYINPUT32), .ZN(new_n787));
  AOI21_X1  g0587(.A(new_n787), .B1(new_n778), .B2(G159), .ZN(new_n788));
  AOI21_X1  g0588(.A(new_n756), .B1(new_n451), .B2(new_n449), .ZN(new_n789));
  INV_X1    g0589(.A(G159), .ZN(new_n790));
  NOR3_X1   g0590(.A1(new_n777), .A2(KEYINPUT32), .A3(new_n790), .ZN(new_n791));
  NOR4_X1   g0591(.A1(new_n788), .A2(new_n789), .A3(new_n791), .A4(new_n282), .ZN(new_n792));
  NAND2_X1  g0592(.A1(new_n786), .A2(new_n792), .ZN(new_n793));
  OAI21_X1  g0593(.A(new_n780), .B1(new_n783), .B2(new_n793), .ZN(new_n794));
  AOI21_X1  g0594(.A(new_n751), .B1(new_n794), .B2(new_n748), .ZN(new_n795));
  INV_X1    g0595(.A(new_n747), .ZN(new_n796));
  OAI21_X1  g0596(.A(new_n795), .B1(new_n673), .B2(new_n796), .ZN(new_n797));
  NAND2_X1  g0597(.A1(new_n673), .A2(G330), .ZN(new_n798));
  OAI21_X1  g0598(.A(new_n798), .B1(new_n730), .B2(new_n733), .ZN(new_n799));
  NOR2_X1   g0599(.A1(new_n673), .A2(G330), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n797), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  XOR2_X1   g0601(.A(new_n801), .B(KEYINPUT102), .Z(new_n802));
  INV_X1    g0602(.A(new_n802), .ZN(G396));
  INV_X1    g0603(.A(new_n748), .ZN(new_n804));
  NAND2_X1  g0604(.A1(new_n804), .A2(new_n746), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n735), .B1(G77), .B2(new_n805), .ZN(new_n806));
  XNOR2_X1  g0606(.A(KEYINPUT103), .B(G283), .ZN(new_n807));
  INV_X1    g0607(.A(new_n807), .ZN(new_n808));
  AOI22_X1  g0608(.A1(new_n766), .A2(new_n808), .B1(new_n774), .B2(G303), .ZN(new_n809));
  OAI21_X1  g0609(.A(new_n809), .B1(new_n436), .B2(new_n759), .ZN(new_n810));
  XOR2_X1   g0610(.A(new_n810), .B(KEYINPUT104), .Z(new_n811));
  NOR2_X1   g0611(.A1(new_n762), .A2(new_n214), .ZN(new_n812));
  NOR3_X1   g0612(.A1(new_n781), .A2(new_n812), .A3(new_n736), .ZN(new_n813));
  AOI22_X1  g0613(.A1(new_n776), .A2(G294), .B1(G311), .B2(new_n778), .ZN(new_n814));
  OAI211_X1 g0614(.A(new_n813), .B(new_n814), .C1(new_n246), .C2(new_n756), .ZN(new_n815));
  AOI22_X1  g0615(.A1(new_n766), .A2(G150), .B1(new_n774), .B2(G137), .ZN(new_n816));
  INV_X1    g0616(.A(new_n776), .ZN(new_n817));
  XNOR2_X1  g0617(.A(KEYINPUT105), .B(G143), .ZN(new_n818));
  OAI221_X1 g0618(.A(new_n816), .B1(new_n790), .B2(new_n759), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  XNOR2_X1  g0619(.A(KEYINPUT106), .B(KEYINPUT34), .ZN(new_n820));
  NAND2_X1  g0620(.A1(new_n819), .A2(new_n820), .ZN(new_n821));
  INV_X1    g0621(.A(G132), .ZN(new_n822));
  NOR2_X1   g0622(.A1(new_n777), .A2(new_n822), .ZN(new_n823));
  NOR2_X1   g0623(.A1(new_n762), .A2(new_n204), .ZN(new_n824));
  INV_X1    g0624(.A(new_n756), .ZN(new_n825));
  AOI211_X1 g0625(.A(new_n823), .B(new_n824), .C1(G50), .C2(new_n825), .ZN(new_n826));
  AOI21_X1  g0626(.A(new_n740), .B1(G58), .B2(new_n771), .ZN(new_n827));
  NAND3_X1  g0627(.A1(new_n821), .A2(new_n826), .A3(new_n827), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n819), .A2(new_n820), .ZN(new_n829));
  OAI22_X1  g0629(.A1(new_n811), .A2(new_n815), .B1(new_n828), .B2(new_n829), .ZN(new_n830));
  AOI21_X1  g0630(.A(new_n806), .B1(new_n830), .B2(new_n748), .ZN(new_n831));
  INV_X1    g0631(.A(KEYINPUT107), .ZN(new_n832));
  OR2_X1    g0632(.A1(new_n418), .A2(new_n660), .ZN(new_n833));
  NOR3_X1   g0633(.A1(new_n423), .A2(new_n832), .A3(new_n833), .ZN(new_n834));
  INV_X1    g0634(.A(new_n834), .ZN(new_n835));
  AND3_X1   g0635(.A1(new_n423), .A2(new_n425), .A3(new_n833), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n832), .B1(new_n423), .B2(new_n833), .ZN(new_n837));
  OAI21_X1  g0637(.A(new_n835), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g0639(.A(new_n831), .B1(new_n839), .B2(new_n746), .ZN(new_n840));
  NAND2_X1  g0640(.A1(new_n710), .A2(new_n838), .ZN(new_n841));
  OAI211_X1 g0641(.A(new_n835), .B(new_n660), .C1(new_n836), .C2(new_n837), .ZN(new_n842));
  INV_X1    g0642(.A(new_n842), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n639), .A2(new_n843), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n841), .A2(new_n844), .ZN(new_n845));
  INV_X1    g0645(.A(new_n709), .ZN(new_n846));
  AOI21_X1  g0646(.A(new_n734), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  INV_X1    g0647(.A(new_n847), .ZN(new_n848));
  NOR2_X1   g0648(.A1(new_n845), .A2(new_n846), .ZN(new_n849));
  OAI21_X1  g0649(.A(new_n840), .B1(new_n848), .B2(new_n849), .ZN(G384));
  OR2_X1    g0650(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n851));
  NAND2_X1  g0651(.A1(new_n535), .A2(KEYINPUT35), .ZN(new_n852));
  NAND4_X1  g0652(.A1(new_n851), .A2(G116), .A3(new_n227), .A4(new_n852), .ZN(new_n853));
  XOR2_X1   g0653(.A(new_n853), .B(KEYINPUT36), .Z(new_n854));
  OAI211_X1 g0654(.A(new_n225), .B(G77), .C1(new_n203), .C2(new_n204), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n201), .A2(G68), .ZN(new_n856));
  AOI211_X1 g0656(.A(new_n208), .B(G13), .C1(new_n855), .C2(new_n856), .ZN(new_n857));
  NOR2_X1   g0657(.A1(new_n854), .A2(new_n857), .ZN(new_n858));
  INV_X1    g0658(.A(KEYINPUT38), .ZN(new_n859));
  INV_X1    g0659(.A(new_n655), .ZN(new_n860));
  AND3_X1   g0660(.A1(new_n402), .A2(new_n387), .A3(new_n860), .ZN(new_n861));
  NAND3_X1  g0661(.A1(new_n391), .A2(new_n395), .A3(new_n365), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n387), .A2(new_n860), .ZN(new_n863));
  NAND3_X1  g0663(.A1(new_n862), .A2(new_n388), .A3(new_n863), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n864), .A2(KEYINPUT37), .ZN(new_n865));
  INV_X1    g0665(.A(KEYINPUT37), .ZN(new_n866));
  NAND4_X1  g0666(.A1(new_n862), .A2(new_n388), .A3(new_n863), .A4(new_n866), .ZN(new_n867));
  AND2_X1   g0667(.A1(new_n865), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g0668(.A(new_n859), .B1(new_n861), .B2(new_n868), .ZN(new_n869));
  INV_X1    g0669(.A(KEYINPUT39), .ZN(new_n870));
  OR2_X1    g0670(.A1(new_n368), .A2(KEYINPUT7), .ZN(new_n871));
  NAND3_X1  g0671(.A1(new_n871), .A2(new_n369), .A3(G68), .ZN(new_n872));
  AOI21_X1  g0672(.A(KEYINPUT16), .B1(new_n872), .B2(new_n367), .ZN(new_n873));
  OAI21_X1  g0673(.A(new_n365), .B1(new_n373), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g0674(.A1(new_n402), .A2(new_n860), .A3(new_n874), .ZN(new_n875));
  NAND2_X1  g0675(.A1(new_n874), .A2(new_n363), .ZN(new_n876));
  NAND2_X1  g0676(.A1(new_n874), .A2(new_n860), .ZN(new_n877));
  AND3_X1   g0677(.A1(new_n862), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  OAI21_X1  g0678(.A(new_n867), .B1(new_n878), .B2(new_n866), .ZN(new_n879));
  NAND3_X1  g0679(.A1(new_n875), .A2(new_n879), .A3(KEYINPUT38), .ZN(new_n880));
  NAND3_X1  g0680(.A1(new_n869), .A2(new_n870), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g0681(.A1(new_n881), .A2(KEYINPUT109), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n881), .A2(KEYINPUT109), .ZN(new_n883));
  INV_X1    g0683(.A(new_n880), .ZN(new_n884));
  AOI21_X1  g0684(.A(KEYINPUT38), .B1(new_n875), .B2(new_n879), .ZN(new_n885));
  OAI21_X1  g0685(.A(KEYINPUT39), .B1(new_n884), .B2(new_n885), .ZN(new_n886));
  AOI21_X1  g0686(.A(new_n882), .B1(new_n883), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g0687(.A1(new_n644), .A2(new_n657), .ZN(new_n888));
  AOI22_X1  g0688(.A1(new_n887), .A2(new_n888), .B1(new_n646), .B2(new_n655), .ZN(new_n889));
  NAND2_X1  g0689(.A1(new_n322), .A2(new_n657), .ZN(new_n890));
  NAND2_X1  g0690(.A1(new_n351), .A2(new_n890), .ZN(new_n891));
  OAI211_X1 g0691(.A(new_n322), .B(new_n657), .C1(new_n350), .C2(new_n344), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g0693(.A1(new_n423), .A2(new_n657), .ZN(new_n894));
  INV_X1    g0694(.A(new_n894), .ZN(new_n895));
  AOI21_X1  g0695(.A(KEYINPUT108), .B1(new_n844), .B2(new_n895), .ZN(new_n896));
  INV_X1    g0696(.A(KEYINPUT108), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n897), .B(new_n894), .C1(new_n639), .C2(new_n843), .ZN(new_n898));
  OAI221_X1 g0698(.A(new_n893), .B1(new_n884), .B2(new_n885), .C1(new_n896), .C2(new_n898), .ZN(new_n899));
  NAND2_X1  g0699(.A1(new_n889), .A2(new_n899), .ZN(new_n900));
  NAND4_X1  g0700(.A1(new_n727), .A2(new_n605), .A3(new_n724), .A4(new_n713), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n901), .A2(new_n648), .ZN(new_n902));
  XNOR2_X1  g0702(.A(new_n900), .B(new_n902), .ZN(new_n903));
  NAND2_X1  g0703(.A1(new_n692), .A2(new_n708), .ZN(new_n904));
  NAND2_X1  g0704(.A1(new_n869), .A2(new_n880), .ZN(new_n905));
  NAND2_X1  g0705(.A1(new_n839), .A2(new_n893), .ZN(new_n906));
  INV_X1    g0706(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g0707(.A1(new_n904), .A2(new_n905), .A3(new_n907), .ZN(new_n908));
  NAND2_X1  g0708(.A1(new_n908), .A2(KEYINPUT40), .ZN(new_n909));
  AOI21_X1  g0709(.A(new_n906), .B1(new_n692), .B2(new_n708), .ZN(new_n910));
  NOR2_X1   g0710(.A1(new_n884), .A2(new_n885), .ZN(new_n911));
  NOR2_X1   g0711(.A1(new_n911), .A2(KEYINPUT40), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n910), .A2(new_n912), .ZN(new_n913));
  NAND2_X1  g0713(.A1(new_n909), .A2(new_n913), .ZN(new_n914));
  AOI21_X1  g0714(.A(new_n428), .B1(new_n692), .B2(new_n708), .ZN(new_n915));
  AOI21_X1  g0715(.A(new_n683), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g0716(.A(new_n916), .B1(new_n915), .B2(new_n914), .ZN(new_n917));
  NAND2_X1  g0717(.A1(new_n903), .A2(new_n917), .ZN(new_n918));
  OAI21_X1  g0718(.A(new_n918), .B1(new_n208), .B2(new_n731), .ZN(new_n919));
  NOR2_X1   g0719(.A1(new_n903), .A2(new_n917), .ZN(new_n920));
  OAI21_X1  g0720(.A(new_n858), .B1(new_n919), .B2(new_n920), .ZN(G367));
  AND2_X1   g0721(.A1(new_n662), .A2(new_n664), .ZN(new_n922));
  OAI21_X1  g0722(.A(new_n637), .B1(new_n538), .B2(new_n660), .ZN(new_n923));
  NAND2_X1  g0723(.A1(new_n613), .A2(new_n657), .ZN(new_n924));
  NAND2_X1  g0724(.A1(new_n923), .A2(new_n924), .ZN(new_n925));
  NAND3_X1  g0725(.A1(new_n922), .A2(KEYINPUT42), .A3(new_n925), .ZN(new_n926));
  INV_X1    g0726(.A(KEYINPUT42), .ZN(new_n927));
  INV_X1    g0727(.A(new_n925), .ZN(new_n928));
  OAI21_X1  g0728(.A(new_n927), .B1(new_n665), .B2(new_n928), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n926), .A2(new_n929), .ZN(new_n930));
  OAI21_X1  g0730(.A(new_n549), .B1(new_n686), .B2(new_n587), .ZN(new_n931));
  NAND2_X1  g0731(.A1(new_n931), .A2(new_n660), .ZN(new_n932));
  NAND2_X1  g0732(.A1(new_n930), .A2(new_n932), .ZN(new_n933));
  INV_X1    g0733(.A(new_n933), .ZN(new_n934));
  NOR2_X1   g0734(.A1(new_n458), .A2(new_n660), .ZN(new_n935));
  NAND2_X1  g0735(.A1(new_n719), .A2(new_n935), .ZN(new_n936));
  OAI21_X1  g0736(.A(new_n936), .B1(new_n614), .B2(new_n935), .ZN(new_n937));
  XOR2_X1   g0737(.A(new_n937), .B(KEYINPUT43), .Z(new_n938));
  INV_X1    g0738(.A(new_n938), .ZN(new_n939));
  OAI21_X1  g0739(.A(KEYINPUT110), .B1(new_n934), .B2(new_n939), .ZN(new_n940));
  OR3_X1    g0740(.A1(new_n933), .A2(KEYINPUT43), .A3(new_n937), .ZN(new_n941));
  INV_X1    g0741(.A(KEYINPUT110), .ZN(new_n942));
  NAND3_X1  g0742(.A1(new_n933), .A2(new_n942), .A3(new_n938), .ZN(new_n943));
  NAND3_X1  g0743(.A1(new_n940), .A2(new_n941), .A3(new_n943), .ZN(new_n944));
  NOR2_X1   g0744(.A1(new_n674), .A2(new_n928), .ZN(new_n945));
  XNOR2_X1  g0745(.A(new_n944), .B(new_n945), .ZN(new_n946));
  XNOR2_X1  g0746(.A(new_n678), .B(KEYINPUT41), .ZN(new_n947));
  XOR2_X1   g0747(.A(KEYINPUT111), .B(KEYINPUT44), .Z(new_n948));
  NAND2_X1  g0748(.A1(new_n667), .A2(new_n928), .ZN(new_n949));
  AOI21_X1  g0749(.A(new_n948), .B1(new_n949), .B2(KEYINPUT112), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n950), .B1(KEYINPUT112), .B2(new_n949), .ZN(new_n951));
  NOR2_X1   g0751(.A1(new_n667), .A2(new_n928), .ZN(new_n952));
  XNOR2_X1  g0752(.A(new_n952), .B(KEYINPUT45), .ZN(new_n953));
  INV_X1    g0753(.A(KEYINPUT112), .ZN(new_n954));
  NAND4_X1  g0754(.A1(new_n667), .A2(new_n954), .A3(new_n928), .A4(new_n948), .ZN(new_n955));
  NAND3_X1  g0755(.A1(new_n951), .A2(new_n953), .A3(new_n955), .ZN(new_n956));
  INV_X1    g0756(.A(new_n674), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NOR2_X1   g0758(.A1(new_n662), .A2(new_n664), .ZN(new_n959));
  NOR2_X1   g0759(.A1(new_n922), .A2(new_n959), .ZN(new_n960));
  XNOR2_X1  g0760(.A(new_n960), .B(new_n798), .ZN(new_n961));
  NAND4_X1  g0761(.A1(new_n951), .A2(new_n953), .A3(new_n674), .A4(new_n955), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n728), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  AOI21_X1  g0763(.A(new_n947), .B1(new_n963), .B2(new_n728), .ZN(new_n964));
  OAI21_X1  g0764(.A(new_n946), .B1(new_n964), .B2(new_n733), .ZN(new_n965));
  INV_X1    g0765(.A(new_n415), .ZN(new_n966));
  OAI221_X1 g0766(.A(new_n749), .B1(new_n229), .B2(new_n966), .C1(new_n741), .C2(new_n241), .ZN(new_n967));
  AND2_X1   g0767(.A1(new_n735), .A2(new_n967), .ZN(new_n968));
  OAI22_X1  g0768(.A1(new_n313), .A2(new_n762), .B1(new_n756), .B2(new_n203), .ZN(new_n969));
  AOI211_X1 g0769(.A(new_n282), .B(new_n969), .C1(G159), .C2(new_n766), .ZN(new_n970));
  INV_X1    g0770(.A(new_n759), .ZN(new_n971));
  AOI22_X1  g0771(.A1(new_n776), .A2(G150), .B1(new_n202), .B2(new_n971), .ZN(new_n972));
  INV_X1    g0772(.A(new_n818), .ZN(new_n973));
  AOI22_X1  g0773(.A1(new_n774), .A2(new_n973), .B1(new_n778), .B2(G137), .ZN(new_n974));
  NOR2_X1   g0774(.A1(new_n770), .A2(new_n204), .ZN(new_n975));
  INV_X1    g0775(.A(new_n975), .ZN(new_n976));
  NAND4_X1  g0776(.A1(new_n970), .A2(new_n972), .A3(new_n974), .A4(new_n976), .ZN(new_n977));
  INV_X1    g0777(.A(new_n568), .ZN(new_n978));
  OAI22_X1  g0778(.A1(new_n817), .A2(new_n978), .B1(new_n759), .B2(new_n807), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n355), .B(new_n979), .C1(G107), .C2(new_n771), .ZN(new_n980));
  NAND3_X1  g0780(.A1(new_n825), .A2(KEYINPUT46), .A3(G116), .ZN(new_n981));
  INV_X1    g0781(.A(KEYINPUT46), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n982), .B1(new_n756), .B2(new_n436), .ZN(new_n983));
  INV_X1    g0783(.A(new_n766), .ZN(new_n984));
  INV_X1    g0784(.A(G294), .ZN(new_n985));
  OAI211_X1 g0785(.A(new_n981), .B(new_n983), .C1(new_n984), .C2(new_n985), .ZN(new_n986));
  INV_X1    g0786(.A(KEYINPUT113), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n986), .A2(new_n987), .ZN(new_n988));
  OAI22_X1  g0788(.A1(new_n760), .A2(new_n773), .B1(new_n762), .B2(new_n248), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n989), .B1(G317), .B2(new_n778), .ZN(new_n990));
  NAND3_X1  g0790(.A1(new_n980), .A2(new_n988), .A3(new_n990), .ZN(new_n991));
  NOR2_X1   g0791(.A1(new_n986), .A2(new_n987), .ZN(new_n992));
  OAI21_X1  g0792(.A(new_n977), .B1(new_n991), .B2(new_n992), .ZN(new_n993));
  XOR2_X1   g0793(.A(new_n993), .B(KEYINPUT47), .Z(new_n994));
  OAI221_X1 g0794(.A(new_n968), .B1(new_n796), .B2(new_n937), .C1(new_n994), .C2(new_n804), .ZN(new_n995));
  NAND2_X1  g0795(.A1(new_n965), .A2(new_n995), .ZN(G387));
  INV_X1    g0796(.A(new_n735), .ZN(new_n997));
  AOI22_X1  g0797(.A1(new_n776), .A2(G317), .B1(new_n568), .B2(new_n971), .ZN(new_n998));
  AOI22_X1  g0798(.A1(new_n766), .A2(G311), .B1(new_n774), .B2(G322), .ZN(new_n999));
  AND2_X1   g0799(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  OR2_X1    g0800(.A1(new_n1000), .A2(KEYINPUT48), .ZN(new_n1001));
  NAND3_X1  g0801(.A1(new_n998), .A2(new_n999), .A3(KEYINPUT48), .ZN(new_n1002));
  AOI22_X1  g0802(.A1(new_n771), .A2(new_n808), .B1(new_n825), .B2(G294), .ZN(new_n1003));
  NAND3_X1  g0803(.A1(new_n1001), .A2(new_n1002), .A3(new_n1003), .ZN(new_n1004));
  INV_X1    g0804(.A(KEYINPUT49), .ZN(new_n1005));
  OR2_X1    g0805(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g0806(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1007));
  AOI22_X1  g0807(.A1(new_n763), .A2(G116), .B1(new_n778), .B2(G326), .ZN(new_n1008));
  NAND4_X1  g0808(.A1(new_n1006), .A2(new_n740), .A3(new_n1007), .A4(new_n1008), .ZN(new_n1009));
  AOI22_X1  g0809(.A1(G159), .A2(new_n774), .B1(new_n971), .B2(G68), .ZN(new_n1010));
  OAI21_X1  g0810(.A(new_n1010), .B1(new_n266), .B2(new_n984), .ZN(new_n1011));
  AOI22_X1  g0811(.A1(G77), .A2(new_n825), .B1(new_n778), .B2(G150), .ZN(new_n1012));
  AOI21_X1  g0812(.A(new_n1011), .B1(KEYINPUT115), .B2(new_n1012), .ZN(new_n1013));
  OAI22_X1  g0813(.A1(new_n817), .A2(new_n315), .B1(new_n762), .B2(new_n248), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n966), .A2(new_n770), .ZN(new_n1015));
  NOR3_X1   g0815(.A1(new_n1014), .A2(new_n1015), .A3(new_n740), .ZN(new_n1016));
  OAI211_X1 g0816(.A(new_n1013), .B(new_n1016), .C1(KEYINPUT115), .C2(new_n1012), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n804), .B1(new_n1009), .B2(new_n1017), .ZN(new_n1018));
  AOI21_X1  g0818(.A(new_n741), .B1(new_n238), .B2(G45), .ZN(new_n1019));
  OAI211_X1 g0819(.A(new_n679), .B(new_n429), .C1(new_n204), .C2(new_n313), .ZN(new_n1020));
  XNOR2_X1  g0820(.A(new_n1020), .B(KEYINPUT114), .ZN(new_n1021));
  NAND2_X1  g0821(.A1(new_n413), .A2(new_n315), .ZN(new_n1022));
  XNOR2_X1  g0822(.A(new_n1022), .B(KEYINPUT50), .ZN(new_n1023));
  OAI21_X1  g0823(.A(new_n1019), .B1(new_n1021), .B2(new_n1023), .ZN(new_n1024));
  OAI221_X1 g0824(.A(new_n1024), .B1(G107), .B2(new_n229), .C1(new_n679), .C2(new_n737), .ZN(new_n1025));
  AOI211_X1 g0825(.A(new_n997), .B(new_n1018), .C1(new_n749), .C2(new_n1025), .ZN(new_n1026));
  OAI21_X1  g0826(.A(new_n1026), .B1(new_n662), .B2(new_n796), .ZN(new_n1027));
  XNOR2_X1  g0827(.A(new_n1027), .B(KEYINPUT116), .ZN(new_n1028));
  AOI21_X1  g0828(.A(new_n1028), .B1(new_n961), .B2(new_n733), .ZN(new_n1029));
  NAND2_X1  g0829(.A1(new_n961), .A2(new_n728), .ZN(new_n1030));
  NAND2_X1  g0830(.A1(new_n1030), .A2(new_n730), .ZN(new_n1031));
  NOR2_X1   g0831(.A1(new_n961), .A2(new_n728), .ZN(new_n1032));
  OAI21_X1  g0832(.A(new_n1029), .B1(new_n1031), .B2(new_n1032), .ZN(G393));
  NAND2_X1  g0833(.A1(new_n958), .A2(new_n962), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n1030), .ZN(new_n1035));
  NAND3_X1  g0835(.A1(new_n1035), .A2(new_n730), .A3(new_n963), .ZN(new_n1036));
  NAND3_X1  g0836(.A1(new_n958), .A2(new_n733), .A3(new_n962), .ZN(new_n1037));
  OAI221_X1 g0837(.A(new_n749), .B1(new_n248), .B2(new_n229), .C1(new_n741), .C2(new_n252), .ZN(new_n1038));
  NAND2_X1  g0838(.A1(new_n735), .A2(new_n1038), .ZN(new_n1039));
  OAI22_X1  g0839(.A1(new_n984), .A2(new_n201), .B1(new_n756), .B2(new_n204), .ZN(new_n1040));
  AOI211_X1 g0840(.A(new_n812), .B(new_n1040), .C1(new_n778), .C2(new_n973), .ZN(new_n1041));
  AOI22_X1  g0841(.A1(new_n776), .A2(G159), .B1(new_n774), .B2(G150), .ZN(new_n1042));
  XOR2_X1   g0842(.A(new_n1042), .B(KEYINPUT51), .Z(new_n1043));
  NAND2_X1  g0843(.A1(new_n413), .A2(new_n971), .ZN(new_n1044));
  NOR2_X1   g0844(.A1(new_n770), .A2(new_n313), .ZN(new_n1045));
  NOR2_X1   g0845(.A1(new_n740), .A2(new_n1045), .ZN(new_n1046));
  NAND4_X1  g0846(.A1(new_n1041), .A2(new_n1043), .A3(new_n1044), .A4(new_n1046), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n825), .A2(new_n808), .B1(new_n778), .B2(G322), .ZN(new_n1048));
  OAI211_X1 g0848(.A(new_n1048), .B(new_n282), .C1(new_n246), .C2(new_n762), .ZN(new_n1049));
  XOR2_X1   g0849(.A(new_n1049), .B(KEYINPUT118), .Z(new_n1050));
  AOI22_X1  g0850(.A1(new_n766), .A2(new_n568), .B1(G294), .B2(new_n971), .ZN(new_n1051));
  OAI211_X1 g0851(.A(new_n1050), .B(new_n1051), .C1(new_n436), .C2(new_n770), .ZN(new_n1052));
  AOI22_X1  g0852(.A1(new_n776), .A2(G311), .B1(new_n774), .B2(G317), .ZN(new_n1053));
  XNOR2_X1  g0853(.A(new_n1053), .B(KEYINPUT117), .ZN(new_n1054));
  XNOR2_X1  g0854(.A(new_n1054), .B(KEYINPUT52), .ZN(new_n1055));
  OAI21_X1  g0855(.A(new_n1047), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1039), .B1(new_n1056), .B2(new_n748), .ZN(new_n1057));
  OAI21_X1  g0857(.A(new_n1057), .B1(new_n925), .B2(new_n796), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1036), .A2(new_n1037), .A3(new_n1058), .ZN(G390));
  NAND2_X1  g0859(.A1(new_n709), .A2(new_n907), .ZN(new_n1060));
  NAND3_X1  g0860(.A1(new_n723), .A2(new_n660), .A3(new_n839), .ZN(new_n1061));
  NAND2_X1  g0861(.A1(new_n1061), .A2(new_n895), .ZN(new_n1062));
  AND3_X1   g0862(.A1(new_n891), .A2(KEYINPUT119), .A3(new_n892), .ZN(new_n1063));
  AOI21_X1  g0863(.A(KEYINPUT119), .B1(new_n891), .B2(new_n892), .ZN(new_n1064));
  NOR2_X1   g0864(.A1(new_n1063), .A2(new_n1064), .ZN(new_n1065));
  INV_X1    g0865(.A(new_n1065), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n1062), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g0867(.A(new_n888), .ZN(new_n1068));
  NAND3_X1  g0868(.A1(new_n1067), .A2(new_n1068), .A3(new_n905), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n844), .A2(new_n895), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n1070), .A2(new_n897), .ZN(new_n1071));
  NAND3_X1  g0871(.A1(new_n844), .A2(KEYINPUT108), .A3(new_n895), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1073));
  AOI21_X1  g0873(.A(new_n888), .B1(new_n1073), .B2(new_n893), .ZN(new_n1074));
  OAI211_X1 g0874(.A(new_n1060), .B(new_n1069), .C1(new_n1074), .C2(new_n887), .ZN(new_n1075));
  INV_X1    g0875(.A(new_n1060), .ZN(new_n1076));
  OAI21_X1  g0876(.A(new_n893), .B1(new_n896), .B2(new_n898), .ZN(new_n1077));
  AOI21_X1  g0877(.A(new_n887), .B1(new_n1077), .B2(new_n1068), .ZN(new_n1078));
  INV_X1    g0878(.A(new_n1069), .ZN(new_n1079));
  OAI21_X1  g0879(.A(new_n1076), .B1(new_n1078), .B2(new_n1079), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1075), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g0881(.A1(new_n605), .A2(new_n709), .ZN(new_n1082));
  AND3_X1   g0882(.A1(new_n901), .A2(new_n648), .A3(new_n1082), .ZN(new_n1083));
  AOI211_X1 g0883(.A(new_n683), .B(new_n838), .C1(new_n692), .C2(new_n708), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n1060), .B1(new_n1084), .B2(new_n893), .ZN(new_n1085));
  NAND2_X1  g0885(.A1(new_n1085), .A2(new_n1073), .ZN(new_n1086));
  AOI21_X1  g0886(.A(new_n1062), .B1(new_n709), .B2(new_n907), .ZN(new_n1087));
  NAND3_X1  g0887(.A1(new_n904), .A2(G330), .A3(new_n839), .ZN(new_n1088));
  NAND2_X1  g0888(.A1(new_n1088), .A2(new_n1065), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n1087), .A2(new_n1089), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n1086), .A2(new_n1090), .ZN(new_n1091));
  NAND2_X1  g0891(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1092));
  NAND2_X1  g0892(.A1(new_n1081), .A2(new_n1092), .ZN(new_n1093));
  AOI22_X1  g0893(.A1(new_n1085), .A2(new_n1073), .B1(new_n1087), .B2(new_n1089), .ZN(new_n1094));
  NAND3_X1  g0894(.A1(new_n901), .A2(new_n1082), .A3(new_n648), .ZN(new_n1095));
  NOR2_X1   g0895(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g0896(.A1(new_n1096), .A2(new_n1075), .A3(new_n1080), .ZN(new_n1097));
  NAND3_X1  g0897(.A1(new_n1093), .A2(new_n730), .A3(new_n1097), .ZN(new_n1098));
  NAND3_X1  g0898(.A1(new_n1075), .A2(new_n1080), .A3(new_n733), .ZN(new_n1099));
  INV_X1    g0899(.A(new_n266), .ZN(new_n1100));
  OAI21_X1  g0900(.A(new_n735), .B1(new_n1100), .B2(new_n805), .ZN(new_n1101));
  NOR2_X1   g0901(.A1(new_n756), .A2(new_n270), .ZN(new_n1102));
  XOR2_X1   g0902(.A(KEYINPUT120), .B(KEYINPUT53), .Z(new_n1103));
  XNOR2_X1  g0903(.A(new_n1102), .B(new_n1103), .ZN(new_n1104));
  NAND2_X1  g0904(.A1(new_n774), .A2(G128), .ZN(new_n1105));
  XOR2_X1   g0905(.A(KEYINPUT54), .B(G143), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n766), .A2(G137), .B1(new_n971), .B2(new_n1106), .ZN(new_n1107));
  NAND3_X1  g0907(.A1(new_n1104), .A2(new_n1105), .A3(new_n1107), .ZN(new_n1108));
  NOR2_X1   g0908(.A1(new_n770), .A2(new_n790), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n736), .B1(new_n201), .B2(new_n762), .ZN(new_n1110));
  INV_X1    g0910(.A(G125), .ZN(new_n1111));
  OAI22_X1  g0911(.A1(new_n817), .A2(new_n822), .B1(new_n777), .B2(new_n1111), .ZN(new_n1112));
  NOR4_X1   g0912(.A1(new_n1108), .A2(new_n1109), .A3(new_n1110), .A4(new_n1112), .ZN(new_n1113));
  INV_X1    g0913(.A(new_n1113), .ZN(new_n1114));
  OR2_X1    g0914(.A1(new_n1114), .A2(KEYINPUT121), .ZN(new_n1115));
  OAI21_X1  g0915(.A(new_n282), .B1(new_n756), .B2(new_n214), .ZN(new_n1116));
  XOR2_X1   g0916(.A(new_n1116), .B(KEYINPUT122), .Z(new_n1117));
  AOI211_X1 g0917(.A(new_n824), .B(new_n1045), .C1(G283), .C2(new_n774), .ZN(new_n1118));
  AOI22_X1  g0918(.A1(new_n766), .A2(G107), .B1(G97), .B2(new_n971), .ZN(new_n1119));
  AOI22_X1  g0919(.A1(new_n776), .A2(G116), .B1(G294), .B2(new_n778), .ZN(new_n1120));
  NAND4_X1  g0920(.A1(new_n1117), .A2(new_n1118), .A3(new_n1119), .A4(new_n1120), .ZN(new_n1121));
  NAND2_X1  g0921(.A1(new_n1114), .A2(KEYINPUT121), .ZN(new_n1122));
  NAND3_X1  g0922(.A1(new_n1115), .A2(new_n1121), .A3(new_n1122), .ZN(new_n1123));
  AOI21_X1  g0923(.A(new_n1101), .B1(new_n1123), .B2(new_n748), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n887), .B2(new_n746), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n1098), .A2(new_n1099), .A3(new_n1125), .ZN(G378));
  XNOR2_X1  g0926(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1127));
  INV_X1    g0927(.A(new_n1127), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n275), .A2(new_n860), .ZN(new_n1129));
  NAND3_X1  g0929(.A1(new_n305), .A2(new_n308), .A3(new_n1129), .ZN(new_n1130));
  INV_X1    g0930(.A(new_n1130), .ZN(new_n1131));
  AOI21_X1  g0931(.A(new_n1129), .B1(new_n305), .B2(new_n308), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1128), .B1(new_n1131), .B2(new_n1132), .ZN(new_n1133));
  INV_X1    g0933(.A(new_n1132), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n1130), .A3(new_n1127), .ZN(new_n1135));
  NAND2_X1  g0935(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n1136), .B1(new_n914), .B2(G330), .ZN(new_n1137));
  AOI22_X1  g0937(.A1(new_n908), .A2(KEYINPUT40), .B1(new_n910), .B2(new_n912), .ZN(new_n1138));
  AND2_X1   g0938(.A1(new_n1133), .A2(new_n1135), .ZN(new_n1139));
  NOR3_X1   g0939(.A1(new_n1138), .A2(new_n1139), .A3(new_n683), .ZN(new_n1140));
  OAI21_X1  g0940(.A(new_n900), .B1(new_n1137), .B2(new_n1140), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n914), .A2(G330), .A3(new_n1136), .ZN(new_n1142));
  OAI21_X1  g0942(.A(new_n1139), .B1(new_n1138), .B2(new_n683), .ZN(new_n1143));
  NAND4_X1  g0943(.A1(new_n1142), .A2(new_n1143), .A3(new_n899), .A4(new_n889), .ZN(new_n1144));
  NAND2_X1  g0944(.A1(new_n1141), .A2(new_n1144), .ZN(new_n1145));
  NAND2_X1  g0945(.A1(new_n1145), .A2(new_n733), .ZN(new_n1146));
  OAI21_X1  g0946(.A(new_n734), .B1(new_n202), .B2(new_n805), .ZN(new_n1147));
  INV_X1    g0947(.A(G137), .ZN(new_n1148));
  OAI22_X1  g0948(.A1(new_n773), .A2(new_n1111), .B1(new_n759), .B2(new_n1148), .ZN(new_n1149));
  AOI22_X1  g0949(.A1(G128), .A2(new_n776), .B1(new_n766), .B2(G132), .ZN(new_n1150));
  OAI21_X1  g0950(.A(new_n1150), .B1(new_n270), .B2(new_n770), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1149), .B(new_n1151), .C1(new_n825), .C2(new_n1106), .ZN(new_n1152));
  INV_X1    g0952(.A(KEYINPUT59), .ZN(new_n1153));
  OR2_X1    g0953(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  NAND2_X1  g0954(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1155));
  OAI211_X1 g0955(.A(new_n267), .B(new_n677), .C1(new_n762), .C2(new_n790), .ZN(new_n1156));
  AOI21_X1  g0956(.A(new_n1156), .B1(G124), .B2(new_n778), .ZN(new_n1157));
  NAND3_X1  g0957(.A1(new_n1154), .A2(new_n1155), .A3(new_n1157), .ZN(new_n1158));
  AOI22_X1  g0958(.A1(new_n763), .A2(G58), .B1(new_n778), .B2(G283), .ZN(new_n1159));
  OAI221_X1 g0959(.A(new_n1159), .B1(new_n313), .B2(new_n756), .C1(new_n246), .C2(new_n817), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n766), .A2(G97), .B1(new_n774), .B2(G116), .ZN(new_n1161));
  OAI21_X1  g0961(.A(new_n1161), .B1(new_n966), .B2(new_n759), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n740), .A2(new_n677), .ZN(new_n1163));
  NOR4_X1   g0963(.A1(new_n1160), .A2(new_n1162), .A3(new_n975), .A4(new_n1163), .ZN(new_n1164));
  OR2_X1    g0964(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1164), .A2(KEYINPUT58), .ZN(new_n1166));
  OAI211_X1 g0966(.A(new_n1163), .B(new_n315), .C1(G33), .C2(G41), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1158), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(new_n1147), .B1(new_n1168), .B2(new_n748), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n1136), .B2(new_n746), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1146), .A2(new_n1170), .ZN(new_n1171));
  INV_X1    g0971(.A(new_n1171), .ZN(new_n1172));
  INV_X1    g0972(.A(KEYINPUT123), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1095), .B(new_n1173), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1097), .A2(new_n1174), .ZN(new_n1175));
  INV_X1    g0975(.A(KEYINPUT57), .ZN(new_n1176));
  AOI21_X1  g0976(.A(new_n1176), .B1(new_n1141), .B2(new_n1144), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1175), .A2(new_n1177), .ZN(new_n1178));
  INV_X1    g0978(.A(KEYINPUT124), .ZN(new_n1179));
  NAND2_X1  g0979(.A1(new_n1178), .A2(new_n1179), .ZN(new_n1180));
  NAND3_X1  g0980(.A1(new_n1175), .A2(KEYINPUT124), .A3(new_n1177), .ZN(new_n1181));
  NAND2_X1  g0981(.A1(new_n1180), .A2(new_n1181), .ZN(new_n1182));
  AOI22_X1  g0982(.A1(new_n1097), .A2(new_n1174), .B1(new_n1144), .B2(new_n1141), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n730), .B1(new_n1183), .B2(KEYINPUT57), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n1172), .B1(new_n1182), .B2(new_n1184), .ZN(G375));
  NAND2_X1  g0985(.A1(new_n1065), .A2(new_n745), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n735), .B1(G68), .B2(new_n805), .ZN(new_n1187));
  OAI22_X1  g0987(.A1(new_n773), .A2(new_n822), .B1(new_n759), .B2(new_n270), .ZN(new_n1188));
  AOI21_X1  g0988(.A(new_n1188), .B1(G137), .B2(new_n776), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n740), .B1(G50), .B2(new_n771), .ZN(new_n1190));
  AOI22_X1  g0990(.A1(new_n766), .A2(new_n1106), .B1(G58), .B2(new_n763), .ZN(new_n1191));
  AOI22_X1  g0991(.A1(G159), .A2(new_n825), .B1(new_n778), .B2(G128), .ZN(new_n1192));
  NAND4_X1  g0992(.A1(new_n1189), .A2(new_n1190), .A3(new_n1191), .A4(new_n1192), .ZN(new_n1193));
  OAI22_X1  g0993(.A1(new_n984), .A2(new_n436), .B1(new_n773), .B2(new_n985), .ZN(new_n1194));
  AOI21_X1  g0994(.A(new_n1194), .B1(G107), .B2(new_n971), .ZN(new_n1195));
  XNOR2_X1  g0995(.A(new_n1195), .B(KEYINPUT125), .ZN(new_n1196));
  AOI21_X1  g0996(.A(new_n1015), .B1(G283), .B2(new_n776), .ZN(new_n1197));
  OR2_X1    g0997(.A1(new_n1197), .A2(KEYINPUT126), .ZN(new_n1198));
  NAND2_X1  g0998(.A1(new_n1197), .A2(KEYINPUT126), .ZN(new_n1199));
  OAI22_X1  g0999(.A1(new_n756), .A2(new_n248), .B1(new_n777), .B2(new_n752), .ZN(new_n1200));
  AOI211_X1 g1000(.A(new_n736), .B(new_n1200), .C1(G77), .C2(new_n763), .ZN(new_n1201));
  NAND3_X1  g1001(.A1(new_n1198), .A2(new_n1199), .A3(new_n1201), .ZN(new_n1202));
  OAI21_X1  g1002(.A(new_n1193), .B1(new_n1196), .B2(new_n1202), .ZN(new_n1203));
  AOI21_X1  g1003(.A(new_n1187), .B1(new_n1203), .B2(new_n748), .ZN(new_n1204));
  AOI22_X1  g1004(.A1(new_n1091), .A2(new_n733), .B1(new_n1186), .B2(new_n1204), .ZN(new_n1205));
  INV_X1    g1005(.A(new_n947), .ZN(new_n1206));
  NAND2_X1  g1006(.A1(new_n1092), .A2(new_n1206), .ZN(new_n1207));
  NOR2_X1   g1007(.A1(new_n1083), .A2(new_n1091), .ZN(new_n1208));
  OAI21_X1  g1008(.A(new_n1205), .B1(new_n1207), .B2(new_n1208), .ZN(G381));
  OR2_X1    g1009(.A1(G393), .A2(G396), .ZN(new_n1210));
  OR4_X1    g1010(.A1(G384), .A2(G390), .A3(new_n1210), .A4(G381), .ZN(new_n1211));
  OR4_X1    g1011(.A1(G387), .A2(new_n1211), .A3(G378), .A4(G375), .ZN(G407));
  INV_X1    g1012(.A(G378), .ZN(new_n1213));
  NAND2_X1  g1013(.A1(new_n656), .A2(G213), .ZN(new_n1214));
  INV_X1    g1014(.A(new_n1214), .ZN(new_n1215));
  NAND2_X1  g1015(.A1(new_n1213), .A2(new_n1215), .ZN(new_n1216));
  OAI211_X1 g1016(.A(G407), .B(G213), .C1(G375), .C2(new_n1216), .ZN(G409));
  INV_X1    g1017(.A(G390), .ZN(new_n1218));
  NAND2_X1  g1018(.A1(G387), .A2(new_n1218), .ZN(new_n1219));
  XNOR2_X1  g1019(.A(G393), .B(new_n802), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(G390), .A2(new_n965), .A3(new_n995), .ZN(new_n1221));
  AND3_X1   g1021(.A1(new_n1219), .A2(new_n1220), .A3(new_n1221), .ZN(new_n1222));
  AOI21_X1  g1022(.A(new_n1220), .B1(new_n1219), .B2(new_n1221), .ZN(new_n1223));
  NOR2_X1   g1023(.A1(new_n1222), .A2(new_n1223), .ZN(new_n1224));
  INV_X1    g1024(.A(KEYINPUT63), .ZN(new_n1225));
  OAI211_X1 g1025(.A(G378), .B(new_n1172), .C1(new_n1182), .C2(new_n1184), .ZN(new_n1226));
  AND2_X1   g1026(.A1(new_n1183), .A2(new_n1206), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1213), .B1(new_n1171), .B2(new_n1227), .ZN(new_n1228));
  NAND2_X1  g1028(.A1(new_n1226), .A2(new_n1228), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1229), .A2(new_n1214), .ZN(new_n1230));
  AOI21_X1  g1030(.A(new_n1208), .B1(KEYINPUT60), .B2(new_n1092), .ZN(new_n1231));
  NAND3_X1  g1031(.A1(new_n1094), .A2(new_n1095), .A3(KEYINPUT60), .ZN(new_n1232));
  NAND2_X1  g1032(.A1(new_n1232), .A2(new_n730), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1205), .B1(new_n1231), .B2(new_n1233), .ZN(new_n1234));
  INV_X1    g1034(.A(G384), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n1234), .A2(new_n1235), .ZN(new_n1236));
  OAI211_X1 g1036(.A(G384), .B(new_n1205), .C1(new_n1231), .C2(new_n1233), .ZN(new_n1237));
  NAND2_X1  g1037(.A1(new_n1236), .A2(new_n1237), .ZN(new_n1238));
  OAI21_X1  g1038(.A(new_n1225), .B1(new_n1230), .B2(new_n1238), .ZN(new_n1239));
  NAND2_X1  g1039(.A1(new_n1215), .A2(KEYINPUT127), .ZN(new_n1240));
  NAND3_X1  g1040(.A1(new_n1236), .A2(new_n1237), .A3(new_n1240), .ZN(new_n1241));
  NAND3_X1  g1041(.A1(new_n1241), .A2(G2897), .A3(new_n1215), .ZN(new_n1242));
  NAND2_X1  g1042(.A1(new_n1215), .A2(G2897), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1236), .A2(new_n1237), .A3(new_n1243), .A4(new_n1240), .ZN(new_n1244));
  AND2_X1   g1044(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1245));
  AOI21_X1  g1045(.A(KEYINPUT61), .B1(new_n1230), .B2(new_n1245), .ZN(new_n1246));
  AOI21_X1  g1046(.A(new_n1215), .B1(new_n1226), .B2(new_n1228), .ZN(new_n1247));
  INV_X1    g1047(.A(new_n1238), .ZN(new_n1248));
  NAND3_X1  g1048(.A1(new_n1247), .A2(KEYINPUT63), .A3(new_n1248), .ZN(new_n1249));
  NAND4_X1  g1049(.A1(new_n1224), .A2(new_n1239), .A3(new_n1246), .A4(new_n1249), .ZN(new_n1250));
  INV_X1    g1050(.A(KEYINPUT62), .ZN(new_n1251));
  AND3_X1   g1051(.A1(new_n1247), .A2(new_n1251), .A3(new_n1248), .ZN(new_n1252));
  INV_X1    g1052(.A(KEYINPUT61), .ZN(new_n1253));
  NAND2_X1  g1053(.A1(new_n1242), .A2(new_n1244), .ZN(new_n1254));
  OAI21_X1  g1054(.A(new_n1253), .B1(new_n1247), .B2(new_n1254), .ZN(new_n1255));
  AOI21_X1  g1055(.A(new_n1251), .B1(new_n1247), .B2(new_n1248), .ZN(new_n1256));
  NOR3_X1   g1056(.A1(new_n1252), .A2(new_n1255), .A3(new_n1256), .ZN(new_n1257));
  OAI21_X1  g1057(.A(new_n1250), .B1(new_n1257), .B2(new_n1224), .ZN(G405));
  NAND2_X1  g1058(.A1(G375), .A2(new_n1213), .ZN(new_n1259));
  NAND3_X1  g1059(.A1(new_n1259), .A2(new_n1238), .A3(new_n1226), .ZN(new_n1260));
  INV_X1    g1060(.A(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1238), .B1(new_n1259), .B2(new_n1226), .ZN(new_n1262));
  NOR2_X1   g1062(.A1(new_n1261), .A2(new_n1262), .ZN(new_n1263));
  XNOR2_X1  g1063(.A(new_n1263), .B(new_n1224), .ZN(G402));
endmodule


