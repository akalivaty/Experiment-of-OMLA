

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588;

  XNOR2_X1 U323 ( .A(n350), .B(n349), .ZN(n355) );
  XNOR2_X1 U324 ( .A(KEYINPUT48), .B(KEYINPUT113), .ZN(n425) );
  XOR2_X1 U325 ( .A(G36GAT), .B(G190GAT), .Z(n339) );
  XNOR2_X1 U326 ( .A(KEYINPUT54), .B(KEYINPUT118), .ZN(n427) );
  XNOR2_X1 U327 ( .A(n348), .B(n386), .ZN(n349) );
  XNOR2_X1 U328 ( .A(n426), .B(n425), .ZN(n535) );
  XNOR2_X1 U329 ( .A(n428), .B(n427), .ZN(n429) );
  XOR2_X1 U330 ( .A(n378), .B(n377), .Z(n567) );
  XNOR2_X1 U331 ( .A(KEYINPUT94), .B(n475), .ZN(n523) );
  XNOR2_X1 U332 ( .A(n461), .B(n460), .ZN(n462) );
  XNOR2_X1 U333 ( .A(n463), .B(n462), .ZN(G1351GAT) );
  XOR2_X1 U334 ( .A(G155GAT), .B(G204GAT), .Z(n292) );
  XNOR2_X1 U335 ( .A(KEYINPUT91), .B(G211GAT), .ZN(n291) );
  XNOR2_X1 U336 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U337 ( .A(n293), .B(G148GAT), .Z(n295) );
  XOR2_X1 U338 ( .A(G106GAT), .B(G78GAT), .Z(n392) );
  XNOR2_X1 U339 ( .A(G22GAT), .B(n392), .ZN(n294) );
  XNOR2_X1 U340 ( .A(n295), .B(n294), .ZN(n300) );
  XNOR2_X1 U341 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n296), .B(KEYINPUT88), .ZN(n325) );
  XOR2_X1 U343 ( .A(G50GAT), .B(G218GAT), .Z(n340) );
  XOR2_X1 U344 ( .A(n325), .B(n340), .Z(n298) );
  NAND2_X1 U345 ( .A1(G228GAT), .A2(G233GAT), .ZN(n297) );
  XNOR2_X1 U346 ( .A(n298), .B(n297), .ZN(n299) );
  XOR2_X1 U347 ( .A(n300), .B(n299), .Z(n308) );
  XOR2_X1 U348 ( .A(KEYINPUT2), .B(G162GAT), .Z(n302) );
  XNOR2_X1 U349 ( .A(KEYINPUT3), .B(KEYINPUT89), .ZN(n301) );
  XNOR2_X1 U350 ( .A(n302), .B(n301), .ZN(n303) );
  XOR2_X1 U351 ( .A(G141GAT), .B(n303), .Z(n313) );
  XOR2_X1 U352 ( .A(KEYINPUT90), .B(KEYINPUT23), .Z(n305) );
  XNOR2_X1 U353 ( .A(KEYINPUT24), .B(KEYINPUT22), .ZN(n304) );
  XNOR2_X1 U354 ( .A(n305), .B(n304), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n313), .B(n306), .ZN(n307) );
  XNOR2_X1 U356 ( .A(n308), .B(n307), .ZN(n478) );
  XOR2_X1 U357 ( .A(G29GAT), .B(G134GAT), .Z(n353) );
  XNOR2_X1 U358 ( .A(G1GAT), .B(G127GAT), .ZN(n309) );
  XNOR2_X1 U359 ( .A(n309), .B(G155GAT), .ZN(n404) );
  XOR2_X1 U360 ( .A(n353), .B(n404), .Z(n311) );
  NAND2_X1 U361 ( .A1(G225GAT), .A2(G233GAT), .ZN(n310) );
  XNOR2_X1 U362 ( .A(n311), .B(n310), .ZN(n312) );
  XNOR2_X1 U363 ( .A(n313), .B(n312), .ZN(n324) );
  XOR2_X1 U364 ( .A(KEYINPUT6), .B(KEYINPUT5), .Z(n315) );
  XNOR2_X1 U365 ( .A(KEYINPUT1), .B(KEYINPUT92), .ZN(n314) );
  XNOR2_X1 U366 ( .A(n315), .B(n314), .ZN(n316) );
  XOR2_X1 U367 ( .A(n316), .B(KEYINPUT93), .Z(n318) );
  XOR2_X1 U368 ( .A(G120GAT), .B(G148GAT), .Z(n385) );
  XNOR2_X1 U369 ( .A(n385), .B(G85GAT), .ZN(n317) );
  XNOR2_X1 U370 ( .A(n318), .B(n317), .ZN(n319) );
  XOR2_X1 U371 ( .A(n319), .B(G57GAT), .Z(n322) );
  XNOR2_X1 U372 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n320) );
  XNOR2_X1 U373 ( .A(n320), .B(KEYINPUT84), .ZN(n439) );
  XNOR2_X1 U374 ( .A(n439), .B(KEYINPUT4), .ZN(n321) );
  XNOR2_X1 U375 ( .A(n322), .B(n321), .ZN(n323) );
  XNOR2_X1 U376 ( .A(n324), .B(n323), .ZN(n475) );
  XNOR2_X1 U377 ( .A(G218GAT), .B(n325), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n326), .B(KEYINPUT95), .ZN(n327) );
  XOR2_X1 U379 ( .A(n339), .B(n327), .Z(n329) );
  NAND2_X1 U380 ( .A1(G226GAT), .A2(G233GAT), .ZN(n328) );
  XNOR2_X1 U381 ( .A(n329), .B(n328), .ZN(n333) );
  XOR2_X1 U382 ( .A(KEYINPUT73), .B(G64GAT), .Z(n331) );
  XNOR2_X1 U383 ( .A(G204GAT), .B(G92GAT), .ZN(n330) );
  XNOR2_X1 U384 ( .A(n331), .B(n330), .ZN(n332) );
  XOR2_X1 U385 ( .A(G176GAT), .B(n332), .Z(n391) );
  XOR2_X1 U386 ( .A(n333), .B(n391), .Z(n338) );
  XOR2_X1 U387 ( .A(KEYINPUT19), .B(KEYINPUT18), .Z(n335) );
  XNOR2_X1 U388 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n334) );
  XNOR2_X1 U389 ( .A(n335), .B(n334), .ZN(n440) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(G183GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n336), .B(G211GAT), .ZN(n403) );
  XNOR2_X1 U392 ( .A(n440), .B(n403), .ZN(n337) );
  XNOR2_X1 U393 ( .A(n338), .B(n337), .ZN(n526) );
  XOR2_X1 U394 ( .A(KEYINPUT11), .B(n339), .Z(n342) );
  XNOR2_X1 U395 ( .A(n340), .B(G106GAT), .ZN(n341) );
  XNOR2_X1 U396 ( .A(n342), .B(n341), .ZN(n344) );
  INV_X1 U397 ( .A(KEYINPUT76), .ZN(n343) );
  XNOR2_X1 U398 ( .A(n344), .B(n343), .ZN(n350) );
  XOR2_X1 U399 ( .A(KEYINPUT75), .B(KEYINPUT78), .Z(n346) );
  XNOR2_X1 U400 ( .A(KEYINPUT9), .B(KEYINPUT77), .ZN(n345) );
  XNOR2_X1 U401 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U402 ( .A(G162GAT), .B(n347), .Z(n348) );
  XOR2_X1 U403 ( .A(G99GAT), .B(G85GAT), .Z(n386) );
  XOR2_X1 U404 ( .A(G43GAT), .B(KEYINPUT7), .Z(n352) );
  XNOR2_X1 U405 ( .A(KEYINPUT8), .B(KEYINPUT67), .ZN(n351) );
  XNOR2_X1 U406 ( .A(n352), .B(n351), .ZN(n370) );
  XNOR2_X1 U407 ( .A(n370), .B(n353), .ZN(n354) );
  XNOR2_X1 U408 ( .A(n355), .B(n354), .ZN(n360) );
  XOR2_X1 U409 ( .A(KEYINPUT10), .B(G92GAT), .Z(n357) );
  NAND2_X1 U410 ( .A1(G232GAT), .A2(G233GAT), .ZN(n356) );
  XNOR2_X1 U411 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U412 ( .A(KEYINPUT64), .B(n358), .Z(n359) );
  XNOR2_X1 U413 ( .A(n360), .B(n359), .ZN(n561) );
  XOR2_X1 U414 ( .A(KEYINPUT69), .B(KEYINPUT65), .Z(n362) );
  XNOR2_X1 U415 ( .A(G113GAT), .B(G1GAT), .ZN(n361) );
  XNOR2_X1 U416 ( .A(n362), .B(n361), .ZN(n378) );
  XOR2_X1 U417 ( .A(G141GAT), .B(G197GAT), .Z(n364) );
  XNOR2_X1 U418 ( .A(G169GAT), .B(G50GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n364), .B(n363), .ZN(n366) );
  XOR2_X1 U420 ( .A(G29GAT), .B(G36GAT), .Z(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n374) );
  XNOR2_X1 U422 ( .A(KEYINPUT29), .B(KEYINPUT66), .ZN(n367) );
  XNOR2_X1 U423 ( .A(n367), .B(G8GAT), .ZN(n368) );
  XOR2_X1 U424 ( .A(n368), .B(KEYINPUT30), .Z(n372) );
  XNOR2_X1 U425 ( .A(G22GAT), .B(G15GAT), .ZN(n369) );
  XNOR2_X1 U426 ( .A(n369), .B(KEYINPUT68), .ZN(n405) );
  XNOR2_X1 U427 ( .A(n370), .B(n405), .ZN(n371) );
  XNOR2_X1 U428 ( .A(n372), .B(n371), .ZN(n373) );
  XNOR2_X1 U429 ( .A(n374), .B(n373), .ZN(n376) );
  NAND2_X1 U430 ( .A1(G229GAT), .A2(G233GAT), .ZN(n375) );
  XNOR2_X1 U431 ( .A(n376), .B(n375), .ZN(n377) );
  XOR2_X1 U432 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n384) );
  XNOR2_X1 U433 ( .A(G71GAT), .B(G57GAT), .ZN(n379) );
  XNOR2_X1 U434 ( .A(n379), .B(KEYINPUT13), .ZN(n402) );
  XOR2_X1 U435 ( .A(KEYINPUT72), .B(KEYINPUT32), .Z(n381) );
  XNOR2_X1 U436 ( .A(KEYINPUT70), .B(KEYINPUT31), .ZN(n380) );
  XNOR2_X1 U437 ( .A(n381), .B(n380), .ZN(n382) );
  XNOR2_X1 U438 ( .A(n402), .B(n382), .ZN(n383) );
  XNOR2_X1 U439 ( .A(n384), .B(n383), .ZN(n390) );
  XOR2_X1 U440 ( .A(n386), .B(n385), .Z(n388) );
  NAND2_X1 U441 ( .A1(G230GAT), .A2(G233GAT), .ZN(n387) );
  XNOR2_X1 U442 ( .A(n388), .B(n387), .ZN(n389) );
  XOR2_X1 U443 ( .A(n390), .B(n389), .Z(n394) );
  XNOR2_X1 U444 ( .A(n392), .B(n391), .ZN(n393) );
  XNOR2_X1 U445 ( .A(n394), .B(n393), .ZN(n576) );
  XNOR2_X1 U446 ( .A(KEYINPUT41), .B(n576), .ZN(n554) );
  NAND2_X1 U447 ( .A1(n567), .A2(n554), .ZN(n395) );
  XNOR2_X1 U448 ( .A(KEYINPUT46), .B(n395), .ZN(n414) );
  XOR2_X1 U449 ( .A(KEYINPUT79), .B(KEYINPUT80), .Z(n397) );
  XNOR2_X1 U450 ( .A(KEYINPUT15), .B(KEYINPUT83), .ZN(n396) );
  XNOR2_X1 U451 ( .A(n397), .B(n396), .ZN(n413) );
  XOR2_X1 U452 ( .A(KEYINPUT81), .B(KEYINPUT12), .Z(n399) );
  XNOR2_X1 U453 ( .A(KEYINPUT82), .B(KEYINPUT14), .ZN(n398) );
  XNOR2_X1 U454 ( .A(n399), .B(n398), .ZN(n401) );
  XOR2_X1 U455 ( .A(G78GAT), .B(G64GAT), .Z(n400) );
  XNOR2_X1 U456 ( .A(n401), .B(n400), .ZN(n409) );
  XOR2_X1 U457 ( .A(n403), .B(n402), .Z(n407) );
  XNOR2_X1 U458 ( .A(n405), .B(n404), .ZN(n406) );
  XNOR2_X1 U459 ( .A(n407), .B(n406), .ZN(n408) );
  XNOR2_X1 U460 ( .A(n409), .B(n408), .ZN(n411) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n410) );
  XNOR2_X1 U462 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U463 ( .A(n413), .B(n412), .ZN(n581) );
  XNOR2_X1 U464 ( .A(KEYINPUT111), .B(n581), .ZN(n543) );
  NAND2_X1 U465 ( .A1(n414), .A2(n543), .ZN(n415) );
  NOR2_X1 U466 ( .A1(n561), .A2(n415), .ZN(n416) );
  XOR2_X1 U467 ( .A(KEYINPUT47), .B(n416), .Z(n424) );
  INV_X1 U468 ( .A(n581), .ZN(n495) );
  XNOR2_X1 U469 ( .A(KEYINPUT36), .B(KEYINPUT103), .ZN(n417) );
  XNOR2_X1 U470 ( .A(n417), .B(n561), .ZN(n586) );
  NOR2_X1 U471 ( .A1(n495), .A2(n586), .ZN(n418) );
  XNOR2_X1 U472 ( .A(KEYINPUT45), .B(n418), .ZN(n421) );
  INV_X1 U473 ( .A(n576), .ZN(n419) );
  NOR2_X1 U474 ( .A1(n567), .A2(n419), .ZN(n420) );
  AND2_X1 U475 ( .A1(n421), .A2(n420), .ZN(n422) );
  XNOR2_X1 U476 ( .A(KEYINPUT112), .B(n422), .ZN(n423) );
  NOR2_X1 U477 ( .A1(n424), .A2(n423), .ZN(n426) );
  NAND2_X1 U478 ( .A1(n526), .A2(n535), .ZN(n428) );
  NOR2_X1 U479 ( .A1(n523), .A2(n429), .ZN(n575) );
  NAND2_X1 U480 ( .A1(n478), .A2(n575), .ZN(n430) );
  XNOR2_X1 U481 ( .A(n430), .B(KEYINPUT55), .ZN(n564) );
  XOR2_X1 U482 ( .A(KEYINPUT20), .B(KEYINPUT86), .Z(n432) );
  XNOR2_X1 U483 ( .A(KEYINPUT85), .B(G71GAT), .ZN(n431) );
  XNOR2_X1 U484 ( .A(n432), .B(n431), .ZN(n448) );
  XOR2_X1 U485 ( .A(G120GAT), .B(G190GAT), .Z(n434) );
  XNOR2_X1 U486 ( .A(G43GAT), .B(G15GAT), .ZN(n433) );
  XNOR2_X1 U487 ( .A(n434), .B(n433), .ZN(n436) );
  XOR2_X1 U488 ( .A(G134GAT), .B(G99GAT), .Z(n435) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n444) );
  XNOR2_X1 U490 ( .A(G183GAT), .B(G127GAT), .ZN(n437) );
  XNOR2_X1 U491 ( .A(n437), .B(G176GAT), .ZN(n438) );
  XOR2_X1 U492 ( .A(n438), .B(KEYINPUT87), .Z(n442) );
  XNOR2_X1 U493 ( .A(n440), .B(n439), .ZN(n441) );
  XNOR2_X1 U494 ( .A(n442), .B(n441), .ZN(n443) );
  XNOR2_X1 U495 ( .A(n444), .B(n443), .ZN(n446) );
  NAND2_X1 U496 ( .A1(G227GAT), .A2(G233GAT), .ZN(n445) );
  XNOR2_X1 U497 ( .A(n446), .B(n445), .ZN(n447) );
  XOR2_X1 U498 ( .A(n448), .B(n447), .Z(n538) );
  NOR2_X1 U499 ( .A1(n543), .A2(n538), .ZN(n449) );
  NAND2_X1 U500 ( .A1(n564), .A2(n449), .ZN(n453) );
  INV_X1 U501 ( .A(G183GAT), .ZN(n451) );
  INV_X1 U502 ( .A(KEYINPUT120), .ZN(n450) );
  XNOR2_X1 U503 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U504 ( .A(n453), .B(n452), .ZN(G1350GAT) );
  INV_X1 U505 ( .A(n538), .ZN(n563) );
  AND2_X1 U506 ( .A1(n563), .A2(n554), .ZN(n454) );
  NAND2_X1 U507 ( .A1(n564), .A2(n454), .ZN(n458) );
  XOR2_X1 U508 ( .A(KEYINPUT57), .B(KEYINPUT119), .Z(n456) );
  XOR2_X1 U509 ( .A(G176GAT), .B(KEYINPUT56), .Z(n455) );
  XNOR2_X1 U510 ( .A(n456), .B(n455), .ZN(n457) );
  XNOR2_X1 U511 ( .A(n458), .B(n457), .ZN(G1349GAT) );
  AND2_X1 U512 ( .A1(n561), .A2(n563), .ZN(n459) );
  NAND2_X1 U513 ( .A1(n564), .A2(n459), .ZN(n463) );
  XOR2_X1 U514 ( .A(KEYINPUT122), .B(KEYINPUT58), .Z(n461) );
  XNOR2_X1 U515 ( .A(G190GAT), .B(KEYINPUT121), .ZN(n460) );
  NAND2_X1 U516 ( .A1(n576), .A2(n567), .ZN(n464) );
  XNOR2_X1 U517 ( .A(n464), .B(KEYINPUT74), .ZN(n498) );
  NOR2_X1 U518 ( .A1(n495), .A2(n561), .ZN(n465) );
  XNOR2_X1 U519 ( .A(n465), .B(KEYINPUT16), .ZN(n484) );
  NAND2_X1 U520 ( .A1(n563), .A2(n526), .ZN(n466) );
  NAND2_X1 U521 ( .A1(n466), .A2(n478), .ZN(n467) );
  XNOR2_X1 U522 ( .A(n467), .B(KEYINPUT99), .ZN(n468) );
  XNOR2_X1 U523 ( .A(n468), .B(KEYINPUT25), .ZN(n472) );
  XNOR2_X1 U524 ( .A(n526), .B(KEYINPUT96), .ZN(n469) );
  XNOR2_X1 U525 ( .A(n469), .B(KEYINPUT27), .ZN(n476) );
  NOR2_X1 U526 ( .A1(n563), .A2(n478), .ZN(n470) );
  XNOR2_X1 U527 ( .A(n470), .B(KEYINPUT26), .ZN(n574) );
  NAND2_X1 U528 ( .A1(n476), .A2(n574), .ZN(n471) );
  NAND2_X1 U529 ( .A1(n472), .A2(n471), .ZN(n473) );
  XOR2_X1 U530 ( .A(KEYINPUT100), .B(n473), .Z(n474) );
  NOR2_X1 U531 ( .A1(n475), .A2(n474), .ZN(n482) );
  NAND2_X1 U532 ( .A1(n523), .A2(n476), .ZN(n477) );
  XNOR2_X1 U533 ( .A(n477), .B(KEYINPUT97), .ZN(n534) );
  XNOR2_X1 U534 ( .A(n478), .B(KEYINPUT28), .ZN(n536) );
  NAND2_X1 U535 ( .A1(n534), .A2(n536), .ZN(n479) );
  NOR2_X1 U536 ( .A1(n563), .A2(n479), .ZN(n480) );
  XNOR2_X1 U537 ( .A(n480), .B(KEYINPUT98), .ZN(n481) );
  NOR2_X1 U538 ( .A1(n482), .A2(n481), .ZN(n494) );
  INV_X1 U539 ( .A(n494), .ZN(n483) );
  NAND2_X1 U540 ( .A1(n484), .A2(n483), .ZN(n512) );
  NOR2_X1 U541 ( .A1(n498), .A2(n512), .ZN(n492) );
  NAND2_X1 U542 ( .A1(n523), .A2(n492), .ZN(n487) );
  XOR2_X1 U543 ( .A(G1GAT), .B(KEYINPUT34), .Z(n485) );
  XNOR2_X1 U544 ( .A(KEYINPUT101), .B(n485), .ZN(n486) );
  XNOR2_X1 U545 ( .A(n487), .B(n486), .ZN(G1324GAT) );
  NAND2_X1 U546 ( .A1(n492), .A2(n526), .ZN(n488) );
  XNOR2_X1 U547 ( .A(n488), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT102), .B(KEYINPUT35), .Z(n490) );
  NAND2_X1 U549 ( .A1(n492), .A2(n563), .ZN(n489) );
  XNOR2_X1 U550 ( .A(n490), .B(n489), .ZN(n491) );
  XNOR2_X1 U551 ( .A(G15GAT), .B(n491), .ZN(G1326GAT) );
  INV_X1 U552 ( .A(n536), .ZN(n529) );
  NAND2_X1 U553 ( .A1(n492), .A2(n529), .ZN(n493) );
  XNOR2_X1 U554 ( .A(n493), .B(G22GAT), .ZN(G1327GAT) );
  XOR2_X1 U555 ( .A(G29GAT), .B(KEYINPUT39), .Z(n502) );
  NOR2_X1 U556 ( .A1(n494), .A2(n586), .ZN(n496) );
  NAND2_X1 U557 ( .A1(n496), .A2(n495), .ZN(n497) );
  XOR2_X1 U558 ( .A(KEYINPUT37), .B(n497), .Z(n522) );
  NOR2_X1 U559 ( .A1(n498), .A2(n522), .ZN(n500) );
  XNOR2_X1 U560 ( .A(KEYINPUT104), .B(KEYINPUT38), .ZN(n499) );
  XNOR2_X1 U561 ( .A(n500), .B(n499), .ZN(n507) );
  NAND2_X1 U562 ( .A1(n507), .A2(n523), .ZN(n501) );
  XNOR2_X1 U563 ( .A(n502), .B(n501), .ZN(G1328GAT) );
  XOR2_X1 U564 ( .A(G36GAT), .B(KEYINPUT105), .Z(n504) );
  NAND2_X1 U565 ( .A1(n507), .A2(n526), .ZN(n503) );
  XNOR2_X1 U566 ( .A(n504), .B(n503), .ZN(G1329GAT) );
  NAND2_X1 U567 ( .A1(n563), .A2(n507), .ZN(n505) );
  XNOR2_X1 U568 ( .A(n505), .B(KEYINPUT40), .ZN(n506) );
  XNOR2_X1 U569 ( .A(G43GAT), .B(n506), .ZN(G1330GAT) );
  XNOR2_X1 U570 ( .A(G50GAT), .B(KEYINPUT106), .ZN(n509) );
  NAND2_X1 U571 ( .A1(n529), .A2(n507), .ZN(n508) );
  XNOR2_X1 U572 ( .A(n509), .B(n508), .ZN(G1331GAT) );
  XNOR2_X1 U573 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n514) );
  INV_X1 U574 ( .A(n567), .ZN(n510) );
  NAND2_X1 U575 ( .A1(n554), .A2(n510), .ZN(n511) );
  XOR2_X1 U576 ( .A(KEYINPUT107), .B(n511), .Z(n521) );
  NOR2_X1 U577 ( .A1(n521), .A2(n512), .ZN(n517) );
  NAND2_X1 U578 ( .A1(n517), .A2(n523), .ZN(n513) );
  XNOR2_X1 U579 ( .A(n514), .B(n513), .ZN(G1332GAT) );
  NAND2_X1 U580 ( .A1(n517), .A2(n526), .ZN(n515) );
  XNOR2_X1 U581 ( .A(n515), .B(G64GAT), .ZN(G1333GAT) );
  NAND2_X1 U582 ( .A1(n563), .A2(n517), .ZN(n516) );
  XNOR2_X1 U583 ( .A(n516), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U584 ( .A(KEYINPUT108), .B(KEYINPUT43), .Z(n519) );
  NAND2_X1 U585 ( .A1(n517), .A2(n529), .ZN(n518) );
  XNOR2_X1 U586 ( .A(n519), .B(n518), .ZN(n520) );
  XNOR2_X1 U587 ( .A(G78GAT), .B(n520), .ZN(G1335GAT) );
  XOR2_X1 U588 ( .A(G85GAT), .B(KEYINPUT109), .Z(n525) );
  NOR2_X1 U589 ( .A1(n522), .A2(n521), .ZN(n530) );
  NAND2_X1 U590 ( .A1(n530), .A2(n523), .ZN(n524) );
  XNOR2_X1 U591 ( .A(n525), .B(n524), .ZN(G1336GAT) );
  NAND2_X1 U592 ( .A1(n530), .A2(n526), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n527), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U594 ( .A1(n563), .A2(n530), .ZN(n528) );
  XNOR2_X1 U595 ( .A(n528), .B(G99GAT), .ZN(G1338GAT) );
  XOR2_X1 U596 ( .A(KEYINPUT44), .B(KEYINPUT110), .Z(n532) );
  NAND2_X1 U597 ( .A1(n530), .A2(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(n533) );
  XOR2_X1 U599 ( .A(G106GAT), .B(n533), .Z(G1339GAT) );
  AND2_X1 U600 ( .A1(n535), .A2(n534), .ZN(n550) );
  NAND2_X1 U601 ( .A1(n550), .A2(n536), .ZN(n537) );
  NOR2_X1 U602 ( .A1(n538), .A2(n537), .ZN(n546) );
  NAND2_X1 U603 ( .A1(n546), .A2(n567), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n539), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U605 ( .A(G120GAT), .B(KEYINPUT49), .Z(n541) );
  NAND2_X1 U606 ( .A1(n546), .A2(n554), .ZN(n540) );
  XNOR2_X1 U607 ( .A(n541), .B(n540), .ZN(G1341GAT) );
  INV_X1 U608 ( .A(n546), .ZN(n542) );
  NOR2_X1 U609 ( .A1(n543), .A2(n542), .ZN(n544) );
  XOR2_X1 U610 ( .A(KEYINPUT50), .B(n544), .Z(n545) );
  XNOR2_X1 U611 ( .A(G127GAT), .B(n545), .ZN(G1342GAT) );
  XOR2_X1 U612 ( .A(KEYINPUT51), .B(KEYINPUT114), .Z(n548) );
  NAND2_X1 U613 ( .A1(n546), .A2(n561), .ZN(n547) );
  XNOR2_X1 U614 ( .A(n548), .B(n547), .ZN(n549) );
  XNOR2_X1 U615 ( .A(G134GAT), .B(n549), .ZN(G1343GAT) );
  NAND2_X1 U616 ( .A1(n550), .A2(n574), .ZN(n551) );
  XNOR2_X1 U617 ( .A(KEYINPUT115), .B(n551), .ZN(n560) );
  NAND2_X1 U618 ( .A1(n560), .A2(n567), .ZN(n552) );
  XNOR2_X1 U619 ( .A(n552), .B(KEYINPUT116), .ZN(n553) );
  XNOR2_X1 U620 ( .A(G141GAT), .B(n553), .ZN(G1344GAT) );
  XOR2_X1 U621 ( .A(KEYINPUT52), .B(KEYINPUT117), .Z(n556) );
  NAND2_X1 U622 ( .A1(n560), .A2(n554), .ZN(n555) );
  XNOR2_X1 U623 ( .A(n556), .B(n555), .ZN(n558) );
  XOR2_X1 U624 ( .A(G148GAT), .B(KEYINPUT53), .Z(n557) );
  XNOR2_X1 U625 ( .A(n558), .B(n557), .ZN(G1345GAT) );
  NAND2_X1 U626 ( .A1(n581), .A2(n560), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n559), .B(G155GAT), .ZN(G1346GAT) );
  NAND2_X1 U628 ( .A1(n561), .A2(n560), .ZN(n562) );
  XNOR2_X1 U629 ( .A(n562), .B(G162GAT), .ZN(G1347GAT) );
  AND2_X1 U630 ( .A1(n564), .A2(n563), .ZN(n565) );
  NAND2_X1 U631 ( .A1(n565), .A2(n567), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n566), .B(G169GAT), .ZN(G1348GAT) );
  AND2_X1 U633 ( .A1(n575), .A2(n574), .ZN(n580) );
  NAND2_X1 U634 ( .A1(n580), .A2(n567), .ZN(n569) );
  XOR2_X1 U635 ( .A(KEYINPUT60), .B(KEYINPUT124), .Z(n568) );
  XNOR2_X1 U636 ( .A(n569), .B(n568), .ZN(n571) );
  INV_X1 U637 ( .A(KEYINPUT59), .ZN(n570) );
  XNOR2_X1 U638 ( .A(n571), .B(n570), .ZN(n573) );
  XNOR2_X1 U639 ( .A(G197GAT), .B(KEYINPUT123), .ZN(n572) );
  XNOR2_X1 U640 ( .A(n573), .B(n572), .ZN(G1352GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT125), .B(KEYINPUT61), .Z(n578) );
  NAND2_X1 U642 ( .A1(n575), .A2(n574), .ZN(n585) );
  OR2_X1 U643 ( .A1(n585), .A2(n576), .ZN(n577) );
  XNOR2_X1 U644 ( .A(n578), .B(n577), .ZN(n579) );
  XOR2_X1 U645 ( .A(G204GAT), .B(n579), .Z(G1353GAT) );
  NAND2_X1 U646 ( .A1(n581), .A2(n580), .ZN(n582) );
  XNOR2_X1 U647 ( .A(n582), .B(G211GAT), .ZN(G1354GAT) );
  XOR2_X1 U648 ( .A(KEYINPUT126), .B(KEYINPUT127), .Z(n584) );
  XNOR2_X1 U649 ( .A(G218GAT), .B(KEYINPUT62), .ZN(n583) );
  XNOR2_X1 U650 ( .A(n584), .B(n583), .ZN(n588) );
  NOR2_X1 U651 ( .A1(n586), .A2(n585), .ZN(n587) );
  XOR2_X1 U652 ( .A(n588), .B(n587), .Z(G1355GAT) );
endmodule

