

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
         n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578,
         n579, n580, n581, n582, n583, n584, n585, n586;

  INV_X1 U325 ( .A(n549), .ZN(n575) );
  XNOR2_X2 U326 ( .A(n405), .B(n404), .ZN(n549) );
  XOR2_X2 U327 ( .A(n442), .B(n441), .Z(n556) );
  NOR2_X1 U328 ( .A1(n515), .A2(n462), .ZN(n568) );
  NAND2_X1 U329 ( .A1(n385), .A2(n384), .ZN(n477) );
  INV_X1 U330 ( .A(KEYINPUT37), .ZN(n407) );
  XOR2_X1 U331 ( .A(n372), .B(n360), .Z(n517) );
  XOR2_X1 U332 ( .A(G204GAT), .B(G211GAT), .Z(n293) );
  XNOR2_X1 U333 ( .A(KEYINPUT89), .B(KEYINPUT25), .ZN(n374) );
  XNOR2_X1 U334 ( .A(n375), .B(n374), .ZN(n378) );
  XNOR2_X1 U335 ( .A(n338), .B(n421), .ZN(n339) );
  XNOR2_X1 U336 ( .A(KEYINPUT64), .B(KEYINPUT48), .ZN(n458) );
  XNOR2_X1 U337 ( .A(n340), .B(n339), .ZN(n341) );
  XNOR2_X1 U338 ( .A(n416), .B(n415), .ZN(n420) );
  XNOR2_X1 U339 ( .A(n459), .B(n458), .ZN(n524) );
  XNOR2_X1 U340 ( .A(n420), .B(n419), .ZN(n424) );
  XOR2_X1 U341 ( .A(n344), .B(n343), .Z(n463) );
  XOR2_X1 U342 ( .A(n372), .B(n371), .Z(n526) );
  XNOR2_X1 U343 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U344 ( .A(n445), .B(G29GAT), .ZN(n446) );
  XNOR2_X1 U345 ( .A(n474), .B(n473), .ZN(G1349GAT) );
  XNOR2_X1 U346 ( .A(n447), .B(n446), .ZN(G1328GAT) );
  XOR2_X1 U347 ( .A(KEYINPUT0), .B(G127GAT), .Z(n362) );
  XOR2_X1 U348 ( .A(n362), .B(G57GAT), .Z(n295) );
  NAND2_X1 U349 ( .A1(G225GAT), .A2(G233GAT), .ZN(n294) );
  XNOR2_X1 U350 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U351 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n297) );
  XNOR2_X1 U352 ( .A(G1GAT), .B(KEYINPUT5), .ZN(n296) );
  XNOR2_X1 U353 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U354 ( .A(n299), .B(n298), .Z(n301) );
  XNOR2_X1 U355 ( .A(G29GAT), .B(G134GAT), .ZN(n300) );
  XNOR2_X1 U356 ( .A(n301), .B(n300), .ZN(n305) );
  XOR2_X1 U357 ( .A(G85GAT), .B(G155GAT), .Z(n303) );
  XNOR2_X1 U358 ( .A(G162GAT), .B(G148GAT), .ZN(n302) );
  XNOR2_X1 U359 ( .A(n303), .B(n302), .ZN(n304) );
  XOR2_X1 U360 ( .A(n305), .B(n304), .Z(n314) );
  XOR2_X1 U361 ( .A(KEYINPUT82), .B(KEYINPUT2), .Z(n307) );
  XNOR2_X1 U362 ( .A(KEYINPUT3), .B(KEYINPUT83), .ZN(n306) );
  XNOR2_X1 U363 ( .A(n307), .B(n306), .ZN(n308) );
  XOR2_X1 U364 ( .A(G141GAT), .B(n308), .Z(n344) );
  INV_X1 U365 ( .A(n344), .ZN(n312) );
  XOR2_X1 U366 ( .A(KEYINPUT4), .B(KEYINPUT86), .Z(n310) );
  XNOR2_X1 U367 ( .A(G113GAT), .B(G120GAT), .ZN(n309) );
  XNOR2_X1 U368 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U369 ( .A(n312), .B(n311), .Z(n313) );
  XNOR2_X1 U370 ( .A(n314), .B(n313), .ZN(n515) );
  XNOR2_X1 U371 ( .A(KEYINPUT97), .B(KEYINPUT38), .ZN(n444) );
  XOR2_X1 U372 ( .A(G50GAT), .B(G162GAT), .Z(n332) );
  XOR2_X1 U373 ( .A(G36GAT), .B(G218GAT), .Z(n357) );
  XNOR2_X1 U374 ( .A(n332), .B(n357), .ZN(n328) );
  XNOR2_X1 U375 ( .A(G43GAT), .B(G190GAT), .ZN(n315) );
  XNOR2_X1 U376 ( .A(n315), .B(G134GAT), .ZN(n361) );
  XOR2_X1 U377 ( .A(KEYINPUT10), .B(n361), .Z(n317) );
  NAND2_X1 U378 ( .A1(G232GAT), .A2(G233GAT), .ZN(n316) );
  XNOR2_X1 U379 ( .A(n317), .B(n316), .ZN(n321) );
  XOR2_X1 U380 ( .A(KEYINPUT72), .B(KEYINPUT9), .Z(n319) );
  XNOR2_X1 U381 ( .A(KEYINPUT65), .B(KEYINPUT11), .ZN(n318) );
  XNOR2_X1 U382 ( .A(n319), .B(n318), .ZN(n320) );
  XNOR2_X1 U383 ( .A(n321), .B(n320), .ZN(n326) );
  XNOR2_X1 U384 ( .A(G29GAT), .B(KEYINPUT8), .ZN(n322) );
  XNOR2_X1 U385 ( .A(n322), .B(KEYINPUT7), .ZN(n432) );
  XOR2_X1 U386 ( .A(G92GAT), .B(G85GAT), .Z(n324) );
  XNOR2_X1 U387 ( .A(G99GAT), .B(G106GAT), .ZN(n323) );
  XNOR2_X1 U388 ( .A(n324), .B(n323), .ZN(n418) );
  XOR2_X1 U389 ( .A(n432), .B(n418), .Z(n325) );
  XNOR2_X1 U390 ( .A(n326), .B(n325), .ZN(n327) );
  XNOR2_X1 U391 ( .A(n328), .B(n327), .ZN(n553) );
  XOR2_X1 U392 ( .A(KEYINPUT73), .B(n553), .Z(n536) );
  XNOR2_X1 U393 ( .A(KEYINPUT36), .B(n536), .ZN(n581) );
  XOR2_X1 U394 ( .A(KEYINPUT23), .B(KEYINPUT24), .Z(n330) );
  XNOR2_X1 U395 ( .A(KEYINPUT84), .B(KEYINPUT22), .ZN(n329) );
  XNOR2_X1 U396 ( .A(n330), .B(n329), .ZN(n342) );
  XNOR2_X1 U397 ( .A(G197GAT), .B(KEYINPUT21), .ZN(n331) );
  XNOR2_X1 U398 ( .A(n293), .B(n331), .ZN(n350) );
  XOR2_X1 U399 ( .A(n332), .B(n350), .Z(n334) );
  NAND2_X1 U400 ( .A1(G228GAT), .A2(G233GAT), .ZN(n333) );
  XNOR2_X1 U401 ( .A(n334), .B(n333), .ZN(n340) );
  XOR2_X1 U402 ( .A(KEYINPUT81), .B(KEYINPUT85), .Z(n336) );
  XNOR2_X1 U403 ( .A(G218GAT), .B(G106GAT), .ZN(n335) );
  XNOR2_X1 U404 ( .A(n336), .B(n335), .ZN(n337) );
  XOR2_X1 U405 ( .A(G22GAT), .B(G155GAT), .Z(n390) );
  XOR2_X1 U406 ( .A(n337), .B(n390), .Z(n338) );
  XOR2_X1 U407 ( .A(G148GAT), .B(G78GAT), .Z(n421) );
  XOR2_X1 U408 ( .A(n342), .B(n341), .Z(n343) );
  XOR2_X1 U409 ( .A(KEYINPUT17), .B(KEYINPUT78), .Z(n346) );
  XNOR2_X1 U410 ( .A(KEYINPUT18), .B(KEYINPUT19), .ZN(n345) );
  XNOR2_X1 U411 ( .A(n346), .B(n345), .ZN(n347) );
  XOR2_X1 U412 ( .A(n347), .B(G183GAT), .Z(n349) );
  XNOR2_X1 U413 ( .A(G169GAT), .B(G176GAT), .ZN(n348) );
  XNOR2_X1 U414 ( .A(n349), .B(n348), .ZN(n372) );
  XOR2_X1 U415 ( .A(KEYINPUT87), .B(n350), .Z(n352) );
  NAND2_X1 U416 ( .A1(G226GAT), .A2(G233GAT), .ZN(n351) );
  XNOR2_X1 U417 ( .A(n352), .B(n351), .ZN(n356) );
  XOR2_X1 U418 ( .A(KEYINPUT88), .B(G64GAT), .Z(n354) );
  XNOR2_X1 U419 ( .A(G190GAT), .B(G92GAT), .ZN(n353) );
  XNOR2_X1 U420 ( .A(n354), .B(n353), .ZN(n355) );
  XOR2_X1 U421 ( .A(n356), .B(n355), .Z(n359) );
  XOR2_X1 U422 ( .A(G8GAT), .B(KEYINPUT74), .Z(n391) );
  XNOR2_X1 U423 ( .A(n357), .B(n391), .ZN(n358) );
  XNOR2_X1 U424 ( .A(n359), .B(n358), .ZN(n360) );
  XOR2_X1 U425 ( .A(n362), .B(n361), .Z(n364) );
  NAND2_X1 U426 ( .A1(G227GAT), .A2(G233GAT), .ZN(n363) );
  XNOR2_X1 U427 ( .A(n364), .B(n363), .ZN(n368) );
  XOR2_X1 U428 ( .A(KEYINPUT79), .B(KEYINPUT77), .Z(n366) );
  XNOR2_X1 U429 ( .A(G99GAT), .B(KEYINPUT20), .ZN(n365) );
  XNOR2_X1 U430 ( .A(n366), .B(n365), .ZN(n367) );
  XOR2_X1 U431 ( .A(n368), .B(n367), .Z(n370) );
  XOR2_X1 U432 ( .A(G113GAT), .B(G15GAT), .Z(n428) );
  XOR2_X1 U433 ( .A(G120GAT), .B(G71GAT), .Z(n422) );
  XNOR2_X1 U434 ( .A(n428), .B(n422), .ZN(n369) );
  XNOR2_X1 U435 ( .A(n370), .B(n369), .ZN(n371) );
  NAND2_X1 U436 ( .A1(n517), .A2(n526), .ZN(n373) );
  NAND2_X1 U437 ( .A1(n463), .A2(n373), .ZN(n375) );
  NOR2_X1 U438 ( .A1(n463), .A2(n526), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n376), .B(KEYINPUT26), .ZN(n567) );
  XNOR2_X1 U440 ( .A(KEYINPUT27), .B(n517), .ZN(n382) );
  NAND2_X1 U441 ( .A1(n567), .A2(n382), .ZN(n377) );
  NAND2_X1 U442 ( .A1(n378), .A2(n377), .ZN(n379) );
  XOR2_X1 U443 ( .A(KEYINPUT90), .B(n379), .Z(n380) );
  NOR2_X1 U444 ( .A1(n515), .A2(n380), .ZN(n381) );
  XNOR2_X1 U445 ( .A(n381), .B(KEYINPUT91), .ZN(n385) );
  XOR2_X1 U446 ( .A(n526), .B(KEYINPUT80), .Z(n383) );
  XOR2_X1 U447 ( .A(n463), .B(KEYINPUT28), .Z(n520) );
  NAND2_X1 U448 ( .A1(n515), .A2(n382), .ZN(n541) );
  NOR2_X1 U449 ( .A1(n520), .A2(n541), .ZN(n525) );
  NAND2_X1 U450 ( .A1(n383), .A2(n525), .ZN(n384) );
  XOR2_X1 U451 ( .A(G127GAT), .B(G71GAT), .Z(n387) );
  XNOR2_X1 U452 ( .A(G15GAT), .B(G183GAT), .ZN(n386) );
  XNOR2_X1 U453 ( .A(n387), .B(n386), .ZN(n405) );
  XOR2_X1 U454 ( .A(KEYINPUT15), .B(KEYINPUT76), .Z(n389) );
  XNOR2_X1 U455 ( .A(G1GAT), .B(KEYINPUT12), .ZN(n388) );
  XNOR2_X1 U456 ( .A(n389), .B(n388), .ZN(n395) );
  XOR2_X1 U457 ( .A(n391), .B(n390), .Z(n393) );
  XNOR2_X1 U458 ( .A(G211GAT), .B(G78GAT), .ZN(n392) );
  XNOR2_X1 U459 ( .A(n393), .B(n392), .ZN(n394) );
  XOR2_X1 U460 ( .A(n395), .B(n394), .Z(n397) );
  NAND2_X1 U461 ( .A1(G231GAT), .A2(G233GAT), .ZN(n396) );
  XNOR2_X1 U462 ( .A(n397), .B(n396), .ZN(n399) );
  INV_X1 U463 ( .A(KEYINPUT14), .ZN(n398) );
  XNOR2_X1 U464 ( .A(n399), .B(n398), .ZN(n403) );
  XOR2_X1 U465 ( .A(G64GAT), .B(KEYINPUT69), .Z(n401) );
  XNOR2_X1 U466 ( .A(G57GAT), .B(KEYINPUT13), .ZN(n400) );
  XNOR2_X1 U467 ( .A(n401), .B(n400), .ZN(n417) );
  XNOR2_X1 U468 ( .A(n417), .B(KEYINPUT75), .ZN(n402) );
  XNOR2_X1 U469 ( .A(n403), .B(n402), .ZN(n404) );
  NAND2_X1 U470 ( .A1(n477), .A2(n549), .ZN(n406) );
  NOR2_X1 U471 ( .A1(n581), .A2(n406), .ZN(n408) );
  XNOR2_X1 U472 ( .A(n408), .B(n407), .ZN(n514) );
  XOR2_X1 U473 ( .A(KEYINPUT31), .B(KEYINPUT70), .Z(n410) );
  NAND2_X1 U474 ( .A1(G230GAT), .A2(G233GAT), .ZN(n409) );
  XNOR2_X1 U475 ( .A(n410), .B(n409), .ZN(n412) );
  INV_X1 U476 ( .A(KEYINPUT32), .ZN(n411) );
  XNOR2_X1 U477 ( .A(n412), .B(n411), .ZN(n416) );
  XOR2_X1 U478 ( .A(KEYINPUT71), .B(KEYINPUT33), .Z(n414) );
  XNOR2_X1 U479 ( .A(G176GAT), .B(G204GAT), .ZN(n413) );
  XNOR2_X1 U480 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U481 ( .A(n418), .B(n417), .ZN(n419) );
  XOR2_X1 U482 ( .A(n422), .B(n421), .Z(n423) );
  XNOR2_X1 U483 ( .A(n424), .B(n423), .ZN(n572) );
  XOR2_X1 U484 ( .A(G197GAT), .B(G50GAT), .Z(n426) );
  XNOR2_X1 U485 ( .A(G43GAT), .B(G36GAT), .ZN(n425) );
  XNOR2_X1 U486 ( .A(n426), .B(n425), .ZN(n427) );
  XOR2_X1 U487 ( .A(n428), .B(n427), .Z(n430) );
  NAND2_X1 U488 ( .A1(G229GAT), .A2(G233GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n431) );
  XOR2_X1 U490 ( .A(n431), .B(KEYINPUT67), .Z(n434) );
  XNOR2_X1 U491 ( .A(n432), .B(KEYINPUT66), .ZN(n433) );
  XNOR2_X1 U492 ( .A(n434), .B(n433), .ZN(n442) );
  XOR2_X1 U493 ( .A(G1GAT), .B(G141GAT), .Z(n436) );
  XNOR2_X1 U494 ( .A(G169GAT), .B(G22GAT), .ZN(n435) );
  XNOR2_X1 U495 ( .A(n436), .B(n435), .ZN(n440) );
  XOR2_X1 U496 ( .A(KEYINPUT30), .B(KEYINPUT29), .Z(n438) );
  XNOR2_X1 U497 ( .A(G8GAT), .B(KEYINPUT68), .ZN(n437) );
  XNOR2_X1 U498 ( .A(n438), .B(n437), .ZN(n439) );
  XOR2_X1 U499 ( .A(n440), .B(n439), .Z(n441) );
  INV_X1 U500 ( .A(n556), .ZN(n569) );
  NOR2_X1 U501 ( .A1(n572), .A2(n569), .ZN(n478) );
  NAND2_X1 U502 ( .A1(n514), .A2(n478), .ZN(n443) );
  XNOR2_X1 U503 ( .A(n444), .B(n443), .ZN(n494) );
  NAND2_X1 U504 ( .A1(n515), .A2(n494), .ZN(n447) );
  XOR2_X1 U505 ( .A(KEYINPUT96), .B(KEYINPUT39), .Z(n445) );
  XOR2_X1 U506 ( .A(n572), .B(KEYINPUT41), .Z(n530) );
  INV_X1 U507 ( .A(KEYINPUT116), .ZN(n468) );
  AND2_X1 U508 ( .A1(n556), .A2(n530), .ZN(n448) );
  XNOR2_X1 U509 ( .A(n448), .B(KEYINPUT46), .ZN(n449) );
  NOR2_X1 U510 ( .A1(n575), .A2(n449), .ZN(n450) );
  XNOR2_X1 U511 ( .A(n450), .B(KEYINPUT108), .ZN(n451) );
  NAND2_X1 U512 ( .A1(n451), .A2(n553), .ZN(n452) );
  XNOR2_X1 U513 ( .A(n452), .B(KEYINPUT47), .ZN(n457) );
  NOR2_X1 U514 ( .A1(n581), .A2(n549), .ZN(n453) );
  XNOR2_X1 U515 ( .A(n453), .B(KEYINPUT45), .ZN(n454) );
  NAND2_X1 U516 ( .A1(n454), .A2(n569), .ZN(n455) );
  NOR2_X1 U517 ( .A1(n455), .A2(n572), .ZN(n456) );
  NOR2_X1 U518 ( .A1(n457), .A2(n456), .ZN(n459) );
  INV_X1 U519 ( .A(n517), .ZN(n460) );
  NOR2_X1 U520 ( .A1(n524), .A2(n460), .ZN(n461) );
  XOR2_X1 U521 ( .A(KEYINPUT54), .B(n461), .Z(n462) );
  NAND2_X1 U522 ( .A1(n568), .A2(n463), .ZN(n465) );
  XOR2_X1 U523 ( .A(KEYINPUT55), .B(KEYINPUT115), .Z(n464) );
  XNOR2_X1 U524 ( .A(n465), .B(n464), .ZN(n466) );
  NAND2_X1 U525 ( .A1(n466), .A2(n526), .ZN(n467) );
  XNOR2_X2 U526 ( .A(n468), .B(n467), .ZN(n561) );
  NAND2_X1 U527 ( .A1(n530), .A2(n561), .ZN(n474) );
  XOR2_X1 U528 ( .A(KEYINPUT120), .B(KEYINPUT119), .Z(n470) );
  XNOR2_X1 U529 ( .A(KEYINPUT118), .B(KEYINPUT57), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(n472) );
  XOR2_X1 U531 ( .A(G176GAT), .B(KEYINPUT56), .Z(n471) );
  XNOR2_X1 U532 ( .A(KEYINPUT93), .B(KEYINPUT34), .ZN(n483) );
  XOR2_X1 U533 ( .A(G1GAT), .B(KEYINPUT94), .Z(n481) );
  NAND2_X1 U534 ( .A1(n536), .A2(n575), .ZN(n475) );
  XOR2_X1 U535 ( .A(KEYINPUT16), .B(n475), .Z(n476) );
  AND2_X1 U536 ( .A1(n477), .A2(n476), .ZN(n498) );
  NAND2_X1 U537 ( .A1(n478), .A2(n498), .ZN(n479) );
  XOR2_X1 U538 ( .A(KEYINPUT92), .B(n479), .Z(n487) );
  NAND2_X1 U539 ( .A1(n515), .A2(n487), .ZN(n480) );
  XNOR2_X1 U540 ( .A(n481), .B(n480), .ZN(n482) );
  XNOR2_X1 U541 ( .A(n483), .B(n482), .ZN(G1324GAT) );
  NAND2_X1 U542 ( .A1(n487), .A2(n517), .ZN(n484) );
  XNOR2_X1 U543 ( .A(n484), .B(G8GAT), .ZN(G1325GAT) );
  XOR2_X1 U544 ( .A(G15GAT), .B(KEYINPUT35), .Z(n486) );
  NAND2_X1 U545 ( .A1(n526), .A2(n487), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n486), .B(n485), .ZN(G1326GAT) );
  XOR2_X1 U547 ( .A(G22GAT), .B(KEYINPUT95), .Z(n489) );
  NAND2_X1 U548 ( .A1(n520), .A2(n487), .ZN(n488) );
  XNOR2_X1 U549 ( .A(n489), .B(n488), .ZN(G1327GAT) );
  NAND2_X1 U550 ( .A1(n494), .A2(n517), .ZN(n490) );
  XNOR2_X1 U551 ( .A(n490), .B(KEYINPUT98), .ZN(n491) );
  XNOR2_X1 U552 ( .A(G36GAT), .B(n491), .ZN(G1329GAT) );
  NAND2_X1 U553 ( .A1(n494), .A2(n526), .ZN(n492) );
  XNOR2_X1 U554 ( .A(n492), .B(KEYINPUT40), .ZN(n493) );
  XNOR2_X1 U555 ( .A(G43GAT), .B(n493), .ZN(G1330GAT) );
  XOR2_X1 U556 ( .A(G50GAT), .B(KEYINPUT99), .Z(n496) );
  NAND2_X1 U557 ( .A1(n520), .A2(n494), .ZN(n495) );
  XNOR2_X1 U558 ( .A(n496), .B(n495), .ZN(G1331GAT) );
  INV_X1 U559 ( .A(n530), .ZN(n546) );
  NOR2_X1 U560 ( .A1(n546), .A2(n556), .ZN(n497) );
  XNOR2_X1 U561 ( .A(n497), .B(KEYINPUT100), .ZN(n513) );
  NAND2_X1 U562 ( .A1(n513), .A2(n498), .ZN(n499) );
  XNOR2_X1 U563 ( .A(n499), .B(KEYINPUT101), .ZN(n509) );
  NAND2_X1 U564 ( .A1(n509), .A2(n515), .ZN(n502) );
  XNOR2_X1 U565 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n500) );
  XNOR2_X1 U566 ( .A(n500), .B(KEYINPUT102), .ZN(n501) );
  XNOR2_X1 U567 ( .A(n502), .B(n501), .ZN(G1332GAT) );
  NAND2_X1 U568 ( .A1(n509), .A2(n517), .ZN(n503) );
  XNOR2_X1 U569 ( .A(n503), .B(G64GAT), .ZN(G1333GAT) );
  XOR2_X1 U570 ( .A(KEYINPUT103), .B(KEYINPUT104), .Z(n505) );
  NAND2_X1 U571 ( .A1(n509), .A2(n526), .ZN(n504) );
  XNOR2_X1 U572 ( .A(n505), .B(n504), .ZN(n506) );
  XNOR2_X1 U573 ( .A(G71GAT), .B(n506), .ZN(G1334GAT) );
  XOR2_X1 U574 ( .A(KEYINPUT107), .B(KEYINPUT106), .Z(n508) );
  XNOR2_X1 U575 ( .A(G78GAT), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U576 ( .A(n508), .B(n507), .ZN(n512) );
  NAND2_X1 U577 ( .A1(n509), .A2(n520), .ZN(n510) );
  XNOR2_X1 U578 ( .A(n510), .B(KEYINPUT105), .ZN(n511) );
  XNOR2_X1 U579 ( .A(n512), .B(n511), .ZN(G1335GAT) );
  AND2_X1 U580 ( .A1(n514), .A2(n513), .ZN(n521) );
  NAND2_X1 U581 ( .A1(n515), .A2(n521), .ZN(n516) );
  XNOR2_X1 U582 ( .A(G85GAT), .B(n516), .ZN(G1336GAT) );
  NAND2_X1 U583 ( .A1(n521), .A2(n517), .ZN(n518) );
  XNOR2_X1 U584 ( .A(n518), .B(G92GAT), .ZN(G1337GAT) );
  NAND2_X1 U585 ( .A1(n521), .A2(n526), .ZN(n519) );
  XNOR2_X1 U586 ( .A(n519), .B(G99GAT), .ZN(G1338GAT) );
  NAND2_X1 U587 ( .A1(n521), .A2(n520), .ZN(n522) );
  XNOR2_X1 U588 ( .A(n522), .B(KEYINPUT44), .ZN(n523) );
  XNOR2_X1 U589 ( .A(G106GAT), .B(n523), .ZN(G1339GAT) );
  XOR2_X1 U590 ( .A(G113GAT), .B(KEYINPUT109), .Z(n529) );
  NAND2_X1 U591 ( .A1(n526), .A2(n525), .ZN(n527) );
  NOR2_X1 U592 ( .A1(n524), .A2(n527), .ZN(n537) );
  NAND2_X1 U593 ( .A1(n537), .A2(n556), .ZN(n528) );
  XNOR2_X1 U594 ( .A(n529), .B(n528), .ZN(G1340GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT110), .B(KEYINPUT49), .Z(n532) );
  NAND2_X1 U596 ( .A1(n537), .A2(n530), .ZN(n531) );
  XNOR2_X1 U597 ( .A(n532), .B(n531), .ZN(n533) );
  XNOR2_X1 U598 ( .A(G120GAT), .B(n533), .ZN(G1341GAT) );
  NAND2_X1 U599 ( .A1(n537), .A2(n575), .ZN(n534) );
  XNOR2_X1 U600 ( .A(n534), .B(KEYINPUT50), .ZN(n535) );
  XNOR2_X1 U601 ( .A(G127GAT), .B(n535), .ZN(G1342GAT) );
  XOR2_X1 U602 ( .A(KEYINPUT51), .B(KEYINPUT111), .Z(n539) );
  INV_X1 U603 ( .A(n536), .ZN(n560) );
  NAND2_X1 U604 ( .A1(n537), .A2(n560), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(n540) );
  XOR2_X1 U606 ( .A(G134GAT), .B(n540), .Z(G1343GAT) );
  NOR2_X1 U607 ( .A1(n524), .A2(n541), .ZN(n542) );
  NAND2_X1 U608 ( .A1(n542), .A2(n567), .ZN(n552) );
  NOR2_X1 U609 ( .A1(n569), .A2(n552), .ZN(n543) );
  XOR2_X1 U610 ( .A(G141GAT), .B(n543), .Z(G1344GAT) );
  XOR2_X1 U611 ( .A(KEYINPUT52), .B(KEYINPUT112), .Z(n545) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n544) );
  XNOR2_X1 U613 ( .A(n545), .B(n544), .ZN(n548) );
  NOR2_X1 U614 ( .A1(n546), .A2(n552), .ZN(n547) );
  XOR2_X1 U615 ( .A(n548), .B(n547), .Z(G1345GAT) );
  NOR2_X1 U616 ( .A1(n549), .A2(n552), .ZN(n551) );
  XNOR2_X1 U617 ( .A(G155GAT), .B(KEYINPUT113), .ZN(n550) );
  XNOR2_X1 U618 ( .A(n551), .B(n550), .ZN(G1346GAT) );
  NOR2_X1 U619 ( .A1(n553), .A2(n552), .ZN(n554) );
  XOR2_X1 U620 ( .A(KEYINPUT114), .B(n554), .Z(n555) );
  XNOR2_X1 U621 ( .A(G162GAT), .B(n555), .ZN(G1347GAT) );
  XOR2_X1 U622 ( .A(G169GAT), .B(KEYINPUT117), .Z(n558) );
  NAND2_X1 U623 ( .A1(n556), .A2(n561), .ZN(n557) );
  XNOR2_X1 U624 ( .A(n558), .B(n557), .ZN(G1348GAT) );
  NAND2_X1 U625 ( .A1(n561), .A2(n575), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n559), .B(G183GAT), .ZN(G1350GAT) );
  NAND2_X1 U627 ( .A1(n561), .A2(n560), .ZN(n563) );
  XOR2_X1 U628 ( .A(KEYINPUT58), .B(KEYINPUT121), .Z(n562) );
  XNOR2_X1 U629 ( .A(n563), .B(n562), .ZN(n564) );
  XNOR2_X1 U630 ( .A(n564), .B(G190GAT), .ZN(G1351GAT) );
  XOR2_X1 U631 ( .A(KEYINPUT122), .B(KEYINPUT59), .Z(n566) );
  XNOR2_X1 U632 ( .A(G197GAT), .B(KEYINPUT60), .ZN(n565) );
  XNOR2_X1 U633 ( .A(n566), .B(n565), .ZN(n571) );
  NAND2_X1 U634 ( .A1(n568), .A2(n567), .ZN(n580) );
  NOR2_X1 U635 ( .A1(n569), .A2(n580), .ZN(n570) );
  XOR2_X1 U636 ( .A(n571), .B(n570), .Z(G1352GAT) );
  XOR2_X1 U637 ( .A(G204GAT), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n580), .ZN(n576) );
  NAND2_X1 U639 ( .A1(n576), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(G1353GAT) );
  XOR2_X1 U641 ( .A(KEYINPUT123), .B(KEYINPUT124), .Z(n578) );
  NAND2_X1 U642 ( .A1(n576), .A2(n575), .ZN(n577) );
  XNOR2_X1 U643 ( .A(n578), .B(n577), .ZN(n579) );
  XNOR2_X1 U644 ( .A(G211GAT), .B(n579), .ZN(G1354GAT) );
  NOR2_X1 U645 ( .A1(n581), .A2(n580), .ZN(n586) );
  XOR2_X1 U646 ( .A(KEYINPUT62), .B(KEYINPUT127), .Z(n583) );
  XNOR2_X1 U647 ( .A(G218GAT), .B(KEYINPUT126), .ZN(n582) );
  XNOR2_X1 U648 ( .A(n583), .B(n582), .ZN(n584) );
  XNOR2_X1 U649 ( .A(KEYINPUT125), .B(n584), .ZN(n585) );
  XNOR2_X1 U650 ( .A(n586), .B(n585), .ZN(G1355GAT) );
endmodule

