

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737;

  XNOR2_X1 U364 ( .A(n341), .B(n525), .ZN(n727) );
  NOR2_X2 U365 ( .A1(n644), .A2(n664), .ZN(n343) );
  OR2_X2 U366 ( .A1(n632), .A2(G902), .ZN(n422) );
  NOR2_X2 U367 ( .A1(n390), .A2(n538), .ZN(n439) );
  XNOR2_X2 U368 ( .A(n387), .B(n403), .ZN(n386) );
  NOR2_X1 U369 ( .A1(n436), .A2(n431), .ZN(n365) );
  NAND2_X1 U370 ( .A1(n344), .A2(n379), .ZN(n644) );
  NOR2_X1 U371 ( .A1(n599), .A2(n673), .ZN(n591) );
  NOR2_X1 U372 ( .A1(n366), .A2(n365), .ZN(n372) );
  XNOR2_X1 U373 ( .A(n511), .B(G137), .ZN(n341) );
  INV_X1 U374 ( .A(G119), .ZN(n443) );
  XNOR2_X1 U375 ( .A(KEYINPUT73), .B(KEYINPUT3), .ZN(n444) );
  OR2_X1 U376 ( .A1(n412), .A2(n411), .ZN(n410) );
  NAND2_X1 U377 ( .A1(n657), .A2(n618), .ZN(n620) );
  AND2_X1 U378 ( .A1(n427), .A2(n579), .ZN(n426) );
  NOR2_X1 U379 ( .A1(n633), .A2(n425), .ZN(n424) );
  XNOR2_X1 U380 ( .A(n346), .B(KEYINPUT71), .ZN(n345) );
  XNOR2_X1 U381 ( .A(n351), .B(n606), .ZN(n350) );
  XNOR2_X1 U382 ( .A(n343), .B(n594), .ZN(n595) );
  INV_X1 U383 ( .A(n653), .ZN(n347) );
  INV_X1 U384 ( .A(n602), .ZN(n344) );
  NOR2_X1 U385 ( .A1(n501), .A2(n585), .ZN(n502) );
  NAND2_X1 U386 ( .A1(n372), .A2(n370), .ZN(n417) );
  XNOR2_X1 U387 ( .A(n592), .B(n543), .ZN(n677) );
  AND2_X1 U388 ( .A1(n433), .A2(n357), .ZN(n371) );
  XNOR2_X1 U389 ( .A(n490), .B(n489), .ZN(n670) );
  OR2_X1 U390 ( .A1(n706), .A2(G902), .ZN(n487) );
  XOR2_X1 U391 ( .A(KEYINPUT59), .B(n621), .Z(n622) );
  XNOR2_X1 U392 ( .A(n447), .B(G953), .ZN(n729) );
  XNOR2_X1 U393 ( .A(n453), .B(G902), .ZN(n618) );
  XNOR2_X1 U394 ( .A(n444), .B(n443), .ZN(n418) );
  INV_X1 U395 ( .A(KEYINPUT75), .ZN(n349) );
  XNOR2_X2 U396 ( .A(n342), .B(G131), .ZN(n511) );
  XNOR2_X2 U397 ( .A(KEYINPUT68), .B(KEYINPUT69), .ZN(n342) );
  NAND2_X1 U398 ( .A1(n350), .A2(n345), .ZN(n609) );
  NAND2_X1 U399 ( .A1(n348), .A2(n347), .ZN(n346) );
  XNOR2_X1 U400 ( .A(n596), .B(n349), .ZN(n348) );
  NAND2_X1 U401 ( .A1(n605), .A2(n604), .ZN(n351) );
  XNOR2_X2 U402 ( .A(n532), .B(KEYINPUT40), .ZN(n605) );
  NOR2_X2 U403 ( .A1(n620), .A2(n656), .ZN(n698) );
  NAND2_X1 U404 ( .A1(n364), .A2(n639), .ZN(n564) );
  XNOR2_X1 U405 ( .A(n381), .B(n380), .ZN(n522) );
  INV_X1 U406 ( .A(KEYINPUT8), .ZN(n380) );
  INV_X1 U407 ( .A(KEYINPUT67), .ZN(n560) );
  OR2_X1 U408 ( .A1(n352), .A2(n618), .ZN(n434) );
  NAND2_X1 U409 ( .A1(n352), .A2(n618), .ZN(n435) );
  NOR2_X1 U410 ( .A1(G953), .A2(G237), .ZN(n503) );
  XOR2_X1 U411 ( .A(KEYINPUT18), .B(KEYINPUT83), .Z(n451) );
  INV_X1 U412 ( .A(n472), .ZN(n403) );
  NOR2_X1 U413 ( .A1(n356), .A2(n430), .ZN(n367) );
  OR2_X1 U414 ( .A1(n588), .A2(n587), .ZN(n440) );
  XNOR2_X1 U415 ( .A(n442), .B(n476), .ZN(n421) );
  XOR2_X1 U416 ( .A(G137), .B(G128), .Z(n442) );
  XOR2_X1 U417 ( .A(KEYINPUT99), .B(KEYINPUT23), .Z(n476) );
  XNOR2_X1 U418 ( .A(n420), .B(n475), .ZN(n419) );
  INV_X1 U419 ( .A(KEYINPUT24), .ZN(n475) );
  XNOR2_X1 U420 ( .A(G119), .B(G110), .ZN(n420) );
  XNOR2_X1 U421 ( .A(KEYINPUT70), .B(G140), .ZN(n478) );
  XNOR2_X1 U422 ( .A(n727), .B(G146), .ZN(n474) );
  BUF_X1 U423 ( .A(n677), .Z(n363) );
  INV_X1 U424 ( .A(KEYINPUT22), .ZN(n541) );
  NAND2_X1 U425 ( .A1(n438), .A2(n670), .ZN(n437) );
  XNOR2_X1 U426 ( .A(n377), .B(n376), .ZN(n382) );
  XNOR2_X1 U427 ( .A(n515), .B(n516), .ZN(n376) );
  OR2_X1 U428 ( .A1(n621), .A2(G902), .ZN(n377) );
  XNOR2_X1 U429 ( .A(n529), .B(n528), .ZN(n556) );
  INV_X1 U430 ( .A(G902), .ZN(n527) );
  INV_X1 U431 ( .A(n382), .ZN(n557) );
  NAND2_X1 U432 ( .A1(n698), .A2(G472), .ZN(n415) );
  INV_X1 U433 ( .A(KEYINPUT64), .ZN(n447) );
  BUF_X1 U434 ( .A(n698), .Z(n705) );
  NAND2_X1 U435 ( .A1(n698), .A2(G210), .ZN(n407) );
  AND2_X1 U436 ( .A1(n375), .A2(n571), .ZN(n664) );
  INV_X1 U437 ( .A(KEYINPUT92), .ZN(n432) );
  NAND2_X1 U438 ( .A1(n429), .A2(n374), .ZN(n373) );
  INV_X1 U439 ( .A(KEYINPUT15), .ZN(n453) );
  NAND2_X1 U440 ( .A1(G234), .A2(G237), .ZN(n491) );
  NOR2_X1 U441 ( .A1(G902), .A2(G237), .ZN(n454) );
  INV_X1 U442 ( .A(n662), .ZN(n438) );
  AND2_X1 U443 ( .A1(n671), .A2(n670), .ZN(n551) );
  XOR2_X1 U444 ( .A(KEYINPUT78), .B(KEYINPUT5), .Z(n459) );
  XNOR2_X1 U445 ( .A(G101), .B(KEYINPUT66), .ZN(n446) );
  XOR2_X1 U446 ( .A(G107), .B(G122), .Z(n519) );
  XNOR2_X1 U447 ( .A(G113), .B(G104), .ZN(n506) );
  XOR2_X1 U448 ( .A(KEYINPUT12), .B(KEYINPUT102), .Z(n507) );
  XOR2_X1 U449 ( .A(KEYINPUT103), .B(KEYINPUT11), .Z(n505) );
  XNOR2_X1 U450 ( .A(n388), .B(n452), .ZN(n385) );
  XNOR2_X1 U451 ( .A(n417), .B(n441), .ZN(n390) );
  XNOR2_X1 U452 ( .A(n393), .B(n392), .ZN(n719) );
  INV_X1 U453 ( .A(G110), .ZN(n392) );
  XNOR2_X1 U454 ( .A(G107), .B(G104), .ZN(n393) );
  XNOR2_X1 U455 ( .A(n421), .B(n419), .ZN(n479) );
  XNOR2_X1 U456 ( .A(n383), .B(KEYINPUT36), .ZN(n600) );
  XNOR2_X1 U457 ( .A(n573), .B(n400), .ZN(n651) );
  XNOR2_X1 U458 ( .A(KEYINPUT31), .B(KEYINPUT101), .ZN(n400) );
  NOR2_X1 U459 ( .A1(n574), .A2(n398), .ZN(n397) );
  INV_X1 U460 ( .A(n570), .ZN(n398) );
  INV_X1 U461 ( .A(n556), .ZN(n531) );
  XNOR2_X1 U462 ( .A(n415), .B(n362), .ZN(n414) );
  XNOR2_X1 U463 ( .A(n402), .B(n401), .ZN(n704) );
  INV_X1 U464 ( .A(n703), .ZN(n401) );
  NAND2_X1 U465 ( .A1(n705), .A2(G478), .ZN(n402) );
  INV_X1 U466 ( .A(KEYINPUT56), .ZN(n428) );
  NAND2_X1 U467 ( .A1(n406), .A2(n624), .ZN(n405) );
  XNOR2_X1 U468 ( .A(n407), .B(n702), .ZN(n406) );
  INV_X1 U469 ( .A(KEYINPUT53), .ZN(n394) );
  NAND2_X1 U470 ( .A1(n410), .A2(n408), .ZN(n395) );
  AND2_X1 U471 ( .A1(n697), .A2(n409), .ZN(n408) );
  AND2_X1 U472 ( .A1(G210), .A2(n466), .ZN(n352) );
  NAND2_X1 U473 ( .A1(n699), .A2(n352), .ZN(n436) );
  XOR2_X1 U474 ( .A(n505), .B(n504), .Z(n353) );
  XNOR2_X1 U475 ( .A(G122), .B(KEYINPUT16), .ZN(n354) );
  OR2_X1 U476 ( .A1(n664), .A2(n578), .ZN(n355) );
  AND2_X1 U477 ( .A1(n429), .A2(n368), .ZN(n356) );
  INV_X1 U478 ( .A(n431), .ZN(n429) );
  NAND2_X1 U479 ( .A1(n659), .A2(n432), .ZN(n431) );
  AND2_X1 U480 ( .A1(n435), .A2(KEYINPUT92), .ZN(n357) );
  AND2_X1 U481 ( .A1(n436), .A2(n435), .ZN(n358) );
  XOR2_X1 U482 ( .A(KEYINPUT35), .B(KEYINPUT87), .Z(n359) );
  XOR2_X1 U483 ( .A(KEYINPUT74), .B(KEYINPUT39), .Z(n360) );
  XOR2_X1 U484 ( .A(KEYINPUT6), .B(KEYINPUT107), .Z(n361) );
  INV_X1 U485 ( .A(n650), .ZN(n375) );
  INV_X1 U486 ( .A(n571), .ZN(n647) );
  XOR2_X1 U487 ( .A(n632), .B(KEYINPUT62), .Z(n362) );
  INV_X1 U488 ( .A(n390), .ZN(n379) );
  AND2_X1 U489 ( .A1(n592), .A2(n551), .ZN(n575) );
  NAND2_X1 U490 ( .A1(n550), .A2(n548), .ZN(n549) );
  XNOR2_X2 U491 ( .A(n542), .B(n541), .ZN(n550) );
  NAND2_X1 U492 ( .A1(n371), .A2(n436), .ZN(n370) );
  INV_X1 U493 ( .A(n567), .ZN(n399) );
  XNOR2_X1 U494 ( .A(n575), .B(KEYINPUT111), .ZN(n498) );
  XNOR2_X1 U495 ( .A(n364), .B(G119), .ZN(G21) );
  XNOR2_X2 U496 ( .A(n549), .B(KEYINPUT32), .ZN(n364) );
  OR2_X2 U497 ( .A1(n699), .A2(n434), .ZN(n433) );
  NAND2_X1 U498 ( .A1(n369), .A2(n367), .ZN(n366) );
  INV_X1 U499 ( .A(n435), .ZN(n368) );
  OR2_X1 U500 ( .A1(n699), .A2(n373), .ZN(n369) );
  INV_X1 U501 ( .A(n434), .ZN(n374) );
  NOR2_X2 U502 ( .A1(n577), .A2(n378), .ZN(n555) );
  NOR2_X1 U503 ( .A1(n693), .A2(n378), .ZN(n694) );
  NOR2_X1 U504 ( .A1(n668), .A2(n378), .ZN(n689) );
  XNOR2_X2 U505 ( .A(n553), .B(n554), .ZN(n378) );
  NAND2_X1 U506 ( .A1(n522), .A2(G217), .ZN(n523) );
  NAND2_X1 U507 ( .A1(n729), .A2(G234), .ZN(n381) );
  NAND2_X1 U508 ( .A1(n382), .A2(n556), .ZN(n571) );
  NAND2_X1 U509 ( .A1(n610), .A2(n384), .ZN(n383) );
  INV_X1 U510 ( .A(n417), .ZN(n384) );
  NOR2_X1 U511 ( .A1(n598), .A2(n599), .ZN(n610) );
  INV_X1 U512 ( .A(n387), .ZN(n404) );
  XNOR2_X2 U513 ( .A(n461), .B(n354), .ZN(n387) );
  XNOR2_X2 U514 ( .A(n418), .B(n445), .ZN(n461) );
  XNOR2_X2 U515 ( .A(n386), .B(n385), .ZN(n699) );
  XNOR2_X1 U516 ( .A(n449), .B(n389), .ZN(n388) );
  XNOR2_X1 U517 ( .A(n448), .B(n457), .ZN(n389) );
  XNOR2_X1 U518 ( .A(n391), .B(n353), .ZN(n514) );
  XNOR2_X1 U519 ( .A(n508), .B(n509), .ZN(n391) );
  NAND2_X1 U520 ( .A1(n426), .A2(n424), .ZN(n423) );
  XNOR2_X1 U521 ( .A(n423), .B(n580), .ZN(n713) );
  NOR2_X1 U522 ( .A1(n713), .A2(n728), .ZN(n619) );
  NOR2_X2 U523 ( .A1(n677), .A2(n676), .ZN(n572) );
  XNOR2_X1 U524 ( .A(n395), .B(n394), .ZN(G75) );
  XNOR2_X2 U525 ( .A(n396), .B(n359), .ZN(n736) );
  NAND2_X1 U526 ( .A1(n559), .A2(n558), .ZN(n396) );
  OR2_X2 U527 ( .A1(n577), .A2(n437), .ZN(n542) );
  NAND2_X1 U528 ( .A1(n399), .A2(n397), .ZN(n639) );
  XNOR2_X1 U529 ( .A(n405), .B(n428), .ZN(G51) );
  OR2_X2 U530 ( .A1(n628), .A2(G902), .ZN(n416) );
  NOR2_X2 U531 ( .A1(n625), .A2(n709), .ZN(n626) );
  XNOR2_X1 U532 ( .A(n404), .B(G101), .ZN(n718) );
  INV_X1 U533 ( .A(G953), .ZN(n409) );
  INV_X1 U534 ( .A(n657), .ZN(n411) );
  XNOR2_X1 U535 ( .A(n656), .B(KEYINPUT86), .ZN(n412) );
  XNOR2_X1 U536 ( .A(n413), .B(KEYINPUT63), .ZN(G57) );
  NAND2_X1 U537 ( .A1(n414), .A2(n624), .ZN(n413) );
  XNOR2_X2 U538 ( .A(n416), .B(G469), .ZN(n592) );
  NAND2_X1 U539 ( .A1(n530), .A2(n647), .ZN(n532) );
  XNOR2_X1 U540 ( .A(n502), .B(n360), .ZN(n530) );
  XNOR2_X1 U541 ( .A(n574), .B(n361), .ZN(n552) );
  XNOR2_X2 U542 ( .A(n422), .B(G472), .ZN(n574) );
  XNOR2_X1 U543 ( .A(n474), .B(n465), .ZN(n632) );
  NOR2_X2 U544 ( .A1(n736), .A2(KEYINPUT44), .ZN(n561) );
  NAND2_X1 U545 ( .A1(n565), .A2(n355), .ZN(n425) );
  NAND2_X1 U546 ( .A1(n563), .A2(n562), .ZN(n427) );
  NAND2_X1 U547 ( .A1(n358), .A2(n433), .ZN(n581) );
  NOR2_X1 U548 ( .A1(n659), .A2(n432), .ZN(n430) );
  XNOR2_X2 U549 ( .A(n439), .B(n539), .ZN(n577) );
  XOR2_X1 U550 ( .A(KEYINPUT19), .B(KEYINPUT80), .Z(n441) );
  INV_X1 U551 ( .A(KEYINPUT47), .ZN(n594) );
  INV_X1 U552 ( .A(n477), .ZN(n448) );
  INV_X1 U553 ( .A(KEYINPUT72), .ZN(n589) );
  INV_X1 U554 ( .A(n462), .ZN(n463) );
  XNOR2_X1 U555 ( .A(n590), .B(n589), .ZN(n599) );
  XNOR2_X1 U556 ( .A(n464), .B(n463), .ZN(n465) );
  INV_X1 U557 ( .A(n582), .ZN(n558) );
  XNOR2_X1 U558 ( .A(n479), .B(n724), .ZN(n481) );
  OR2_X1 U559 ( .A1(n729), .A2(G952), .ZN(n624) );
  INV_X1 U560 ( .A(n624), .ZN(n709) );
  XOR2_X1 U561 ( .A(G113), .B(G116), .Z(n445) );
  XNOR2_X1 U562 ( .A(n446), .B(KEYINPUT4), .ZN(n462) );
  XNOR2_X1 U563 ( .A(n719), .B(n462), .ZN(n472) );
  NAND2_X1 U564 ( .A1(n729), .A2(G224), .ZN(n449) );
  XNOR2_X2 U565 ( .A(G146), .B(G125), .ZN(n477) );
  XNOR2_X1 U566 ( .A(G143), .B(G128), .ZN(n457) );
  XNOR2_X1 U567 ( .A(KEYINPUT17), .B(KEYINPUT84), .ZN(n450) );
  XNOR2_X1 U568 ( .A(n451), .B(n450), .ZN(n452) );
  XNOR2_X1 U569 ( .A(n454), .B(KEYINPUT77), .ZN(n466) );
  INV_X1 U570 ( .A(KEYINPUT76), .ZN(n455) );
  XNOR2_X1 U571 ( .A(n455), .B(KEYINPUT38), .ZN(n456) );
  XNOR2_X1 U572 ( .A(n581), .B(n456), .ZN(n658) );
  XNOR2_X1 U573 ( .A(n457), .B(G134), .ZN(n525) );
  NAND2_X1 U574 ( .A1(n503), .A2(G210), .ZN(n458) );
  XNOR2_X1 U575 ( .A(n459), .B(n458), .ZN(n460) );
  XNOR2_X1 U576 ( .A(n461), .B(n460), .ZN(n464) );
  NAND2_X1 U577 ( .A1(G214), .A2(n466), .ZN(n659) );
  AND2_X1 U578 ( .A1(n574), .A2(n659), .ZN(n467) );
  XNOR2_X1 U579 ( .A(n467), .B(KEYINPUT30), .ZN(n584) );
  NAND2_X1 U580 ( .A1(n658), .A2(n584), .ZN(n501) );
  XNOR2_X1 U581 ( .A(KEYINPUT81), .B(KEYINPUT82), .ZN(n468) );
  XNOR2_X1 U582 ( .A(n478), .B(n468), .ZN(n470) );
  NAND2_X1 U583 ( .A1(n729), .A2(G227), .ZN(n469) );
  XNOR2_X1 U584 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U585 ( .A(n472), .B(n471), .ZN(n473) );
  XNOR2_X1 U586 ( .A(n474), .B(n473), .ZN(n628) );
  XNOR2_X1 U587 ( .A(KEYINPUT10), .B(n477), .ZN(n509) );
  XNOR2_X1 U588 ( .A(n509), .B(n478), .ZN(n724) );
  NAND2_X1 U589 ( .A1(G221), .A2(n522), .ZN(n480) );
  XNOR2_X1 U590 ( .A(n481), .B(n480), .ZN(n706) );
  XOR2_X1 U591 ( .A(KEYINPUT100), .B(KEYINPUT25), .Z(n485) );
  INV_X1 U592 ( .A(n618), .ZN(n482) );
  NAND2_X1 U593 ( .A1(G234), .A2(n482), .ZN(n483) );
  XNOR2_X1 U594 ( .A(KEYINPUT20), .B(n483), .ZN(n488) );
  NAND2_X1 U595 ( .A1(n488), .A2(G217), .ZN(n484) );
  XNOR2_X1 U596 ( .A(n485), .B(n484), .ZN(n486) );
  XNOR2_X2 U597 ( .A(n487), .B(n486), .ZN(n671) );
  NAND2_X1 U598 ( .A1(n488), .A2(G221), .ZN(n490) );
  INV_X1 U599 ( .A(KEYINPUT21), .ZN(n489) );
  XNOR2_X1 U600 ( .A(n491), .B(KEYINPUT94), .ZN(n492) );
  XNOR2_X1 U601 ( .A(KEYINPUT14), .B(n492), .ZN(n494) );
  NAND2_X1 U602 ( .A1(n494), .A2(G952), .ZN(n493) );
  XOR2_X1 U603 ( .A(KEYINPUT95), .B(n493), .Z(n692) );
  NOR2_X1 U604 ( .A1(n692), .A2(G953), .ZN(n537) );
  NAND2_X1 U605 ( .A1(n494), .A2(G902), .ZN(n495) );
  XOR2_X1 U606 ( .A(n495), .B(KEYINPUT97), .Z(n534) );
  OR2_X1 U607 ( .A1(n729), .A2(G900), .ZN(n496) );
  NOR2_X1 U608 ( .A1(n534), .A2(n496), .ZN(n497) );
  NOR2_X1 U609 ( .A1(n537), .A2(n497), .ZN(n588) );
  OR2_X1 U610 ( .A1(n498), .A2(n588), .ZN(n500) );
  INV_X1 U611 ( .A(KEYINPUT79), .ZN(n499) );
  XNOR2_X1 U612 ( .A(n500), .B(n499), .ZN(n585) );
  NAND2_X1 U613 ( .A1(G214), .A2(n503), .ZN(n504) );
  XNOR2_X1 U614 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U615 ( .A(G143), .B(G122), .ZN(n510) );
  XNOR2_X1 U616 ( .A(n510), .B(G140), .ZN(n512) );
  XNOR2_X1 U617 ( .A(n511), .B(n512), .ZN(n513) );
  XNOR2_X1 U618 ( .A(n514), .B(n513), .ZN(n621) );
  XNOR2_X1 U619 ( .A(KEYINPUT104), .B(KEYINPUT13), .ZN(n515) );
  INV_X1 U620 ( .A(G475), .ZN(n516) );
  XNOR2_X1 U621 ( .A(G116), .B(KEYINPUT105), .ZN(n517) );
  XNOR2_X1 U622 ( .A(n517), .B(KEYINPUT7), .ZN(n521) );
  XNOR2_X1 U623 ( .A(KEYINPUT106), .B(KEYINPUT9), .ZN(n518) );
  XNOR2_X1 U624 ( .A(n519), .B(n518), .ZN(n520) );
  XOR2_X1 U625 ( .A(n521), .B(n520), .Z(n524) );
  XNOR2_X1 U626 ( .A(n524), .B(n523), .ZN(n526) );
  XNOR2_X1 U627 ( .A(n526), .B(n525), .ZN(n703) );
  NAND2_X1 U628 ( .A1(n703), .A2(n527), .ZN(n529) );
  INV_X1 U629 ( .A(G478), .ZN(n528) );
  AND2_X1 U630 ( .A1(n557), .A2(n531), .ZN(n650) );
  AND2_X1 U631 ( .A1(n530), .A2(n650), .ZN(n615) );
  XOR2_X1 U632 ( .A(G134), .B(n615), .Z(G36) );
  XOR2_X1 U633 ( .A(G131), .B(KEYINPUT126), .Z(n533) );
  XOR2_X1 U634 ( .A(n533), .B(n605), .Z(G33) );
  XOR2_X1 U635 ( .A(G898), .B(KEYINPUT96), .Z(n712) );
  NAND2_X1 U636 ( .A1(G953), .A2(n712), .ZN(n721) );
  NOR2_X1 U637 ( .A1(n534), .A2(n721), .ZN(n535) );
  XNOR2_X1 U638 ( .A(n535), .B(KEYINPUT98), .ZN(n536) );
  NOR2_X1 U639 ( .A1(n537), .A2(n536), .ZN(n538) );
  XNOR2_X1 U640 ( .A(KEYINPUT65), .B(KEYINPUT0), .ZN(n539) );
  NAND2_X1 U641 ( .A1(n556), .A2(n557), .ZN(n540) );
  XNOR2_X1 U642 ( .A(n540), .B(KEYINPUT108), .ZN(n662) );
  INV_X1 U643 ( .A(KEYINPUT1), .ZN(n543) );
  INV_X1 U644 ( .A(n677), .ZN(n544) );
  INV_X1 U645 ( .A(n671), .ZN(n570) );
  NAND2_X1 U646 ( .A1(n544), .A2(n570), .ZN(n545) );
  XNOR2_X1 U647 ( .A(n545), .B(KEYINPUT109), .ZN(n546) );
  NAND2_X1 U648 ( .A1(n546), .A2(n552), .ZN(n547) );
  XNOR2_X1 U649 ( .A(n547), .B(KEYINPUT85), .ZN(n548) );
  NAND2_X1 U650 ( .A1(n550), .A2(n363), .ZN(n567) );
  XNOR2_X1 U651 ( .A(n564), .B(KEYINPUT91), .ZN(n563) );
  XOR2_X1 U652 ( .A(KEYINPUT110), .B(KEYINPUT33), .Z(n554) );
  INV_X1 U653 ( .A(n551), .ZN(n676) );
  INV_X1 U654 ( .A(n552), .ZN(n597) );
  NAND2_X1 U655 ( .A1(n572), .A2(n597), .ZN(n553) );
  XNOR2_X1 U656 ( .A(n555), .B(KEYINPUT34), .ZN(n559) );
  OR2_X1 U657 ( .A1(n557), .A2(n556), .ZN(n582) );
  XNOR2_X1 U658 ( .A(n561), .B(n560), .ZN(n562) );
  NAND2_X1 U659 ( .A1(n564), .A2(KEYINPUT44), .ZN(n565) );
  NAND2_X1 U660 ( .A1(KEYINPUT44), .A2(n736), .ZN(n566) );
  XNOR2_X1 U661 ( .A(n566), .B(KEYINPUT90), .ZN(n579) );
  NOR2_X1 U662 ( .A1(n597), .A2(n567), .ZN(n568) );
  XNOR2_X1 U663 ( .A(n568), .B(KEYINPUT89), .ZN(n569) );
  NOR2_X1 U664 ( .A1(n570), .A2(n569), .ZN(n633) );
  NAND2_X1 U665 ( .A1(n574), .A2(n572), .ZN(n682) );
  NOR2_X1 U666 ( .A1(n577), .A2(n682), .ZN(n573) );
  INV_X1 U667 ( .A(n574), .ZN(n673) );
  NAND2_X1 U668 ( .A1(n575), .A2(n673), .ZN(n576) );
  NOR2_X1 U669 ( .A1(n577), .A2(n576), .ZN(n635) );
  NOR2_X1 U670 ( .A1(n651), .A2(n635), .ZN(n578) );
  INV_X1 U671 ( .A(KEYINPUT45), .ZN(n580) );
  INV_X1 U672 ( .A(n581), .ZN(n613) );
  NOR2_X1 U673 ( .A1(n613), .A2(n582), .ZN(n583) );
  NAND2_X1 U674 ( .A1(n584), .A2(n583), .ZN(n586) );
  NOR2_X1 U675 ( .A1(n586), .A2(n585), .ZN(n643) );
  INV_X1 U676 ( .A(n670), .ZN(n587) );
  NOR2_X1 U677 ( .A1(n671), .A2(n440), .ZN(n590) );
  XNOR2_X1 U678 ( .A(n591), .B(KEYINPUT28), .ZN(n593) );
  NAND2_X1 U679 ( .A1(n593), .A2(n592), .ZN(n602) );
  NOR2_X1 U680 ( .A1(n643), .A2(n595), .ZN(n596) );
  NAND2_X1 U681 ( .A1(n647), .A2(n597), .ZN(n598) );
  NOR2_X1 U682 ( .A1(n600), .A2(n363), .ZN(n653) );
  NAND2_X1 U683 ( .A1(n659), .A2(n658), .ZN(n665) );
  NOR2_X1 U684 ( .A1(n665), .A2(n662), .ZN(n601) );
  XNOR2_X1 U685 ( .A(n601), .B(KEYINPUT41), .ZN(n693) );
  NOR2_X1 U686 ( .A1(n693), .A2(n602), .ZN(n603) );
  XNOR2_X1 U687 ( .A(n603), .B(KEYINPUT42), .ZN(n737) );
  INV_X1 U688 ( .A(n737), .ZN(n604) );
  INV_X1 U689 ( .A(KEYINPUT46), .ZN(n606) );
  INV_X1 U690 ( .A(KEYINPUT88), .ZN(n607) );
  XNOR2_X1 U691 ( .A(n607), .B(KEYINPUT48), .ZN(n608) );
  XNOR2_X1 U692 ( .A(n609), .B(n608), .ZN(n617) );
  AND2_X1 U693 ( .A1(n610), .A2(n659), .ZN(n611) );
  NAND2_X1 U694 ( .A1(n611), .A2(n363), .ZN(n612) );
  XNOR2_X1 U695 ( .A(n612), .B(KEYINPUT43), .ZN(n614) );
  AND2_X1 U696 ( .A1(n614), .A2(n613), .ZN(n655) );
  NOR2_X1 U697 ( .A1(n615), .A2(n655), .ZN(n616) );
  NAND2_X1 U698 ( .A1(n617), .A2(n616), .ZN(n728) );
  NAND2_X1 U699 ( .A1(n619), .A2(KEYINPUT2), .ZN(n657) );
  NOR2_X1 U700 ( .A1(n619), .A2(KEYINPUT2), .ZN(n656) );
  NAND2_X1 U701 ( .A1(n698), .A2(G475), .ZN(n623) );
  XNOR2_X1 U702 ( .A(n623), .B(n622), .ZN(n625) );
  XNOR2_X1 U703 ( .A(n626), .B(KEYINPUT60), .ZN(G60) );
  NAND2_X1 U704 ( .A1(n705), .A2(G469), .ZN(n630) );
  XOR2_X1 U705 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n627) );
  XNOR2_X1 U706 ( .A(n628), .B(n627), .ZN(n629) );
  XNOR2_X1 U707 ( .A(n630), .B(n629), .ZN(n631) );
  NOR2_X1 U708 ( .A1(n631), .A2(n709), .ZN(G54) );
  XOR2_X1 U709 ( .A(n633), .B(G101), .Z(G3) );
  NAND2_X1 U710 ( .A1(n635), .A2(n647), .ZN(n634) );
  XNOR2_X1 U711 ( .A(n634), .B(G104), .ZN(G6) );
  XOR2_X1 U712 ( .A(KEYINPUT27), .B(KEYINPUT26), .Z(n637) );
  NAND2_X1 U713 ( .A1(n635), .A2(n650), .ZN(n636) );
  XNOR2_X1 U714 ( .A(n637), .B(n636), .ZN(n638) );
  XNOR2_X1 U715 ( .A(G107), .B(n638), .ZN(G9) );
  XNOR2_X1 U716 ( .A(n639), .B(G110), .ZN(G12) );
  NOR2_X1 U717 ( .A1(n375), .A2(n644), .ZN(n641) );
  XNOR2_X1 U718 ( .A(KEYINPUT112), .B(KEYINPUT29), .ZN(n640) );
  XNOR2_X1 U719 ( .A(n641), .B(n640), .ZN(n642) );
  XNOR2_X1 U720 ( .A(G128), .B(n642), .ZN(G30) );
  XOR2_X1 U721 ( .A(G143), .B(n643), .Z(G45) );
  NOR2_X1 U722 ( .A1(n571), .A2(n644), .ZN(n646) );
  XNOR2_X1 U723 ( .A(G146), .B(KEYINPUT113), .ZN(n645) );
  XNOR2_X1 U724 ( .A(n646), .B(n645), .ZN(G48) );
  NAND2_X1 U725 ( .A1(n651), .A2(n647), .ZN(n648) );
  XNOR2_X1 U726 ( .A(n648), .B(KEYINPUT114), .ZN(n649) );
  XNOR2_X1 U727 ( .A(G113), .B(n649), .ZN(G15) );
  NAND2_X1 U728 ( .A1(n651), .A2(n650), .ZN(n652) );
  XNOR2_X1 U729 ( .A(n652), .B(G116), .ZN(G18) );
  XNOR2_X1 U730 ( .A(G125), .B(n653), .ZN(n654) );
  XNOR2_X1 U731 ( .A(n654), .B(KEYINPUT37), .ZN(G27) );
  XOR2_X1 U732 ( .A(G140), .B(n655), .Z(G42) );
  NOR2_X1 U733 ( .A1(n659), .A2(n658), .ZN(n660) );
  XNOR2_X1 U734 ( .A(n660), .B(KEYINPUT120), .ZN(n661) );
  NOR2_X1 U735 ( .A1(n662), .A2(n661), .ZN(n663) );
  XOR2_X1 U736 ( .A(KEYINPUT121), .B(n663), .Z(n667) );
  NOR2_X1 U737 ( .A1(n665), .A2(n664), .ZN(n666) );
  NOR2_X1 U738 ( .A1(n667), .A2(n666), .ZN(n668) );
  XNOR2_X1 U739 ( .A(KEYINPUT117), .B(KEYINPUT118), .ZN(n669) );
  XNOR2_X1 U740 ( .A(n669), .B(KEYINPUT51), .ZN(n685) );
  NOR2_X1 U741 ( .A1(n671), .A2(n670), .ZN(n672) );
  XNOR2_X1 U742 ( .A(n672), .B(KEYINPUT49), .ZN(n674) );
  NAND2_X1 U743 ( .A1(n674), .A2(n673), .ZN(n675) );
  XNOR2_X1 U744 ( .A(KEYINPUT115), .B(n675), .ZN(n680) );
  NAND2_X1 U745 ( .A1(n363), .A2(n676), .ZN(n678) );
  XNOR2_X1 U746 ( .A(KEYINPUT50), .B(n678), .ZN(n679) );
  NAND2_X1 U747 ( .A1(n680), .A2(n679), .ZN(n681) );
  XNOR2_X1 U748 ( .A(n681), .B(KEYINPUT116), .ZN(n683) );
  NAND2_X1 U749 ( .A1(n683), .A2(n682), .ZN(n684) );
  XOR2_X1 U750 ( .A(n685), .B(n684), .Z(n686) );
  NOR2_X1 U751 ( .A1(n693), .A2(n686), .ZN(n687) );
  XOR2_X1 U752 ( .A(KEYINPUT119), .B(n687), .Z(n688) );
  NOR2_X1 U753 ( .A1(n689), .A2(n688), .ZN(n690) );
  XNOR2_X1 U754 ( .A(n690), .B(KEYINPUT52), .ZN(n691) );
  NOR2_X1 U755 ( .A1(n692), .A2(n691), .ZN(n695) );
  NOR2_X1 U756 ( .A1(n695), .A2(n694), .ZN(n696) );
  XNOR2_X1 U757 ( .A(n696), .B(KEYINPUT122), .ZN(n697) );
  XOR2_X1 U758 ( .A(KEYINPUT54), .B(KEYINPUT55), .Z(n701) );
  XNOR2_X1 U759 ( .A(n699), .B(KEYINPUT93), .ZN(n700) );
  XNOR2_X1 U760 ( .A(n701), .B(n700), .ZN(n702) );
  NOR2_X1 U761 ( .A1(n709), .A2(n704), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n705), .A2(G217), .ZN(n707) );
  XNOR2_X1 U763 ( .A(n707), .B(n706), .ZN(n708) );
  NOR2_X1 U764 ( .A1(n709), .A2(n708), .ZN(G66) );
  NAND2_X1 U765 ( .A1(G953), .A2(G224), .ZN(n710) );
  XOR2_X1 U766 ( .A(KEYINPUT61), .B(n710), .Z(n711) );
  NOR2_X1 U767 ( .A1(n712), .A2(n711), .ZN(n716) );
  NOR2_X1 U768 ( .A1(G953), .A2(n713), .ZN(n714) );
  XOR2_X1 U769 ( .A(KEYINPUT123), .B(n714), .Z(n715) );
  NOR2_X1 U770 ( .A1(n716), .A2(n715), .ZN(n717) );
  XOR2_X1 U771 ( .A(KEYINPUT124), .B(n717), .Z(n723) );
  XNOR2_X1 U772 ( .A(n719), .B(n718), .ZN(n720) );
  NAND2_X1 U773 ( .A1(n721), .A2(n720), .ZN(n722) );
  XOR2_X1 U774 ( .A(n723), .B(n722), .Z(G69) );
  XNOR2_X1 U775 ( .A(n724), .B(KEYINPUT125), .ZN(n725) );
  XNOR2_X1 U776 ( .A(n725), .B(KEYINPUT4), .ZN(n726) );
  XOR2_X1 U777 ( .A(n727), .B(n726), .Z(n731) );
  XNOR2_X1 U778 ( .A(n728), .B(n731), .ZN(n730) );
  NAND2_X1 U779 ( .A1(n730), .A2(n729), .ZN(n735) );
  XNOR2_X1 U780 ( .A(G227), .B(n731), .ZN(n732) );
  NAND2_X1 U781 ( .A1(n732), .A2(G900), .ZN(n733) );
  NAND2_X1 U782 ( .A1(n733), .A2(G953), .ZN(n734) );
  NAND2_X1 U783 ( .A1(n735), .A2(n734), .ZN(G72) );
  XOR2_X1 U784 ( .A(n736), .B(G122), .Z(G24) );
  XOR2_X1 U785 ( .A(G137), .B(n737), .Z(G39) );
endmodule

