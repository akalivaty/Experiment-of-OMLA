//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 1 1 0 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 0 0 1 1 1 0 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 1 1 0 1 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n698, new_n699,
    new_n700, new_n701, new_n702, new_n703, new_n704, new_n705, new_n707,
    new_n708, new_n709, new_n710, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n790, new_n791,
    new_n792, new_n793, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n800, new_n802, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n812, new_n813, new_n814, new_n815, new_n816,
    new_n817, new_n818, new_n819, new_n821, new_n822, new_n823, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n867, new_n868, new_n870,
    new_n871, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n919, new_n920, new_n922, new_n923, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n981,
    new_n982, new_n983;
  INV_X1    g000(.A(KEYINPUT80), .ZN(new_n202));
  INV_X1    g001(.A(G141gat), .ZN(new_n203));
  NAND2_X1  g002(.A1(new_n203), .A2(G148gat), .ZN(new_n204));
  INV_X1    g003(.A(G148gat), .ZN(new_n205));
  NAND2_X1  g004(.A1(new_n205), .A2(G141gat), .ZN(new_n206));
  NAND2_X1  g005(.A1(new_n204), .A2(new_n206), .ZN(new_n207));
  XNOR2_X1  g006(.A(G155gat), .B(G162gat), .ZN(new_n208));
  INV_X1    g007(.A(G155gat), .ZN(new_n209));
  INV_X1    g008(.A(G162gat), .ZN(new_n210));
  OAI21_X1  g009(.A(KEYINPUT2), .B1(new_n209), .B2(new_n210), .ZN(new_n211));
  AND3_X1   g010(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n212));
  AOI21_X1  g011(.A(new_n208), .B1(new_n211), .B2(new_n207), .ZN(new_n213));
  OAI21_X1  g012(.A(new_n202), .B1(new_n212), .B2(new_n213), .ZN(new_n214));
  AND2_X1   g013(.A1(G155gat), .A2(G162gat), .ZN(new_n215));
  NOR2_X1   g014(.A1(G155gat), .A2(G162gat), .ZN(new_n216));
  NOR2_X1   g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  XNOR2_X1  g016(.A(G141gat), .B(G148gat), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT2), .ZN(new_n219));
  AOI21_X1  g018(.A(new_n219), .B1(G155gat), .B2(G162gat), .ZN(new_n220));
  OAI21_X1  g019(.A(new_n217), .B1(new_n218), .B2(new_n220), .ZN(new_n221));
  NAND3_X1  g020(.A1(new_n207), .A2(new_n208), .A3(new_n211), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n221), .A2(new_n222), .A3(KEYINPUT80), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n214), .A2(new_n223), .ZN(new_n224));
  AND2_X1   g023(.A1(G211gat), .A2(G218gat), .ZN(new_n225));
  NOR2_X1   g024(.A1(G211gat), .A2(G218gat), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT77), .ZN(new_n227));
  OR3_X1    g026(.A1(new_n225), .A2(new_n226), .A3(new_n227), .ZN(new_n228));
  OAI21_X1  g027(.A(new_n227), .B1(new_n225), .B2(new_n226), .ZN(new_n229));
  NAND2_X1  g028(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  INV_X1    g029(.A(G197gat), .ZN(new_n231));
  INV_X1    g030(.A(G204gat), .ZN(new_n232));
  NAND2_X1  g031(.A1(new_n231), .A2(new_n232), .ZN(new_n233));
  NAND2_X1  g032(.A1(G197gat), .A2(G204gat), .ZN(new_n234));
  INV_X1    g033(.A(KEYINPUT22), .ZN(new_n235));
  NAND2_X1  g034(.A1(G211gat), .A2(G218gat), .ZN(new_n236));
  AOI22_X1  g035(.A1(new_n233), .A2(new_n234), .B1(new_n235), .B2(new_n236), .ZN(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n230), .A2(new_n238), .ZN(new_n239));
  INV_X1    g038(.A(KEYINPUT29), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n228), .A2(new_n229), .A3(new_n237), .ZN(new_n241));
  NAND3_X1  g040(.A1(new_n239), .A2(new_n240), .A3(new_n241), .ZN(new_n242));
  AOI21_X1  g041(.A(KEYINPUT3), .B1(new_n242), .B2(KEYINPUT87), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT87), .ZN(new_n244));
  NAND4_X1  g043(.A1(new_n239), .A2(new_n244), .A3(new_n240), .A4(new_n241), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n224), .B1(new_n243), .B2(new_n245), .ZN(new_n246));
  INV_X1    g045(.A(G228gat), .ZN(new_n247));
  INV_X1    g046(.A(G233gat), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT76), .ZN(new_n250));
  OAI21_X1  g049(.A(new_n237), .B1(new_n230), .B2(new_n250), .ZN(new_n251));
  NAND4_X1  g050(.A1(new_n238), .A2(KEYINPUT76), .A3(new_n228), .A4(new_n229), .ZN(new_n252));
  NAND2_X1  g051(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n221), .A2(new_n222), .ZN(new_n254));
  OR2_X1    g053(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n255));
  AOI21_X1  g054(.A(new_n253), .B1(new_n240), .B2(new_n255), .ZN(new_n256));
  OR3_X1    g055(.A1(new_n246), .A2(new_n249), .A3(new_n256), .ZN(new_n257));
  INV_X1    g056(.A(G22gat), .ZN(new_n258));
  AOI21_X1  g057(.A(KEYINPUT29), .B1(new_n251), .B2(new_n252), .ZN(new_n259));
  OAI21_X1  g058(.A(new_n254), .B1(new_n259), .B2(KEYINPUT3), .ZN(new_n260));
  INV_X1    g059(.A(new_n253), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n255), .A2(new_n240), .ZN(new_n262));
  NAND2_X1  g061(.A1(new_n261), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n260), .A2(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n264), .A2(new_n249), .ZN(new_n265));
  NAND3_X1  g064(.A1(new_n257), .A2(new_n258), .A3(new_n265), .ZN(new_n266));
  NOR3_X1   g065(.A1(new_n246), .A2(new_n249), .A3(new_n256), .ZN(new_n267));
  AOI211_X1 g066(.A(new_n247), .B(new_n248), .C1(new_n260), .C2(new_n263), .ZN(new_n268));
  OAI21_X1  g067(.A(G22gat), .B1(new_n267), .B2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT86), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n269), .A3(new_n270), .ZN(new_n271));
  XNOR2_X1  g070(.A(G78gat), .B(G106gat), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  XNOR2_X1  g072(.A(KEYINPUT85), .B(KEYINPUT31), .ZN(new_n274));
  INV_X1    g073(.A(G50gat), .ZN(new_n275));
  XNOR2_X1  g074(.A(new_n274), .B(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n272), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n266), .A2(new_n269), .A3(new_n270), .A4(new_n277), .ZN(new_n278));
  AND3_X1   g077(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n276), .B1(new_n273), .B2(new_n278), .ZN(new_n280));
  NOR2_X1   g079(.A1(new_n279), .A2(new_n280), .ZN(new_n281));
  NAND2_X1  g080(.A1(G169gat), .A2(G176gat), .ZN(new_n282));
  NOR2_X1   g081(.A1(G169gat), .A2(G176gat), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n282), .B1(new_n283), .B2(KEYINPUT23), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n283), .A2(KEYINPUT23), .ZN(new_n286));
  AOI21_X1  g085(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n287));
  XNOR2_X1  g086(.A(new_n287), .B(KEYINPUT65), .ZN(new_n288));
  NAND3_X1  g087(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n289));
  OAI21_X1  g088(.A(new_n289), .B1(G183gat), .B2(G190gat), .ZN(new_n290));
  OAI211_X1 g089(.A(new_n285), .B(new_n286), .C1(new_n288), .C2(new_n290), .ZN(new_n291));
  XNOR2_X1  g090(.A(KEYINPUT64), .B(G176gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G169gat), .ZN(new_n293));
  AOI21_X1  g092(.A(new_n284), .B1(new_n293), .B2(KEYINPUT23), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n290), .A2(new_n287), .ZN(new_n295));
  NOR2_X1   g094(.A1(new_n295), .A2(KEYINPUT25), .ZN(new_n296));
  AOI22_X1  g095(.A1(new_n291), .A2(KEYINPUT25), .B1(new_n294), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT66), .ZN(new_n298));
  INV_X1    g097(.A(G183gat), .ZN(new_n299));
  OAI21_X1  g098(.A(KEYINPUT27), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT28), .ZN(new_n301));
  INV_X1    g100(.A(G190gat), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT27), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n303), .A2(KEYINPUT66), .A3(G183gat), .ZN(new_n304));
  NAND4_X1  g103(.A1(new_n300), .A2(new_n301), .A3(new_n302), .A4(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  XNOR2_X1  g105(.A(KEYINPUT27), .B(G183gat), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n301), .B1(new_n307), .B2(new_n302), .ZN(new_n308));
  OAI21_X1  g107(.A(KEYINPUT67), .B1(new_n306), .B2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(KEYINPUT67), .ZN(new_n310));
  AND2_X1   g109(.A1(new_n307), .A2(new_n302), .ZN(new_n311));
  OAI211_X1 g110(.A(new_n310), .B(new_n305), .C1(new_n311), .C2(new_n301), .ZN(new_n312));
  INV_X1    g111(.A(new_n283), .ZN(new_n313));
  OR2_X1    g112(.A1(new_n313), .A2(KEYINPUT26), .ZN(new_n314));
  INV_X1    g113(.A(new_n282), .ZN(new_n315));
  AOI21_X1  g114(.A(new_n315), .B1(new_n313), .B2(KEYINPUT26), .ZN(new_n316));
  AOI22_X1  g115(.A1(new_n314), .A2(new_n316), .B1(G183gat), .B2(G190gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n309), .A2(new_n312), .A3(new_n317), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n297), .A2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT1), .ZN(new_n320));
  INV_X1    g119(.A(G113gat), .ZN(new_n321));
  NOR2_X1   g120(.A1(new_n321), .A2(G120gat), .ZN(new_n322));
  INV_X1    g121(.A(G120gat), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n323), .A2(G113gat), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n320), .B1(new_n322), .B2(new_n324), .ZN(new_n325));
  INV_X1    g124(.A(G127gat), .ZN(new_n326));
  NAND2_X1  g125(.A1(new_n326), .A2(G134gat), .ZN(new_n327));
  INV_X1    g126(.A(G134gat), .ZN(new_n328));
  NAND2_X1  g127(.A1(new_n328), .A2(G127gat), .ZN(new_n329));
  NAND2_X1  g128(.A1(new_n327), .A2(new_n329), .ZN(new_n330));
  NOR2_X1   g129(.A1(new_n325), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n327), .A2(new_n329), .A3(KEYINPUT68), .ZN(new_n333));
  OR3_X1    g132(.A1(new_n328), .A2(KEYINPUT68), .A3(G127gat), .ZN(new_n334));
  XNOR2_X1  g133(.A(G113gat), .B(G120gat), .ZN(new_n335));
  OAI211_X1 g134(.A(new_n333), .B(new_n334), .C1(KEYINPUT1), .C2(new_n335), .ZN(new_n336));
  AND2_X1   g135(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT69), .ZN(new_n338));
  NAND4_X1  g137(.A1(new_n325), .A2(new_n338), .A3(new_n334), .A4(new_n333), .ZN(new_n339));
  INV_X1    g138(.A(new_n339), .ZN(new_n340));
  OAI21_X1  g139(.A(new_n332), .B1(new_n337), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n319), .A2(new_n341), .ZN(new_n342));
  INV_X1    g141(.A(G227gat), .ZN(new_n343));
  NOR2_X1   g142(.A1(new_n343), .A2(new_n248), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n336), .A2(KEYINPUT69), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n331), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n346), .B1(new_n297), .B2(new_n318), .ZN(new_n347));
  NOR3_X1   g146(.A1(new_n342), .A2(new_n344), .A3(new_n347), .ZN(new_n348));
  AND2_X1   g147(.A1(KEYINPUT72), .A2(KEYINPUT34), .ZN(new_n349));
  NAND2_X1  g148(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  XNOR2_X1  g149(.A(KEYINPUT72), .B(KEYINPUT34), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n350), .B1(new_n348), .B2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n352), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n344), .B1(new_n342), .B2(new_n347), .ZN(new_n354));
  INV_X1    g153(.A(KEYINPUT70), .ZN(new_n355));
  OR2_X1    g154(.A1(new_n355), .A2(KEYINPUT33), .ZN(new_n356));
  NAND2_X1  g155(.A1(new_n355), .A2(KEYINPUT33), .ZN(new_n357));
  NAND3_X1  g156(.A1(new_n354), .A2(new_n356), .A3(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n354), .A2(KEYINPUT32), .ZN(new_n359));
  XNOR2_X1  g158(.A(G15gat), .B(G43gat), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n360), .B(G99gat), .ZN(new_n361));
  XNOR2_X1  g160(.A(KEYINPUT71), .B(G71gat), .ZN(new_n362));
  XNOR2_X1  g161(.A(new_n361), .B(new_n362), .ZN(new_n363));
  AND3_X1   g162(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n359), .B1(new_n358), .B2(new_n363), .ZN(new_n365));
  OAI21_X1  g164(.A(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(KEYINPUT73), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT73), .ZN(new_n368));
  OAI211_X1 g167(.A(new_n353), .B(new_n368), .C1(new_n364), .C2(new_n365), .ZN(new_n369));
  INV_X1    g168(.A(KEYINPUT74), .ZN(new_n370));
  NOR2_X1   g169(.A1(new_n364), .A2(new_n365), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n370), .B1(new_n371), .B2(new_n352), .ZN(new_n372));
  NAND2_X1  g171(.A1(new_n358), .A2(new_n363), .ZN(new_n373));
  INV_X1    g172(.A(new_n359), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n363), .ZN(new_n376));
  AND4_X1   g175(.A1(new_n370), .A2(new_n375), .A3(new_n376), .A4(new_n352), .ZN(new_n377));
  OAI211_X1 g176(.A(new_n367), .B(new_n369), .C1(new_n372), .C2(new_n377), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n281), .A2(new_n378), .ZN(new_n379));
  AOI21_X1  g178(.A(KEYINPUT29), .B1(new_n297), .B2(new_n318), .ZN(new_n380));
  NAND2_X1  g179(.A1(G226gat), .A2(G233gat), .ZN(new_n381));
  XOR2_X1   g180(.A(new_n381), .B(KEYINPUT78), .Z(new_n382));
  INV_X1    g181(.A(new_n319), .ZN(new_n383));
  OAI221_X1 g182(.A(new_n261), .B1(new_n380), .B2(new_n382), .C1(new_n381), .C2(new_n383), .ZN(new_n384));
  AND2_X1   g183(.A1(new_n319), .A2(new_n382), .ZN(new_n385));
  INV_X1    g184(.A(new_n381), .ZN(new_n386));
  AOI21_X1  g185(.A(new_n386), .B1(new_n319), .B2(new_n240), .ZN(new_n387));
  OAI21_X1  g186(.A(new_n253), .B1(new_n385), .B2(new_n387), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n384), .A2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G8gat), .B(G36gat), .ZN(new_n390));
  INV_X1    g189(.A(G64gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  INV_X1    g191(.A(G92gat), .ZN(new_n393));
  XNOR2_X1  g192(.A(new_n392), .B(new_n393), .ZN(new_n394));
  INV_X1    g193(.A(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n389), .A2(new_n395), .ZN(new_n396));
  NAND2_X1  g195(.A1(new_n396), .A2(KEYINPUT79), .ZN(new_n397));
  INV_X1    g196(.A(KEYINPUT30), .ZN(new_n398));
  INV_X1    g197(.A(KEYINPUT79), .ZN(new_n399));
  NAND3_X1  g198(.A1(new_n389), .A2(new_n399), .A3(new_n395), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n397), .A2(new_n398), .A3(new_n400), .ZN(new_n401));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n388), .A3(new_n394), .ZN(new_n402));
  NAND3_X1  g201(.A1(new_n389), .A2(KEYINPUT30), .A3(new_n395), .ZN(new_n403));
  NAND3_X1  g202(.A1(new_n401), .A2(new_n402), .A3(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(G225gat), .A2(G233gat), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n254), .A2(KEYINPUT3), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n255), .A2(new_n407), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n406), .B1(new_n408), .B2(new_n346), .ZN(new_n409));
  INV_X1    g208(.A(new_n409), .ZN(new_n410));
  INV_X1    g209(.A(new_n254), .ZN(new_n411));
  OAI211_X1 g210(.A(new_n332), .B(new_n411), .C1(new_n337), .C2(new_n340), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT83), .ZN(new_n413));
  NAND3_X1  g212(.A1(new_n412), .A2(new_n413), .A3(KEYINPUT4), .ZN(new_n414));
  INV_X1    g213(.A(KEYINPUT4), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n346), .A2(new_n224), .A3(new_n415), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AOI21_X1  g216(.A(new_n413), .B1(new_n412), .B2(KEYINPUT4), .ZN(new_n418));
  OAI211_X1 g217(.A(new_n405), .B(new_n410), .C1(new_n417), .C2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(new_n419), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT82), .ZN(new_n421));
  NAND2_X1  g220(.A1(new_n341), .A2(new_n254), .ZN(new_n422));
  AOI21_X1  g221(.A(KEYINPUT81), .B1(new_n346), .B2(new_n411), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(new_n406), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n341), .A2(KEYINPUT81), .A3(new_n254), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n346), .A2(new_n224), .A3(KEYINPUT4), .ZN(new_n428));
  AOI211_X1 g227(.A(new_n331), .B(new_n254), .C1(new_n345), .C2(new_n339), .ZN(new_n429));
  OAI21_X1  g228(.A(new_n428), .B1(KEYINPUT4), .B2(new_n429), .ZN(new_n430));
  OAI21_X1  g229(.A(KEYINPUT5), .B1(new_n430), .B2(new_n409), .ZN(new_n431));
  OAI21_X1  g230(.A(new_n421), .B1(new_n427), .B2(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n424), .A2(new_n425), .A3(new_n426), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n341), .A2(new_n255), .A3(new_n407), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n412), .A2(new_n415), .ZN(new_n435));
  NAND4_X1  g234(.A1(new_n434), .A2(new_n435), .A3(new_n406), .A4(new_n428), .ZN(new_n436));
  NAND4_X1  g235(.A1(new_n433), .A2(KEYINPUT82), .A3(new_n436), .A4(KEYINPUT5), .ZN(new_n437));
  AOI21_X1  g236(.A(new_n420), .B1(new_n432), .B2(new_n437), .ZN(new_n438));
  XNOR2_X1  g237(.A(KEYINPUT0), .B(G57gat), .ZN(new_n439));
  XNOR2_X1  g238(.A(new_n439), .B(G85gat), .ZN(new_n440));
  XNOR2_X1  g239(.A(G1gat), .B(G29gat), .ZN(new_n441));
  XOR2_X1   g240(.A(new_n440), .B(new_n441), .Z(new_n442));
  XOR2_X1   g241(.A(KEYINPUT84), .B(KEYINPUT6), .Z(new_n443));
  INV_X1    g242(.A(new_n443), .ZN(new_n444));
  NOR3_X1   g243(.A1(new_n438), .A2(new_n442), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(new_n445), .ZN(new_n446));
  AND2_X1   g245(.A1(new_n435), .A2(new_n428), .ZN(new_n447));
  AOI21_X1  g246(.A(new_n405), .B1(new_n447), .B2(new_n410), .ZN(new_n448));
  AOI21_X1  g247(.A(KEYINPUT82), .B1(new_n448), .B2(new_n433), .ZN(new_n449));
  INV_X1    g248(.A(new_n437), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n419), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n442), .ZN(new_n452));
  NAND2_X1  g251(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  NAND2_X1  g252(.A1(new_n438), .A2(new_n442), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n453), .A2(new_n444), .A3(new_n454), .ZN(new_n455));
  AOI21_X1  g254(.A(new_n404), .B1(new_n446), .B2(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n379), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(KEYINPUT35), .ZN(new_n458));
  INV_X1    g257(.A(new_n280), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n273), .A2(new_n276), .A3(new_n278), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g260(.A(new_n366), .ZN(new_n462));
  NAND3_X1  g261(.A1(new_n371), .A2(new_n370), .A3(new_n352), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n375), .A2(new_n376), .A3(new_n352), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(KEYINPUT74), .ZN(new_n465));
  AOI21_X1  g264(.A(new_n462), .B1(new_n463), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n461), .A2(new_n466), .ZN(new_n467));
  INV_X1    g266(.A(new_n467), .ZN(new_n468));
  AOI211_X1 g267(.A(new_n452), .B(new_n420), .C1(new_n432), .C2(new_n437), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n432), .A2(new_n437), .ZN(new_n470));
  AOI21_X1  g269(.A(new_n442), .B1(new_n470), .B2(new_n419), .ZN(new_n471));
  NOR3_X1   g270(.A1(new_n469), .A2(new_n471), .A3(new_n443), .ZN(new_n472));
  OAI21_X1  g271(.A(KEYINPUT89), .B1(new_n472), .B2(new_n445), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT89), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n455), .A2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n404), .B1(new_n473), .B2(new_n475), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n468), .B1(new_n476), .B2(KEYINPUT91), .ZN(new_n477));
  INV_X1    g276(.A(new_n404), .ZN(new_n478));
  AOI21_X1  g277(.A(new_n474), .B1(new_n455), .B2(new_n446), .ZN(new_n479));
  NOR2_X1   g278(.A1(new_n469), .A2(new_n471), .ZN(new_n480));
  AOI21_X1  g279(.A(KEYINPUT89), .B1(new_n480), .B2(new_n444), .ZN(new_n481));
  OAI211_X1 g280(.A(KEYINPUT91), .B(new_n478), .C1(new_n479), .C2(new_n481), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT35), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n482), .A2(new_n483), .ZN(new_n484));
  OAI21_X1  g283(.A(new_n458), .B1(new_n477), .B2(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(KEYINPUT90), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n397), .A2(new_n400), .ZN(new_n487));
  INV_X1    g286(.A(KEYINPUT37), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n389), .A2(new_n488), .ZN(new_n489));
  NAND2_X1  g288(.A1(new_n489), .A2(new_n394), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n389), .A2(new_n488), .ZN(new_n491));
  OAI21_X1  g290(.A(KEYINPUT38), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  OAI22_X1  g291(.A1(new_n383), .A2(new_n381), .B1(new_n380), .B2(new_n382), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(new_n253), .ZN(new_n494));
  OR2_X1    g293(.A1(new_n385), .A2(new_n387), .ZN(new_n495));
  OAI211_X1 g294(.A(KEYINPUT37), .B(new_n494), .C1(new_n495), .C2(new_n253), .ZN(new_n496));
  INV_X1    g295(.A(KEYINPUT38), .ZN(new_n497));
  NAND4_X1  g296(.A1(new_n489), .A2(new_n496), .A3(new_n497), .A4(new_n394), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n487), .A2(new_n492), .A3(new_n498), .ZN(new_n499));
  NOR3_X1   g298(.A1(new_n479), .A2(new_n481), .A3(new_n499), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT83), .B1(new_n429), .B2(new_n415), .ZN(new_n501));
  NAND3_X1  g300(.A1(new_n501), .A2(new_n416), .A3(new_n414), .ZN(new_n502));
  AOI21_X1  g301(.A(new_n406), .B1(new_n502), .B2(new_n434), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(KEYINPUT88), .ZN(new_n505));
  AND2_X1   g304(.A1(new_n424), .A2(new_n426), .ZN(new_n506));
  OAI211_X1 g305(.A(new_n505), .B(KEYINPUT39), .C1(new_n506), .C2(new_n425), .ZN(new_n507));
  AOI21_X1  g306(.A(new_n425), .B1(new_n424), .B2(new_n426), .ZN(new_n508));
  INV_X1    g307(.A(KEYINPUT39), .ZN(new_n509));
  OAI21_X1  g308(.A(KEYINPUT88), .B1(new_n508), .B2(new_n509), .ZN(new_n510));
  NAND3_X1  g309(.A1(new_n504), .A2(new_n507), .A3(new_n510), .ZN(new_n511));
  AOI21_X1  g310(.A(new_n452), .B1(new_n503), .B2(new_n509), .ZN(new_n512));
  AND3_X1   g311(.A1(new_n511), .A2(KEYINPUT40), .A3(new_n512), .ZN(new_n513));
  AOI21_X1  g312(.A(KEYINPUT40), .B1(new_n511), .B2(new_n512), .ZN(new_n514));
  NOR3_X1   g313(.A1(new_n513), .A2(new_n514), .A3(new_n471), .ZN(new_n515));
  NAND2_X1  g314(.A1(new_n515), .A2(new_n404), .ZN(new_n516));
  NAND2_X1  g315(.A1(new_n461), .A2(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n486), .B1(new_n500), .B2(new_n517), .ZN(new_n518));
  INV_X1    g317(.A(new_n466), .ZN(new_n519));
  XOR2_X1   g318(.A(KEYINPUT75), .B(KEYINPUT36), .Z(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n463), .A2(new_n465), .ZN(new_n522));
  NAND4_X1  g321(.A1(new_n522), .A2(KEYINPUT36), .A3(new_n367), .A4(new_n369), .ZN(new_n523));
  INV_X1    g322(.A(new_n456), .ZN(new_n524));
  AOI22_X1  g323(.A1(new_n521), .A2(new_n523), .B1(new_n524), .B2(new_n281), .ZN(new_n525));
  INV_X1    g324(.A(new_n499), .ZN(new_n526));
  AOI21_X1  g325(.A(new_n445), .B1(new_n480), .B2(new_n444), .ZN(new_n527));
  OAI211_X1 g326(.A(new_n475), .B(new_n526), .C1(new_n527), .C2(new_n474), .ZN(new_n528));
  AOI22_X1  g327(.A1(new_n460), .A2(new_n459), .B1(new_n515), .B2(new_n404), .ZN(new_n529));
  NAND3_X1  g328(.A1(new_n528), .A2(KEYINPUT90), .A3(new_n529), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n518), .A2(new_n525), .A3(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n485), .A2(new_n531), .ZN(new_n532));
  INV_X1    g331(.A(G29gat), .ZN(new_n533));
  INV_X1    g332(.A(G36gat), .ZN(new_n534));
  OAI21_X1  g333(.A(KEYINPUT92), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g334(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n536));
  INV_X1    g335(.A(KEYINPUT14), .ZN(new_n537));
  NAND3_X1  g336(.A1(new_n537), .A2(new_n533), .A3(new_n534), .ZN(new_n538));
  AOI21_X1  g337(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT15), .ZN(new_n540));
  XNOR2_X1  g339(.A(G43gat), .B(G50gat), .ZN(new_n541));
  INV_X1    g340(.A(new_n541), .ZN(new_n542));
  OR3_X1    g341(.A1(new_n539), .A2(new_n540), .A3(new_n542), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n542), .A2(new_n540), .ZN(new_n544));
  NAND2_X1  g343(.A1(new_n541), .A2(KEYINPUT15), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n544), .A2(new_n539), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n543), .A2(new_n546), .ZN(new_n547));
  INV_X1    g346(.A(KEYINPUT17), .ZN(new_n548));
  NAND2_X1  g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT93), .ZN(new_n550));
  XNOR2_X1  g349(.A(G15gat), .B(G22gat), .ZN(new_n551));
  INV_X1    g350(.A(G1gat), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n552), .A2(KEYINPUT16), .ZN(new_n553));
  NAND2_X1  g352(.A1(new_n551), .A2(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n554), .B1(G1gat), .B2(new_n551), .ZN(new_n555));
  INV_X1    g354(.A(G8gat), .ZN(new_n556));
  XNOR2_X1  g355(.A(new_n555), .B(new_n556), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n543), .A2(KEYINPUT17), .A3(new_n546), .ZN(new_n558));
  NAND4_X1  g357(.A1(new_n549), .A2(new_n550), .A3(new_n557), .A4(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n549), .A2(new_n558), .ZN(new_n560));
  INV_X1    g359(.A(new_n557), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  NAND2_X1  g361(.A1(new_n561), .A2(new_n547), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n563), .A2(KEYINPUT93), .ZN(new_n564));
  OAI21_X1  g363(.A(new_n559), .B1(new_n562), .B2(new_n564), .ZN(new_n565));
  NAND2_X1  g364(.A1(G229gat), .A2(G233gat), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  INV_X1    g366(.A(KEYINPUT18), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  XOR2_X1   g368(.A(new_n557), .B(new_n547), .Z(new_n570));
  INV_X1    g369(.A(new_n570), .ZN(new_n571));
  XNOR2_X1  g370(.A(new_n566), .B(KEYINPUT13), .ZN(new_n572));
  OR2_X1    g371(.A1(new_n571), .A2(new_n572), .ZN(new_n573));
  NAND3_X1  g372(.A1(new_n565), .A2(KEYINPUT18), .A3(new_n566), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n573), .A3(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n569), .A2(KEYINPUT94), .ZN(new_n576));
  XNOR2_X1  g375(.A(KEYINPUT11), .B(G169gat), .ZN(new_n577));
  XNOR2_X1  g376(.A(new_n577), .B(new_n231), .ZN(new_n578));
  XOR2_X1   g377(.A(G113gat), .B(G141gat), .Z(new_n579));
  XNOR2_X1  g378(.A(new_n578), .B(new_n579), .ZN(new_n580));
  XNOR2_X1  g379(.A(new_n580), .B(KEYINPUT12), .ZN(new_n581));
  NAND3_X1  g380(.A1(new_n575), .A2(new_n576), .A3(new_n581), .ZN(new_n582));
  AOI21_X1  g381(.A(KEYINPUT18), .B1(new_n565), .B2(new_n566), .ZN(new_n583));
  INV_X1    g382(.A(KEYINPUT94), .ZN(new_n584));
  OAI21_X1  g383(.A(new_n581), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND4_X1  g384(.A1(new_n585), .A2(new_n569), .A3(new_n573), .A4(new_n574), .ZN(new_n586));
  NAND2_X1  g385(.A1(new_n582), .A2(new_n586), .ZN(new_n587));
  AOI21_X1  g386(.A(KEYINPUT95), .B1(new_n532), .B2(new_n587), .ZN(new_n588));
  INV_X1    g387(.A(KEYINPUT95), .ZN(new_n589));
  AND2_X1   g388(.A1(new_n582), .A2(new_n586), .ZN(new_n590));
  AOI211_X1 g389(.A(new_n589), .B(new_n590), .C1(new_n485), .C2(new_n531), .ZN(new_n591));
  NOR2_X1   g390(.A1(new_n588), .A2(new_n591), .ZN(new_n592));
  XNOR2_X1  g391(.A(G127gat), .B(G155gat), .ZN(new_n593));
  INV_X1    g392(.A(G211gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT21), .ZN(new_n596));
  XNOR2_X1  g395(.A(KEYINPUT97), .B(G64gat), .ZN(new_n597));
  INV_X1    g396(.A(G57gat), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n597), .A2(new_n598), .ZN(new_n599));
  INV_X1    g398(.A(KEYINPUT9), .ZN(new_n600));
  INV_X1    g399(.A(G71gat), .ZN(new_n601));
  INV_X1    g400(.A(G78gat), .ZN(new_n602));
  OAI21_X1  g401(.A(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  OR2_X1    g402(.A1(KEYINPUT97), .A2(G64gat), .ZN(new_n604));
  NAND2_X1  g403(.A1(KEYINPUT97), .A2(G64gat), .ZN(new_n605));
  NAND3_X1  g404(.A1(new_n604), .A2(G57gat), .A3(new_n605), .ZN(new_n606));
  NAND3_X1  g405(.A1(new_n599), .A2(new_n603), .A3(new_n606), .ZN(new_n607));
  XNOR2_X1  g406(.A(G71gat), .B(G78gat), .ZN(new_n608));
  INV_X1    g407(.A(KEYINPUT96), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  OAI21_X1  g409(.A(KEYINPUT96), .B1(new_n601), .B2(new_n602), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n607), .A2(new_n610), .A3(new_n611), .ZN(new_n612));
  OR3_X1    g411(.A1(new_n598), .A2(new_n391), .A3(KEYINPUT98), .ZN(new_n613));
  OAI21_X1  g412(.A(new_n391), .B1(new_n598), .B2(KEYINPUT98), .ZN(new_n614));
  NAND4_X1  g413(.A1(new_n613), .A2(new_n608), .A3(new_n603), .A4(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n612), .A2(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n557), .B1(new_n596), .B2(new_n616), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(new_n299), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT99), .ZN(new_n619));
  OR2_X1    g418(.A1(new_n618), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g419(.A1(G231gat), .A2(G233gat), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n618), .A2(new_n619), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n620), .A2(new_n622), .A3(new_n623), .ZN(new_n624));
  INV_X1    g423(.A(new_n624), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n622), .B1(new_n620), .B2(new_n623), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n595), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  INV_X1    g426(.A(new_n626), .ZN(new_n628));
  INV_X1    g427(.A(new_n595), .ZN(new_n629));
  NAND3_X1  g428(.A1(new_n628), .A2(new_n624), .A3(new_n629), .ZN(new_n630));
  NAND2_X1  g429(.A1(new_n627), .A2(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n616), .A2(new_n596), .ZN(new_n632));
  XNOR2_X1  g431(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n633));
  XOR2_X1   g432(.A(new_n632), .B(new_n633), .Z(new_n634));
  INV_X1    g433(.A(new_n634), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n631), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g435(.A1(new_n627), .A2(new_n630), .A3(new_n634), .ZN(new_n637));
  NAND2_X1  g436(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND2_X1  g438(.A1(G99gat), .A2(G106gat), .ZN(new_n640));
  INV_X1    g439(.A(G85gat), .ZN(new_n641));
  AOI22_X1  g440(.A1(KEYINPUT8), .A2(new_n640), .B1(new_n641), .B2(new_n393), .ZN(new_n642));
  INV_X1    g441(.A(KEYINPUT7), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n643), .B1(new_n641), .B2(new_n393), .ZN(new_n644));
  NAND3_X1  g443(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n645));
  NAND3_X1  g444(.A1(new_n642), .A2(new_n644), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g445(.A(G99gat), .B(G106gat), .Z(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n646), .B(new_n648), .ZN(new_n649));
  AND2_X1   g448(.A1(G232gat), .A2(G233gat), .ZN(new_n650));
  AOI22_X1  g449(.A1(new_n547), .A2(new_n649), .B1(KEYINPUT41), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g450(.A(new_n651), .B1(new_n560), .B2(new_n649), .ZN(new_n652));
  XOR2_X1   g451(.A(G134gat), .B(G162gat), .Z(new_n653));
  XNOR2_X1  g452(.A(new_n652), .B(new_n653), .ZN(new_n654));
  NOR2_X1   g453(.A1(new_n650), .A2(KEYINPUT41), .ZN(new_n655));
  XNOR2_X1  g454(.A(G190gat), .B(G218gat), .ZN(new_n656));
  XNOR2_X1  g455(.A(new_n655), .B(new_n656), .ZN(new_n657));
  XOR2_X1   g456(.A(new_n654), .B(new_n657), .Z(new_n658));
  XNOR2_X1  g457(.A(G120gat), .B(G148gat), .ZN(new_n659));
  INV_X1    g458(.A(G176gat), .ZN(new_n660));
  XNOR2_X1  g459(.A(new_n659), .B(new_n660), .ZN(new_n661));
  XNOR2_X1  g460(.A(new_n661), .B(new_n232), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n649), .A2(KEYINPUT10), .A3(new_n612), .A4(new_n615), .ZN(new_n664));
  INV_X1    g463(.A(KEYINPUT102), .ZN(new_n665));
  XNOR2_X1  g464(.A(new_n664), .B(new_n665), .ZN(new_n666));
  INV_X1    g465(.A(KEYINPUT101), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n616), .A2(new_n649), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n646), .A2(KEYINPUT100), .ZN(new_n669));
  NAND2_X1  g468(.A1(new_n669), .A2(new_n647), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n646), .A2(new_n648), .A3(KEYINPUT100), .ZN(new_n671));
  NAND4_X1  g470(.A1(new_n612), .A2(new_n670), .A3(new_n615), .A4(new_n671), .ZN(new_n672));
  NAND2_X1  g471(.A1(new_n668), .A2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(KEYINPUT10), .ZN(new_n674));
  AOI21_X1  g473(.A(new_n667), .B1(new_n673), .B2(new_n674), .ZN(new_n675));
  AOI211_X1 g474(.A(KEYINPUT101), .B(KEYINPUT10), .C1(new_n668), .C2(new_n672), .ZN(new_n676));
  OAI21_X1  g475(.A(new_n666), .B1(new_n675), .B2(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(G230gat), .A2(G233gat), .ZN(new_n678));
  XOR2_X1   g477(.A(new_n678), .B(KEYINPUT103), .Z(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  NAND2_X1  g479(.A1(new_n677), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g480(.A1(new_n668), .A2(new_n679), .A3(new_n672), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n663), .B1(new_n681), .B2(new_n682), .ZN(new_n683));
  XNOR2_X1  g482(.A(new_n683), .B(KEYINPUT105), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n681), .A2(new_n682), .A3(new_n663), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT104), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n684), .A2(new_n686), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NAND4_X1  g487(.A1(new_n639), .A2(KEYINPUT106), .A3(new_n658), .A4(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(KEYINPUT106), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n636), .A2(new_n637), .A3(new_n658), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n690), .B1(new_n691), .B2(new_n687), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n689), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n592), .A2(new_n693), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n694), .A2(new_n527), .ZN(new_n695));
  XNOR2_X1  g494(.A(KEYINPUT107), .B(G1gat), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n695), .B(new_n696), .ZN(G1324gat));
  NOR3_X1   g496(.A1(new_n592), .A2(new_n478), .A3(new_n693), .ZN(new_n698));
  NAND2_X1  g497(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n699));
  OR2_X1    g498(.A1(KEYINPUT16), .A2(G8gat), .ZN(new_n700));
  NAND3_X1  g499(.A1(new_n698), .A2(new_n699), .A3(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT42), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n701), .A2(new_n702), .ZN(new_n703));
  OR2_X1    g502(.A1(new_n698), .A2(new_n556), .ZN(new_n704));
  NAND2_X1  g503(.A1(new_n701), .A2(new_n702), .ZN(new_n705));
  NAND3_X1  g504(.A1(new_n703), .A2(new_n704), .A3(new_n705), .ZN(G1325gat));
  AOI21_X1  g505(.A(G15gat), .B1(new_n694), .B2(new_n466), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n521), .A2(new_n523), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  AND2_X1   g508(.A1(new_n709), .A2(G15gat), .ZN(new_n710));
  AOI21_X1  g509(.A(new_n707), .B1(new_n694), .B2(new_n710), .ZN(G1326gat));
  NAND2_X1  g510(.A1(new_n694), .A2(new_n281), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  XNOR2_X1  g512(.A(new_n712), .B(new_n713), .ZN(G1327gat));
  INV_X1    g513(.A(new_n658), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n528), .A2(KEYINPUT90), .A3(new_n529), .ZN(new_n716));
  AOI21_X1  g515(.A(KEYINPUT90), .B1(new_n528), .B2(new_n529), .ZN(new_n717));
  NOR2_X1   g516(.A1(new_n372), .A2(new_n377), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n367), .A2(new_n369), .ZN(new_n719));
  INV_X1    g518(.A(KEYINPUT36), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n718), .A2(new_n719), .A3(new_n720), .ZN(new_n721));
  INV_X1    g520(.A(new_n520), .ZN(new_n722));
  NOR2_X1   g521(.A1(new_n466), .A2(new_n722), .ZN(new_n723));
  OAI22_X1  g522(.A1(new_n721), .A2(new_n723), .B1(new_n456), .B2(new_n461), .ZN(new_n724));
  NOR3_X1   g523(.A1(new_n716), .A2(new_n717), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n483), .B1(new_n379), .B2(new_n456), .ZN(new_n726));
  AND2_X1   g525(.A1(new_n482), .A2(new_n483), .ZN(new_n727));
  OAI21_X1  g526(.A(new_n478), .B1(new_n479), .B2(new_n481), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT91), .ZN(new_n729));
  AOI21_X1  g528(.A(new_n467), .B1(new_n728), .B2(new_n729), .ZN(new_n730));
  AOI21_X1  g529(.A(new_n726), .B1(new_n727), .B2(new_n730), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n715), .B1(new_n725), .B2(new_n731), .ZN(new_n732));
  INV_X1    g531(.A(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  NAND3_X1  g533(.A1(new_n532), .A2(KEYINPUT44), .A3(new_n715), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n638), .A2(new_n688), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n736), .A2(new_n590), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n734), .A2(new_n735), .A3(new_n737), .ZN(new_n738));
  NAND2_X1  g537(.A1(new_n455), .A2(new_n446), .ZN(new_n739));
  OAI21_X1  g538(.A(G29gat), .B1(new_n738), .B2(new_n739), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n587), .B1(new_n725), .B2(new_n731), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(new_n589), .ZN(new_n742));
  NAND3_X1  g541(.A1(new_n532), .A2(KEYINPUT95), .A3(new_n587), .ZN(new_n743));
  NAND2_X1  g542(.A1(new_n742), .A2(new_n743), .ZN(new_n744));
  NOR2_X1   g543(.A1(new_n736), .A2(new_n658), .ZN(new_n745));
  AND2_X1   g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  NAND3_X1  g545(.A1(new_n746), .A2(new_n533), .A3(new_n527), .ZN(new_n747));
  AND2_X1   g546(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n748));
  NOR2_X1   g547(.A1(new_n747), .A2(KEYINPUT45), .ZN(new_n749));
  OAI21_X1  g548(.A(new_n740), .B1(new_n748), .B2(new_n749), .ZN(G1328gat));
  NAND3_X1  g549(.A1(new_n746), .A2(new_n534), .A3(new_n404), .ZN(new_n751));
  XNOR2_X1  g550(.A(KEYINPUT108), .B(KEYINPUT46), .ZN(new_n752));
  OR2_X1    g551(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI21_X1  g552(.A(G36gat), .B1(new_n738), .B2(new_n478), .ZN(new_n754));
  NAND2_X1  g553(.A1(new_n751), .A2(new_n752), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(G1329gat));
  NAND4_X1  g555(.A1(new_n734), .A2(new_n709), .A3(new_n735), .A4(new_n737), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(G43gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n519), .A2(G43gat), .ZN(new_n759));
  OAI211_X1 g558(.A(new_n745), .B(new_n759), .C1(new_n588), .C2(new_n591), .ZN(new_n760));
  NAND3_X1  g559(.A1(new_n758), .A2(KEYINPUT47), .A3(new_n760), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(KEYINPUT111), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT111), .ZN(new_n763));
  NAND4_X1  g562(.A1(new_n758), .A2(new_n763), .A3(KEYINPUT47), .A4(new_n760), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n762), .A2(new_n764), .ZN(new_n765));
  NAND2_X1  g564(.A1(new_n760), .A2(KEYINPUT109), .ZN(new_n766));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n767));
  NAND4_X1  g566(.A1(new_n744), .A2(new_n767), .A3(new_n745), .A4(new_n759), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n766), .A2(new_n758), .A3(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT110), .ZN(new_n770));
  INV_X1    g569(.A(KEYINPUT47), .ZN(new_n771));
  AND3_X1   g570(.A1(new_n769), .A2(new_n770), .A3(new_n771), .ZN(new_n772));
  AOI21_X1  g571(.A(new_n770), .B1(new_n769), .B2(new_n771), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n765), .B1(new_n772), .B2(new_n773), .ZN(G1330gat));
  OAI21_X1  g573(.A(G50gat), .B1(new_n738), .B2(new_n461), .ZN(new_n775));
  NAND4_X1  g574(.A1(new_n744), .A2(new_n275), .A3(new_n281), .A4(new_n745), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT112), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT48), .ZN(new_n778));
  OAI211_X1 g577(.A(new_n777), .B(new_n778), .C1(KEYINPUT112), .C2(new_n775), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n775), .A2(new_n776), .A3(KEYINPUT48), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT113), .ZN(new_n781));
  AND2_X1   g580(.A1(new_n780), .A2(new_n781), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n780), .A2(new_n781), .ZN(new_n783));
  OAI21_X1  g582(.A(new_n779), .B1(new_n782), .B2(new_n783), .ZN(G1331gat));
  AOI21_X1  g583(.A(new_n691), .B1(new_n485), .B2(new_n531), .ZN(new_n785));
  NOR2_X1   g584(.A1(new_n688), .A2(new_n587), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n785), .A2(new_n786), .ZN(new_n787));
  NOR2_X1   g586(.A1(new_n787), .A2(new_n739), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n788), .B(new_n598), .ZN(G1332gat));
  NOR2_X1   g588(.A1(new_n787), .A2(new_n478), .ZN(new_n790));
  NOR2_X1   g589(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n791));
  AND2_X1   g590(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n792));
  OAI21_X1  g591(.A(new_n790), .B1(new_n791), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g592(.A(new_n793), .B1(new_n790), .B2(new_n791), .ZN(G1333gat));
  OR3_X1    g593(.A1(new_n787), .A2(KEYINPUT115), .A3(new_n519), .ZN(new_n795));
  OAI21_X1  g594(.A(KEYINPUT115), .B1(new_n787), .B2(new_n519), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n795), .A2(new_n601), .A3(new_n796), .ZN(new_n797));
  NAND4_X1  g596(.A1(new_n785), .A2(G71gat), .A3(new_n709), .A4(new_n786), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n798), .B(KEYINPUT114), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n797), .A2(new_n799), .ZN(new_n800));
  XNOR2_X1  g599(.A(new_n800), .B(KEYINPUT50), .ZN(G1334gat));
  NOR2_X1   g600(.A1(new_n787), .A2(new_n461), .ZN(new_n802));
  XNOR2_X1  g601(.A(new_n802), .B(new_n602), .ZN(G1335gat));
  NAND4_X1  g602(.A1(new_n734), .A2(new_n638), .A3(new_n735), .A4(new_n786), .ZN(new_n804));
  NOR3_X1   g603(.A1(new_n804), .A2(new_n641), .A3(new_n739), .ZN(new_n805));
  AOI211_X1 g604(.A(new_n587), .B(new_n658), .C1(new_n485), .C2(new_n531), .ZN(new_n806));
  AND3_X1   g605(.A1(new_n806), .A2(KEYINPUT51), .A3(new_n638), .ZN(new_n807));
  AOI21_X1  g606(.A(KEYINPUT51), .B1(new_n806), .B2(new_n638), .ZN(new_n808));
  OR2_X1    g607(.A1(new_n807), .A2(new_n808), .ZN(new_n809));
  NAND3_X1  g608(.A1(new_n809), .A2(new_n527), .A3(new_n687), .ZN(new_n810));
  AOI21_X1  g609(.A(new_n805), .B1(new_n810), .B2(new_n641), .ZN(G1336gat));
  INV_X1    g610(.A(KEYINPUT52), .ZN(new_n812));
  OAI21_X1  g611(.A(G92gat), .B1(new_n804), .B2(new_n478), .ZN(new_n813));
  INV_X1    g612(.A(KEYINPUT117), .ZN(new_n814));
  AOI21_X1  g613(.A(new_n812), .B1(new_n813), .B2(new_n814), .ZN(new_n815));
  NAND3_X1  g614(.A1(new_n687), .A2(new_n393), .A3(new_n404), .ZN(new_n816));
  XOR2_X1   g615(.A(new_n816), .B(KEYINPUT116), .Z(new_n817));
  OAI21_X1  g616(.A(new_n817), .B1(new_n807), .B2(new_n808), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n813), .A2(new_n818), .ZN(new_n819));
  XNOR2_X1  g618(.A(new_n815), .B(new_n819), .ZN(G1337gat));
  OR3_X1    g619(.A1(new_n804), .A2(KEYINPUT118), .A3(new_n708), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT118), .B1(new_n804), .B2(new_n708), .ZN(new_n822));
  NAND3_X1  g621(.A1(new_n821), .A2(G99gat), .A3(new_n822), .ZN(new_n823));
  NOR2_X1   g622(.A1(new_n519), .A2(G99gat), .ZN(new_n824));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n687), .A3(new_n824), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n823), .A2(new_n825), .ZN(G1338gat));
  NOR2_X1   g625(.A1(new_n461), .A2(G106gat), .ZN(new_n827));
  OAI211_X1 g626(.A(new_n687), .B(new_n827), .C1(new_n807), .C2(new_n808), .ZN(new_n828));
  OAI21_X1  g627(.A(G106gat), .B1(new_n804), .B2(new_n461), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  XNOR2_X1  g629(.A(new_n830), .B(KEYINPUT53), .ZN(G1339gat));
  NOR2_X1   g630(.A1(new_n575), .A2(new_n581), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n565), .A2(new_n566), .ZN(new_n833));
  AOI21_X1  g632(.A(new_n833), .B1(new_n571), .B2(new_n572), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n834), .A2(new_n580), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n832), .A2(new_n835), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n687), .A2(new_n836), .ZN(new_n837));
  OAI211_X1 g636(.A(new_n679), .B(new_n666), .C1(new_n675), .C2(new_n676), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n681), .A2(KEYINPUT54), .A3(new_n838), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n839), .A2(KEYINPUT119), .ZN(new_n840));
  INV_X1    g639(.A(KEYINPUT119), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n681), .A2(new_n841), .A3(KEYINPUT54), .A4(new_n838), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n840), .A2(new_n842), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n662), .B1(new_n681), .B2(KEYINPUT54), .ZN(new_n844));
  INV_X1    g643(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n843), .A2(new_n845), .ZN(new_n846));
  INV_X1    g645(.A(KEYINPUT55), .ZN(new_n847));
  OAI211_X1 g646(.A(new_n587), .B(new_n686), .C1(new_n846), .C2(new_n847), .ZN(new_n848));
  AOI21_X1  g647(.A(new_n844), .B1(new_n840), .B2(new_n842), .ZN(new_n849));
  NOR2_X1   g648(.A1(new_n849), .A2(KEYINPUT55), .ZN(new_n850));
  OAI21_X1  g649(.A(new_n837), .B1(new_n848), .B2(new_n850), .ZN(new_n851));
  NAND2_X1  g650(.A1(new_n851), .A2(new_n658), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n686), .B1(new_n846), .B2(new_n847), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n715), .ZN(new_n854));
  OR3_X1    g653(.A1(new_n853), .A2(new_n854), .A3(new_n850), .ZN(new_n855));
  AOI21_X1  g654(.A(new_n639), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  NOR3_X1   g655(.A1(new_n691), .A2(new_n587), .A3(new_n687), .ZN(new_n857));
  OR2_X1    g656(.A1(new_n856), .A2(new_n857), .ZN(new_n858));
  AND2_X1   g657(.A1(new_n858), .A2(new_n379), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n739), .A2(new_n404), .ZN(new_n860));
  AND2_X1   g659(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n861), .A2(new_n321), .A3(new_n587), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n858), .A2(new_n468), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n863), .A2(new_n860), .ZN(new_n864));
  OAI21_X1  g663(.A(G113gat), .B1(new_n864), .B2(new_n590), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n862), .A2(new_n865), .ZN(G1340gat));
  NAND3_X1  g665(.A1(new_n861), .A2(new_n323), .A3(new_n687), .ZN(new_n867));
  OAI21_X1  g666(.A(G120gat), .B1(new_n864), .B2(new_n688), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n867), .A2(new_n868), .ZN(G1341gat));
  AOI21_X1  g668(.A(G127gat), .B1(new_n861), .B2(new_n639), .ZN(new_n870));
  NOR3_X1   g669(.A1(new_n864), .A2(new_n326), .A3(new_n638), .ZN(new_n871));
  NOR2_X1   g670(.A1(new_n870), .A2(new_n871), .ZN(G1342gat));
  NAND3_X1  g671(.A1(new_n861), .A2(new_n328), .A3(new_n715), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  OAI21_X1  g673(.A(G134gat), .B1(new_n864), .B2(new_n658), .ZN(new_n875));
  NAND2_X1  g674(.A1(new_n874), .A2(new_n875), .ZN(G1343gat));
  INV_X1    g675(.A(new_n848), .ZN(new_n877));
  NOR2_X1   g676(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT121), .ZN(new_n879));
  AOI211_X1 g678(.A(new_n879), .B(new_n844), .C1(new_n840), .C2(new_n842), .ZN(new_n880));
  NOR3_X1   g679(.A1(new_n878), .A2(new_n880), .A3(KEYINPUT55), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n877), .B1(new_n881), .B2(KEYINPUT122), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n846), .A2(new_n879), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n849), .A2(KEYINPUT121), .ZN(new_n884));
  NAND3_X1  g683(.A1(new_n883), .A2(new_n847), .A3(new_n884), .ZN(new_n885));
  INV_X1    g684(.A(KEYINPUT122), .ZN(new_n886));
  NOR2_X1   g685(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  OAI21_X1  g686(.A(new_n837), .B1(new_n882), .B2(new_n887), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n888), .A2(new_n658), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n639), .B1(new_n889), .B2(new_n855), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n281), .B1(new_n890), .B2(new_n857), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n891), .A2(KEYINPUT57), .ZN(new_n892));
  OAI21_X1  g691(.A(new_n281), .B1(new_n856), .B2(new_n857), .ZN(new_n893));
  OR2_X1    g692(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n894));
  AND2_X1   g693(.A1(new_n708), .A2(new_n860), .ZN(new_n895));
  XNOR2_X1  g694(.A(new_n895), .B(KEYINPUT120), .ZN(new_n896));
  NAND4_X1  g695(.A1(new_n892), .A2(new_n894), .A3(new_n587), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n897), .A2(G141gat), .ZN(new_n898));
  AND3_X1   g697(.A1(new_n858), .A2(new_n281), .A3(new_n895), .ZN(new_n899));
  NAND3_X1  g698(.A1(new_n899), .A2(new_n203), .A3(new_n587), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n898), .A2(new_n900), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n901), .A2(KEYINPUT58), .ZN(new_n902));
  INV_X1    g701(.A(KEYINPUT58), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n898), .A2(new_n903), .A3(new_n900), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n902), .A2(new_n904), .ZN(G1344gat));
  INV_X1    g704(.A(KEYINPUT59), .ZN(new_n906));
  NAND3_X1  g705(.A1(new_n892), .A2(new_n896), .A3(new_n894), .ZN(new_n907));
  OAI211_X1 g706(.A(new_n906), .B(G148gat), .C1(new_n907), .C2(new_n688), .ZN(new_n908));
  NOR2_X1   g707(.A1(new_n461), .A2(KEYINPUT57), .ZN(new_n909));
  AND3_X1   g708(.A1(new_n689), .A2(new_n590), .A3(new_n692), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n909), .B1(new_n890), .B2(new_n910), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n893), .A2(KEYINPUT57), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AND2_X1   g712(.A1(new_n896), .A2(new_n687), .ZN(new_n914));
  AOI21_X1  g713(.A(new_n205), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g714(.A(new_n908), .B1(new_n906), .B2(new_n915), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n899), .A2(new_n205), .A3(new_n687), .ZN(new_n917));
  NAND2_X1  g716(.A1(new_n916), .A2(new_n917), .ZN(G1345gat));
  AOI21_X1  g717(.A(G155gat), .B1(new_n899), .B2(new_n639), .ZN(new_n919));
  NOR2_X1   g718(.A1(new_n907), .A2(new_n209), .ZN(new_n920));
  AOI21_X1  g719(.A(new_n919), .B1(new_n920), .B2(new_n639), .ZN(G1346gat));
  AOI21_X1  g720(.A(G162gat), .B1(new_n899), .B2(new_n715), .ZN(new_n922));
  NOR2_X1   g721(.A1(new_n907), .A2(new_n658), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(G162gat), .ZN(G1347gat));
  NOR2_X1   g723(.A1(new_n527), .A2(new_n478), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n859), .A2(new_n925), .ZN(new_n926));
  XOR2_X1   g725(.A(new_n926), .B(KEYINPUT123), .Z(new_n927));
  INV_X1    g726(.A(G169gat), .ZN(new_n928));
  NAND3_X1  g727(.A1(new_n927), .A2(new_n928), .A3(new_n587), .ZN(new_n929));
  XOR2_X1   g728(.A(new_n925), .B(KEYINPUT124), .Z(new_n930));
  NAND2_X1  g729(.A1(new_n863), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G169gat), .B1(new_n931), .B2(new_n590), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(G1348gat));
  INV_X1    g732(.A(new_n292), .ZN(new_n934));
  NOR3_X1   g733(.A1(new_n931), .A2(new_n934), .A3(new_n688), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n927), .A2(new_n687), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n935), .B1(new_n936), .B2(new_n660), .ZN(G1349gat));
  OAI21_X1  g736(.A(G183gat), .B1(new_n931), .B2(new_n638), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n859), .A2(new_n307), .A3(new_n925), .ZN(new_n939));
  OAI21_X1  g738(.A(new_n938), .B1(new_n638), .B2(new_n939), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g740(.A1(new_n927), .A2(new_n302), .A3(new_n715), .ZN(new_n942));
  OAI21_X1  g741(.A(G190gat), .B1(new_n931), .B2(new_n658), .ZN(new_n943));
  NOR2_X1   g742(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n944));
  AND2_X1   g743(.A1(new_n943), .A2(KEYINPUT61), .ZN(new_n945));
  OAI21_X1  g744(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(G1351gat));
  AND2_X1   g745(.A1(new_n930), .A2(new_n708), .ZN(new_n947));
  AOI21_X1  g746(.A(new_n848), .B1(new_n885), .B2(new_n886), .ZN(new_n948));
  NAND2_X1  g747(.A1(new_n881), .A2(KEYINPUT122), .ZN(new_n949));
  AOI22_X1  g748(.A1(new_n948), .A2(new_n949), .B1(new_n687), .B2(new_n836), .ZN(new_n950));
  OAI21_X1  g749(.A(new_n855), .B1(new_n950), .B2(new_n715), .ZN(new_n951));
  AOI21_X1  g750(.A(new_n910), .B1(new_n951), .B2(new_n638), .ZN(new_n952));
  INV_X1    g751(.A(new_n909), .ZN(new_n953));
  OAI211_X1 g752(.A(new_n912), .B(new_n947), .C1(new_n952), .C2(new_n953), .ZN(new_n954));
  OAI21_X1  g753(.A(G197gat), .B1(new_n954), .B2(new_n590), .ZN(new_n955));
  NOR2_X1   g754(.A1(new_n893), .A2(new_n709), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n925), .ZN(new_n957));
  INV_X1    g756(.A(new_n957), .ZN(new_n958));
  NAND3_X1  g757(.A1(new_n958), .A2(new_n231), .A3(new_n587), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n955), .A2(new_n959), .ZN(G1352gat));
  INV_X1    g759(.A(new_n954), .ZN(new_n961));
  NAND3_X1  g760(.A1(new_n961), .A2(KEYINPUT125), .A3(new_n687), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT125), .ZN(new_n963));
  OAI21_X1  g762(.A(new_n963), .B1(new_n954), .B2(new_n688), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n962), .A2(G204gat), .A3(new_n964), .ZN(new_n965));
  NOR2_X1   g764(.A1(new_n688), .A2(G204gat), .ZN(new_n966));
  INV_X1    g765(.A(new_n966), .ZN(new_n967));
  OAI21_X1  g766(.A(KEYINPUT62), .B1(new_n957), .B2(new_n967), .ZN(new_n968));
  OR3_X1    g767(.A1(new_n957), .A2(KEYINPUT62), .A3(new_n967), .ZN(new_n969));
  NAND3_X1  g768(.A1(new_n965), .A2(new_n968), .A3(new_n969), .ZN(G1353gat));
  NAND3_X1  g769(.A1(new_n958), .A2(new_n594), .A3(new_n639), .ZN(new_n971));
  OAI211_X1 g770(.A(KEYINPUT63), .B(G211gat), .C1(new_n954), .C2(new_n638), .ZN(new_n972));
  INV_X1    g771(.A(new_n972), .ZN(new_n973));
  NAND4_X1  g772(.A1(new_n911), .A2(new_n639), .A3(new_n912), .A4(new_n947), .ZN(new_n974));
  AOI21_X1  g773(.A(KEYINPUT63), .B1(new_n974), .B2(G211gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n971), .B1(new_n973), .B2(new_n975), .ZN(new_n976));
  INV_X1    g775(.A(KEYINPUT126), .ZN(new_n977));
  NAND2_X1  g776(.A1(new_n976), .A2(new_n977), .ZN(new_n978));
  OAI211_X1 g777(.A(KEYINPUT126), .B(new_n971), .C1(new_n973), .C2(new_n975), .ZN(new_n979));
  NAND2_X1  g778(.A1(new_n978), .A2(new_n979), .ZN(G1354gat));
  AOI21_X1  g779(.A(G218gat), .B1(new_n958), .B2(new_n715), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n715), .A2(G218gat), .ZN(new_n982));
  XOR2_X1   g781(.A(new_n982), .B(KEYINPUT127), .Z(new_n983));
  AOI21_X1  g782(.A(new_n981), .B1(new_n961), .B2(new_n983), .ZN(G1355gat));
endmodule


