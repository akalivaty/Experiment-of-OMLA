

module locked_locked_c1908 ( G101, G104, G107, G110, G113, G116, G119, G122, 
        G125, G128, G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, 
        G224, G227, G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, 
        G953, G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, 
        G36, G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G101, G104, G107, G110, G113, G116, G119, G122, G125, G128, G131, G134,
         G137, G140, G143, G146, G210, G214, G217, G221, G224, G227, G234,
         G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
         KEYINPUT63, KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59,
         KEYINPUT58, KEYINPUT57, KEYINPUT56, KEYINPUT55, KEYINPUT54,
         KEYINPUT53, KEYINPUT52, KEYINPUT51, KEYINPUT50, KEYINPUT49,
         KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, KEYINPUT44,
         KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39,
         KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34,
         KEYINPUT33, KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29,
         KEYINPUT28, KEYINPUT27, KEYINPUT26, KEYINPUT25, KEYINPUT24,
         KEYINPUT23, KEYINPUT22, KEYINPUT21, KEYINPUT20, KEYINPUT19,
         KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, KEYINPUT14,
         KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, KEYINPUT8,
         KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, KEYINPUT2,
         KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125,
         KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120,
         KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115,
         KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110,
         KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105,
         KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100,
         KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95,
         KEYINPUT94, KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90,
         KEYINPUT89, KEYINPUT88, KEYINPUT87, KEYINPUT86, KEYINPUT85,
         KEYINPUT84, KEYINPUT83, KEYINPUT82, KEYINPUT81, KEYINPUT80,
         KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, KEYINPUT75,
         KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70,
         KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65,
         KEYINPUT64;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
         G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire   n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738;

  NOR2_X1 U372 ( .A1(G902), .A2(n710), .ZN(n414) );
  NOR2_X1 U373 ( .A1(n737), .A2(n736), .ZN(n532) );
  XNOR2_X1 U374 ( .A(n455), .B(KEYINPUT4), .ZN(n492) );
  NOR2_X1 U375 ( .A1(n572), .A2(n668), .ZN(n573) );
  XNOR2_X1 U376 ( .A(n368), .B(KEYINPUT87), .ZN(n600) );
  XNOR2_X2 U377 ( .A(n505), .B(n504), .ZN(n574) );
  OR2_X2 U378 ( .A1(n539), .A2(n536), .ZN(n538) );
  XNOR2_X2 U379 ( .A(n444), .B(KEYINPUT0), .ZN(n539) );
  XNOR2_X2 U380 ( .A(KEYINPUT67), .B(G101), .ZN(n424) );
  INV_X4 U381 ( .A(G953), .ZN(n423) );
  AND2_X1 U382 ( .A1(n366), .A2(n600), .ZN(n365) );
  AND2_X1 U383 ( .A1(n392), .A2(n390), .ZN(n583) );
  INV_X1 U384 ( .A(KEYINPUT48), .ZN(n386) );
  NAND2_X1 U385 ( .A1(n397), .A2(n597), .ZN(n604) );
  NAND2_X1 U386 ( .A1(n603), .A2(n602), .ZN(n695) );
  NAND2_X1 U387 ( .A1(n385), .A2(n654), .ZN(n368) );
  XNOR2_X1 U388 ( .A(n387), .B(n386), .ZN(n385) );
  NOR2_X1 U389 ( .A1(n738), .A2(n735), .ZN(n590) );
  NOR2_X1 U390 ( .A1(n526), .A2(n523), .ZN(n524) );
  NOR2_X1 U391 ( .A1(n526), .A2(n525), .ZN(n528) );
  XNOR2_X1 U392 ( .A(n584), .B(KEYINPUT39), .ZN(n595) );
  XNOR2_X1 U393 ( .A(n538), .B(n537), .ZN(n648) );
  NOR2_X1 U394 ( .A1(n568), .A2(n569), .ZN(n392) );
  XNOR2_X1 U395 ( .A(n574), .B(KEYINPUT1), .ZN(n662) );
  XNOR2_X1 U396 ( .A(n399), .B(n351), .ZN(n542) );
  XNOR2_X1 U397 ( .A(n427), .B(n405), .ZN(n725) );
  AND2_X1 U398 ( .A1(n604), .A2(n695), .ZN(n350) );
  AND2_X2 U399 ( .A1(n604), .A2(n695), .ZN(n708) );
  XNOR2_X1 U400 ( .A(G119), .B(G128), .ZN(n406) );
  XNOR2_X1 U401 ( .A(n484), .B(G125), .ZN(n427) );
  INV_X2 U402 ( .A(G146), .ZN(n484) );
  XNOR2_X1 U403 ( .A(n510), .B(n509), .ZN(n663) );
  NOR2_X2 U404 ( .A1(n689), .A2(n539), .ZN(n516) );
  XNOR2_X2 U405 ( .A(n515), .B(n514), .ZN(n689) );
  INV_X1 U406 ( .A(KEYINPUT10), .ZN(n405) );
  NAND2_X1 U407 ( .A1(n626), .A2(n552), .ZN(n372) );
  NAND2_X1 U408 ( .A1(n374), .A2(n373), .ZN(n380) );
  NOR2_X1 U409 ( .A1(n656), .A2(KEYINPUT104), .ZN(n373) );
  INV_X1 U410 ( .A(n540), .ZN(n374) );
  AND2_X1 U411 ( .A1(n648), .A2(n383), .ZN(n377) );
  XNOR2_X1 U412 ( .A(n492), .B(n491), .ZN(n496) );
  NAND2_X1 U413 ( .A1(n541), .A2(n472), .ZN(n678) );
  INV_X1 U414 ( .A(KEYINPUT95), .ZN(n418) );
  XNOR2_X1 U415 ( .A(G140), .B(G137), .ZN(n495) );
  XNOR2_X1 U416 ( .A(n401), .B(KEYINPUT71), .ZN(n358) );
  XNOR2_X1 U417 ( .A(n370), .B(n369), .ZN(n384) );
  XNOR2_X1 U418 ( .A(KEYINPUT79), .B(G110), .ZN(n369) );
  XNOR2_X1 U419 ( .A(n406), .B(n371), .ZN(n370) );
  INV_X1 U420 ( .A(KEYINPUT24), .ZN(n371) );
  XNOR2_X1 U421 ( .A(n471), .B(n400), .ZN(n617) );
  XNOR2_X1 U422 ( .A(n470), .B(n353), .ZN(n400) );
  XNOR2_X1 U423 ( .A(n496), .B(n495), .ZN(n726) );
  NAND2_X1 U424 ( .A1(n583), .A2(n675), .ZN(n584) );
  XNOR2_X1 U425 ( .A(n436), .B(n435), .ZN(n577) );
  XNOR2_X1 U426 ( .A(KEYINPUT77), .B(KEYINPUT19), .ZN(n435) );
  AND2_X1 U427 ( .A1(n380), .A2(n382), .ZN(n379) );
  INV_X1 U428 ( .A(n680), .ZN(n382) );
  NOR2_X1 U429 ( .A1(G237), .A2(G953), .ZN(n463) );
  NAND2_X1 U430 ( .A1(G234), .A2(G237), .ZN(n437) );
  NOR2_X1 U431 ( .A1(n580), .A2(n640), .ZN(n361) );
  INV_X1 U432 ( .A(G902), .ZN(n503) );
  XNOR2_X1 U433 ( .A(KEYINPUT102), .B(KEYINPUT5), .ZN(n478) );
  XOR2_X1 U434 ( .A(G137), .B(G116), .Z(n479) );
  XNOR2_X1 U435 ( .A(KEYINPUT69), .B(KEYINPUT3), .ZN(n419) );
  XOR2_X1 U436 ( .A(G140), .B(G143), .Z(n462) );
  OR2_X1 U437 ( .A1(G237), .A2(G902), .ZN(n434) );
  XOR2_X1 U438 ( .A(G116), .B(G107), .Z(n448) );
  NAND2_X1 U439 ( .A1(n552), .A2(KEYINPUT86), .ZN(n363) );
  XNOR2_X1 U440 ( .A(n567), .B(n391), .ZN(n390) );
  INV_X1 U441 ( .A(KEYINPUT30), .ZN(n391) );
  OR2_X1 U442 ( .A1(n617), .A2(G902), .ZN(n399) );
  BUF_X1 U443 ( .A(n662), .Z(n359) );
  OR2_X1 U444 ( .A1(n539), .A2(n568), .ZN(n540) );
  XNOR2_X1 U445 ( .A(n384), .B(n725), .ZN(n407) );
  XNOR2_X1 U446 ( .A(n358), .B(n495), .ZN(n404) );
  XNOR2_X1 U447 ( .A(n726), .B(n502), .ZN(n701) );
  XNOR2_X1 U448 ( .A(G110), .B(G107), .ZN(n498) );
  XNOR2_X1 U449 ( .A(n715), .B(n432), .ZN(n626) );
  XNOR2_X1 U450 ( .A(n610), .B(n609), .ZN(n714) );
  NOR2_X1 U451 ( .A1(n577), .A2(n587), .ZN(n578) );
  NOR2_X1 U452 ( .A1(n540), .A2(n656), .ZN(n632) );
  XNOR2_X1 U453 ( .A(n394), .B(n393), .ZN(n697) );
  INV_X1 U454 ( .A(KEYINPUT123), .ZN(n393) );
  INV_X1 U455 ( .A(KEYINPUT86), .ZN(n398) );
  XOR2_X1 U456 ( .A(KEYINPUT13), .B(G475), .Z(n351) );
  XOR2_X1 U457 ( .A(n433), .B(KEYINPUT82), .Z(n352) );
  XOR2_X1 U458 ( .A(n462), .B(n461), .Z(n353) );
  XOR2_X1 U459 ( .A(KEYINPUT97), .B(n443), .Z(n354) );
  AND2_X1 U460 ( .A1(n653), .A2(n363), .ZN(n355) );
  AND2_X1 U461 ( .A1(n364), .A2(n355), .ZN(n356) );
  INV_X1 U462 ( .A(KEYINPUT104), .ZN(n383) );
  AND2_X1 U463 ( .A1(n596), .A2(n398), .ZN(n357) );
  NOR2_X1 U464 ( .A1(n508), .A2(n658), .ZN(n510) );
  XNOR2_X2 U465 ( .A(n414), .B(n413), .ZN(n508) );
  XNOR2_X1 U466 ( .A(n404), .B(n403), .ZN(n408) );
  XNOR2_X1 U467 ( .A(n475), .B(KEYINPUT22), .ZN(n522) );
  NAND2_X1 U468 ( .A1(n360), .A2(n354), .ZN(n444) );
  INV_X1 U469 ( .A(n577), .ZN(n360) );
  AND2_X1 U470 ( .A1(n361), .A2(n581), .ZN(n389) );
  XNOR2_X1 U471 ( .A(n362), .B(n489), .ZN(n605) );
  XNOR2_X1 U472 ( .A(n488), .B(n496), .ZN(n362) );
  XNOR2_X1 U473 ( .A(n481), .B(n480), .ZN(n483) );
  NOR2_X2 U474 ( .A1(n663), .A2(n662), .ZN(n512) );
  OR2_X1 U475 ( .A1(n663), .A2(n574), .ZN(n568) );
  AND2_X1 U476 ( .A1(n600), .A2(n653), .ZN(n728) );
  NAND2_X1 U477 ( .A1(n365), .A2(n356), .ZN(n397) );
  NAND2_X1 U478 ( .A1(n601), .A2(n357), .ZN(n364) );
  NAND2_X1 U479 ( .A1(n367), .A2(KEYINPUT86), .ZN(n366) );
  INV_X1 U480 ( .A(n601), .ZN(n367) );
  XNOR2_X2 U481 ( .A(n551), .B(KEYINPUT45), .ZN(n601) );
  INV_X1 U482 ( .A(n553), .ZN(n593) );
  XNOR2_X2 U483 ( .A(n372), .B(n352), .ZN(n553) );
  INV_X1 U484 ( .A(n424), .ZN(n485) );
  NAND2_X1 U485 ( .A1(n376), .A2(n375), .ZN(n381) );
  NOR2_X1 U486 ( .A1(n632), .A2(n383), .ZN(n375) );
  INV_X1 U487 ( .A(n648), .ZN(n376) );
  NOR2_X1 U488 ( .A1(n378), .A2(n377), .ZN(n545) );
  NAND2_X1 U489 ( .A1(n381), .A2(n379), .ZN(n378) );
  XNOR2_X2 U490 ( .A(n485), .B(n484), .ZN(n501) );
  NAND2_X1 U491 ( .A1(n389), .A2(n388), .ZN(n387) );
  XNOR2_X1 U492 ( .A(n590), .B(KEYINPUT46), .ZN(n388) );
  NAND2_X1 U493 ( .A1(n395), .A2(n696), .ZN(n394) );
  NAND2_X1 U494 ( .A1(n396), .A2(n695), .ZN(n395) );
  NAND2_X1 U495 ( .A1(n694), .A2(n693), .ZN(n396) );
  INV_X1 U496 ( .A(n535), .ZN(n529) );
  XNOR2_X1 U497 ( .A(n710), .B(n709), .ZN(n711) );
  XOR2_X2 U498 ( .A(G122), .B(G104), .Z(n469) );
  INV_X1 U499 ( .A(KEYINPUT101), .ZN(n486) );
  XNOR2_X1 U500 ( .A(n487), .B(n486), .ZN(n488) );
  INV_X1 U501 ( .A(KEYINPUT23), .ZN(n401) );
  INV_X1 U502 ( .A(KEYINPUT75), .ZN(n511) );
  XNOR2_X1 U503 ( .A(n712), .B(n711), .ZN(n713) );
  NAND2_X1 U504 ( .A1(G234), .A2(n423), .ZN(n402) );
  XOR2_X1 U505 ( .A(KEYINPUT8), .B(n402), .Z(n449) );
  NAND2_X1 U506 ( .A1(G221), .A2(n449), .ZN(n403) );
  XNOR2_X1 U507 ( .A(n408), .B(n407), .ZN(n710) );
  XOR2_X1 U508 ( .A(KEYINPUT25), .B(KEYINPUT78), .Z(n411) );
  XNOR2_X2 U509 ( .A(G902), .B(KEYINPUT15), .ZN(n552) );
  NAND2_X1 U510 ( .A1(n552), .A2(G234), .ZN(n409) );
  XNOR2_X1 U511 ( .A(n409), .B(KEYINPUT20), .ZN(n445) );
  NAND2_X1 U512 ( .A1(G217), .A2(n445), .ZN(n410) );
  XNOR2_X1 U513 ( .A(n411), .B(n410), .ZN(n412) );
  XNOR2_X1 U514 ( .A(KEYINPUT98), .B(n412), .ZN(n413) );
  XOR2_X1 U515 ( .A(G110), .B(KEYINPUT16), .Z(n415) );
  XNOR2_X1 U516 ( .A(n469), .B(n415), .ZN(n416) );
  XNOR2_X1 U517 ( .A(n416), .B(n448), .ZN(n422) );
  XNOR2_X1 U518 ( .A(G119), .B(KEYINPUT70), .ZN(n417) );
  XNOR2_X1 U519 ( .A(n417), .B(G113), .ZN(n421) );
  XNOR2_X1 U520 ( .A(n419), .B(n418), .ZN(n420) );
  XNOR2_X1 U521 ( .A(n421), .B(n420), .ZN(n482) );
  XNOR2_X1 U522 ( .A(n422), .B(n482), .ZN(n715) );
  XNOR2_X2 U523 ( .A(G143), .B(G128), .ZN(n455) );
  NAND2_X1 U524 ( .A1(G224), .A2(n423), .ZN(n425) );
  XNOR2_X1 U525 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U526 ( .A(n492), .B(n426), .ZN(n431) );
  XOR2_X1 U527 ( .A(KEYINPUT17), .B(KEYINPUT18), .Z(n429) );
  INV_X1 U528 ( .A(n427), .ZN(n428) );
  XOR2_X1 U529 ( .A(n429), .B(n428), .Z(n430) );
  XNOR2_X1 U530 ( .A(n431), .B(n430), .ZN(n432) );
  NAND2_X1 U531 ( .A1(G210), .A2(n434), .ZN(n433) );
  NAND2_X1 U532 ( .A1(G214), .A2(n434), .ZN(n674) );
  NAND2_X1 U533 ( .A1(n553), .A2(n674), .ZN(n436) );
  XOR2_X1 U534 ( .A(KEYINPUT73), .B(KEYINPUT14), .Z(n438) );
  XNOR2_X1 U535 ( .A(n438), .B(n437), .ZN(n439) );
  NAND2_X1 U536 ( .A1(G952), .A2(n439), .ZN(n688) );
  NOR2_X1 U537 ( .A1(G953), .A2(n688), .ZN(n558) );
  INV_X1 U538 ( .A(n558), .ZN(n442) );
  NOR2_X1 U539 ( .A1(G898), .A2(n423), .ZN(n717) );
  NAND2_X1 U540 ( .A1(n439), .A2(G902), .ZN(n440) );
  XOR2_X1 U541 ( .A(KEYINPUT96), .B(n440), .Z(n554) );
  NAND2_X1 U542 ( .A1(n717), .A2(n554), .ZN(n441) );
  NAND2_X1 U543 ( .A1(n442), .A2(n441), .ZN(n443) );
  XOR2_X1 U544 ( .A(KEYINPUT99), .B(KEYINPUT21), .Z(n447) );
  NAND2_X1 U545 ( .A1(G221), .A2(n445), .ZN(n446) );
  XNOR2_X1 U546 ( .A(n447), .B(n446), .ZN(n658) );
  XOR2_X1 U547 ( .A(n448), .B(KEYINPUT9), .Z(n451) );
  NAND2_X1 U548 ( .A1(G217), .A2(n449), .ZN(n450) );
  XNOR2_X1 U549 ( .A(n451), .B(n450), .ZN(n452) );
  XOR2_X1 U550 ( .A(n452), .B(G122), .Z(n459) );
  XOR2_X1 U551 ( .A(KEYINPUT109), .B(KEYINPUT108), .Z(n454) );
  XNOR2_X1 U552 ( .A(KEYINPUT110), .B(KEYINPUT7), .ZN(n453) );
  XNOR2_X1 U553 ( .A(n454), .B(n453), .ZN(n457) );
  XOR2_X1 U554 ( .A(n455), .B(G134), .Z(n456) );
  XNOR2_X1 U555 ( .A(n457), .B(n456), .ZN(n458) );
  XNOR2_X1 U556 ( .A(n459), .B(n458), .ZN(n705) );
  NOR2_X1 U557 ( .A1(G902), .A2(n705), .ZN(n460) );
  XNOR2_X1 U558 ( .A(G478), .B(n460), .ZN(n541) );
  XNOR2_X1 U559 ( .A(G113), .B(G131), .ZN(n461) );
  XNOR2_X1 U560 ( .A(n463), .B(KEYINPUT76), .ZN(n477) );
  NAND2_X1 U561 ( .A1(n477), .A2(G214), .ZN(n467) );
  XOR2_X1 U562 ( .A(KEYINPUT106), .B(KEYINPUT107), .Z(n465) );
  XNOR2_X1 U563 ( .A(KEYINPUT11), .B(KEYINPUT12), .ZN(n464) );
  XNOR2_X1 U564 ( .A(n465), .B(n464), .ZN(n466) );
  XNOR2_X1 U565 ( .A(n467), .B(n466), .ZN(n468) );
  XOR2_X1 U566 ( .A(n468), .B(KEYINPUT105), .Z(n471) );
  XNOR2_X1 U567 ( .A(n469), .B(n725), .ZN(n470) );
  INV_X1 U568 ( .A(n542), .ZN(n472) );
  NOR2_X1 U569 ( .A1(n658), .A2(n678), .ZN(n473) );
  XNOR2_X1 U570 ( .A(n473), .B(KEYINPUT111), .ZN(n474) );
  NOR2_X1 U571 ( .A1(n539), .A2(n474), .ZN(n475) );
  INV_X1 U572 ( .A(n522), .ZN(n476) );
  NOR2_X1 U573 ( .A1(n508), .A2(n476), .ZN(n507) );
  AND2_X1 U574 ( .A1(G210), .A2(n477), .ZN(n481) );
  XNOR2_X1 U575 ( .A(n479), .B(n478), .ZN(n480) );
  XNOR2_X1 U576 ( .A(n483), .B(n482), .ZN(n489) );
  XNOR2_X1 U577 ( .A(n501), .B(KEYINPUT100), .ZN(n487) );
  INV_X1 U578 ( .A(G131), .ZN(n490) );
  XNOR2_X1 U579 ( .A(n490), .B(G134), .ZN(n491) );
  NAND2_X1 U580 ( .A1(n605), .A2(n503), .ZN(n493) );
  XNOR2_X2 U581 ( .A(n493), .B(G472), .ZN(n566) );
  INV_X1 U582 ( .A(KEYINPUT6), .ZN(n494) );
  XNOR2_X1 U583 ( .A(n566), .B(n494), .ZN(n560) );
  NAND2_X1 U584 ( .A1(n423), .A2(G227), .ZN(n497) );
  XNOR2_X1 U585 ( .A(n497), .B(G104), .ZN(n499) );
  XNOR2_X1 U586 ( .A(n499), .B(n498), .ZN(n500) );
  XNOR2_X1 U587 ( .A(n501), .B(n500), .ZN(n502) );
  NAND2_X1 U588 ( .A1(n701), .A2(n503), .ZN(n505) );
  INV_X1 U589 ( .A(G469), .ZN(n504) );
  INV_X1 U590 ( .A(n359), .ZN(n564) );
  NOR2_X1 U591 ( .A1(n560), .A2(n564), .ZN(n506) );
  AND2_X1 U592 ( .A1(n507), .A2(n506), .ZN(n544) );
  XOR2_X1 U593 ( .A(G101), .B(n544), .Z(G3) );
  INV_X1 U594 ( .A(KEYINPUT68), .ZN(n509) );
  XNOR2_X2 U595 ( .A(n512), .B(n511), .ZN(n655) );
  NAND2_X1 U596 ( .A1(n655), .A2(n560), .ZN(n515) );
  INV_X1 U597 ( .A(KEYINPUT72), .ZN(n513) );
  XNOR2_X1 U598 ( .A(n513), .B(KEYINPUT33), .ZN(n514) );
  XNOR2_X1 U599 ( .A(n516), .B(KEYINPUT34), .ZN(n519) );
  INV_X1 U600 ( .A(n541), .ZN(n517) );
  NAND2_X1 U601 ( .A1(n542), .A2(n517), .ZN(n571) );
  INV_X1 U602 ( .A(n571), .ZN(n518) );
  NAND2_X1 U603 ( .A1(n519), .A2(n518), .ZN(n521) );
  XNOR2_X1 U604 ( .A(KEYINPUT80), .B(KEYINPUT35), .ZN(n520) );
  XNOR2_X2 U605 ( .A(n521), .B(n520), .ZN(n535) );
  XOR2_X1 U606 ( .A(n535), .B(G122), .Z(G24) );
  NAND2_X1 U607 ( .A1(n508), .A2(n522), .ZN(n526) );
  INV_X1 U608 ( .A(n566), .ZN(n668) );
  NAND2_X1 U609 ( .A1(n668), .A2(n359), .ZN(n523) );
  XNOR2_X1 U610 ( .A(n524), .B(KEYINPUT112), .ZN(n737) );
  OR2_X1 U611 ( .A1(n560), .A2(n359), .ZN(n525) );
  XNOR2_X1 U612 ( .A(KEYINPUT64), .B(KEYINPUT32), .ZN(n527) );
  XNOR2_X1 U613 ( .A(n528), .B(n527), .ZN(n736) );
  NAND2_X1 U614 ( .A1(n532), .A2(n529), .ZN(n531) );
  INV_X1 U615 ( .A(KEYINPUT44), .ZN(n530) );
  NAND2_X1 U616 ( .A1(n531), .A2(n530), .ZN(n534) );
  NAND2_X1 U617 ( .A1(n532), .A2(KEYINPUT44), .ZN(n533) );
  NAND2_X1 U618 ( .A1(n534), .A2(n533), .ZN(n550) );
  NAND2_X1 U619 ( .A1(n535), .A2(KEYINPUT44), .ZN(n547) );
  INV_X1 U620 ( .A(n668), .ZN(n656) );
  NAND2_X1 U621 ( .A1(n655), .A2(n656), .ZN(n536) );
  XOR2_X1 U622 ( .A(KEYINPUT31), .B(KEYINPUT103), .Z(n537) );
  NAND2_X1 U623 ( .A1(n541), .A2(n542), .ZN(n642) );
  INV_X1 U624 ( .A(n642), .ZN(n644) );
  OR2_X1 U625 ( .A1(n542), .A2(n541), .ZN(n543) );
  INV_X1 U626 ( .A(n543), .ZN(n647) );
  NOR2_X1 U627 ( .A1(n644), .A2(n647), .ZN(n680) );
  NOR2_X1 U628 ( .A1(n545), .A2(n544), .ZN(n546) );
  NAND2_X1 U629 ( .A1(n547), .A2(n546), .ZN(n548) );
  XNOR2_X1 U630 ( .A(n548), .B(KEYINPUT89), .ZN(n549) );
  NAND2_X1 U631 ( .A1(n550), .A2(n549), .ZN(n551) );
  INV_X1 U632 ( .A(n552), .ZN(n596) );
  NAND2_X1 U633 ( .A1(G953), .A2(n554), .ZN(n555) );
  NOR2_X1 U634 ( .A1(G900), .A2(n555), .ZN(n556) );
  XOR2_X1 U635 ( .A(KEYINPUT113), .B(n556), .Z(n557) );
  NOR2_X1 U636 ( .A1(n558), .A2(n557), .ZN(n569) );
  NOR2_X1 U637 ( .A1(n658), .A2(n569), .ZN(n559) );
  NAND2_X1 U638 ( .A1(n508), .A2(n559), .ZN(n572) );
  NAND2_X1 U639 ( .A1(n560), .A2(n674), .ZN(n561) );
  OR2_X1 U640 ( .A1(n642), .A2(n561), .ZN(n562) );
  NOR2_X1 U641 ( .A1(n572), .A2(n562), .ZN(n591) );
  AND2_X1 U642 ( .A1(n553), .A2(n591), .ZN(n563) );
  XNOR2_X1 U643 ( .A(n563), .B(KEYINPUT36), .ZN(n565) );
  NAND2_X1 U644 ( .A1(n565), .A2(n564), .ZN(n651) );
  XNOR2_X1 U645 ( .A(n651), .B(KEYINPUT88), .ZN(n581) );
  NAND2_X1 U646 ( .A1(n566), .A2(n674), .ZN(n567) );
  NAND2_X1 U647 ( .A1(n583), .A2(n553), .ZN(n570) );
  NOR2_X1 U648 ( .A1(n571), .A2(n570), .ZN(n640) );
  XNOR2_X1 U649 ( .A(KEYINPUT28), .B(n573), .ZN(n576) );
  INV_X1 U650 ( .A(n574), .ZN(n575) );
  NAND2_X1 U651 ( .A1(n576), .A2(n575), .ZN(n587) );
  XNOR2_X1 U652 ( .A(n578), .B(KEYINPUT81), .ZN(n641) );
  NOR2_X1 U653 ( .A1(n641), .A2(n680), .ZN(n579) );
  XOR2_X1 U654 ( .A(KEYINPUT47), .B(n579), .Z(n580) );
  XNOR2_X1 U655 ( .A(KEYINPUT74), .B(KEYINPUT38), .ZN(n582) );
  XOR2_X1 U656 ( .A(n582), .B(n553), .Z(n675) );
  AND2_X1 U657 ( .A1(n595), .A2(n644), .ZN(n585) );
  XNOR2_X1 U658 ( .A(n585), .B(KEYINPUT40), .ZN(n738) );
  NAND2_X1 U659 ( .A1(n675), .A2(n674), .ZN(n679) );
  NOR2_X1 U660 ( .A1(n679), .A2(n678), .ZN(n586) );
  XNOR2_X1 U661 ( .A(n586), .B(KEYINPUT41), .ZN(n690) );
  NOR2_X1 U662 ( .A1(n690), .A2(n587), .ZN(n589) );
  XNOR2_X1 U663 ( .A(KEYINPUT114), .B(KEYINPUT42), .ZN(n588) );
  XNOR2_X1 U664 ( .A(n589), .B(n588), .ZN(n735) );
  NAND2_X1 U665 ( .A1(n591), .A2(n359), .ZN(n592) );
  XNOR2_X1 U666 ( .A(n592), .B(KEYINPUT43), .ZN(n594) );
  NAND2_X1 U667 ( .A1(n594), .A2(n593), .ZN(n654) );
  NAND2_X1 U668 ( .A1(n595), .A2(n647), .ZN(n653) );
  NAND2_X1 U669 ( .A1(n596), .A2(KEYINPUT2), .ZN(n597) );
  NAND2_X1 U670 ( .A1(n653), .A2(KEYINPUT2), .ZN(n598) );
  XNOR2_X1 U671 ( .A(n598), .B(KEYINPUT83), .ZN(n599) );
  AND2_X1 U672 ( .A1(n600), .A2(n599), .ZN(n603) );
  BUF_X1 U673 ( .A(n601), .Z(n602) );
  NAND2_X1 U674 ( .A1(n708), .A2(G472), .ZN(n607) );
  XOR2_X1 U675 ( .A(KEYINPUT62), .B(n605), .Z(n606) );
  XNOR2_X1 U676 ( .A(n607), .B(n606), .ZN(n611) );
  INV_X1 U677 ( .A(G952), .ZN(n608) );
  NAND2_X1 U678 ( .A1(n608), .A2(G953), .ZN(n610) );
  INV_X1 U679 ( .A(KEYINPUT94), .ZN(n609) );
  NOR2_X2 U680 ( .A1(n611), .A2(n714), .ZN(n614) );
  XNOR2_X1 U681 ( .A(KEYINPUT93), .B(KEYINPUT63), .ZN(n612) );
  XNOR2_X1 U682 ( .A(n612), .B(KEYINPUT90), .ZN(n613) );
  XNOR2_X1 U683 ( .A(n614), .B(n613), .ZN(G57) );
  NAND2_X1 U684 ( .A1(n708), .A2(G475), .ZN(n619) );
  XNOR2_X1 U685 ( .A(KEYINPUT65), .B(KEYINPUT92), .ZN(n615) );
  XNOR2_X1 U686 ( .A(n615), .B(KEYINPUT59), .ZN(n616) );
  XNOR2_X1 U687 ( .A(n617), .B(n616), .ZN(n618) );
  XNOR2_X1 U688 ( .A(n619), .B(n618), .ZN(n620) );
  NOR2_X2 U689 ( .A1(n620), .A2(n714), .ZN(n622) );
  XNOR2_X1 U690 ( .A(KEYINPUT66), .B(KEYINPUT60), .ZN(n621) );
  XNOR2_X1 U691 ( .A(n622), .B(n621), .ZN(G60) );
  NAND2_X1 U692 ( .A1(n708), .A2(G210), .ZN(n628) );
  XOR2_X1 U693 ( .A(KEYINPUT91), .B(KEYINPUT54), .Z(n624) );
  XNOR2_X1 U694 ( .A(KEYINPUT55), .B(KEYINPUT84), .ZN(n623) );
  XNOR2_X1 U695 ( .A(n624), .B(n623), .ZN(n625) );
  XNOR2_X1 U696 ( .A(n626), .B(n625), .ZN(n627) );
  XNOR2_X1 U697 ( .A(n628), .B(n627), .ZN(n629) );
  NOR2_X2 U698 ( .A1(n629), .A2(n714), .ZN(n630) );
  XNOR2_X1 U699 ( .A(n630), .B(KEYINPUT56), .ZN(G51) );
  NAND2_X1 U700 ( .A1(n632), .A2(n644), .ZN(n631) );
  XNOR2_X1 U701 ( .A(n631), .B(G104), .ZN(G6) );
  XOR2_X1 U702 ( .A(KEYINPUT115), .B(KEYINPUT27), .Z(n634) );
  NAND2_X1 U703 ( .A1(n632), .A2(n647), .ZN(n633) );
  XNOR2_X1 U704 ( .A(n634), .B(n633), .ZN(n636) );
  XOR2_X1 U705 ( .A(G107), .B(KEYINPUT26), .Z(n635) );
  XNOR2_X1 U706 ( .A(n636), .B(n635), .ZN(G9) );
  NOR2_X1 U707 ( .A1(n543), .A2(n641), .ZN(n638) );
  XNOR2_X1 U708 ( .A(KEYINPUT116), .B(KEYINPUT29), .ZN(n637) );
  XNOR2_X1 U709 ( .A(n638), .B(n637), .ZN(n639) );
  XNOR2_X1 U710 ( .A(G128), .B(n639), .ZN(G30) );
  XOR2_X1 U711 ( .A(G143), .B(n640), .Z(G45) );
  NOR2_X1 U712 ( .A1(n642), .A2(n641), .ZN(n643) );
  XOR2_X1 U713 ( .A(G146), .B(n643), .Z(G48) );
  XOR2_X1 U714 ( .A(G113), .B(KEYINPUT117), .Z(n646) );
  NAND2_X1 U715 ( .A1(n648), .A2(n644), .ZN(n645) );
  XNOR2_X1 U716 ( .A(n646), .B(n645), .ZN(G15) );
  NAND2_X1 U717 ( .A1(n648), .A2(n647), .ZN(n649) );
  XNOR2_X1 U718 ( .A(n649), .B(G116), .ZN(G18) );
  XOR2_X1 U719 ( .A(KEYINPUT37), .B(KEYINPUT118), .Z(n650) );
  XNOR2_X1 U720 ( .A(n651), .B(n650), .ZN(n652) );
  XNOR2_X1 U721 ( .A(G125), .B(n652), .ZN(G27) );
  XNOR2_X1 U722 ( .A(G134), .B(n653), .ZN(G36) );
  XNOR2_X1 U723 ( .A(G140), .B(n654), .ZN(G42) );
  INV_X1 U724 ( .A(n655), .ZN(n657) );
  NAND2_X1 U725 ( .A1(n657), .A2(n656), .ZN(n671) );
  NAND2_X1 U726 ( .A1(n508), .A2(n658), .ZN(n661) );
  XNOR2_X1 U727 ( .A(KEYINPUT120), .B(KEYINPUT49), .ZN(n659) );
  XNOR2_X1 U728 ( .A(n659), .B(KEYINPUT119), .ZN(n660) );
  XNOR2_X1 U729 ( .A(n661), .B(n660), .ZN(n667) );
  NAND2_X1 U730 ( .A1(n663), .A2(n359), .ZN(n665) );
  XOR2_X1 U731 ( .A(KEYINPUT121), .B(KEYINPUT50), .Z(n664) );
  XNOR2_X1 U732 ( .A(n665), .B(n664), .ZN(n666) );
  NAND2_X1 U733 ( .A1(n667), .A2(n666), .ZN(n669) );
  NAND2_X1 U734 ( .A1(n669), .A2(n668), .ZN(n670) );
  NAND2_X1 U735 ( .A1(n671), .A2(n670), .ZN(n672) );
  XOR2_X1 U736 ( .A(KEYINPUT51), .B(n672), .Z(n673) );
  NOR2_X1 U737 ( .A1(n690), .A2(n673), .ZN(n685) );
  NOR2_X1 U738 ( .A1(n675), .A2(n674), .ZN(n676) );
  XNOR2_X1 U739 ( .A(n676), .B(KEYINPUT122), .ZN(n677) );
  NOR2_X1 U740 ( .A1(n678), .A2(n677), .ZN(n682) );
  NOR2_X1 U741 ( .A1(n680), .A2(n679), .ZN(n681) );
  NOR2_X1 U742 ( .A1(n682), .A2(n681), .ZN(n683) );
  NOR2_X1 U743 ( .A1(n689), .A2(n683), .ZN(n684) );
  NOR2_X1 U744 ( .A1(n685), .A2(n684), .ZN(n686) );
  XNOR2_X1 U745 ( .A(n686), .B(KEYINPUT52), .ZN(n687) );
  NOR2_X1 U746 ( .A1(n688), .A2(n687), .ZN(n692) );
  NOR2_X1 U747 ( .A1(n690), .A2(n689), .ZN(n691) );
  NOR2_X1 U748 ( .A1(n692), .A2(n691), .ZN(n696) );
  NAND2_X1 U749 ( .A1(n728), .A2(n602), .ZN(n694) );
  XNOR2_X1 U750 ( .A(KEYINPUT85), .B(KEYINPUT2), .ZN(n693) );
  NOR2_X1 U751 ( .A1(G953), .A2(n697), .ZN(n698) );
  XNOR2_X1 U752 ( .A(KEYINPUT53), .B(n698), .ZN(G75) );
  NAND2_X1 U753 ( .A1(n350), .A2(G469), .ZN(n703) );
  XOR2_X1 U754 ( .A(KEYINPUT57), .B(KEYINPUT58), .Z(n699) );
  XOR2_X1 U755 ( .A(n699), .B(KEYINPUT124), .Z(n700) );
  XNOR2_X1 U756 ( .A(n701), .B(n700), .ZN(n702) );
  XNOR2_X1 U757 ( .A(n703), .B(n702), .ZN(n704) );
  NOR2_X1 U758 ( .A1(n714), .A2(n704), .ZN(G54) );
  NAND2_X1 U759 ( .A1(n350), .A2(G478), .ZN(n706) );
  XNOR2_X1 U760 ( .A(n706), .B(n705), .ZN(n707) );
  NOR2_X1 U761 ( .A1(n714), .A2(n707), .ZN(G63) );
  NAND2_X1 U762 ( .A1(n350), .A2(G217), .ZN(n712) );
  INV_X1 U763 ( .A(KEYINPUT125), .ZN(n709) );
  NOR2_X1 U764 ( .A1(n714), .A2(n713), .ZN(G66) );
  XNOR2_X1 U765 ( .A(G101), .B(n715), .ZN(n716) );
  NOR2_X1 U766 ( .A1(n717), .A2(n716), .ZN(n724) );
  NAND2_X1 U767 ( .A1(n602), .A2(n423), .ZN(n718) );
  XNOR2_X1 U768 ( .A(n718), .B(KEYINPUT126), .ZN(n722) );
  NAND2_X1 U769 ( .A1(G953), .A2(G224), .ZN(n719) );
  XNOR2_X1 U770 ( .A(KEYINPUT61), .B(n719), .ZN(n720) );
  NAND2_X1 U771 ( .A1(n720), .A2(G898), .ZN(n721) );
  NAND2_X1 U772 ( .A1(n722), .A2(n721), .ZN(n723) );
  XNOR2_X1 U773 ( .A(n724), .B(n723), .ZN(G69) );
  XOR2_X1 U774 ( .A(n725), .B(KEYINPUT127), .Z(n727) );
  XNOR2_X1 U775 ( .A(n727), .B(n726), .ZN(n730) );
  XOR2_X1 U776 ( .A(n730), .B(n728), .Z(n729) );
  NAND2_X1 U777 ( .A1(n729), .A2(n423), .ZN(n734) );
  XNOR2_X1 U778 ( .A(G227), .B(n730), .ZN(n731) );
  NAND2_X1 U779 ( .A1(n731), .A2(G900), .ZN(n732) );
  NAND2_X1 U780 ( .A1(n732), .A2(G953), .ZN(n733) );
  NAND2_X1 U781 ( .A1(n734), .A2(n733), .ZN(G72) );
  XOR2_X1 U782 ( .A(G137), .B(n735), .Z(G39) );
  XOR2_X1 U783 ( .A(n736), .B(G119), .Z(G21) );
  XOR2_X1 U784 ( .A(G110), .B(n737), .Z(G12) );
  XOR2_X1 U785 ( .A(n738), .B(G131), .Z(G33) );
endmodule

