//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 0 0 0 0 1 1 0 0 0 1 1 0 0 0 0 0 1 1 1 1 0 0 1 1 0 0 0 1 1 0 1 1 0 0 0 1 0 1 0 1 1 0 1 1 1 1 0 1 1 0 1 0 0 1 1 0 1 0 1 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:30:02 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n448, new_n450, new_n452, new_n453,
    new_n456, new_n457, new_n458, new_n461, new_n462, new_n463, new_n464,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n522, new_n523, new_n524, new_n525, new_n526,
    new_n527, new_n528, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n552, new_n553, new_n554, new_n555, new_n556,
    new_n557, new_n558, new_n559, new_n560, new_n561, new_n564, new_n565,
    new_n567, new_n568, new_n569, new_n570, new_n571, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n581, new_n582, new_n583, new_n584, new_n585, new_n586, new_n587,
    new_n588, new_n589, new_n590, new_n591, new_n593, new_n594, new_n595,
    new_n597, new_n598, new_n599, new_n600, new_n601, new_n602, new_n604,
    new_n605, new_n606, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n615, new_n616, new_n617, new_n618, new_n619, new_n620,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n649, new_n651, new_n652, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n672, new_n673, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n912, new_n913, new_n914, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n920, new_n921, new_n922, new_n923,
    new_n924, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n957, new_n958, new_n959, new_n960,
    new_n961, new_n962, new_n963, new_n964, new_n965, new_n966, new_n967,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1193;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  XNOR2_X1  g008(.A(KEYINPUT64), .B(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  XNOR2_X1  g011(.A(KEYINPUT65), .B(G96), .ZN(G221));
  XNOR2_X1  g012(.A(KEYINPUT66), .B(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  NAND2_X1  g022(.A1(G94), .A2(G452), .ZN(new_n448));
  XNOR2_X1  g023(.A(new_n448), .B(KEYINPUT67), .ZN(G173));
  NAND2_X1  g024(.A1(G7), .A2(G661), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT1), .Z(G223));
  INV_X1    g026(.A(G567), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n450), .A2(new_n452), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT68), .ZN(G234));
  NAND3_X1  g029(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  OR4_X1    g030(.A1(G219), .A2(G218), .A3(G220), .A4(G221), .ZN(new_n456));
  XOR2_X1   g031(.A(new_n456), .B(KEYINPUT2), .Z(new_n457));
  NOR4_X1   g032(.A1(G235), .A2(G237), .A3(G238), .A4(G236), .ZN(new_n458));
  NAND2_X1  g033(.A1(new_n457), .A2(new_n458), .ZN(G261));
  INV_X1    g034(.A(G261), .ZN(G325));
  INV_X1    g035(.A(new_n457), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G2106), .ZN(new_n462));
  OR2_X1    g037(.A1(new_n458), .A2(new_n452), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(new_n464), .ZN(G319));
  AND2_X1   g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NOR2_X1   g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  OR2_X1    g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  AND2_X1   g043(.A1(new_n468), .A2(G125), .ZN(new_n469));
  AND2_X1   g044(.A1(G113), .A2(G2104), .ZN(new_n470));
  OAI21_X1  g045(.A(G2105), .B1(new_n469), .B2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n466), .A2(new_n467), .ZN(new_n472));
  NOR2_X1   g047(.A1(new_n472), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(G2105), .ZN(new_n474));
  AND2_X1   g049(.A1(new_n474), .A2(G2104), .ZN(new_n475));
  AOI22_X1  g050(.A1(new_n473), .A2(G137), .B1(G101), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n471), .A2(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NAND2_X1  g053(.A1(new_n473), .A2(G136), .ZN(new_n479));
  NOR2_X1   g054(.A1(new_n472), .A2(new_n474), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n480), .A2(G124), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n474), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND2_X1  g060(.A1(new_n468), .A2(G2105), .ZN(new_n486));
  INV_X1    g061(.A(G126), .ZN(new_n487));
  NOR2_X1   g062(.A1(new_n474), .A2(G114), .ZN(new_n488));
  OAI21_X1  g063(.A(G2104), .B1(G102), .B2(G2105), .ZN(new_n489));
  OAI22_X1  g064(.A1(new_n486), .A2(new_n487), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n468), .A2(new_n474), .ZN(new_n491));
  INV_X1    g066(.A(G138), .ZN(new_n492));
  OAI21_X1  g067(.A(KEYINPUT4), .B1(new_n491), .B2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n473), .A2(new_n494), .A3(G138), .ZN(new_n495));
  AOI21_X1  g070(.A(new_n490), .B1(new_n493), .B2(new_n495), .ZN(G164));
  NAND2_X1  g071(.A1(G75), .A2(G543), .ZN(new_n497));
  AND2_X1   g072(.A1(KEYINPUT5), .A2(G543), .ZN(new_n498));
  NOR2_X1   g073(.A1(KEYINPUT5), .A2(G543), .ZN(new_n499));
  NOR2_X1   g074(.A1(new_n498), .A2(new_n499), .ZN(new_n500));
  INV_X1    g075(.A(G62), .ZN(new_n501));
  OAI21_X1  g076(.A(new_n497), .B1(new_n500), .B2(new_n501), .ZN(new_n502));
  NAND2_X1  g077(.A1(new_n502), .A2(G651), .ZN(new_n503));
  OR2_X1    g078(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  OR2_X1    g080(.A1(KEYINPUT6), .A2(G651), .ZN(new_n506));
  NAND2_X1  g081(.A1(KEYINPUT6), .A2(G651), .ZN(new_n507));
  AOI21_X1  g082(.A(new_n505), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n508), .A2(KEYINPUT69), .A3(G50), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT69), .ZN(new_n510));
  AND2_X1   g085(.A1(KEYINPUT6), .A2(G651), .ZN(new_n511));
  NOR2_X1   g086(.A1(KEYINPUT6), .A2(G651), .ZN(new_n512));
  OAI21_X1  g087(.A(G543), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  INV_X1    g088(.A(G50), .ZN(new_n514));
  OAI21_X1  g089(.A(new_n510), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  OAI22_X1  g090(.A1(new_n512), .A2(new_n511), .B1(new_n498), .B2(new_n499), .ZN(new_n516));
  INV_X1    g091(.A(new_n516), .ZN(new_n517));
  AOI22_X1  g092(.A1(new_n509), .A2(new_n515), .B1(new_n517), .B2(G88), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n503), .A2(KEYINPUT70), .ZN(new_n519));
  NAND3_X1  g094(.A1(new_n504), .A2(new_n518), .A3(new_n519), .ZN(G303));
  INV_X1    g095(.A(G303), .ZN(G166));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n522));
  NAND3_X1  g097(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n523));
  NAND2_X1  g098(.A1(new_n523), .A2(KEYINPUT7), .ZN(new_n524));
  INV_X1    g099(.A(KEYINPUT7), .ZN(new_n525));
  NAND4_X1  g100(.A1(new_n525), .A2(G76), .A3(G543), .A4(G651), .ZN(new_n526));
  NAND2_X1  g101(.A1(new_n524), .A2(new_n526), .ZN(new_n527));
  INV_X1    g102(.A(G89), .ZN(new_n528));
  OAI211_X1 g103(.A(new_n522), .B(new_n527), .C1(new_n516), .C2(new_n528), .ZN(new_n529));
  INV_X1    g104(.A(KEYINPUT5), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n530), .A2(new_n505), .ZN(new_n531));
  NAND2_X1  g106(.A1(KEYINPUT5), .A2(G543), .ZN(new_n532));
  NAND2_X1  g107(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  AND2_X1   g108(.A1(G63), .A2(G651), .ZN(new_n534));
  AOI22_X1  g109(.A1(new_n508), .A2(G51), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g110(.A1(new_n529), .A2(new_n535), .ZN(new_n536));
  XNOR2_X1  g111(.A(KEYINPUT6), .B(G651), .ZN(new_n537));
  NAND3_X1  g112(.A1(new_n533), .A2(new_n537), .A3(G89), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n522), .B1(new_n538), .B2(new_n527), .ZN(new_n539));
  NOR2_X1   g114(.A1(new_n536), .A2(new_n539), .ZN(G168));
  OAI21_X1  g115(.A(G64), .B1(new_n498), .B2(new_n499), .ZN(new_n541));
  NAND2_X1  g116(.A1(G77), .A2(G543), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g118(.A(KEYINPUT72), .B1(new_n543), .B2(G651), .ZN(new_n544));
  INV_X1    g119(.A(KEYINPUT72), .ZN(new_n545));
  INV_X1    g120(.A(G651), .ZN(new_n546));
  AOI211_X1 g121(.A(new_n545), .B(new_n546), .C1(new_n541), .C2(new_n542), .ZN(new_n547));
  INV_X1    g122(.A(G90), .ZN(new_n548));
  XNOR2_X1  g123(.A(KEYINPUT73), .B(G52), .ZN(new_n549));
  OAI22_X1  g124(.A1(new_n516), .A2(new_n548), .B1(new_n513), .B2(new_n549), .ZN(new_n550));
  NOR3_X1   g125(.A1(new_n544), .A2(new_n547), .A3(new_n550), .ZN(G171));
  NAND2_X1  g126(.A1(new_n533), .A2(G56), .ZN(new_n552));
  NAND2_X1  g127(.A1(G68), .A2(G543), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n552), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g129(.A1(new_n554), .A2(G651), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  INV_X1    g131(.A(KEYINPUT74), .ZN(new_n557));
  NAND3_X1  g132(.A1(new_n554), .A2(new_n557), .A3(G651), .ZN(new_n558));
  AOI22_X1  g133(.A1(new_n517), .A2(G81), .B1(G43), .B2(new_n508), .ZN(new_n559));
  NAND3_X1  g134(.A1(new_n556), .A2(new_n558), .A3(new_n559), .ZN(new_n560));
  INV_X1    g135(.A(new_n560), .ZN(new_n561));
  NAND2_X1  g136(.A1(new_n561), .A2(G860), .ZN(G153));
  NAND4_X1  g137(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g138(.A1(G1), .A2(G3), .ZN(new_n564));
  XNOR2_X1  g139(.A(new_n564), .B(KEYINPUT8), .ZN(new_n565));
  NAND4_X1  g140(.A1(G319), .A2(G483), .A3(G661), .A4(new_n565), .ZN(G188));
  NAND3_X1  g141(.A1(new_n537), .A2(G53), .A3(G543), .ZN(new_n567));
  INV_X1    g142(.A(KEYINPUT75), .ZN(new_n568));
  OAI21_X1  g143(.A(KEYINPUT9), .B1(new_n567), .B2(new_n568), .ZN(new_n569));
  NAND2_X1  g144(.A1(new_n567), .A2(new_n568), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  NAND3_X1  g146(.A1(new_n567), .A2(new_n568), .A3(KEYINPUT9), .ZN(new_n572));
  AOI22_X1  g147(.A1(new_n571), .A2(new_n572), .B1(G91), .B2(new_n517), .ZN(new_n573));
  AND2_X1   g148(.A1(G78), .A2(G543), .ZN(new_n574));
  OAI21_X1  g149(.A(KEYINPUT76), .B1(new_n498), .B2(new_n499), .ZN(new_n575));
  INV_X1    g150(.A(KEYINPUT76), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n531), .A2(new_n576), .A3(new_n532), .ZN(new_n577));
  NAND2_X1  g152(.A1(new_n575), .A2(new_n577), .ZN(new_n578));
  AOI21_X1  g153(.A(new_n574), .B1(new_n578), .B2(G65), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n546), .B1(new_n579), .B2(KEYINPUT77), .ZN(new_n580));
  INV_X1    g155(.A(KEYINPUT77), .ZN(new_n581));
  INV_X1    g156(.A(G65), .ZN(new_n582));
  AOI21_X1  g157(.A(new_n582), .B1(new_n575), .B2(new_n577), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n581), .B1(new_n583), .B2(new_n574), .ZN(new_n584));
  AOI21_X1  g159(.A(KEYINPUT78), .B1(new_n580), .B2(new_n584), .ZN(new_n585));
  NOR3_X1   g160(.A1(new_n498), .A2(new_n499), .A3(KEYINPUT76), .ZN(new_n586));
  AOI21_X1  g161(.A(new_n576), .B1(new_n531), .B2(new_n532), .ZN(new_n587));
  OAI21_X1  g162(.A(G65), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n574), .ZN(new_n589));
  NAND3_X1  g164(.A1(new_n588), .A2(KEYINPUT77), .A3(new_n589), .ZN(new_n590));
  AND4_X1   g165(.A1(KEYINPUT78), .A2(new_n590), .A3(new_n584), .A4(G651), .ZN(new_n591));
  OAI21_X1  g166(.A(new_n573), .B1(new_n585), .B2(new_n591), .ZN(G299));
  INV_X1    g167(.A(new_n544), .ZN(new_n593));
  INV_X1    g168(.A(new_n547), .ZN(new_n594));
  INV_X1    g169(.A(new_n550), .ZN(new_n595));
  NAND3_X1  g170(.A1(new_n593), .A2(new_n594), .A3(new_n595), .ZN(G301));
  OAI21_X1  g171(.A(KEYINPUT79), .B1(new_n536), .B2(new_n539), .ZN(new_n597));
  OAI21_X1  g172(.A(new_n527), .B1(new_n516), .B2(new_n528), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(KEYINPUT71), .ZN(new_n599));
  INV_X1    g174(.A(KEYINPUT79), .ZN(new_n600));
  NAND4_X1  g175(.A1(new_n599), .A2(new_n600), .A3(new_n529), .A4(new_n535), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n597), .A2(new_n601), .ZN(new_n602));
  INV_X1    g177(.A(new_n602), .ZN(G286));
  OR2_X1    g178(.A1(new_n533), .A2(G74), .ZN(new_n604));
  AOI22_X1  g179(.A1(new_n604), .A2(G651), .B1(new_n508), .B2(G49), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n517), .A2(G87), .ZN(new_n606));
  NAND2_X1  g181(.A1(new_n605), .A2(new_n606), .ZN(G288));
  AOI22_X1  g182(.A1(new_n533), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n608), .A2(new_n546), .ZN(new_n609));
  INV_X1    g184(.A(G86), .ZN(new_n610));
  INV_X1    g185(.A(G48), .ZN(new_n611));
  OAI22_X1  g186(.A1(new_n516), .A2(new_n610), .B1(new_n513), .B2(new_n611), .ZN(new_n612));
  NOR2_X1   g187(.A1(new_n609), .A2(new_n612), .ZN(new_n613));
  INV_X1    g188(.A(new_n613), .ZN(G305));
  AOI22_X1  g189(.A1(new_n533), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n615));
  NOR2_X1   g190(.A1(new_n615), .A2(new_n546), .ZN(new_n616));
  INV_X1    g191(.A(G85), .ZN(new_n617));
  INV_X1    g192(.A(G47), .ZN(new_n618));
  OAI22_X1  g193(.A1(new_n516), .A2(new_n617), .B1(new_n513), .B2(new_n618), .ZN(new_n619));
  NOR2_X1   g194(.A1(new_n616), .A2(new_n619), .ZN(new_n620));
  INV_X1    g195(.A(new_n620), .ZN(G290));
  NAND2_X1  g196(.A1(G301), .A2(G868), .ZN(new_n622));
  INV_X1    g197(.A(G92), .ZN(new_n623));
  NOR2_X1   g198(.A1(new_n516), .A2(new_n623), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(KEYINPUT10), .ZN(new_n625));
  AND2_X1   g200(.A1(new_n578), .A2(G66), .ZN(new_n626));
  AND2_X1   g201(.A1(G79), .A2(G543), .ZN(new_n627));
  OAI21_X1  g202(.A(G651), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  INV_X1    g203(.A(G54), .ZN(new_n629));
  INV_X1    g204(.A(KEYINPUT80), .ZN(new_n630));
  AOI21_X1  g205(.A(new_n629), .B1(new_n513), .B2(new_n630), .ZN(new_n631));
  OAI21_X1  g206(.A(new_n631), .B1(new_n630), .B2(new_n513), .ZN(new_n632));
  NAND3_X1  g207(.A1(new_n625), .A2(new_n628), .A3(new_n632), .ZN(new_n633));
  INV_X1    g208(.A(new_n633), .ZN(new_n634));
  OAI21_X1  g209(.A(new_n622), .B1(new_n634), .B2(G868), .ZN(G284));
  OAI21_X1  g210(.A(new_n622), .B1(new_n634), .B2(G868), .ZN(G321));
  INV_X1    g211(.A(G868), .ZN(new_n637));
  NOR2_X1   g212(.A1(G286), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n571), .A2(new_n572), .ZN(new_n639));
  NAND2_X1  g214(.A1(new_n517), .A2(G91), .ZN(new_n640));
  NAND2_X1  g215(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND3_X1  g216(.A1(new_n590), .A2(new_n584), .A3(G651), .ZN(new_n642));
  INV_X1    g217(.A(KEYINPUT78), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  NAND3_X1  g219(.A1(new_n580), .A2(KEYINPUT78), .A3(new_n584), .ZN(new_n645));
  AOI21_X1  g220(.A(new_n641), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  AOI21_X1  g221(.A(new_n638), .B1(new_n637), .B2(new_n646), .ZN(G297));
  AOI21_X1  g222(.A(new_n638), .B1(new_n637), .B2(new_n646), .ZN(G280));
  INV_X1    g223(.A(G559), .ZN(new_n649));
  OAI21_X1  g224(.A(new_n634), .B1(new_n649), .B2(G860), .ZN(G148));
  NAND2_X1  g225(.A1(new_n560), .A2(new_n637), .ZN(new_n651));
  NOR2_X1   g226(.A1(new_n633), .A2(G559), .ZN(new_n652));
  OAI21_X1  g227(.A(new_n651), .B1(new_n652), .B2(new_n637), .ZN(G323));
  XNOR2_X1  g228(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g229(.A1(new_n468), .A2(new_n475), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n655), .B(KEYINPUT12), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT13), .ZN(new_n657));
  INV_X1    g232(.A(G2100), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT82), .Z(new_n660));
  NOR2_X1   g235(.A1(new_n657), .A2(new_n658), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT81), .ZN(new_n662));
  NAND2_X1  g237(.A1(new_n480), .A2(G123), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n663), .B(KEYINPUT83), .ZN(new_n664));
  OAI21_X1  g239(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n665));
  INV_X1    g240(.A(G111), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n666), .B2(G2105), .ZN(new_n667));
  AOI21_X1  g242(.A(new_n667), .B1(new_n473), .B2(G135), .ZN(new_n668));
  AND2_X1   g243(.A1(new_n664), .A2(new_n668), .ZN(new_n669));
  XNOR2_X1  g244(.A(new_n669), .B(G2096), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n660), .A2(new_n662), .A3(new_n670), .ZN(G156));
  XNOR2_X1  g246(.A(G2427), .B(G2438), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2430), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT15), .B(G2435), .ZN(new_n674));
  OR2_X1    g249(.A1(new_n673), .A2(new_n674), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n673), .A2(new_n674), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n675), .A2(KEYINPUT14), .A3(new_n676), .ZN(new_n677));
  XNOR2_X1  g252(.A(G2451), .B(G2454), .ZN(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT16), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n677), .B(new_n679), .ZN(new_n680));
  XNOR2_X1  g255(.A(G2443), .B(G2446), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XNOR2_X1  g257(.A(G1341), .B(G1348), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  XOR2_X1   g259(.A(new_n684), .B(KEYINPUT84), .Z(new_n685));
  OAI21_X1  g260(.A(G14), .B1(new_n682), .B2(new_n683), .ZN(new_n686));
  NOR2_X1   g261(.A1(new_n685), .A2(new_n686), .ZN(G401));
  XNOR2_X1  g262(.A(G2067), .B(G2678), .ZN(new_n688));
  NOR2_X1   g263(.A1(G2072), .A2(G2078), .ZN(new_n689));
  NOR2_X1   g264(.A1(new_n444), .A2(new_n689), .ZN(new_n690));
  INV_X1    g265(.A(new_n690), .ZN(new_n691));
  AOI21_X1  g266(.A(new_n688), .B1(new_n691), .B2(KEYINPUT85), .ZN(new_n692));
  OAI21_X1  g267(.A(new_n692), .B1(KEYINPUT85), .B2(new_n691), .ZN(new_n693));
  XOR2_X1   g268(.A(G2084), .B(G2090), .Z(new_n694));
  INV_X1    g269(.A(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n690), .B(KEYINPUT17), .ZN(new_n696));
  INV_X1    g271(.A(new_n688), .ZN(new_n697));
  OAI211_X1 g272(.A(new_n693), .B(new_n695), .C1(new_n696), .C2(new_n697), .ZN(new_n698));
  NOR3_X1   g273(.A1(new_n695), .A2(new_n690), .A3(new_n697), .ZN(new_n699));
  XNOR2_X1  g274(.A(new_n699), .B(KEYINPUT18), .ZN(new_n700));
  NAND3_X1  g275(.A1(new_n696), .A2(new_n697), .A3(new_n694), .ZN(new_n701));
  NAND3_X1  g276(.A1(new_n698), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  XOR2_X1   g277(.A(G2096), .B(G2100), .Z(new_n703));
  XNOR2_X1  g278(.A(new_n702), .B(new_n703), .ZN(G227));
  XOR2_X1   g279(.A(KEYINPUT86), .B(KEYINPUT19), .Z(new_n705));
  XNOR2_X1  g280(.A(G1971), .B(G1976), .ZN(new_n706));
  XNOR2_X1  g281(.A(new_n705), .B(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(G1956), .B(G2474), .ZN(new_n708));
  XNOR2_X1  g283(.A(G1961), .B(G1966), .ZN(new_n709));
  NOR2_X1   g284(.A1(new_n708), .A2(new_n709), .ZN(new_n710));
  NAND2_X1  g285(.A1(new_n707), .A2(new_n710), .ZN(new_n711));
  XOR2_X1   g286(.A(new_n711), .B(KEYINPUT20), .Z(new_n712));
  AND2_X1   g287(.A1(new_n708), .A2(new_n709), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n707), .A2(new_n713), .ZN(new_n714));
  XNOR2_X1  g289(.A(new_n714), .B(KEYINPUT87), .ZN(new_n715));
  NOR3_X1   g290(.A1(new_n707), .A2(new_n710), .A3(new_n713), .ZN(new_n716));
  NOR3_X1   g291(.A1(new_n712), .A2(new_n715), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT88), .ZN(new_n719));
  XNOR2_X1  g294(.A(new_n717), .B(new_n719), .ZN(new_n720));
  XNOR2_X1  g295(.A(G1991), .B(G1996), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(G1981), .B(G1986), .ZN(new_n723));
  XNOR2_X1  g298(.A(new_n722), .B(new_n723), .ZN(new_n724));
  INV_X1    g299(.A(new_n724), .ZN(G229));
  INV_X1    g300(.A(G29), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G32), .ZN(new_n727));
  NAND3_X1  g302(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT26), .Z(new_n729));
  INV_X1    g304(.A(G129), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n729), .B1(new_n486), .B2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n475), .A2(G105), .ZN(new_n732));
  INV_X1    g307(.A(G141), .ZN(new_n733));
  OAI21_X1  g308(.A(new_n732), .B1(new_n491), .B2(new_n733), .ZN(new_n734));
  NOR2_X1   g309(.A1(new_n731), .A2(new_n734), .ZN(new_n735));
  OAI21_X1  g310(.A(new_n727), .B1(new_n735), .B2(new_n726), .ZN(new_n736));
  XNOR2_X1  g311(.A(KEYINPUT27), .B(G1996), .ZN(new_n737));
  INV_X1    g312(.A(new_n737), .ZN(new_n738));
  NOR2_X1   g313(.A1(new_n736), .A2(new_n738), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(KEYINPUT95), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G27), .ZN(new_n741));
  OAI21_X1  g316(.A(new_n741), .B1(G164), .B2(new_n726), .ZN(new_n742));
  XNOR2_X1  g317(.A(new_n742), .B(new_n443), .ZN(new_n743));
  AND2_X1   g318(.A1(new_n740), .A2(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n726), .A2(G35), .ZN(new_n745));
  OAI21_X1  g320(.A(new_n745), .B1(G162), .B2(new_n726), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT29), .Z(new_n747));
  INV_X1    g322(.A(G2090), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n747), .A2(new_n748), .ZN(new_n749));
  NAND2_X1  g324(.A1(new_n468), .A2(G127), .ZN(new_n750));
  NAND2_X1  g325(.A1(G115), .A2(G2104), .ZN(new_n751));
  AOI21_X1  g326(.A(new_n474), .B1(new_n750), .B2(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n473), .A2(G139), .ZN(new_n753));
  INV_X1    g328(.A(new_n753), .ZN(new_n754));
  NAND3_X1  g329(.A1(new_n474), .A2(G103), .A3(G2104), .ZN(new_n755));
  XNOR2_X1  g330(.A(new_n755), .B(KEYINPUT25), .ZN(new_n756));
  NOR3_X1   g331(.A1(new_n752), .A2(new_n754), .A3(new_n756), .ZN(new_n757));
  XNOR2_X1  g332(.A(new_n757), .B(KEYINPUT94), .ZN(new_n758));
  NOR2_X1   g333(.A1(new_n758), .A2(new_n726), .ZN(new_n759));
  AOI21_X1  g334(.A(new_n759), .B1(new_n726), .B2(G33), .ZN(new_n760));
  OAI211_X1 g335(.A(new_n744), .B(new_n749), .C1(new_n442), .C2(new_n760), .ZN(new_n761));
  NOR2_X1   g336(.A1(new_n747), .A2(new_n748), .ZN(new_n762));
  XOR2_X1   g337(.A(new_n762), .B(KEYINPUT99), .Z(new_n763));
  NOR2_X1   g338(.A1(G16), .A2(G19), .ZN(new_n764));
  AOI21_X1  g339(.A(new_n764), .B1(new_n561), .B2(G16), .ZN(new_n765));
  XOR2_X1   g340(.A(new_n765), .B(G1341), .Z(new_n766));
  INV_X1    g341(.A(G1961), .ZN(new_n767));
  INV_X1    g342(.A(G16), .ZN(new_n768));
  NOR2_X1   g343(.A1(G171), .A2(new_n768), .ZN(new_n769));
  AOI21_X1  g344(.A(new_n769), .B1(G5), .B2(new_n768), .ZN(new_n770));
  NAND2_X1  g345(.A1(new_n768), .A2(G21), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n771), .B1(G168), .B2(new_n768), .ZN(new_n772));
  XNOR2_X1  g347(.A(KEYINPUT96), .B(G1966), .ZN(new_n773));
  INV_X1    g348(.A(new_n773), .ZN(new_n774));
  OAI221_X1 g349(.A(new_n766), .B1(new_n767), .B2(new_n770), .C1(new_n772), .C2(new_n774), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n761), .A2(new_n763), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n770), .A2(new_n767), .ZN(new_n777));
  INV_X1    g352(.A(G2084), .ZN(new_n778));
  INV_X1    g353(.A(G34), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n779), .B2(KEYINPUT24), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT24), .B2(new_n779), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(new_n477), .B2(new_n726), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n778), .A2(new_n782), .B1(new_n736), .B2(new_n738), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n777), .A2(new_n783), .ZN(new_n784));
  XOR2_X1   g359(.A(new_n784), .B(KEYINPUT98), .Z(new_n785));
  NAND2_X1  g360(.A1(new_n669), .A2(G29), .ZN(new_n786));
  XOR2_X1   g361(.A(new_n786), .B(KEYINPUT97), .Z(new_n787));
  NAND2_X1  g362(.A1(new_n726), .A2(G26), .ZN(new_n788));
  XOR2_X1   g363(.A(new_n788), .B(KEYINPUT28), .Z(new_n789));
  OR2_X1    g364(.A1(G104), .A2(G2105), .ZN(new_n790));
  OAI211_X1 g365(.A(new_n790), .B(G2104), .C1(G116), .C2(new_n474), .ZN(new_n791));
  XOR2_X1   g366(.A(new_n791), .B(KEYINPUT93), .Z(new_n792));
  AOI22_X1  g367(.A1(G128), .A2(new_n480), .B1(new_n473), .B2(G140), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n792), .A2(new_n793), .ZN(new_n794));
  AOI21_X1  g369(.A(new_n789), .B1(new_n794), .B2(G29), .ZN(new_n795));
  INV_X1    g370(.A(G2067), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n795), .B(new_n796), .ZN(new_n797));
  XNOR2_X1  g372(.A(KEYINPUT30), .B(G28), .ZN(new_n798));
  OR2_X1    g373(.A1(KEYINPUT31), .A2(G11), .ZN(new_n799));
  NAND2_X1  g374(.A1(KEYINPUT31), .A2(G11), .ZN(new_n800));
  AOI22_X1  g375(.A1(new_n798), .A2(new_n726), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(new_n782), .B2(new_n778), .ZN(new_n802));
  NOR3_X1   g377(.A1(new_n787), .A2(new_n797), .A3(new_n802), .ZN(new_n803));
  NAND2_X1  g378(.A1(new_n768), .A2(G4), .ZN(new_n804));
  OAI21_X1  g379(.A(new_n804), .B1(new_n634), .B2(new_n768), .ZN(new_n805));
  INV_X1    g380(.A(G1348), .ZN(new_n806));
  XNOR2_X1  g381(.A(new_n805), .B(new_n806), .ZN(new_n807));
  AOI22_X1  g382(.A1(new_n760), .A2(new_n442), .B1(new_n772), .B2(new_n774), .ZN(new_n808));
  AND4_X1   g383(.A1(new_n785), .A2(new_n803), .A3(new_n807), .A4(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n768), .A2(G20), .ZN(new_n810));
  XNOR2_X1  g385(.A(new_n810), .B(KEYINPUT23), .ZN(new_n811));
  OAI21_X1  g386(.A(new_n811), .B1(new_n646), .B2(new_n768), .ZN(new_n812));
  INV_X1    g387(.A(G1956), .ZN(new_n813));
  XNOR2_X1  g388(.A(new_n812), .B(new_n813), .ZN(new_n814));
  NAND3_X1  g389(.A1(new_n776), .A2(new_n809), .A3(new_n814), .ZN(new_n815));
  XNOR2_X1  g390(.A(new_n815), .B(KEYINPUT100), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n768), .A2(G24), .ZN(new_n817));
  OAI21_X1  g392(.A(new_n817), .B1(new_n620), .B2(new_n768), .ZN(new_n818));
  INV_X1    g393(.A(G1986), .ZN(new_n819));
  XNOR2_X1  g394(.A(new_n818), .B(new_n819), .ZN(new_n820));
  NAND2_X1  g395(.A1(new_n473), .A2(G131), .ZN(new_n821));
  NAND2_X1  g396(.A1(new_n480), .A2(G119), .ZN(new_n822));
  NOR2_X1   g397(.A1(new_n474), .A2(G107), .ZN(new_n823));
  OAI21_X1  g398(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n824));
  OAI211_X1 g399(.A(new_n821), .B(new_n822), .C1(new_n823), .C2(new_n824), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(KEYINPUT89), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n826), .B(KEYINPUT90), .ZN(new_n827));
  MUX2_X1   g402(.A(G25), .B(new_n827), .S(G29), .Z(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT35), .B(G1991), .ZN(new_n829));
  XOR2_X1   g404(.A(new_n829), .B(KEYINPUT91), .Z(new_n830));
  OAI21_X1  g405(.A(new_n820), .B1(new_n828), .B2(new_n830), .ZN(new_n831));
  AOI21_X1  g406(.A(new_n831), .B1(new_n828), .B2(new_n830), .ZN(new_n832));
  NOR2_X1   g407(.A1(G6), .A2(G16), .ZN(new_n833));
  AOI21_X1  g408(.A(new_n833), .B1(new_n613), .B2(G16), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT32), .ZN(new_n835));
  INV_X1    g410(.A(G1981), .ZN(new_n836));
  XNOR2_X1  g411(.A(new_n835), .B(new_n836), .ZN(new_n837));
  NAND2_X1  g412(.A1(G166), .A2(G16), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(G16), .B2(G22), .ZN(new_n839));
  INV_X1    g414(.A(G1971), .ZN(new_n840));
  NAND2_X1  g415(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OR2_X1    g416(.A1(new_n839), .A2(new_n840), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n768), .A2(G23), .ZN(new_n843));
  INV_X1    g418(.A(G288), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n843), .B1(new_n844), .B2(new_n768), .ZN(new_n845));
  XNOR2_X1  g420(.A(KEYINPUT33), .B(G1976), .ZN(new_n846));
  XNOR2_X1  g421(.A(new_n845), .B(new_n846), .ZN(new_n847));
  NAND4_X1  g422(.A1(new_n837), .A2(new_n841), .A3(new_n842), .A4(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n849));
  NAND2_X1  g424(.A1(new_n848), .A2(KEYINPUT34), .ZN(new_n850));
  NAND3_X1  g425(.A1(new_n832), .A2(new_n849), .A3(new_n850), .ZN(new_n851));
  XOR2_X1   g426(.A(KEYINPUT92), .B(KEYINPUT36), .Z(new_n852));
  XNOR2_X1  g427(.A(new_n851), .B(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n816), .A2(new_n853), .ZN(G150));
  INV_X1    g429(.A(G150), .ZN(G311));
  NAND2_X1  g430(.A1(new_n533), .A2(G67), .ZN(new_n856));
  NAND2_X1  g431(.A1(G80), .A2(G543), .ZN(new_n857));
  AOI21_X1  g432(.A(new_n546), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g433(.A(G93), .ZN(new_n859));
  XNOR2_X1  g434(.A(KEYINPUT101), .B(G55), .ZN(new_n860));
  OAI22_X1  g435(.A1(new_n516), .A2(new_n859), .B1(new_n513), .B2(new_n860), .ZN(new_n861));
  NOR2_X1   g436(.A1(new_n858), .A2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(G860), .ZN(new_n863));
  NOR2_X1   g438(.A1(new_n862), .A2(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT37), .ZN(new_n865));
  NAND2_X1  g440(.A1(new_n634), .A2(G559), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT38), .ZN(new_n867));
  INV_X1    g442(.A(new_n862), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n560), .A2(new_n868), .ZN(new_n869));
  NAND4_X1  g444(.A1(new_n556), .A2(new_n862), .A3(new_n558), .A4(new_n559), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n869), .A2(new_n870), .ZN(new_n871));
  XNOR2_X1  g446(.A(new_n867), .B(new_n871), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT39), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT102), .Z(new_n875));
  OAI21_X1  g450(.A(new_n863), .B1(new_n873), .B2(KEYINPUT39), .ZN(new_n876));
  OAI21_X1  g451(.A(new_n865), .B1(new_n875), .B2(new_n876), .ZN(G145));
  NAND2_X1  g452(.A1(new_n493), .A2(new_n495), .ZN(new_n878));
  INV_X1    g453(.A(new_n490), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  XNOR2_X1  g455(.A(new_n880), .B(new_n794), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(new_n735), .ZN(new_n882));
  NOR2_X1   g457(.A1(new_n882), .A2(new_n757), .ZN(new_n883));
  AOI21_X1  g458(.A(new_n883), .B1(new_n758), .B2(new_n882), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n480), .A2(G130), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n474), .A2(G118), .ZN(new_n886));
  OAI21_X1  g461(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n887));
  OAI21_X1  g462(.A(new_n885), .B1(new_n886), .B2(new_n887), .ZN(new_n888));
  AOI21_X1  g463(.A(new_n888), .B1(G142), .B2(new_n473), .ZN(new_n889));
  XNOR2_X1  g464(.A(new_n889), .B(new_n656), .ZN(new_n890));
  XOR2_X1   g465(.A(new_n890), .B(new_n826), .Z(new_n891));
  INV_X1    g466(.A(new_n891), .ZN(new_n892));
  OR2_X1    g467(.A1(new_n884), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n884), .A2(new_n892), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  XNOR2_X1  g470(.A(new_n477), .B(new_n484), .ZN(new_n896));
  XOR2_X1   g471(.A(new_n896), .B(new_n669), .Z(new_n897));
  AOI21_X1  g472(.A(G37), .B1(new_n895), .B2(new_n897), .ZN(new_n898));
  OAI21_X1  g473(.A(new_n898), .B1(new_n897), .B2(new_n895), .ZN(new_n899));
  XNOR2_X1  g474(.A(new_n899), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g475(.A1(new_n868), .A2(new_n637), .ZN(new_n901));
  XNOR2_X1  g476(.A(new_n871), .B(new_n652), .ZN(new_n902));
  OAI211_X1 g477(.A(new_n573), .B(new_n633), .C1(new_n585), .C2(new_n591), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n903), .A2(KEYINPUT41), .ZN(new_n904));
  INV_X1    g479(.A(KEYINPUT103), .ZN(new_n905));
  OAI21_X1  g480(.A(new_n905), .B1(new_n646), .B2(new_n633), .ZN(new_n906));
  NAND3_X1  g481(.A1(G299), .A2(KEYINPUT103), .A3(new_n634), .ZN(new_n907));
  AOI21_X1  g482(.A(new_n904), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  NAND2_X1  g483(.A1(G299), .A2(new_n634), .ZN(new_n909));
  AOI21_X1  g484(.A(KEYINPUT41), .B1(new_n909), .B2(new_n903), .ZN(new_n910));
  OAI21_X1  g485(.A(new_n902), .B1(new_n908), .B2(new_n910), .ZN(new_n911));
  INV_X1    g486(.A(new_n903), .ZN(new_n912));
  AOI21_X1  g487(.A(new_n912), .B1(new_n906), .B2(new_n907), .ZN(new_n913));
  OAI21_X1  g488(.A(new_n911), .B1(new_n902), .B2(new_n913), .ZN(new_n914));
  XNOR2_X1  g489(.A(G303), .B(G290), .ZN(new_n915));
  XNOR2_X1  g490(.A(G288), .B(new_n613), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n915), .A2(new_n917), .ZN(new_n918));
  NOR2_X1   g493(.A1(G166), .A2(G290), .ZN(new_n919));
  NOR2_X1   g494(.A1(G303), .A2(new_n620), .ZN(new_n920));
  OAI21_X1  g495(.A(new_n916), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g496(.A1(new_n918), .A2(new_n921), .ZN(new_n922));
  XNOR2_X1  g497(.A(new_n922), .B(KEYINPUT42), .ZN(new_n923));
  XNOR2_X1  g498(.A(new_n914), .B(new_n923), .ZN(new_n924));
  OAI21_X1  g499(.A(new_n901), .B1(new_n924), .B2(new_n637), .ZN(G295));
  OAI21_X1  g500(.A(new_n901), .B1(new_n924), .B2(new_n637), .ZN(G331));
  INV_X1    g501(.A(KEYINPUT44), .ZN(new_n927));
  NAND3_X1  g502(.A1(new_n597), .A2(G171), .A3(new_n601), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n599), .A2(new_n529), .A3(new_n535), .ZN(new_n929));
  OAI21_X1  g504(.A(KEYINPUT105), .B1(G171), .B2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(KEYINPUT105), .ZN(new_n931));
  NAND3_X1  g506(.A1(G301), .A2(G168), .A3(new_n931), .ZN(new_n932));
  NAND3_X1  g507(.A1(new_n928), .A2(new_n930), .A3(new_n932), .ZN(new_n933));
  XNOR2_X1  g508(.A(new_n933), .B(new_n871), .ZN(new_n934));
  NOR3_X1   g509(.A1(new_n908), .A2(new_n934), .A3(new_n910), .ZN(new_n935));
  AND2_X1   g510(.A1(new_n913), .A2(new_n934), .ZN(new_n936));
  OAI21_X1  g511(.A(new_n922), .B1(new_n935), .B2(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(KEYINPUT41), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n933), .A2(new_n869), .A3(new_n870), .ZN(new_n939));
  NAND4_X1  g514(.A1(new_n871), .A2(new_n928), .A3(new_n932), .A4(new_n930), .ZN(new_n940));
  AOI21_X1  g515(.A(new_n938), .B1(new_n939), .B2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n909), .A2(new_n903), .ZN(new_n942));
  AOI21_X1  g517(.A(new_n922), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  OAI21_X1  g518(.A(new_n913), .B1(new_n934), .B2(new_n938), .ZN(new_n944));
  AOI21_X1  g519(.A(G37), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n937), .A2(new_n945), .ZN(new_n946));
  AOI21_X1  g521(.A(new_n927), .B1(new_n946), .B2(KEYINPUT43), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n938), .B1(new_n646), .B2(new_n633), .ZN(new_n948));
  NOR3_X1   g523(.A1(new_n646), .A2(new_n905), .A3(new_n633), .ZN(new_n949));
  AOI21_X1  g524(.A(KEYINPUT103), .B1(G299), .B2(new_n634), .ZN(new_n950));
  OAI21_X1  g525(.A(new_n948), .B1(new_n949), .B2(new_n950), .ZN(new_n951));
  NAND2_X1  g526(.A1(new_n942), .A2(new_n938), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n939), .A2(new_n940), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n952), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(new_n922), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n913), .A2(new_n934), .ZN(new_n956));
  NAND3_X1  g531(.A1(new_n954), .A2(new_n955), .A3(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT106), .ZN(new_n958));
  INV_X1    g533(.A(G37), .ZN(new_n959));
  NAND3_X1  g534(.A1(new_n957), .A2(new_n958), .A3(new_n959), .ZN(new_n960));
  NAND2_X1  g535(.A1(new_n960), .A2(new_n937), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n958), .B1(new_n957), .B2(new_n959), .ZN(new_n962));
  OR2_X1    g537(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  XOR2_X1   g538(.A(KEYINPUT104), .B(KEYINPUT43), .Z(new_n964));
  INV_X1    g539(.A(new_n964), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n947), .B1(new_n963), .B2(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT108), .ZN(new_n967));
  NAND3_X1  g542(.A1(new_n937), .A2(new_n964), .A3(new_n945), .ZN(new_n968));
  INV_X1    g543(.A(KEYINPUT107), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n968), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g545(.A1(new_n937), .A2(KEYINPUT107), .A3(new_n945), .A4(new_n964), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  OAI21_X1  g547(.A(new_n965), .B1(new_n961), .B2(new_n962), .ZN(new_n973));
  AOI211_X1 g548(.A(new_n967), .B(KEYINPUT44), .C1(new_n972), .C2(new_n973), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n973), .A2(new_n970), .A3(new_n971), .ZN(new_n975));
  AOI21_X1  g550(.A(KEYINPUT108), .B1(new_n975), .B2(new_n927), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n966), .B1(new_n974), .B2(new_n976), .ZN(G397));
  AOI21_X1  g552(.A(G1384), .B1(new_n878), .B2(new_n879), .ZN(new_n978));
  NOR2_X1   g553(.A1(new_n978), .A2(KEYINPUT45), .ZN(new_n979));
  AND3_X1   g554(.A1(new_n471), .A2(G40), .A3(new_n476), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n979), .A2(new_n980), .ZN(new_n981));
  XNOR2_X1  g556(.A(new_n794), .B(new_n796), .ZN(new_n982));
  OAI21_X1  g557(.A(G1996), .B1(new_n731), .B2(new_n734), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n981), .B1(new_n982), .B2(new_n983), .ZN(new_n984));
  NOR2_X1   g559(.A1(new_n981), .A2(G1996), .ZN(new_n985));
  XNOR2_X1  g560(.A(new_n985), .B(KEYINPUT109), .ZN(new_n986));
  AOI21_X1  g561(.A(new_n984), .B1(new_n986), .B2(new_n735), .ZN(new_n987));
  XOR2_X1   g562(.A(new_n826), .B(new_n829), .Z(new_n988));
  OAI21_X1  g563(.A(new_n987), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n620), .A2(new_n819), .ZN(new_n990));
  NAND2_X1  g565(.A1(G290), .A2(G1986), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n981), .B1(new_n990), .B2(new_n991), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n989), .A2(new_n992), .ZN(new_n993));
  INV_X1    g568(.A(G8), .ZN(new_n994));
  AOI21_X1  g569(.A(new_n994), .B1(new_n978), .B2(new_n980), .ZN(new_n995));
  NAND2_X1  g570(.A1(G305), .A2(G1981), .ZN(new_n996));
  NAND2_X1  g571(.A1(new_n613), .A2(new_n836), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(KEYINPUT114), .A3(new_n997), .ZN(new_n998));
  OR3_X1    g573(.A1(new_n613), .A2(KEYINPUT114), .A3(new_n836), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  INV_X1    g575(.A(KEYINPUT49), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n1001), .A2(KEYINPUT115), .ZN(new_n1002));
  NAND2_X1  g577(.A1(new_n1000), .A2(new_n1002), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n998), .A2(KEYINPUT115), .A3(new_n1001), .A4(new_n999), .ZN(new_n1004));
  NAND3_X1  g579(.A1(new_n1003), .A2(new_n1004), .A3(new_n995), .ZN(new_n1005));
  NOR2_X1   g580(.A1(G288), .A2(G1976), .ZN(new_n1006));
  AND2_X1   g581(.A1(new_n1005), .A2(new_n1006), .ZN(new_n1007));
  INV_X1    g582(.A(new_n997), .ZN(new_n1008));
  OAI21_X1  g583(.A(new_n995), .B1(new_n1007), .B2(new_n1008), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n844), .A2(G1976), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT52), .B1(new_n995), .B2(new_n1010), .ZN(new_n1011));
  AOI21_X1  g586(.A(KEYINPUT113), .B1(new_n844), .B2(G1976), .ZN(new_n1012));
  NAND2_X1  g587(.A1(new_n995), .A2(new_n1012), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1011), .A2(new_n1013), .ZN(new_n1014));
  OAI211_X1 g589(.A(new_n995), .B(new_n1012), .C1(KEYINPUT52), .C2(new_n1010), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1016), .A2(new_n1005), .ZN(new_n1017));
  NAND3_X1  g592(.A1(new_n471), .A2(G40), .A3(new_n476), .ZN(new_n1018));
  AOI21_X1  g593(.A(new_n1018), .B1(new_n978), .B2(KEYINPUT45), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT45), .ZN(new_n1020));
  OAI21_X1  g595(.A(new_n1020), .B1(G164), .B2(G1384), .ZN(new_n1021));
  NOR2_X1   g596(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1022));
  INV_X1    g597(.A(KEYINPUT110), .ZN(new_n1023));
  INV_X1    g598(.A(G1384), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n880), .A2(new_n1024), .ZN(new_n1025));
  AOI21_X1  g600(.A(new_n1023), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1026));
  OAI21_X1  g601(.A(new_n1019), .B1(new_n1022), .B2(new_n1026), .ZN(new_n1027));
  NAND2_X1  g602(.A1(new_n1027), .A2(new_n840), .ZN(new_n1028));
  XOR2_X1   g603(.A(KEYINPUT111), .B(KEYINPUT50), .Z(new_n1029));
  AOI21_X1  g604(.A(new_n1018), .B1(new_n978), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n1031));
  AND2_X1   g606(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1032));
  NAND2_X1  g607(.A1(new_n1032), .A2(new_n748), .ZN(new_n1033));
  AOI21_X1  g608(.A(new_n994), .B1(new_n1028), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(G303), .A2(G8), .ZN(new_n1035));
  XNOR2_X1  g610(.A(new_n1035), .B(KEYINPUT55), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT112), .ZN(new_n1037));
  XNOR2_X1  g612(.A(new_n1036), .B(new_n1037), .ZN(new_n1038));
  NAND2_X1  g613(.A1(new_n1034), .A2(new_n1038), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1009), .B1(new_n1017), .B2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT63), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1021), .A2(KEYINPUT110), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1025), .A2(new_n1023), .A3(new_n1020), .ZN(new_n1043));
  NAND2_X1  g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  AOI21_X1  g619(.A(G1971), .B1(new_n1044), .B2(new_n1019), .ZN(new_n1045));
  INV_X1    g620(.A(KEYINPUT50), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n978), .A2(new_n1046), .ZN(new_n1047));
  OAI211_X1 g622(.A(new_n1047), .B(new_n980), .C1(new_n978), .C2(new_n1029), .ZN(new_n1048));
  NOR2_X1   g623(.A1(new_n1048), .A2(G2090), .ZN(new_n1049));
  OAI21_X1  g624(.A(G8), .B1(new_n1045), .B2(new_n1049), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1050), .A2(new_n1036), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  NAND3_X1  g627(.A1(new_n1016), .A2(new_n1005), .A3(new_n1052), .ZN(new_n1053));
  INV_X1    g628(.A(new_n1053), .ZN(new_n1054));
  AOI21_X1  g629(.A(new_n1052), .B1(new_n1016), .B2(new_n1005), .ZN(new_n1055));
  OAI211_X1 g630(.A(new_n1039), .B(new_n1051), .C1(new_n1054), .C2(new_n1055), .ZN(new_n1056));
  OAI21_X1  g631(.A(new_n980), .B1(new_n1025), .B2(new_n1020), .ZN(new_n1057));
  OAI21_X1  g632(.A(new_n773), .B1(new_n1057), .B2(new_n979), .ZN(new_n1058));
  NAND3_X1  g633(.A1(new_n1030), .A2(new_n778), .A3(new_n1031), .ZN(new_n1059));
  AOI21_X1  g634(.A(new_n994), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(new_n602), .ZN(new_n1061));
  OAI21_X1  g636(.A(new_n1041), .B1(new_n1056), .B2(new_n1061), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1017), .A2(new_n1061), .A3(new_n1041), .ZN(new_n1063));
  INV_X1    g638(.A(new_n1036), .ZN(new_n1064));
  OAI211_X1 g639(.A(new_n1063), .B(new_n1039), .C1(new_n1034), .C2(new_n1064), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n1040), .B1(new_n1062), .B2(new_n1065), .ZN(new_n1066));
  AOI21_X1  g641(.A(G1348), .B1(new_n1030), .B2(new_n1031), .ZN(new_n1067));
  NAND2_X1  g642(.A1(new_n978), .A2(new_n980), .ZN(new_n1068));
  NOR2_X1   g643(.A1(new_n1068), .A2(G2067), .ZN(new_n1069));
  OAI21_X1  g644(.A(KEYINPUT118), .B1(new_n1067), .B2(new_n1069), .ZN(new_n1070));
  INV_X1    g645(.A(new_n1070), .ZN(new_n1071));
  NOR3_X1   g646(.A1(new_n1067), .A2(KEYINPUT118), .A3(new_n1069), .ZN(new_n1072));
  OAI21_X1  g647(.A(KEYINPUT60), .B1(new_n1071), .B2(new_n1072), .ZN(new_n1073));
  INV_X1    g648(.A(new_n1072), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT60), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1074), .A2(new_n1075), .A3(new_n1070), .ZN(new_n1076));
  NAND3_X1  g651(.A1(new_n1073), .A2(new_n1076), .A3(new_n634), .ZN(new_n1077));
  INV_X1    g652(.A(G1996), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1044), .A2(new_n1078), .A3(new_n1019), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  NAND2_X1  g655(.A1(new_n1068), .A2(new_n1080), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g657(.A(KEYINPUT59), .B1(new_n1082), .B2(new_n561), .ZN(new_n1083));
  INV_X1    g658(.A(KEYINPUT59), .ZN(new_n1084));
  AOI211_X1 g659(.A(new_n1084), .B(new_n560), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1085));
  NOR2_X1   g660(.A1(new_n1083), .A2(new_n1085), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1057), .B1(new_n1042), .B2(new_n1043), .ZN(new_n1087));
  XNOR2_X1  g662(.A(KEYINPUT56), .B(G2072), .ZN(new_n1088));
  AOI22_X1  g663(.A1(new_n1087), .A2(new_n1088), .B1(new_n813), .B2(new_n1048), .ZN(new_n1089));
  XNOR2_X1  g664(.A(new_n646), .B(KEYINPUT57), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1089), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(new_n1090), .ZN(new_n1092));
  NAND2_X1  g667(.A1(new_n1048), .A2(new_n813), .ZN(new_n1093));
  INV_X1    g668(.A(new_n1088), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1093), .B1(new_n1027), .B2(new_n1094), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1092), .A2(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1091), .A2(new_n1096), .A3(KEYINPUT61), .ZN(new_n1097));
  OAI211_X1 g672(.A(KEYINPUT60), .B(new_n633), .C1(new_n1071), .C2(new_n1072), .ZN(new_n1098));
  AND4_X1   g673(.A1(new_n1077), .A2(new_n1086), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  NOR2_X1   g674(.A1(new_n1091), .A2(KEYINPUT117), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT117), .ZN(new_n1101));
  AOI21_X1  g676(.A(new_n1101), .B1(new_n1089), .B2(new_n1090), .ZN(new_n1102));
  OAI21_X1  g677(.A(new_n1096), .B1(new_n1100), .B2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT61), .ZN(new_n1104));
  NAND2_X1  g679(.A1(new_n1103), .A2(new_n1104), .ZN(new_n1105));
  OR2_X1    g680(.A1(new_n1100), .A2(new_n1102), .ZN(new_n1106));
  NAND3_X1  g681(.A1(new_n1074), .A2(new_n634), .A3(new_n1070), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1107), .A2(new_n1096), .ZN(new_n1108));
  AOI22_X1  g683(.A1(new_n1099), .A2(new_n1105), .B1(new_n1106), .B2(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT54), .ZN(new_n1110));
  INV_X1    g685(.A(KEYINPUT121), .ZN(new_n1111));
  NAND3_X1  g686(.A1(new_n1044), .A2(new_n443), .A3(new_n1019), .ZN(new_n1112));
  INV_X1    g687(.A(KEYINPUT53), .ZN(new_n1113));
  NAND2_X1  g688(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  NOR2_X1   g689(.A1(new_n1057), .A2(new_n979), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(G2078), .ZN(new_n1116));
  NAND2_X1  g691(.A1(new_n1030), .A2(new_n1031), .ZN(new_n1117));
  AOI22_X1  g692(.A1(new_n1115), .A2(new_n1116), .B1(new_n1117), .B2(new_n767), .ZN(new_n1118));
  NAND2_X1  g693(.A1(new_n1114), .A2(new_n1118), .ZN(new_n1119));
  AOI21_X1  g694(.A(new_n1111), .B1(new_n1119), .B2(G171), .ZN(new_n1120));
  AOI211_X1 g695(.A(KEYINPUT121), .B(G301), .C1(new_n1114), .C2(new_n1118), .ZN(new_n1121));
  NOR2_X1   g696(.A1(new_n1120), .A2(new_n1121), .ZN(new_n1122));
  NAND3_X1  g697(.A1(new_n1019), .A2(new_n1021), .A3(new_n1116), .ZN(new_n1123));
  OAI21_X1  g698(.A(new_n1123), .B1(new_n1032), .B2(G1961), .ZN(new_n1124));
  AOI21_X1  g699(.A(new_n1124), .B1(new_n1113), .B2(new_n1112), .ZN(new_n1125));
  INV_X1    g700(.A(KEYINPUT122), .ZN(new_n1126));
  NAND3_X1  g701(.A1(new_n1125), .A2(new_n1126), .A3(G301), .ZN(new_n1127));
  NAND3_X1  g702(.A1(new_n1114), .A2(G301), .A3(new_n1118), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1128), .A2(KEYINPUT122), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1127), .A2(new_n1129), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1110), .B1(new_n1122), .B2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1119), .A2(G171), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1132), .A2(KEYINPUT54), .A3(new_n1128), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1017), .A2(KEYINPUT116), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1134), .A2(new_n1053), .ZN(new_n1135));
  AOI22_X1  g710(.A1(new_n1034), .A2(new_n1038), .B1(new_n1050), .B2(new_n1036), .ZN(new_n1136));
  AND3_X1   g711(.A1(new_n1133), .A2(new_n1135), .A3(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n929), .A2(G8), .ZN(new_n1138));
  XOR2_X1   g713(.A(new_n1138), .B(KEYINPUT119), .Z(new_n1139));
  AOI21_X1  g714(.A(new_n1139), .B1(new_n1058), .B2(new_n1059), .ZN(new_n1140));
  INV_X1    g715(.A(KEYINPUT120), .ZN(new_n1141));
  INV_X1    g716(.A(new_n1059), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n774), .B1(new_n1019), .B2(new_n1021), .ZN(new_n1143));
  OAI21_X1  g718(.A(G8), .B1(new_n1142), .B2(new_n1143), .ZN(new_n1144));
  AOI21_X1  g719(.A(new_n1141), .B1(new_n1144), .B2(new_n1139), .ZN(new_n1145));
  INV_X1    g720(.A(KEYINPUT51), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1140), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  INV_X1    g722(.A(new_n1139), .ZN(new_n1148));
  OAI21_X1  g723(.A(KEYINPUT120), .B1(new_n1060), .B2(new_n1148), .ZN(new_n1149));
  NAND3_X1  g724(.A1(new_n1144), .A2(new_n1141), .A3(new_n1139), .ZN(new_n1150));
  NAND3_X1  g725(.A1(new_n1149), .A2(new_n1150), .A3(KEYINPUT51), .ZN(new_n1151));
  NAND2_X1  g726(.A1(new_n1147), .A2(new_n1151), .ZN(new_n1152));
  NAND3_X1  g727(.A1(new_n1131), .A2(new_n1137), .A3(new_n1152), .ZN(new_n1153));
  OAI21_X1  g728(.A(new_n1066), .B1(new_n1109), .B2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT62), .ZN(new_n1155));
  AND3_X1   g730(.A1(new_n1147), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1156));
  OAI21_X1  g731(.A(KEYINPUT121), .B1(new_n1125), .B2(G301), .ZN(new_n1157));
  NAND3_X1  g732(.A1(new_n1119), .A2(new_n1111), .A3(G171), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1135), .A2(new_n1136), .A3(new_n1157), .A4(new_n1158), .ZN(new_n1159));
  OAI21_X1  g734(.A(KEYINPUT123), .B1(new_n1156), .B2(new_n1159), .ZN(new_n1160));
  INV_X1    g735(.A(new_n1056), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT123), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n1147), .A2(new_n1151), .A3(new_n1155), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1161), .A2(new_n1162), .A3(new_n1163), .A4(new_n1122), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1152), .A2(KEYINPUT62), .ZN(new_n1165));
  AND3_X1   g740(.A1(new_n1160), .A2(new_n1164), .A3(new_n1165), .ZN(new_n1166));
  OAI21_X1  g741(.A(new_n993), .B1(new_n1154), .B2(new_n1166), .ZN(new_n1167));
  OR2_X1    g742(.A1(new_n989), .A2(KEYINPUT125), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n989), .A2(KEYINPUT125), .ZN(new_n1169));
  NOR2_X1   g744(.A1(new_n981), .A2(new_n990), .ZN(new_n1170));
  XOR2_X1   g745(.A(KEYINPUT126), .B(KEYINPUT48), .Z(new_n1171));
  XNOR2_X1  g746(.A(new_n1171), .B(KEYINPUT127), .ZN(new_n1172));
  XNOR2_X1  g747(.A(new_n1170), .B(new_n1172), .ZN(new_n1173));
  NAND3_X1  g748(.A1(new_n1168), .A2(new_n1169), .A3(new_n1173), .ZN(new_n1174));
  INV_X1    g749(.A(KEYINPUT46), .ZN(new_n1175));
  XNOR2_X1  g750(.A(new_n986), .B(new_n1175), .ZN(new_n1176));
  AOI21_X1  g751(.A(new_n981), .B1(new_n982), .B2(new_n735), .ZN(new_n1177));
  INV_X1    g752(.A(new_n1177), .ZN(new_n1178));
  NAND2_X1  g753(.A1(new_n1176), .A2(new_n1178), .ZN(new_n1179));
  INV_X1    g754(.A(KEYINPUT124), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1179), .A2(new_n1180), .ZN(new_n1181));
  NAND3_X1  g756(.A1(new_n1176), .A2(KEYINPUT124), .A3(new_n1178), .ZN(new_n1182));
  NAND3_X1  g757(.A1(new_n1181), .A2(new_n1182), .A3(KEYINPUT47), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1174), .A2(new_n1183), .ZN(new_n1184));
  AOI21_X1  g759(.A(KEYINPUT47), .B1(new_n1181), .B2(new_n1182), .ZN(new_n1185));
  NOR2_X1   g760(.A1(new_n794), .A2(G2067), .ZN(new_n1186));
  NOR2_X1   g761(.A1(new_n827), .A2(new_n829), .ZN(new_n1187));
  AOI21_X1  g762(.A(new_n1186), .B1(new_n987), .B2(new_n1187), .ZN(new_n1188));
  NOR2_X1   g763(.A1(new_n1188), .A2(new_n981), .ZN(new_n1189));
  NOR3_X1   g764(.A1(new_n1184), .A2(new_n1185), .A3(new_n1189), .ZN(new_n1190));
  NAND2_X1  g765(.A1(new_n1167), .A2(new_n1190), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g766(.A1(G401), .A2(new_n464), .A3(G227), .ZN(new_n1193));
  NAND4_X1  g767(.A1(new_n899), .A2(new_n975), .A3(new_n724), .A4(new_n1193), .ZN(G225));
  INV_X1    g768(.A(G225), .ZN(G308));
endmodule


