//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 1 0 1 1 1 1 1 1 0 0 0 0 1 1 1 1 1 1 1 1 1 0 1 0 0 0 0 0 1 0 1 0 0 1 1 0 1 0 1 1 0 1 0 1 1 0 0 1 0 0 1 0 0 1 0 1 0 1 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:39 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n639, new_n640, new_n641, new_n642, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n671, new_n672, new_n673, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n731,
    new_n732, new_n733, new_n734, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n894, new_n895, new_n896, new_n897, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n904, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n915, new_n916, new_n917, new_n918, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n953, new_n954, new_n955, new_n956, new_n957, new_n958, new_n959,
    new_n960, new_n961, new_n962, new_n963;
  INV_X1    g000(.A(G237), .ZN(new_n187));
  NAND2_X1  g001(.A1(new_n187), .A2(KEYINPUT67), .ZN(new_n188));
  INV_X1    g002(.A(KEYINPUT67), .ZN(new_n189));
  NAND2_X1  g003(.A1(new_n189), .A2(G237), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n188), .A2(new_n190), .ZN(new_n191));
  INV_X1    g005(.A(G953), .ZN(new_n192));
  INV_X1    g006(.A(G214), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  AOI21_X1  g008(.A(new_n193), .B1(KEYINPUT86), .B2(new_n194), .ZN(new_n195));
  NAND3_X1  g009(.A1(new_n191), .A2(new_n192), .A3(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(new_n194), .A2(KEYINPUT86), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n196), .A2(new_n197), .ZN(new_n198));
  AOI21_X1  g012(.A(G953), .B1(new_n188), .B2(new_n190), .ZN(new_n199));
  INV_X1    g013(.A(new_n197), .ZN(new_n200));
  NAND3_X1  g014(.A1(new_n199), .A2(new_n195), .A3(new_n200), .ZN(new_n201));
  AOI21_X1  g015(.A(G131), .B1(new_n198), .B2(new_n201), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n198), .A2(G131), .A3(new_n201), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(KEYINPUT87), .ZN(new_n204));
  INV_X1    g018(.A(KEYINPUT87), .ZN(new_n205));
  NAND4_X1  g019(.A1(new_n198), .A2(new_n205), .A3(G131), .A4(new_n201), .ZN(new_n206));
  AOI21_X1  g020(.A(new_n202), .B1(new_n204), .B2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  XNOR2_X1  g022(.A(G125), .B(G140), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(KEYINPUT16), .ZN(new_n210));
  INV_X1    g024(.A(G125), .ZN(new_n211));
  OR3_X1    g025(.A1(new_n211), .A2(KEYINPUT16), .A3(G140), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n210), .A2(G146), .A3(new_n212), .ZN(new_n213));
  NAND2_X1  g027(.A1(new_n213), .A2(KEYINPUT75), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT75), .ZN(new_n215));
  NAND4_X1  g029(.A1(new_n210), .A2(new_n215), .A3(G146), .A4(new_n212), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n214), .A2(new_n216), .ZN(new_n217));
  INV_X1    g031(.A(new_n217), .ZN(new_n218));
  XOR2_X1   g032(.A(new_n209), .B(KEYINPUT19), .Z(new_n219));
  OAI211_X1 g033(.A(new_n208), .B(new_n218), .C1(G146), .C2(new_n219), .ZN(new_n220));
  XNOR2_X1  g034(.A(G113), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  INV_X1    g037(.A(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(KEYINPUT18), .ZN(new_n225));
  OR2_X1    g039(.A1(new_n203), .A2(new_n225), .ZN(new_n226));
  NAND2_X1  g040(.A1(new_n198), .A2(new_n201), .ZN(new_n227));
  INV_X1    g041(.A(G131), .ZN(new_n228));
  OAI21_X1  g042(.A(new_n227), .B1(new_n225), .B2(new_n228), .ZN(new_n229));
  INV_X1    g043(.A(G146), .ZN(new_n230));
  XNOR2_X1  g044(.A(new_n209), .B(new_n230), .ZN(new_n231));
  NAND3_X1  g045(.A1(new_n226), .A2(new_n229), .A3(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n220), .A2(new_n224), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(G475), .A2(G902), .ZN(new_n234));
  INV_X1    g048(.A(new_n232), .ZN(new_n235));
  INV_X1    g049(.A(KEYINPUT89), .ZN(new_n236));
  NAND2_X1  g050(.A1(new_n204), .A2(new_n206), .ZN(new_n237));
  INV_X1    g051(.A(KEYINPUT17), .ZN(new_n238));
  INV_X1    g052(.A(new_n202), .ZN(new_n239));
  AND4_X1   g053(.A1(new_n236), .A2(new_n237), .A3(new_n238), .A4(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(new_n236), .B1(new_n207), .B2(new_n238), .ZN(new_n241));
  NOR2_X1   g055(.A1(new_n240), .A2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n210), .A2(new_n212), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n243), .A2(new_n230), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(new_n213), .ZN(new_n245));
  INV_X1    g059(.A(KEYINPUT88), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n246), .B1(new_n237), .B2(new_n238), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n204), .A2(KEYINPUT88), .A3(KEYINPUT17), .A4(new_n206), .ZN(new_n248));
  AOI21_X1  g062(.A(new_n245), .B1(new_n247), .B2(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n235), .B1(new_n242), .B2(new_n249), .ZN(new_n250));
  OAI211_X1 g064(.A(new_n233), .B(new_n234), .C1(new_n250), .C2(new_n224), .ZN(new_n251));
  OAI21_X1  g065(.A(KEYINPUT90), .B1(new_n251), .B2(KEYINPUT20), .ZN(new_n252));
  AND3_X1   g066(.A1(new_n220), .A2(new_n224), .A3(new_n232), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n247), .A2(new_n248), .ZN(new_n254));
  NAND3_X1  g068(.A1(new_n237), .A2(new_n238), .A3(new_n239), .ZN(new_n255));
  NAND2_X1  g069(.A1(new_n255), .A2(KEYINPUT89), .ZN(new_n256));
  INV_X1    g070(.A(new_n245), .ZN(new_n257));
  NAND3_X1  g071(.A1(new_n207), .A2(new_n236), .A3(new_n238), .ZN(new_n258));
  NAND4_X1  g072(.A1(new_n254), .A2(new_n256), .A3(new_n257), .A4(new_n258), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n259), .A2(new_n232), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n253), .B1(new_n260), .B2(new_n223), .ZN(new_n261));
  INV_X1    g075(.A(KEYINPUT90), .ZN(new_n262));
  INV_X1    g076(.A(KEYINPUT20), .ZN(new_n263));
  NAND4_X1  g077(.A1(new_n261), .A2(new_n262), .A3(new_n263), .A4(new_n234), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n251), .A2(KEYINPUT20), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n252), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G478), .ZN(new_n267));
  NOR2_X1   g081(.A1(new_n267), .A2(KEYINPUT15), .ZN(new_n268));
  INV_X1    g082(.A(G902), .ZN(new_n269));
  XNOR2_X1  g083(.A(G128), .B(G143), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(KEYINPUT13), .ZN(new_n271));
  INV_X1    g085(.A(G128), .ZN(new_n272));
  NOR3_X1   g086(.A1(new_n272), .A2(KEYINPUT13), .A3(G143), .ZN(new_n273));
  INV_X1    g087(.A(G134), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  AOI22_X1  g089(.A1(new_n271), .A2(new_n275), .B1(new_n274), .B2(new_n270), .ZN(new_n276));
  INV_X1    g090(.A(G122), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n277), .A2(G116), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT92), .ZN(new_n279));
  XNOR2_X1  g093(.A(new_n278), .B(new_n279), .ZN(new_n280));
  INV_X1    g094(.A(G107), .ZN(new_n281));
  INV_X1    g095(.A(G116), .ZN(new_n282));
  NAND2_X1  g096(.A1(new_n282), .A2(G122), .ZN(new_n283));
  NAND3_X1  g097(.A1(new_n280), .A2(new_n281), .A3(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n281), .B1(new_n280), .B2(new_n283), .ZN(new_n286));
  OAI21_X1  g100(.A(new_n276), .B1(new_n285), .B2(new_n286), .ZN(new_n287));
  XNOR2_X1  g101(.A(new_n278), .B(KEYINPUT92), .ZN(new_n288));
  XNOR2_X1  g102(.A(new_n283), .B(KEYINPUT14), .ZN(new_n289));
  OAI21_X1  g103(.A(G107), .B1(new_n288), .B2(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(new_n270), .B(new_n274), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n284), .A3(new_n291), .ZN(new_n292));
  XOR2_X1   g106(.A(KEYINPUT72), .B(G217), .Z(new_n293));
  XNOR2_X1  g107(.A(KEYINPUT9), .B(G234), .ZN(new_n294));
  NOR3_X1   g108(.A1(new_n293), .A2(G953), .A3(new_n294), .ZN(new_n295));
  AND3_X1   g109(.A1(new_n287), .A2(new_n292), .A3(new_n295), .ZN(new_n296));
  AOI21_X1  g110(.A(new_n295), .B1(new_n287), .B2(new_n292), .ZN(new_n297));
  OAI21_X1  g111(.A(new_n269), .B1(new_n296), .B2(new_n297), .ZN(new_n298));
  AOI21_X1  g112(.A(new_n268), .B1(new_n298), .B2(KEYINPUT93), .ZN(new_n299));
  XNOR2_X1  g113(.A(new_n298), .B(KEYINPUT93), .ZN(new_n300));
  AOI21_X1  g114(.A(new_n299), .B1(new_n300), .B2(new_n268), .ZN(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(G952), .ZN(new_n303));
  AOI211_X1 g117(.A(G953), .B(new_n303), .C1(G234), .C2(G237), .ZN(new_n304));
  AOI211_X1 g118(.A(new_n269), .B(new_n192), .C1(G234), .C2(G237), .ZN(new_n305));
  XNOR2_X1  g119(.A(KEYINPUT21), .B(G898), .ZN(new_n306));
  AOI21_X1  g120(.A(new_n304), .B1(new_n305), .B2(new_n306), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n302), .A2(new_n307), .ZN(new_n308));
  NOR2_X1   g122(.A1(new_n223), .A2(KEYINPUT91), .ZN(new_n309));
  INV_X1    g123(.A(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n260), .A2(new_n310), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n259), .A2(new_n309), .A3(new_n232), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n311), .A2(new_n269), .A3(new_n312), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n313), .A2(G475), .ZN(new_n314));
  NAND3_X1  g128(.A1(new_n266), .A2(new_n308), .A3(new_n314), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(KEYINPUT94), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT94), .ZN(new_n317));
  NAND4_X1  g131(.A1(new_n266), .A2(new_n308), .A3(new_n317), .A4(new_n314), .ZN(new_n318));
  NAND2_X1  g132(.A1(new_n316), .A2(new_n318), .ZN(new_n319));
  XOR2_X1   g133(.A(KEYINPUT2), .B(G113), .Z(new_n320));
  XNOR2_X1  g134(.A(G116), .B(G119), .ZN(new_n321));
  XOR2_X1   g135(.A(new_n320), .B(new_n321), .Z(new_n322));
  OAI21_X1  g136(.A(KEYINPUT1), .B1(new_n194), .B2(G146), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n323), .A2(G128), .ZN(new_n324));
  NAND2_X1  g138(.A1(new_n230), .A2(G143), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n194), .A2(G146), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n324), .A2(new_n327), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT1), .ZN(new_n329));
  NAND4_X1  g143(.A1(new_n325), .A2(new_n326), .A3(new_n329), .A4(G128), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(KEYINPUT11), .B1(new_n274), .B2(G137), .ZN(new_n332));
  INV_X1    g146(.A(KEYINPUT11), .ZN(new_n333));
  INV_X1    g147(.A(G137), .ZN(new_n334));
  NAND3_X1  g148(.A1(new_n333), .A2(new_n334), .A3(G134), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n332), .A2(new_n335), .ZN(new_n336));
  OAI21_X1  g150(.A(KEYINPUT66), .B1(new_n334), .B2(G134), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT66), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n338), .A2(new_n274), .A3(G137), .ZN(new_n339));
  NAND4_X1  g153(.A1(new_n336), .A2(new_n228), .A3(new_n337), .A4(new_n339), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n274), .A2(G137), .ZN(new_n341));
  NOR2_X1   g155(.A1(new_n334), .A2(G134), .ZN(new_n342));
  OAI21_X1  g156(.A(G131), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  NAND3_X1  g157(.A1(new_n331), .A2(new_n340), .A3(new_n343), .ZN(new_n344));
  AND2_X1   g158(.A1(new_n332), .A2(new_n335), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n337), .A2(new_n339), .ZN(new_n346));
  OAI21_X1  g160(.A(G131), .B1(new_n345), .B2(new_n346), .ZN(new_n347));
  AND2_X1   g161(.A1(new_n347), .A2(new_n340), .ZN(new_n348));
  AND2_X1   g162(.A1(KEYINPUT0), .A2(G128), .ZN(new_n349));
  AOI21_X1  g163(.A(new_n349), .B1(new_n325), .B2(new_n326), .ZN(new_n350));
  INV_X1    g164(.A(KEYINPUT0), .ZN(new_n351));
  NAND3_X1  g165(.A1(new_n351), .A2(new_n272), .A3(KEYINPUT64), .ZN(new_n352));
  INV_X1    g166(.A(KEYINPUT64), .ZN(new_n353));
  OAI21_X1  g167(.A(new_n353), .B1(KEYINPUT0), .B2(G128), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n352), .A2(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n350), .A2(new_n355), .ZN(new_n356));
  INV_X1    g170(.A(KEYINPUT65), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  NAND3_X1  g172(.A1(new_n350), .A2(new_n355), .A3(KEYINPUT65), .ZN(new_n359));
  NAND3_X1  g173(.A1(new_n325), .A2(new_n326), .A3(new_n349), .ZN(new_n360));
  NAND3_X1  g174(.A1(new_n358), .A2(new_n359), .A3(new_n360), .ZN(new_n361));
  OAI211_X1 g175(.A(new_n322), .B(new_n344), .C1(new_n348), .C2(new_n361), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT28), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n362), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT70), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n364), .A2(new_n365), .ZN(new_n366));
  NAND3_X1  g180(.A1(new_n362), .A2(KEYINPUT70), .A3(new_n363), .ZN(new_n367));
  AND2_X1   g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n199), .A2(G210), .ZN(new_n369));
  XNOR2_X1  g183(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n370));
  XNOR2_X1  g184(.A(new_n369), .B(new_n370), .ZN(new_n371));
  XNOR2_X1  g185(.A(KEYINPUT26), .B(G101), .ZN(new_n372));
  XNOR2_X1  g186(.A(new_n371), .B(new_n372), .ZN(new_n373));
  INV_X1    g187(.A(new_n362), .ZN(new_n374));
  NAND2_X1  g188(.A1(new_n347), .A2(new_n340), .ZN(new_n375));
  AND2_X1   g189(.A1(new_n359), .A2(new_n360), .ZN(new_n376));
  NAND3_X1  g190(.A1(new_n375), .A2(new_n376), .A3(new_n358), .ZN(new_n377));
  AOI21_X1  g191(.A(new_n322), .B1(new_n377), .B2(new_n344), .ZN(new_n378));
  OAI21_X1  g192(.A(KEYINPUT28), .B1(new_n374), .B2(new_n378), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n368), .A2(KEYINPUT71), .A3(new_n373), .A4(new_n379), .ZN(new_n380));
  INV_X1    g194(.A(new_n322), .ZN(new_n381));
  INV_X1    g195(.A(KEYINPUT30), .ZN(new_n382));
  OAI211_X1 g196(.A(new_n382), .B(new_n344), .C1(new_n348), .C2(new_n361), .ZN(new_n383));
  INV_X1    g197(.A(new_n383), .ZN(new_n384));
  AOI21_X1  g198(.A(new_n382), .B1(new_n377), .B2(new_n344), .ZN(new_n385));
  OAI21_X1  g199(.A(new_n381), .B1(new_n384), .B2(new_n385), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(new_n362), .ZN(new_n387));
  INV_X1    g201(.A(new_n373), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n387), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n379), .A2(new_n366), .A3(new_n373), .A4(new_n367), .ZN(new_n390));
  INV_X1    g204(.A(KEYINPUT71), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  INV_X1    g206(.A(KEYINPUT29), .ZN(new_n393));
  NAND4_X1  g207(.A1(new_n380), .A2(new_n389), .A3(new_n392), .A4(new_n393), .ZN(new_n394));
  NOR2_X1   g208(.A1(new_n390), .A2(new_n393), .ZN(new_n395));
  NOR2_X1   g209(.A1(new_n395), .A2(G902), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n394), .A2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(G472), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT32), .ZN(new_n399));
  NAND3_X1  g213(.A1(new_n386), .A2(new_n362), .A3(new_n373), .ZN(new_n400));
  INV_X1    g214(.A(KEYINPUT69), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n400), .A2(new_n401), .ZN(new_n402));
  NAND4_X1  g216(.A1(new_n386), .A2(KEYINPUT69), .A3(new_n362), .A4(new_n373), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n402), .A2(KEYINPUT31), .A3(new_n403), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n344), .B1(new_n348), .B2(new_n361), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n405), .A2(KEYINPUT30), .ZN(new_n406));
  AOI21_X1  g220(.A(new_n322), .B1(new_n406), .B2(new_n383), .ZN(new_n407));
  NOR3_X1   g221(.A1(new_n407), .A2(new_n374), .A3(new_n388), .ZN(new_n408));
  INV_X1    g222(.A(KEYINPUT31), .ZN(new_n409));
  NAND3_X1  g223(.A1(new_n379), .A2(new_n366), .A3(new_n367), .ZN(new_n410));
  AOI22_X1  g224(.A1(new_n408), .A2(new_n409), .B1(new_n410), .B2(new_n388), .ZN(new_n411));
  NAND2_X1  g225(.A1(new_n404), .A2(new_n411), .ZN(new_n412));
  NOR2_X1   g226(.A1(G472), .A2(G902), .ZN(new_n413));
  AOI21_X1  g227(.A(new_n399), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n413), .ZN(new_n415));
  AOI211_X1 g229(.A(KEYINPUT32), .B(new_n415), .C1(new_n404), .C2(new_n411), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n398), .B1(new_n414), .B2(new_n416), .ZN(new_n417));
  AOI21_X1  g231(.A(new_n293), .B1(G234), .B2(new_n269), .ZN(new_n418));
  INV_X1    g232(.A(new_n418), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n209), .A2(new_n230), .ZN(new_n420));
  INV_X1    g234(.A(KEYINPUT23), .ZN(new_n421));
  INV_X1    g235(.A(G119), .ZN(new_n422));
  OAI21_X1  g236(.A(new_n421), .B1(new_n422), .B2(G128), .ZN(new_n423));
  NAND3_X1  g237(.A1(new_n272), .A2(KEYINPUT23), .A3(G119), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n423), .B(new_n424), .C1(G119), .C2(new_n272), .ZN(new_n425));
  XOR2_X1   g239(.A(KEYINPUT74), .B(G110), .Z(new_n426));
  XNOR2_X1  g240(.A(G119), .B(G128), .ZN(new_n427));
  XOR2_X1   g241(.A(KEYINPUT24), .B(G110), .Z(new_n428));
  OAI22_X1  g242(.A1(new_n425), .A2(new_n426), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  NAND4_X1  g243(.A1(new_n214), .A2(new_n216), .A3(new_n420), .A4(new_n429), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT22), .B(G137), .ZN(new_n431));
  NAND3_X1  g245(.A1(new_n192), .A2(G221), .A3(G234), .ZN(new_n432));
  XNOR2_X1  g246(.A(new_n431), .B(new_n432), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n428), .A2(new_n427), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n245), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g249(.A1(new_n425), .A2(G110), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT73), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND3_X1  g252(.A1(new_n425), .A2(KEYINPUT73), .A3(G110), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g254(.A(new_n430), .B(new_n433), .C1(new_n435), .C2(new_n440), .ZN(new_n441));
  AND2_X1   g255(.A1(new_n429), .A2(new_n420), .ZN(new_n442));
  AOI22_X1  g256(.A1(new_n244), .A2(new_n213), .B1(new_n427), .B2(new_n428), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n438), .A2(new_n439), .ZN(new_n444));
  AOI22_X1  g258(.A1(new_n218), .A2(new_n442), .B1(new_n443), .B2(new_n444), .ZN(new_n445));
  XOR2_X1   g259(.A(new_n433), .B(KEYINPUT76), .Z(new_n446));
  OAI211_X1 g260(.A(new_n441), .B(new_n269), .C1(new_n445), .C2(new_n446), .ZN(new_n447));
  INV_X1    g261(.A(KEYINPUT25), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n447), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(new_n446), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n430), .B1(new_n435), .B2(new_n440), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n450), .A2(new_n451), .ZN(new_n452));
  NAND4_X1  g266(.A1(new_n452), .A2(KEYINPUT25), .A3(new_n269), .A4(new_n441), .ZN(new_n453));
  AOI21_X1  g267(.A(new_n419), .B1(new_n449), .B2(new_n453), .ZN(new_n454));
  AND2_X1   g268(.A1(new_n452), .A2(new_n441), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n418), .A2(G902), .ZN(new_n456));
  AND2_X1   g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n454), .A2(new_n457), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n417), .A2(new_n458), .ZN(new_n459));
  INV_X1    g273(.A(new_n459), .ZN(new_n460));
  OAI21_X1  g274(.A(G221), .B1(new_n294), .B2(G902), .ZN(new_n461));
  INV_X1    g275(.A(new_n461), .ZN(new_n462));
  XNOR2_X1  g276(.A(G110), .B(G140), .ZN(new_n463));
  INV_X1    g277(.A(G227), .ZN(new_n464));
  NOR2_X1   g278(.A1(new_n464), .A2(G953), .ZN(new_n465));
  XNOR2_X1  g279(.A(new_n463), .B(new_n465), .ZN(new_n466));
  OAI21_X1  g280(.A(KEYINPUT3), .B1(new_n222), .B2(G107), .ZN(new_n467));
  INV_X1    g281(.A(KEYINPUT3), .ZN(new_n468));
  NAND3_X1  g282(.A1(new_n468), .A2(new_n281), .A3(G104), .ZN(new_n469));
  INV_X1    g283(.A(G101), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n222), .A2(G107), .ZN(new_n471));
  NAND4_X1  g285(.A1(new_n467), .A2(new_n469), .A3(new_n470), .A4(new_n471), .ZN(new_n472));
  NOR2_X1   g286(.A1(new_n222), .A2(G107), .ZN(new_n473));
  NOR2_X1   g287(.A1(new_n281), .A2(G104), .ZN(new_n474));
  OAI21_X1  g288(.A(G101), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g289(.A(new_n330), .ZN(new_n476));
  AOI22_X1  g290(.A1(new_n323), .A2(G128), .B1(new_n325), .B2(new_n326), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n472), .B(new_n475), .C1(new_n476), .C2(new_n477), .ZN(new_n478));
  INV_X1    g292(.A(KEYINPUT10), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n478), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n472), .A2(new_n475), .ZN(new_n481));
  INV_X1    g295(.A(new_n481), .ZN(new_n482));
  NAND3_X1  g296(.A1(new_n482), .A2(new_n331), .A3(KEYINPUT10), .ZN(new_n483));
  NAND2_X1  g297(.A1(new_n480), .A2(new_n483), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n472), .A2(KEYINPUT4), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n467), .A2(new_n469), .A3(new_n471), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT77), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n470), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  NAND4_X1  g302(.A1(new_n467), .A2(new_n469), .A3(KEYINPUT77), .A4(new_n471), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n485), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n486), .A2(new_n487), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT4), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n491), .A2(new_n492), .A3(G101), .A4(new_n489), .ZN(new_n493));
  NAND2_X1  g307(.A1(new_n493), .A2(KEYINPUT78), .ZN(new_n494));
  INV_X1    g308(.A(KEYINPUT78), .ZN(new_n495));
  NAND4_X1  g309(.A1(new_n488), .A2(new_n495), .A3(new_n492), .A4(new_n489), .ZN(new_n496));
  AOI21_X1  g310(.A(new_n490), .B1(new_n494), .B2(new_n496), .ZN(new_n497));
  INV_X1    g311(.A(new_n361), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n484), .B1(new_n497), .B2(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(new_n466), .B1(new_n499), .B2(new_n348), .ZN(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n348), .B2(new_n499), .ZN(new_n501));
  NAND2_X1  g315(.A1(new_n494), .A2(new_n496), .ZN(new_n502));
  INV_X1    g316(.A(new_n490), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n502), .A2(new_n498), .A3(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(new_n484), .ZN(new_n505));
  NAND3_X1  g319(.A1(new_n504), .A2(new_n348), .A3(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(KEYINPUT12), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n481), .A2(new_n330), .A3(new_n328), .ZN(new_n509));
  AOI221_X4 g323(.A(new_n508), .B1(new_n347), .B2(new_n340), .C1(new_n509), .C2(new_n478), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n509), .A2(new_n478), .ZN(new_n511));
  AOI21_X1  g325(.A(KEYINPUT12), .B1(new_n511), .B2(new_n375), .ZN(new_n512));
  NOR2_X1   g326(.A1(new_n510), .A2(new_n512), .ZN(new_n513));
  OAI21_X1  g327(.A(new_n466), .B1(new_n507), .B2(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n501), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(new_n515), .ZN(new_n516));
  OAI21_X1  g330(.A(G469), .B1(new_n516), .B2(G902), .ZN(new_n517));
  NAND2_X1  g331(.A1(new_n511), .A2(new_n375), .ZN(new_n518));
  NAND2_X1  g332(.A1(new_n518), .A2(new_n508), .ZN(new_n519));
  NAND3_X1  g333(.A1(new_n511), .A2(KEYINPUT12), .A3(new_n375), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n519), .A2(KEYINPUT79), .A3(new_n520), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT79), .ZN(new_n522));
  OAI21_X1  g336(.A(new_n522), .B1(new_n510), .B2(new_n512), .ZN(new_n523));
  INV_X1    g337(.A(new_n466), .ZN(new_n524));
  NAND4_X1  g338(.A1(new_n506), .A2(new_n521), .A3(new_n523), .A4(new_n524), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT80), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n500), .A2(KEYINPUT80), .A3(new_n523), .A4(new_n521), .ZN(new_n528));
  AOI21_X1  g342(.A(new_n348), .B1(new_n504), .B2(new_n505), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n466), .B1(new_n507), .B2(new_n529), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n527), .A2(new_n528), .A3(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G469), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n269), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n462), .B1(new_n517), .B2(new_n533), .ZN(new_n534));
  OAI21_X1  g348(.A(G214), .B1(G237), .B2(G902), .ZN(new_n535));
  OAI21_X1  g349(.A(G210), .B1(G237), .B2(G902), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n359), .A2(new_n360), .ZN(new_n537));
  AOI21_X1  g351(.A(KEYINPUT65), .B1(new_n350), .B2(new_n355), .ZN(new_n538));
  OAI21_X1  g352(.A(G125), .B1(new_n537), .B2(new_n538), .ZN(new_n539));
  INV_X1    g353(.A(KEYINPUT82), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n539), .A2(new_n540), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n361), .A2(KEYINPUT82), .A3(G125), .ZN(new_n542));
  NAND3_X1  g356(.A1(new_n328), .A2(new_n211), .A3(new_n330), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n541), .A2(new_n542), .A3(new_n543), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n192), .A2(G224), .ZN(new_n545));
  XOR2_X1   g359(.A(new_n544), .B(new_n545), .Z(new_n546));
  NAND3_X1  g360(.A1(new_n502), .A2(new_n381), .A3(new_n503), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n321), .A2(KEYINPUT5), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n422), .A2(G116), .ZN(new_n549));
  OAI211_X1 g363(.A(new_n548), .B(G113), .C1(KEYINPUT5), .C2(new_n549), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n320), .A2(new_n321), .ZN(new_n551));
  NAND2_X1  g365(.A1(new_n550), .A2(new_n551), .ZN(new_n552));
  NOR2_X1   g366(.A1(new_n552), .A2(new_n481), .ZN(new_n553));
  INV_X1    g367(.A(new_n553), .ZN(new_n554));
  XNOR2_X1  g368(.A(G110), .B(G122), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n547), .A2(new_n554), .A3(new_n555), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n547), .A2(new_n554), .ZN(new_n557));
  XOR2_X1   g371(.A(new_n555), .B(KEYINPUT81), .Z(new_n558));
  AOI22_X1  g372(.A1(new_n556), .A2(KEYINPUT6), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  AOI211_X1 g373(.A(new_n322), .B(new_n490), .C1(new_n494), .C2(new_n496), .ZN(new_n560));
  OAI21_X1  g374(.A(new_n558), .B1(new_n560), .B2(new_n553), .ZN(new_n561));
  INV_X1    g375(.A(KEYINPUT6), .ZN(new_n562));
  NOR2_X1   g376(.A1(new_n561), .A2(new_n562), .ZN(new_n563));
  OAI21_X1  g377(.A(new_n546), .B1(new_n559), .B2(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n545), .A2(KEYINPUT7), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n544), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(new_n565), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n541), .A2(new_n542), .A3(new_n543), .A4(new_n567), .ZN(new_n568));
  INV_X1    g382(.A(KEYINPUT84), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n569), .B1(new_n482), .B2(KEYINPUT83), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n570), .A2(new_n551), .A3(new_n550), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n555), .B(KEYINPUT8), .ZN(new_n572));
  OAI21_X1  g386(.A(new_n552), .B1(KEYINPUT84), .B2(new_n481), .ZN(new_n573));
  OAI211_X1 g387(.A(new_n571), .B(new_n572), .C1(new_n573), .C2(new_n570), .ZN(new_n574));
  NAND4_X1  g388(.A1(new_n556), .A2(new_n566), .A3(new_n568), .A4(new_n574), .ZN(new_n575));
  AND2_X1   g389(.A1(new_n575), .A2(new_n269), .ZN(new_n576));
  AOI21_X1  g390(.A(new_n536), .B1(new_n564), .B2(new_n576), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT85), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n577), .A2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(new_n536), .ZN(new_n580));
  XNOR2_X1  g394(.A(new_n544), .B(new_n545), .ZN(new_n581));
  INV_X1    g395(.A(new_n555), .ZN(new_n582));
  AOI211_X1 g396(.A(new_n553), .B(new_n582), .C1(new_n497), .C2(new_n381), .ZN(new_n583));
  OAI21_X1  g397(.A(new_n561), .B1(new_n583), .B2(new_n562), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n557), .A2(KEYINPUT6), .A3(new_n558), .ZN(new_n585));
  AOI21_X1  g399(.A(new_n581), .B1(new_n584), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n575), .A2(new_n269), .ZN(new_n587));
  OAI21_X1  g401(.A(new_n580), .B1(new_n586), .B2(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n564), .A2(new_n536), .A3(new_n576), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n588), .A2(new_n589), .A3(KEYINPUT85), .ZN(new_n590));
  NAND4_X1  g404(.A1(new_n534), .A2(new_n535), .A3(new_n579), .A4(new_n590), .ZN(new_n591));
  INV_X1    g405(.A(new_n591), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n319), .A2(new_n460), .A3(new_n592), .ZN(new_n593));
  XNOR2_X1  g407(.A(KEYINPUT95), .B(G101), .ZN(new_n594));
  XNOR2_X1  g408(.A(new_n593), .B(new_n594), .ZN(G3));
  NAND2_X1  g409(.A1(new_n266), .A2(new_n314), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n588), .A2(new_n589), .ZN(new_n597));
  NAND2_X1  g411(.A1(new_n597), .A2(new_n535), .ZN(new_n598));
  NOR2_X1   g412(.A1(new_n598), .A2(new_n307), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n298), .A2(new_n267), .ZN(new_n600));
  XOR2_X1   g414(.A(new_n600), .B(KEYINPUT96), .Z(new_n601));
  NOR2_X1   g415(.A1(new_n296), .A2(new_n297), .ZN(new_n602));
  XOR2_X1   g416(.A(new_n602), .B(KEYINPUT33), .Z(new_n603));
  NAND3_X1  g417(.A1(new_n603), .A2(G478), .A3(new_n269), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n601), .A2(new_n604), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n596), .A2(new_n599), .A3(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n412), .A2(new_n269), .ZN(new_n607));
  NAND2_X1  g421(.A1(new_n607), .A2(G472), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n412), .A2(new_n413), .ZN(new_n609));
  NAND4_X1  g423(.A1(new_n534), .A2(new_n608), .A3(new_n609), .A4(new_n458), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n606), .A2(new_n610), .ZN(new_n611));
  XNOR2_X1  g425(.A(KEYINPUT34), .B(G104), .ZN(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND3_X1  g427(.A1(new_n261), .A2(new_n263), .A3(new_n234), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n614), .A2(new_n265), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n301), .B1(new_n313), .B2(G475), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n615), .A2(new_n616), .ZN(new_n617));
  NOR4_X1   g431(.A1(new_n610), .A2(new_n307), .A3(new_n617), .A4(new_n598), .ZN(new_n618));
  XNOR2_X1  g432(.A(KEYINPUT35), .B(G107), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n618), .B(new_n619), .ZN(G9));
  NAND2_X1  g434(.A1(new_n608), .A2(new_n609), .ZN(new_n621));
  INV_X1    g435(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n449), .A2(new_n453), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n418), .ZN(new_n624));
  NOR2_X1   g438(.A1(new_n450), .A2(KEYINPUT36), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(new_n451), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(new_n456), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n624), .A2(new_n627), .ZN(new_n628));
  AOI21_X1  g442(.A(KEYINPUT97), .B1(new_n622), .B2(new_n628), .ZN(new_n629));
  INV_X1    g443(.A(KEYINPUT97), .ZN(new_n630));
  INV_X1    g444(.A(new_n628), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n621), .A2(new_n630), .A3(new_n631), .ZN(new_n632));
  NOR2_X1   g446(.A1(new_n629), .A2(new_n632), .ZN(new_n633));
  AOI21_X1  g447(.A(new_n591), .B1(new_n316), .B2(new_n318), .ZN(new_n634));
  NAND2_X1  g448(.A1(new_n633), .A2(new_n634), .ZN(new_n635));
  XOR2_X1   g449(.A(KEYINPUT37), .B(G110), .Z(new_n636));
  XNOR2_X1  g450(.A(new_n636), .B(KEYINPUT98), .ZN(new_n637));
  XNOR2_X1  g451(.A(new_n635), .B(new_n637), .ZN(G12));
  INV_X1    g452(.A(new_n598), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n417), .A2(new_n534), .A3(new_n639), .A4(new_n628), .ZN(new_n640));
  INV_X1    g454(.A(G900), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n305), .A2(new_n641), .ZN(new_n642));
  INV_X1    g456(.A(new_n304), .ZN(new_n643));
  NAND2_X1  g457(.A1(new_n642), .A2(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NOR2_X1   g459(.A1(new_n617), .A2(new_n645), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n640), .A2(new_n646), .ZN(new_n647));
  XNOR2_X1  g461(.A(new_n647), .B(G128), .ZN(G30));
  NAND2_X1  g462(.A1(new_n590), .A2(new_n579), .ZN(new_n649));
  XOR2_X1   g463(.A(new_n649), .B(KEYINPUT38), .Z(new_n650));
  XNOR2_X1  g464(.A(new_n644), .B(KEYINPUT39), .ZN(new_n651));
  NAND2_X1  g465(.A1(new_n534), .A2(new_n651), .ZN(new_n652));
  XOR2_X1   g466(.A(new_n652), .B(KEYINPUT40), .Z(new_n653));
  INV_X1    g467(.A(new_n596), .ZN(new_n654));
  NOR2_X1   g468(.A1(new_n654), .A2(new_n301), .ZN(new_n655));
  INV_X1    g469(.A(G472), .ZN(new_n656));
  AND2_X1   g470(.A1(new_n402), .A2(new_n403), .ZN(new_n657));
  OAI21_X1  g471(.A(new_n388), .B1(new_n374), .B2(new_n378), .ZN(new_n658));
  AOI21_X1  g472(.A(G902), .B1(new_n657), .B2(new_n658), .ZN(new_n659));
  OAI22_X1  g473(.A1(new_n414), .A2(new_n416), .B1(new_n656), .B2(new_n659), .ZN(new_n660));
  AND3_X1   g474(.A1(new_n660), .A2(new_n535), .A3(new_n631), .ZN(new_n661));
  AND4_X1   g475(.A1(new_n650), .A2(new_n653), .A3(new_n655), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(new_n194), .ZN(G45));
  NAND3_X1  g477(.A1(new_n596), .A2(new_n605), .A3(new_n644), .ZN(new_n664));
  NAND2_X1  g478(.A1(new_n664), .A2(KEYINPUT99), .ZN(new_n665));
  AOI22_X1  g479(.A1(new_n266), .A2(new_n314), .B1(new_n601), .B2(new_n604), .ZN(new_n666));
  INV_X1    g480(.A(KEYINPUT99), .ZN(new_n667));
  NAND3_X1  g481(.A1(new_n666), .A2(new_n667), .A3(new_n644), .ZN(new_n668));
  NAND3_X1  g482(.A1(new_n665), .A2(new_n640), .A3(new_n668), .ZN(new_n669));
  INV_X1    g483(.A(KEYINPUT100), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n669), .A2(new_n670), .ZN(new_n671));
  NAND4_X1  g485(.A1(new_n665), .A2(KEYINPUT100), .A3(new_n668), .A4(new_n640), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(new_n673), .B(G146), .ZN(G48));
  INV_X1    g488(.A(new_n533), .ZN(new_n675));
  AOI21_X1  g489(.A(new_n532), .B1(new_n531), .B2(new_n269), .ZN(new_n676));
  NOR3_X1   g490(.A1(new_n675), .A2(new_n676), .A3(new_n462), .ZN(new_n677));
  NAND3_X1  g491(.A1(new_n417), .A2(new_n458), .A3(new_n677), .ZN(new_n678));
  NOR2_X1   g492(.A1(new_n606), .A2(new_n678), .ZN(new_n679));
  XOR2_X1   g493(.A(KEYINPUT41), .B(G113), .Z(new_n680));
  XNOR2_X1  g494(.A(new_n679), .B(new_n680), .ZN(G15));
  NOR3_X1   g495(.A1(new_n454), .A2(new_n457), .A3(new_n307), .ZN(new_n682));
  AND3_X1   g496(.A1(new_n615), .A2(new_n616), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g497(.A1(new_n531), .A2(new_n269), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  NAND3_X1  g499(.A1(new_n685), .A2(new_n461), .A3(new_n533), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n686), .A2(new_n598), .ZN(new_n687));
  NAND3_X1  g501(.A1(new_n683), .A2(new_n687), .A3(new_n417), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G116), .ZN(G18));
  NAND4_X1  g503(.A1(new_n417), .A2(new_n639), .A3(new_n628), .A4(new_n677), .ZN(new_n690));
  AOI21_X1  g504(.A(new_n690), .B1(new_n318), .B2(new_n316), .ZN(new_n691));
  XNOR2_X1  g505(.A(new_n691), .B(new_n422), .ZN(G21));
  AOI211_X1 g506(.A(new_n301), .B(new_n598), .C1(new_n266), .C2(new_n314), .ZN(new_n693));
  INV_X1    g507(.A(KEYINPUT102), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n455), .A2(new_n456), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n624), .A2(new_n694), .A3(new_n695), .ZN(new_n696));
  OAI21_X1  g510(.A(KEYINPUT102), .B1(new_n454), .B2(new_n457), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n696), .A2(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n413), .B(KEYINPUT101), .ZN(new_n699));
  NAND2_X1  g513(.A1(new_n412), .A2(new_n699), .ZN(new_n700));
  AOI21_X1  g514(.A(G902), .B1(new_n404), .B2(new_n411), .ZN(new_n701));
  OAI211_X1 g515(.A(new_n698), .B(new_n700), .C1(new_n656), .C2(new_n701), .ZN(new_n702));
  INV_X1    g516(.A(KEYINPUT103), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n702), .A2(new_n703), .ZN(new_n704));
  NAND4_X1  g518(.A1(new_n608), .A2(KEYINPUT103), .A3(new_n698), .A4(new_n700), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NOR2_X1   g520(.A1(new_n686), .A2(new_n307), .ZN(new_n707));
  AND3_X1   g521(.A1(new_n693), .A2(new_n706), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(new_n277), .ZN(G24));
  INV_X1    g523(.A(new_n687), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n608), .A2(new_n628), .A3(new_n700), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n665), .A2(new_n712), .A3(new_n668), .ZN(new_n713));
  XNOR2_X1  g527(.A(new_n713), .B(G125), .ZN(G27));
  AND2_X1   g528(.A1(new_n417), .A2(new_n698), .ZN(new_n715));
  NAND3_X1  g529(.A1(new_n665), .A2(new_n668), .A3(new_n715), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n649), .A2(new_n535), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(KEYINPUT104), .ZN(new_n718));
  INV_X1    g532(.A(KEYINPUT104), .ZN(new_n719));
  NAND3_X1  g533(.A1(new_n649), .A2(new_n719), .A3(new_n535), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n718), .A2(new_n534), .A3(new_n720), .ZN(new_n721));
  OAI21_X1  g535(.A(KEYINPUT42), .B1(new_n716), .B2(new_n721), .ZN(new_n722));
  NOR2_X1   g536(.A1(new_n721), .A2(new_n459), .ZN(new_n723));
  INV_X1    g537(.A(KEYINPUT42), .ZN(new_n724));
  NAND4_X1  g538(.A1(new_n723), .A2(new_n724), .A3(new_n668), .A4(new_n665), .ZN(new_n725));
  AND2_X1   g539(.A1(new_n722), .A2(new_n725), .ZN(new_n726));
  XOR2_X1   g540(.A(KEYINPUT105), .B(G131), .Z(new_n727));
  XNOR2_X1  g541(.A(new_n726), .B(new_n727), .ZN(G33));
  AOI21_X1  g542(.A(new_n719), .B1(new_n649), .B2(new_n535), .ZN(new_n729));
  INV_X1    g543(.A(new_n535), .ZN(new_n730));
  AOI211_X1 g544(.A(KEYINPUT104), .B(new_n730), .C1(new_n590), .C2(new_n579), .ZN(new_n731));
  INV_X1    g545(.A(new_n534), .ZN(new_n732));
  NOR3_X1   g546(.A1(new_n729), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n733), .A2(new_n460), .A3(new_n646), .ZN(new_n734));
  XNOR2_X1  g548(.A(new_n734), .B(G134), .ZN(G36));
  INV_X1    g549(.A(KEYINPUT45), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n532), .B1(new_n515), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n736), .B2(new_n515), .ZN(new_n738));
  NAND2_X1  g552(.A1(G469), .A2(G902), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n738), .A2(new_n739), .ZN(new_n740));
  INV_X1    g554(.A(KEYINPUT46), .ZN(new_n741));
  NAND2_X1  g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  NAND2_X1  g556(.A1(new_n742), .A2(new_n533), .ZN(new_n743));
  NOR2_X1   g557(.A1(new_n740), .A2(new_n741), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n461), .B(new_n651), .C1(new_n743), .C2(new_n744), .ZN(new_n745));
  NOR2_X1   g559(.A1(new_n729), .A2(new_n731), .ZN(new_n746));
  INV_X1    g560(.A(new_n746), .ZN(new_n747));
  NOR2_X1   g561(.A1(new_n745), .A2(new_n747), .ZN(new_n748));
  INV_X1    g562(.A(KEYINPUT43), .ZN(new_n749));
  NAND2_X1  g563(.A1(new_n749), .A2(KEYINPUT106), .ZN(new_n750));
  XOR2_X1   g564(.A(KEYINPUT106), .B(KEYINPUT43), .Z(new_n751));
  NAND2_X1  g565(.A1(new_n654), .A2(new_n605), .ZN(new_n752));
  MUX2_X1   g566(.A(new_n750), .B(new_n751), .S(new_n752), .Z(new_n753));
  NOR2_X1   g567(.A1(new_n622), .A2(new_n631), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n753), .A2(new_n754), .ZN(new_n755));
  AND2_X1   g569(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n756));
  NOR2_X1   g570(.A1(new_n755), .A2(KEYINPUT44), .ZN(new_n757));
  OAI21_X1  g571(.A(new_n748), .B1(new_n756), .B2(new_n757), .ZN(new_n758));
  XNOR2_X1  g572(.A(new_n758), .B(G137), .ZN(G39));
  OAI21_X1  g573(.A(new_n461), .B1(new_n743), .B2(new_n744), .ZN(new_n760));
  XNOR2_X1  g574(.A(KEYINPUT107), .B(KEYINPUT47), .ZN(new_n761));
  XNOR2_X1  g575(.A(new_n760), .B(new_n761), .ZN(new_n762));
  INV_X1    g576(.A(new_n762), .ZN(new_n763));
  NOR3_X1   g577(.A1(new_n763), .A2(new_n417), .A3(new_n458), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n764), .A2(new_n668), .A3(new_n665), .A4(new_n746), .ZN(new_n765));
  XNOR2_X1  g579(.A(new_n765), .B(G140), .ZN(G42));
  NOR2_X1   g580(.A1(new_n675), .A2(new_n676), .ZN(new_n767));
  INV_X1    g581(.A(KEYINPUT49), .ZN(new_n768));
  NOR2_X1   g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g583(.A1(new_n698), .A2(new_n535), .A3(new_n461), .ZN(new_n770));
  NOR3_X1   g584(.A1(new_n752), .A2(new_n769), .A3(new_n770), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT108), .ZN(new_n772));
  OR2_X1    g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  AOI211_X1 g587(.A(new_n660), .B(new_n650), .C1(new_n768), .C2(new_n767), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND3_X1  g589(.A1(new_n773), .A2(new_n774), .A3(new_n775), .ZN(new_n776));
  NOR2_X1   g590(.A1(new_n711), .A2(new_n732), .ZN(new_n777));
  NAND4_X1  g591(.A1(new_n665), .A2(new_n668), .A3(new_n746), .A4(new_n777), .ZN(new_n778));
  AND2_X1   g592(.A1(new_n778), .A2(new_n734), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT110), .ZN(new_n780));
  NOR3_X1   g594(.A1(new_n302), .A2(new_n631), .A3(new_n645), .ZN(new_n781));
  AND4_X1   g595(.A1(new_n417), .A2(new_n314), .A3(new_n615), .A4(new_n781), .ZN(new_n782));
  AND4_X1   g596(.A1(new_n780), .A2(new_n782), .A3(new_n746), .A4(new_n534), .ZN(new_n783));
  AOI21_X1  g597(.A(new_n780), .B1(new_n733), .B2(new_n782), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g599(.A1(new_n779), .A2(new_n785), .A3(new_n722), .A4(new_n725), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n591), .B(new_n459), .C1(new_n316), .C2(new_n318), .ZN(new_n787));
  INV_X1    g601(.A(new_n307), .ZN(new_n788));
  NAND4_X1  g602(.A1(new_n590), .A2(new_n579), .A3(new_n788), .A4(new_n535), .ZN(new_n789));
  NOR2_X1   g603(.A1(new_n610), .A2(new_n789), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n790), .A2(new_n666), .ZN(new_n791));
  INV_X1    g605(.A(new_n791), .ZN(new_n792));
  OAI21_X1  g606(.A(KEYINPUT109), .B1(new_n787), .B2(new_n792), .ZN(new_n793));
  OAI21_X1  g607(.A(new_n688), .B1(new_n606), .B2(new_n678), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n708), .A2(new_n691), .A3(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT109), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n593), .A2(new_n796), .A3(new_n791), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n596), .A2(new_n301), .ZN(new_n798));
  AOI22_X1  g612(.A1(new_n633), .A2(new_n634), .B1(new_n790), .B2(new_n798), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n793), .A2(new_n795), .A3(new_n797), .A4(new_n799), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n786), .A2(new_n800), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n713), .A2(new_n647), .ZN(new_n802));
  AOI21_X1  g616(.A(new_n802), .B1(new_n671), .B2(new_n672), .ZN(new_n803));
  NAND3_X1  g617(.A1(new_n534), .A2(new_n631), .A3(new_n644), .ZN(new_n804));
  XNOR2_X1  g618(.A(new_n804), .B(KEYINPUT111), .ZN(new_n805));
  NAND3_X1  g619(.A1(new_n805), .A2(new_n660), .A3(new_n693), .ZN(new_n806));
  AOI21_X1  g620(.A(KEYINPUT52), .B1(new_n803), .B2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n802), .ZN(new_n808));
  AND4_X1   g622(.A1(KEYINPUT52), .A2(new_n673), .A3(new_n808), .A4(new_n806), .ZN(new_n809));
  OAI21_X1  g623(.A(new_n801), .B1(new_n807), .B2(new_n809), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT53), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT53), .ZN(new_n812));
  NAND3_X1  g626(.A1(new_n673), .A2(new_n808), .A3(new_n806), .ZN(new_n813));
  XNOR2_X1  g627(.A(KEYINPUT113), .B(KEYINPUT52), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n813), .A2(KEYINPUT112), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n814), .B1(new_n813), .B2(KEYINPUT112), .ZN(new_n816));
  OAI211_X1 g630(.A(new_n812), .B(new_n801), .C1(new_n815), .C2(new_n816), .ZN(new_n817));
  AND2_X1   g631(.A1(new_n811), .A2(new_n817), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n818), .A2(KEYINPUT54), .ZN(new_n819));
  INV_X1    g633(.A(KEYINPUT115), .ZN(new_n820));
  OR2_X1    g634(.A1(new_n795), .A2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n795), .A2(new_n820), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n821), .A2(KEYINPUT53), .A3(new_n822), .ZN(new_n823));
  NAND3_X1  g637(.A1(new_n793), .A2(new_n797), .A3(new_n799), .ZN(new_n824));
  NOR3_X1   g638(.A1(new_n823), .A2(new_n824), .A3(new_n786), .ZN(new_n825));
  OAI21_X1  g639(.A(new_n825), .B1(new_n816), .B2(new_n815), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT114), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT52), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n813), .A2(new_n828), .ZN(new_n829));
  NAND3_X1  g643(.A1(new_n803), .A2(KEYINPUT52), .A3(new_n806), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AOI211_X1 g645(.A(new_n827), .B(KEYINPUT53), .C1(new_n831), .C2(new_n801), .ZN(new_n832));
  AOI21_X1  g646(.A(KEYINPUT114), .B1(new_n810), .B2(new_n812), .ZN(new_n833));
  OAI21_X1  g647(.A(new_n826), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  OAI21_X1  g648(.A(new_n819), .B1(new_n834), .B2(KEYINPUT54), .ZN(new_n835));
  XOR2_X1   g649(.A(KEYINPUT116), .B(KEYINPUT51), .Z(new_n836));
  AND2_X1   g650(.A1(new_n753), .A2(new_n304), .ZN(new_n837));
  NOR3_X1   g651(.A1(new_n650), .A2(new_n535), .A3(new_n686), .ZN(new_n838));
  NAND3_X1  g652(.A1(new_n837), .A2(new_n706), .A3(new_n838), .ZN(new_n839));
  XOR2_X1   g653(.A(new_n839), .B(KEYINPUT50), .Z(new_n840));
  NAND2_X1  g654(.A1(new_n458), .A2(new_n304), .ZN(new_n841));
  OR4_X1    g655(.A1(new_n660), .A2(new_n747), .A3(new_n686), .A4(new_n841), .ZN(new_n842));
  NOR3_X1   g656(.A1(new_n842), .A2(new_n596), .A3(new_n605), .ZN(new_n843));
  NOR2_X1   g657(.A1(new_n747), .A2(new_n686), .ZN(new_n844));
  AND2_X1   g658(.A1(new_n837), .A2(new_n844), .ZN(new_n845));
  INV_X1    g659(.A(new_n711), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n843), .B1(new_n845), .B2(new_n846), .ZN(new_n847));
  NAND2_X1  g661(.A1(new_n840), .A2(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(new_n848), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n837), .A2(new_n706), .ZN(new_n850));
  NOR2_X1   g664(.A1(new_n850), .A2(new_n747), .ZN(new_n851));
  NOR2_X1   g665(.A1(new_n763), .A2(KEYINPUT117), .ZN(new_n852));
  NAND2_X1  g666(.A1(new_n767), .A2(new_n462), .ZN(new_n853));
  INV_X1    g667(.A(KEYINPUT117), .ZN(new_n854));
  OAI21_X1  g668(.A(new_n853), .B1(new_n762), .B2(new_n854), .ZN(new_n855));
  OAI21_X1  g669(.A(new_n851), .B1(new_n852), .B2(new_n855), .ZN(new_n856));
  AOI21_X1  g670(.A(new_n836), .B1(new_n849), .B2(new_n856), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n303), .A2(G953), .ZN(new_n858));
  INV_X1    g672(.A(new_n666), .ZN(new_n859));
  OAI221_X1 g673(.A(new_n858), .B1(new_n859), .B2(new_n842), .C1(new_n850), .C2(new_n710), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n845), .A2(new_n715), .ZN(new_n861));
  OR2_X1    g675(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n862));
  NAND2_X1  g676(.A1(new_n861), .A2(KEYINPUT48), .ZN(new_n863));
  AOI21_X1  g677(.A(new_n860), .B1(new_n862), .B2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n763), .A2(new_n853), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n851), .A2(new_n865), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n866), .A2(KEYINPUT51), .ZN(new_n867));
  OAI21_X1  g681(.A(new_n864), .B1(new_n848), .B2(new_n867), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n835), .A2(new_n857), .A3(new_n868), .ZN(new_n869));
  NOR2_X1   g683(.A1(G952), .A2(G953), .ZN(new_n870));
  OAI21_X1  g684(.A(new_n776), .B1(new_n869), .B2(new_n870), .ZN(G75));
  NAND2_X1  g685(.A1(new_n303), .A2(G953), .ZN(new_n872));
  XOR2_X1   g686(.A(new_n872), .B(KEYINPUT119), .Z(new_n873));
  INV_X1    g687(.A(new_n873), .ZN(new_n874));
  INV_X1    g688(.A(KEYINPUT56), .ZN(new_n875));
  NAND2_X1  g689(.A1(new_n834), .A2(G902), .ZN(new_n876));
  INV_X1    g690(.A(G210), .ZN(new_n877));
  OAI21_X1  g691(.A(new_n875), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n559), .A2(new_n563), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n879), .A2(new_n581), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(new_n564), .ZN(new_n881));
  XNOR2_X1  g695(.A(new_n881), .B(KEYINPUT55), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  AOI21_X1  g697(.A(new_n882), .B1(new_n883), .B2(new_n875), .ZN(new_n884));
  OR2_X1    g698(.A1(new_n878), .A2(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n878), .A2(new_n884), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n874), .B1(new_n885), .B2(new_n886), .ZN(G51));
  INV_X1    g701(.A(KEYINPUT54), .ZN(new_n888));
  XNOR2_X1  g702(.A(new_n834), .B(new_n888), .ZN(new_n889));
  XNOR2_X1  g703(.A(new_n739), .B(KEYINPUT57), .ZN(new_n890));
  OAI21_X1  g704(.A(new_n531), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  OR2_X1    g705(.A1(new_n876), .A2(new_n738), .ZN(new_n892));
  AOI21_X1  g706(.A(new_n874), .B1(new_n891), .B2(new_n892), .ZN(G54));
  AND4_X1   g707(.A1(KEYINPUT58), .A2(new_n834), .A3(G475), .A4(G902), .ZN(new_n894));
  INV_X1    g708(.A(new_n261), .ZN(new_n895));
  OR2_X1    g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND2_X1  g710(.A1(new_n894), .A2(new_n895), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n874), .B1(new_n896), .B2(new_n897), .ZN(G60));
  XNOR2_X1  g712(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n899));
  NAND2_X1  g713(.A1(G478), .A2(G902), .ZN(new_n900));
  XNOR2_X1  g714(.A(new_n899), .B(new_n900), .ZN(new_n901));
  NAND2_X1  g715(.A1(new_n603), .A2(new_n901), .ZN(new_n902));
  OAI21_X1  g716(.A(new_n873), .B1(new_n889), .B2(new_n902), .ZN(new_n903));
  AOI21_X1  g717(.A(new_n603), .B1(new_n835), .B2(new_n901), .ZN(new_n904));
  NOR2_X1   g718(.A1(new_n903), .A2(new_n904), .ZN(G63));
  NAND2_X1  g719(.A1(G217), .A2(G902), .ZN(new_n906));
  XNOR2_X1  g720(.A(new_n906), .B(KEYINPUT60), .ZN(new_n907));
  INV_X1    g721(.A(new_n907), .ZN(new_n908));
  NAND3_X1  g722(.A1(new_n834), .A2(new_n626), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n810), .A2(new_n812), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n910), .A2(new_n827), .ZN(new_n911));
  NAND3_X1  g725(.A1(new_n810), .A2(KEYINPUT114), .A3(new_n812), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  AOI21_X1  g727(.A(new_n907), .B1(new_n913), .B2(new_n826), .ZN(new_n914));
  OAI211_X1 g728(.A(new_n873), .B(new_n909), .C1(new_n914), .C2(new_n455), .ZN(new_n915));
  INV_X1    g729(.A(KEYINPUT121), .ZN(new_n916));
  AND3_X1   g730(.A1(new_n915), .A2(new_n916), .A3(KEYINPUT61), .ZN(new_n917));
  AOI21_X1  g731(.A(KEYINPUT61), .B1(new_n915), .B2(new_n916), .ZN(new_n918));
  NOR2_X1   g732(.A1(new_n917), .A2(new_n918), .ZN(G66));
  INV_X1    g733(.A(G224), .ZN(new_n920));
  OAI21_X1  g734(.A(G953), .B1(new_n306), .B2(new_n920), .ZN(new_n921));
  INV_X1    g735(.A(new_n800), .ZN(new_n922));
  OAI21_X1  g736(.A(new_n921), .B1(new_n922), .B2(G953), .ZN(new_n923));
  OAI21_X1  g737(.A(new_n879), .B1(G898), .B2(new_n192), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT122), .ZN(new_n925));
  XNOR2_X1  g739(.A(new_n923), .B(new_n925), .ZN(G69));
  NOR2_X1   g740(.A1(new_n384), .A2(new_n385), .ZN(new_n927));
  XNOR2_X1  g741(.A(new_n219), .B(KEYINPUT123), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n927), .B(new_n928), .ZN(new_n929));
  AND2_X1   g743(.A1(new_n758), .A2(new_n765), .ZN(new_n930));
  INV_X1    g744(.A(new_n662), .ZN(new_n931));
  NAND2_X1  g745(.A1(new_n803), .A2(new_n931), .ZN(new_n932));
  XOR2_X1   g746(.A(new_n932), .B(KEYINPUT62), .Z(new_n933));
  OAI211_X1 g747(.A(new_n723), .B(new_n651), .C1(new_n666), .C2(new_n798), .ZN(new_n934));
  AND3_X1   g748(.A1(new_n930), .A2(new_n933), .A3(new_n934), .ZN(new_n935));
  OAI21_X1  g749(.A(new_n929), .B1(new_n935), .B2(G953), .ZN(new_n936));
  NOR2_X1   g750(.A1(new_n192), .A2(G900), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n693), .A2(new_n715), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n745), .A2(new_n938), .ZN(new_n939));
  AOI21_X1  g753(.A(new_n939), .B1(new_n646), .B2(new_n723), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n726), .A2(new_n940), .ZN(new_n941));
  INV_X1    g755(.A(new_n941), .ZN(new_n942));
  NAND4_X1  g756(.A1(new_n930), .A2(KEYINPUT125), .A3(new_n803), .A4(new_n942), .ZN(new_n943));
  INV_X1    g757(.A(KEYINPUT125), .ZN(new_n944));
  NAND3_X1  g758(.A1(new_n758), .A2(new_n765), .A3(new_n803), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n944), .B1(new_n945), .B2(new_n941), .ZN(new_n946));
  NAND2_X1  g760(.A1(new_n943), .A2(new_n946), .ZN(new_n947));
  AOI21_X1  g761(.A(new_n937), .B1(new_n947), .B2(new_n192), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n936), .B1(new_n948), .B2(new_n929), .ZN(new_n949));
  OAI21_X1  g763(.A(G953), .B1(new_n464), .B2(new_n641), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT124), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n949), .B(new_n951), .ZN(G72));
  XNOR2_X1  g766(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n656), .A2(new_n269), .ZN(new_n954));
  XOR2_X1   g768(.A(new_n953), .B(new_n954), .Z(new_n955));
  INV_X1    g769(.A(new_n955), .ZN(new_n956));
  AOI21_X1  g770(.A(new_n956), .B1(new_n657), .B2(new_n389), .ZN(new_n957));
  NAND2_X1  g771(.A1(new_n818), .A2(new_n957), .ZN(new_n958));
  XOR2_X1   g772(.A(new_n958), .B(KEYINPUT127), .Z(new_n959));
  OAI21_X1  g773(.A(new_n955), .B1(new_n947), .B2(new_n800), .ZN(new_n960));
  NAND4_X1  g774(.A1(new_n960), .A2(new_n362), .A3(new_n386), .A4(new_n388), .ZN(new_n961));
  AND2_X1   g775(.A1(new_n935), .A2(new_n922), .ZN(new_n962));
  OAI211_X1 g776(.A(new_n387), .B(new_n373), .C1(new_n962), .C2(new_n956), .ZN(new_n963));
  AND4_X1   g777(.A1(new_n873), .A2(new_n959), .A3(new_n961), .A4(new_n963), .ZN(G57));
endmodule


