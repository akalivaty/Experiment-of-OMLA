//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 0 0 1 1 0 0 1 1 0 1 0 1 0 1 0 0 0 1 0 0 1 1 0 1 0 0 0 1 1 1 1 1 0 0 1 0 1 1 1 0 0 1 0 0 1 0 1 1 1 1 0 0 0 1 0 1 1 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:27:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n625, new_n626, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n655, new_n656, new_n657, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n674, new_n675,
    new_n676, new_n677, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n685, new_n686, new_n688, new_n689, new_n691, new_n692,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n745,
    new_n746, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n780, new_n781, new_n782,
    new_n783, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n901, new_n902, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n928, new_n929, new_n930, new_n931, new_n932, new_n933, new_n934,
    new_n935, new_n936, new_n937, new_n938, new_n939, new_n940, new_n942,
    new_n943, new_n944, new_n945, new_n946, new_n947, new_n948, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n974, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n986, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n992, new_n993, new_n994;
  NOR2_X1   g000(.A1(G472), .A2(G902), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  INV_X1    g003(.A(G143), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G146), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n189), .A2(new_n191), .ZN(new_n192));
  NOR2_X1   g006(.A1(KEYINPUT0), .A2(G128), .ZN(new_n193));
  INV_X1    g007(.A(KEYINPUT0), .ZN(new_n194));
  INV_X1    g008(.A(G128), .ZN(new_n195));
  NOR2_X1   g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  OAI21_X1  g010(.A(new_n192), .B1(new_n193), .B2(new_n196), .ZN(new_n197));
  OAI211_X1 g011(.A(new_n189), .B(new_n191), .C1(new_n194), .C2(new_n195), .ZN(new_n198));
  NAND2_X1  g012(.A1(new_n197), .A2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(G134), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(G137), .ZN(new_n201));
  INV_X1    g015(.A(G137), .ZN(new_n202));
  AOI21_X1  g016(.A(KEYINPUT64), .B1(new_n202), .B2(G134), .ZN(new_n203));
  INV_X1    g017(.A(KEYINPUT11), .ZN(new_n204));
  OAI21_X1  g018(.A(new_n201), .B1(new_n203), .B2(new_n204), .ZN(new_n205));
  INV_X1    g019(.A(KEYINPUT64), .ZN(new_n206));
  OAI211_X1 g020(.A(new_n206), .B(new_n204), .C1(new_n200), .C2(G137), .ZN(new_n207));
  INV_X1    g021(.A(new_n207), .ZN(new_n208));
  NOR3_X1   g022(.A1(new_n205), .A2(new_n208), .A3(G131), .ZN(new_n209));
  INV_X1    g023(.A(G131), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n202), .A2(G134), .ZN(new_n211));
  OAI21_X1  g025(.A(new_n206), .B1(new_n200), .B2(G137), .ZN(new_n212));
  AOI21_X1  g026(.A(new_n211), .B1(new_n212), .B2(KEYINPUT11), .ZN(new_n213));
  AOI21_X1  g027(.A(new_n210), .B1(new_n213), .B2(new_n207), .ZN(new_n214));
  OAI21_X1  g028(.A(new_n199), .B1(new_n209), .B2(new_n214), .ZN(new_n215));
  INV_X1    g029(.A(G119), .ZN(new_n216));
  OAI21_X1  g030(.A(KEYINPUT66), .B1(new_n216), .B2(G116), .ZN(new_n217));
  INV_X1    g031(.A(KEYINPUT66), .ZN(new_n218));
  INV_X1    g032(.A(G116), .ZN(new_n219));
  NAND3_X1  g033(.A1(new_n218), .A2(new_n219), .A3(G119), .ZN(new_n220));
  AOI22_X1  g034(.A1(new_n217), .A2(new_n220), .B1(G116), .B2(new_n216), .ZN(new_n221));
  NOR2_X1   g035(.A1(KEYINPUT2), .A2(G113), .ZN(new_n222));
  NAND2_X1  g036(.A1(KEYINPUT2), .A2(G113), .ZN(new_n223));
  INV_X1    g037(.A(KEYINPUT65), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND3_X1  g039(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n226));
  AOI21_X1  g040(.A(new_n222), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  AND2_X1   g041(.A1(new_n221), .A2(new_n227), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n221), .A2(new_n227), .ZN(new_n229));
  NOR2_X1   g043(.A1(new_n228), .A2(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(new_n212), .A2(KEYINPUT11), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n231), .A2(new_n210), .A3(new_n207), .A4(new_n201), .ZN(new_n232));
  NOR2_X1   g046(.A1(new_n195), .A2(KEYINPUT1), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n233), .A2(new_n189), .A3(new_n191), .ZN(new_n234));
  OAI211_X1 g048(.A(new_n190), .B(G146), .C1(new_n195), .C2(KEYINPUT1), .ZN(new_n235));
  NAND3_X1  g049(.A1(new_n195), .A2(new_n188), .A3(G143), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n234), .A2(new_n235), .A3(new_n236), .ZN(new_n237));
  NOR2_X1   g051(.A1(new_n200), .A2(G137), .ZN(new_n238));
  OAI21_X1  g052(.A(G131), .B1(new_n238), .B2(new_n211), .ZN(new_n239));
  NAND3_X1  g053(.A1(new_n232), .A2(new_n237), .A3(new_n239), .ZN(new_n240));
  NAND3_X1  g054(.A1(new_n215), .A2(new_n230), .A3(new_n240), .ZN(new_n241));
  NAND2_X1  g055(.A1(new_n241), .A2(KEYINPUT67), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT67), .ZN(new_n243));
  NAND4_X1  g057(.A1(new_n215), .A2(new_n230), .A3(new_n243), .A4(new_n240), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT26), .B(G101), .ZN(new_n245));
  NOR2_X1   g059(.A1(G237), .A2(G953), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n246), .A2(G210), .ZN(new_n247));
  XNOR2_X1  g061(.A(new_n245), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g062(.A(KEYINPUT68), .B(KEYINPUT27), .ZN(new_n249));
  XOR2_X1   g063(.A(new_n248), .B(new_n249), .Z(new_n250));
  NAND3_X1  g064(.A1(new_n242), .A2(new_n244), .A3(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(KEYINPUT69), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n251), .A2(new_n252), .ZN(new_n253));
  NAND4_X1  g067(.A1(new_n242), .A2(KEYINPUT69), .A3(new_n244), .A4(new_n250), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT30), .ZN(new_n255));
  OAI21_X1  g069(.A(G131), .B1(new_n205), .B2(new_n208), .ZN(new_n256));
  AOI22_X1  g070(.A1(new_n256), .A2(new_n232), .B1(new_n197), .B2(new_n198), .ZN(new_n257));
  INV_X1    g071(.A(new_n240), .ZN(new_n258));
  OAI21_X1  g072(.A(new_n255), .B1(new_n257), .B2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n215), .A2(KEYINPUT30), .A3(new_n240), .ZN(new_n260));
  XNOR2_X1  g074(.A(new_n221), .B(new_n227), .ZN(new_n261));
  AND3_X1   g075(.A1(new_n259), .A2(new_n260), .A3(new_n261), .ZN(new_n262));
  INV_X1    g076(.A(new_n262), .ZN(new_n263));
  NAND3_X1  g077(.A1(new_n253), .A2(new_n254), .A3(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT31), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n262), .B1(new_n251), .B2(new_n252), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT31), .A3(new_n254), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n266), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g083(.A1(new_n215), .A2(new_n240), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n270), .A2(new_n261), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n242), .A2(new_n271), .A3(new_n244), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(KEYINPUT28), .ZN(new_n273));
  INV_X1    g087(.A(new_n241), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n274), .A2(KEYINPUT28), .ZN(new_n275));
  INV_X1    g089(.A(new_n275), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n250), .B1(new_n273), .B2(new_n276), .ZN(new_n277));
  INV_X1    g091(.A(new_n277), .ZN(new_n278));
  AOI21_X1  g092(.A(KEYINPUT70), .B1(new_n269), .B2(new_n278), .ZN(new_n279));
  INV_X1    g093(.A(KEYINPUT70), .ZN(new_n280));
  AOI211_X1 g094(.A(new_n280), .B(new_n277), .C1(new_n266), .C2(new_n268), .ZN(new_n281));
  OAI21_X1  g095(.A(new_n187), .B1(new_n279), .B2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(KEYINPUT71), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n282), .A2(new_n283), .ZN(new_n284));
  INV_X1    g098(.A(KEYINPUT32), .ZN(new_n285));
  AND4_X1   g099(.A1(KEYINPUT31), .A2(new_n253), .A3(new_n254), .A4(new_n263), .ZN(new_n286));
  AOI21_X1  g100(.A(KEYINPUT31), .B1(new_n267), .B2(new_n254), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n278), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  NAND2_X1  g102(.A1(new_n288), .A2(new_n280), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n269), .A2(KEYINPUT70), .A3(new_n278), .ZN(new_n290));
  NAND2_X1  g104(.A1(new_n289), .A2(new_n290), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n291), .A2(KEYINPUT71), .A3(new_n187), .ZN(new_n292));
  NAND3_X1  g106(.A1(new_n284), .A2(new_n285), .A3(new_n292), .ZN(new_n293));
  INV_X1    g107(.A(new_n187), .ZN(new_n294));
  AOI21_X1  g108(.A(new_n294), .B1(new_n289), .B2(new_n290), .ZN(new_n295));
  NAND4_X1  g109(.A1(new_n273), .A2(new_n276), .A3(KEYINPUT29), .A4(new_n250), .ZN(new_n296));
  INV_X1    g110(.A(KEYINPUT72), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  INV_X1    g112(.A(G902), .ZN(new_n299));
  AOI21_X1  g113(.A(new_n275), .B1(new_n272), .B2(KEYINPUT28), .ZN(new_n300));
  NAND4_X1  g114(.A1(new_n300), .A2(KEYINPUT72), .A3(KEYINPUT29), .A4(new_n250), .ZN(new_n301));
  NAND3_X1  g115(.A1(new_n298), .A2(new_n299), .A3(new_n301), .ZN(new_n302));
  INV_X1    g116(.A(KEYINPUT73), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n302), .A2(new_n303), .ZN(new_n304));
  NAND4_X1  g118(.A1(new_n298), .A2(KEYINPUT73), .A3(new_n301), .A4(new_n299), .ZN(new_n305));
  NAND3_X1  g119(.A1(new_n263), .A2(new_n242), .A3(new_n244), .ZN(new_n306));
  INV_X1    g120(.A(new_n250), .ZN(new_n307));
  NAND2_X1  g121(.A1(new_n306), .A2(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT29), .ZN(new_n309));
  INV_X1    g123(.A(new_n300), .ZN(new_n310));
  OAI211_X1 g124(.A(new_n308), .B(new_n309), .C1(new_n310), .C2(new_n307), .ZN(new_n311));
  NAND3_X1  g125(.A1(new_n304), .A2(new_n305), .A3(new_n311), .ZN(new_n312));
  AOI22_X1  g126(.A1(new_n295), .A2(KEYINPUT32), .B1(new_n312), .B2(G472), .ZN(new_n313));
  NAND2_X1  g127(.A1(new_n293), .A2(new_n313), .ZN(new_n314));
  INV_X1    g128(.A(G140), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n315), .A2(G125), .ZN(new_n316));
  NOR2_X1   g130(.A1(new_n316), .A2(KEYINPUT16), .ZN(new_n317));
  INV_X1    g131(.A(new_n317), .ZN(new_n318));
  NOR3_X1   g132(.A1(new_n315), .A2(KEYINPUT75), .A3(G125), .ZN(new_n319));
  XNOR2_X1  g133(.A(G125), .B(G140), .ZN(new_n320));
  AOI21_X1  g134(.A(new_n319), .B1(new_n320), .B2(KEYINPUT75), .ZN(new_n321));
  INV_X1    g135(.A(KEYINPUT16), .ZN(new_n322));
  OAI211_X1 g136(.A(G146), .B(new_n318), .C1(new_n321), .C2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n320), .A2(new_n188), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT23), .ZN(new_n325));
  OAI21_X1  g139(.A(new_n325), .B1(new_n216), .B2(G128), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n216), .A2(G128), .ZN(new_n327));
  NAND3_X1  g141(.A1(new_n195), .A2(KEYINPUT23), .A3(G119), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n326), .A2(new_n327), .A3(new_n328), .ZN(new_n329));
  NOR2_X1   g143(.A1(new_n329), .A2(G110), .ZN(new_n330));
  NAND2_X1  g144(.A1(new_n195), .A2(G119), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n331), .A2(new_n327), .ZN(new_n332));
  XNOR2_X1  g146(.A(KEYINPUT24), .B(G110), .ZN(new_n333));
  AND2_X1   g147(.A1(new_n332), .A2(new_n333), .ZN(new_n334));
  OAI211_X1 g148(.A(new_n323), .B(new_n324), .C1(new_n330), .C2(new_n334), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n329), .A2(G110), .ZN(new_n336));
  OAI21_X1  g150(.A(new_n336), .B1(new_n332), .B2(new_n333), .ZN(new_n337));
  INV_X1    g151(.A(G125), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(G140), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n339), .A2(new_n316), .A3(KEYINPUT75), .ZN(new_n340));
  OR3_X1    g154(.A1(new_n315), .A2(KEYINPUT75), .A3(G125), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n322), .B1(new_n340), .B2(new_n341), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n188), .B1(new_n342), .B2(new_n317), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n337), .B1(new_n343), .B2(new_n323), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n345));
  NOR2_X1   g159(.A1(new_n344), .A2(new_n345), .ZN(new_n346));
  AOI211_X1 g160(.A(KEYINPUT76), .B(new_n337), .C1(new_n343), .C2(new_n323), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n335), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  XNOR2_X1  g162(.A(KEYINPUT22), .B(G137), .ZN(new_n349));
  XNOR2_X1  g163(.A(new_n349), .B(KEYINPUT77), .ZN(new_n350));
  INV_X1    g164(.A(G221), .ZN(new_n351));
  INV_X1    g165(.A(G234), .ZN(new_n352));
  NOR3_X1   g166(.A1(new_n351), .A2(new_n352), .A3(G953), .ZN(new_n353));
  XOR2_X1   g167(.A(new_n350), .B(new_n353), .Z(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n348), .A2(new_n355), .ZN(new_n356));
  OAI211_X1 g170(.A(new_n335), .B(new_n354), .C1(new_n346), .C2(new_n347), .ZN(new_n357));
  NAND2_X1  g171(.A1(new_n356), .A2(new_n357), .ZN(new_n358));
  AOI21_X1  g172(.A(G902), .B1(new_n352), .B2(G217), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  OAI21_X1  g174(.A(G217), .B1(new_n352), .B2(G902), .ZN(new_n361));
  XOR2_X1   g175(.A(new_n361), .B(KEYINPUT74), .Z(new_n362));
  INV_X1    g176(.A(new_n362), .ZN(new_n363));
  AOI21_X1  g177(.A(G902), .B1(new_n356), .B2(new_n357), .ZN(new_n364));
  INV_X1    g178(.A(KEYINPUT25), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n363), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  AOI211_X1 g180(.A(KEYINPUT25), .B(G902), .C1(new_n356), .C2(new_n357), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n360), .B1(new_n366), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(KEYINPUT78), .ZN(new_n369));
  INV_X1    g183(.A(KEYINPUT78), .ZN(new_n370));
  OAI211_X1 g184(.A(new_n360), .B(new_n370), .C1(new_n366), .C2(new_n367), .ZN(new_n371));
  NAND2_X1  g185(.A1(new_n369), .A2(new_n371), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  XNOR2_X1  g187(.A(KEYINPUT9), .B(G234), .ZN(new_n374));
  INV_X1    g188(.A(new_n374), .ZN(new_n375));
  AOI21_X1  g189(.A(new_n351), .B1(new_n375), .B2(new_n299), .ZN(new_n376));
  INV_X1    g190(.A(KEYINPUT10), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n235), .A2(new_n236), .ZN(new_n378));
  INV_X1    g192(.A(KEYINPUT81), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n235), .A2(KEYINPUT81), .A3(new_n236), .ZN(new_n381));
  AND3_X1   g195(.A1(new_n380), .A2(new_n234), .A3(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT80), .ZN(new_n383));
  INV_X1    g197(.A(G107), .ZN(new_n384));
  OAI21_X1  g198(.A(new_n383), .B1(new_n384), .B2(G104), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(G104), .ZN(new_n386));
  INV_X1    g200(.A(G104), .ZN(new_n387));
  NAND3_X1  g201(.A1(new_n387), .A2(KEYINPUT80), .A3(G107), .ZN(new_n388));
  NAND3_X1  g202(.A1(new_n385), .A2(new_n386), .A3(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G101), .ZN(new_n390));
  XNOR2_X1  g204(.A(KEYINPUT79), .B(G101), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n386), .A2(KEYINPUT3), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n387), .A2(G107), .ZN(new_n393));
  INV_X1    g207(.A(KEYINPUT3), .ZN(new_n394));
  NAND3_X1  g208(.A1(new_n394), .A2(new_n384), .A3(G104), .ZN(new_n395));
  NAND4_X1  g209(.A1(new_n391), .A2(new_n392), .A3(new_n393), .A4(new_n395), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n390), .A2(new_n396), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n377), .B1(new_n382), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n392), .A2(new_n395), .A3(new_n393), .ZN(new_n399));
  NAND2_X1  g213(.A1(new_n399), .A2(G101), .ZN(new_n400));
  NAND3_X1  g214(.A1(new_n400), .A2(KEYINPUT4), .A3(new_n396), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT4), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n399), .A2(new_n402), .A3(G101), .ZN(new_n403));
  NAND3_X1  g217(.A1(new_n401), .A2(new_n199), .A3(new_n403), .ZN(new_n404));
  INV_X1    g218(.A(new_n237), .ZN(new_n405));
  NOR2_X1   g219(.A1(new_n405), .A2(new_n377), .ZN(new_n406));
  AND2_X1   g220(.A1(new_n390), .A2(new_n396), .ZN(new_n407));
  NAND2_X1  g221(.A1(new_n406), .A2(new_n407), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n209), .A2(new_n214), .ZN(new_n409));
  NAND4_X1  g223(.A1(new_n398), .A2(new_n404), .A3(new_n408), .A4(new_n409), .ZN(new_n410));
  XNOR2_X1  g224(.A(G110), .B(G140), .ZN(new_n411));
  INV_X1    g225(.A(G227), .ZN(new_n412));
  NOR2_X1   g226(.A1(new_n412), .A2(G953), .ZN(new_n413));
  XNOR2_X1  g227(.A(new_n411), .B(new_n413), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  AND2_X1   g229(.A1(new_n410), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n380), .A2(new_n234), .A3(new_n381), .ZN(new_n417));
  NAND2_X1  g231(.A1(new_n407), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g232(.A1(new_n397), .A2(new_n405), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n418), .A2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n409), .ZN(new_n421));
  NAND4_X1  g235(.A1(new_n420), .A2(KEYINPUT82), .A3(KEYINPUT12), .A4(new_n421), .ZN(new_n422));
  INV_X1    g236(.A(KEYINPUT12), .ZN(new_n423));
  AOI21_X1  g237(.A(new_n237), .B1(new_n396), .B2(new_n390), .ZN(new_n424));
  AOI21_X1  g238(.A(new_n424), .B1(new_n407), .B2(new_n417), .ZN(new_n425));
  OAI21_X1  g239(.A(new_n423), .B1(new_n425), .B2(new_n409), .ZN(new_n426));
  NAND2_X1  g240(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n409), .B1(new_n418), .B2(new_n419), .ZN(new_n428));
  AOI21_X1  g242(.A(KEYINPUT82), .B1(new_n428), .B2(KEYINPUT12), .ZN(new_n429));
  OAI21_X1  g243(.A(new_n416), .B1(new_n427), .B2(new_n429), .ZN(new_n430));
  NAND3_X1  g244(.A1(new_n398), .A2(new_n404), .A3(new_n408), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(new_n421), .ZN(new_n432));
  NAND2_X1  g246(.A1(new_n432), .A2(new_n410), .ZN(new_n433));
  NAND2_X1  g247(.A1(new_n433), .A2(new_n414), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n430), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G469), .ZN(new_n436));
  NAND3_X1  g250(.A1(new_n435), .A2(new_n436), .A3(new_n299), .ZN(new_n437));
  INV_X1    g251(.A(KEYINPUT83), .ZN(new_n438));
  NAND2_X1  g252(.A1(new_n437), .A2(new_n438), .ZN(new_n439));
  AOI21_X1  g253(.A(G902), .B1(new_n430), .B2(new_n434), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n440), .A2(KEYINPUT83), .A3(new_n436), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n439), .A2(new_n441), .ZN(new_n442));
  AND3_X1   g256(.A1(new_n432), .A2(new_n410), .A3(new_n415), .ZN(new_n443));
  NAND3_X1  g257(.A1(new_n420), .A2(KEYINPUT12), .A3(new_n421), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT82), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g260(.A1(new_n446), .A2(new_n426), .A3(new_n422), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n447), .A2(new_n410), .ZN(new_n448));
  AOI21_X1  g262(.A(new_n443), .B1(new_n448), .B2(new_n414), .ZN(new_n449));
  OAI21_X1  g263(.A(G469), .B1(new_n449), .B2(G902), .ZN(new_n450));
  AOI21_X1  g264(.A(new_n376), .B1(new_n442), .B2(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  OAI21_X1  g266(.A(G214), .B1(G237), .B2(G902), .ZN(new_n453));
  XNOR2_X1  g267(.A(new_n453), .B(KEYINPUT84), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n199), .A2(G125), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n237), .A2(new_n338), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  XNOR2_X1  g271(.A(new_n457), .B(KEYINPUT86), .ZN(new_n458));
  INV_X1    g272(.A(G953), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n459), .A2(G224), .ZN(new_n460));
  XNOR2_X1  g274(.A(new_n458), .B(new_n460), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n261), .A2(new_n401), .A3(new_n403), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n462), .A2(KEYINPUT85), .ZN(new_n463));
  INV_X1    g277(.A(KEYINPUT85), .ZN(new_n464));
  NAND4_X1  g278(.A1(new_n261), .A2(new_n401), .A3(new_n464), .A4(new_n403), .ZN(new_n465));
  NAND2_X1  g279(.A1(new_n221), .A2(KEYINPUT5), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n216), .A2(G116), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n466), .B(G113), .C1(KEYINPUT5), .C2(new_n467), .ZN(new_n468));
  INV_X1    g282(.A(new_n228), .ZN(new_n469));
  NAND3_X1  g283(.A1(new_n468), .A2(new_n469), .A3(new_n407), .ZN(new_n470));
  NAND3_X1  g284(.A1(new_n463), .A2(new_n465), .A3(new_n470), .ZN(new_n471));
  XNOR2_X1  g285(.A(G110), .B(G122), .ZN(new_n472));
  INV_X1    g286(.A(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n471), .A2(new_n473), .ZN(new_n474));
  NAND4_X1  g288(.A1(new_n463), .A2(new_n472), .A3(new_n465), .A4(new_n470), .ZN(new_n475));
  NAND3_X1  g289(.A1(new_n474), .A2(KEYINPUT6), .A3(new_n475), .ZN(new_n476));
  INV_X1    g290(.A(KEYINPUT6), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n471), .A2(new_n477), .A3(new_n473), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n461), .A2(new_n476), .A3(new_n478), .ZN(new_n479));
  AND2_X1   g293(.A1(new_n460), .A2(KEYINPUT7), .ZN(new_n480));
  XNOR2_X1  g294(.A(new_n457), .B(new_n480), .ZN(new_n481));
  NAND2_X1  g295(.A1(new_n470), .A2(KEYINPUT87), .ZN(new_n482));
  INV_X1    g296(.A(KEYINPUT87), .ZN(new_n483));
  NAND4_X1  g297(.A1(new_n468), .A2(new_n483), .A3(new_n469), .A4(new_n407), .ZN(new_n484));
  AND2_X1   g298(.A1(new_n468), .A2(new_n469), .ZN(new_n485));
  OAI211_X1 g299(.A(new_n482), .B(new_n484), .C1(new_n407), .C2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n472), .B(KEYINPUT8), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n481), .B1(new_n486), .B2(new_n487), .ZN(new_n488));
  AOI21_X1  g302(.A(G902), .B1(new_n488), .B2(new_n475), .ZN(new_n489));
  OAI21_X1  g303(.A(G210), .B1(G237), .B2(G902), .ZN(new_n490));
  INV_X1    g304(.A(new_n490), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT88), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n479), .A2(new_n489), .A3(new_n493), .ZN(new_n494));
  AOI21_X1  g308(.A(new_n493), .B1(new_n479), .B2(new_n489), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(G475), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n299), .ZN(new_n498));
  XNOR2_X1  g312(.A(new_n498), .B(KEYINPUT92), .ZN(new_n499));
  INV_X1    g313(.A(new_n499), .ZN(new_n500));
  NAND3_X1  g314(.A1(new_n246), .A2(G143), .A3(G214), .ZN(new_n501));
  INV_X1    g315(.A(new_n501), .ZN(new_n502));
  AOI21_X1  g316(.A(G143), .B1(new_n246), .B2(G214), .ZN(new_n503));
  OAI211_X1 g317(.A(KEYINPUT17), .B(G131), .C1(new_n502), .C2(new_n503), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT91), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  INV_X1    g320(.A(G237), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n507), .A2(new_n459), .A3(G214), .ZN(new_n508));
  NAND2_X1  g322(.A1(new_n508), .A2(new_n190), .ZN(new_n509));
  AOI21_X1  g323(.A(new_n210), .B1(new_n509), .B2(new_n501), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n510), .A2(KEYINPUT91), .A3(KEYINPUT17), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n506), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(new_n510), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT17), .ZN(new_n514));
  NAND3_X1  g328(.A1(new_n509), .A2(new_n210), .A3(new_n501), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n513), .A2(new_n514), .A3(new_n515), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n512), .A2(new_n516), .A3(new_n343), .A4(new_n323), .ZN(new_n517));
  XNOR2_X1  g331(.A(G113), .B(G122), .ZN(new_n518));
  XNOR2_X1  g332(.A(new_n518), .B(new_n387), .ZN(new_n519));
  INV_X1    g333(.A(KEYINPUT89), .ZN(new_n520));
  NAND2_X1  g334(.A1(new_n340), .A2(new_n341), .ZN(new_n521));
  OAI21_X1  g335(.A(new_n520), .B1(new_n521), .B2(new_n188), .ZN(new_n522));
  NAND3_X1  g336(.A1(new_n321), .A2(KEYINPUT89), .A3(G146), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n522), .A2(new_n523), .A3(new_n324), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT18), .ZN(new_n525));
  OAI211_X1 g339(.A(new_n509), .B(new_n501), .C1(new_n525), .C2(new_n210), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT90), .ZN(new_n527));
  OR2_X1    g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NAND2_X1  g342(.A1(new_n526), .A2(new_n527), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n510), .A2(KEYINPUT18), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n524), .A2(new_n528), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n517), .A2(new_n519), .A3(new_n531), .ZN(new_n532));
  AND2_X1   g346(.A1(new_n521), .A2(KEYINPUT19), .ZN(new_n533));
  NOR2_X1   g347(.A1(new_n320), .A2(KEYINPUT19), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n188), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n513), .A2(new_n515), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n535), .A2(new_n323), .A3(new_n536), .ZN(new_n537));
  AOI21_X1  g351(.A(new_n519), .B1(new_n537), .B2(new_n531), .ZN(new_n538));
  OAI21_X1  g352(.A(new_n500), .B1(new_n532), .B2(new_n538), .ZN(new_n539));
  NAND2_X1  g353(.A1(new_n539), .A2(KEYINPUT20), .ZN(new_n540));
  NAND2_X1  g354(.A1(new_n537), .A2(new_n531), .ZN(new_n541));
  INV_X1    g355(.A(new_n519), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  NAND3_X1  g357(.A1(new_n517), .A2(new_n531), .A3(new_n519), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(KEYINPUT20), .ZN(new_n546));
  NAND3_X1  g360(.A1(new_n545), .A2(new_n546), .A3(new_n500), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n540), .A2(new_n547), .ZN(new_n548));
  XNOR2_X1  g362(.A(G128), .B(G143), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n549), .A2(KEYINPUT13), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n190), .A2(G128), .ZN(new_n551));
  OAI211_X1 g365(.A(new_n550), .B(G134), .C1(KEYINPUT13), .C2(new_n551), .ZN(new_n552));
  XOR2_X1   g366(.A(G116), .B(G122), .Z(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(G107), .ZN(new_n554));
  XNOR2_X1  g368(.A(G116), .B(G122), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(new_n384), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n554), .A2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n549), .A2(new_n200), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n552), .A2(new_n557), .A3(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(new_n549), .B(new_n200), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n219), .A2(KEYINPUT14), .A3(G122), .ZN(new_n561));
  OAI211_X1 g375(.A(G107), .B(new_n561), .C1(new_n553), .C2(KEYINPUT14), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n560), .A2(new_n556), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  NAND3_X1  g378(.A1(new_n375), .A2(G217), .A3(new_n459), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT93), .ZN(new_n567));
  INV_X1    g381(.A(new_n565), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n559), .A2(new_n563), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n566), .A2(new_n567), .A3(new_n569), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n564), .A2(KEYINPUT93), .A3(new_n565), .ZN(new_n571));
  NAND3_X1  g385(.A1(new_n570), .A2(new_n299), .A3(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(G478), .ZN(new_n573));
  NOR2_X1   g387(.A1(new_n573), .A2(KEYINPUT15), .ZN(new_n574));
  INV_X1    g388(.A(new_n574), .ZN(new_n575));
  XNOR2_X1  g389(.A(new_n572), .B(new_n575), .ZN(new_n576));
  AND2_X1   g390(.A1(new_n459), .A2(G952), .ZN(new_n577));
  OAI21_X1  g391(.A(new_n577), .B1(new_n352), .B2(new_n507), .ZN(new_n578));
  INV_X1    g392(.A(new_n578), .ZN(new_n579));
  AOI211_X1 g393(.A(new_n299), .B(new_n459), .C1(G234), .C2(G237), .ZN(new_n580));
  XNOR2_X1  g394(.A(KEYINPUT21), .B(G898), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n579), .B1(new_n580), .B2(new_n581), .ZN(new_n582));
  INV_X1    g396(.A(new_n582), .ZN(new_n583));
  AOI21_X1  g397(.A(new_n519), .B1(new_n517), .B2(new_n531), .ZN(new_n584));
  OAI21_X1  g398(.A(new_n299), .B1(new_n532), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n585), .A2(G475), .ZN(new_n586));
  NAND4_X1  g400(.A1(new_n548), .A2(new_n576), .A3(new_n583), .A4(new_n586), .ZN(new_n587));
  NOR4_X1   g401(.A1(new_n452), .A2(new_n454), .A3(new_n496), .A4(new_n587), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n314), .A2(new_n373), .A3(new_n588), .ZN(new_n589));
  XNOR2_X1  g403(.A(new_n589), .B(KEYINPUT94), .ZN(new_n590));
  XNOR2_X1  g404(.A(new_n590), .B(new_n391), .ZN(G3));
  AOI22_X1  g405(.A1(new_n447), .A2(new_n416), .B1(new_n433), .B2(new_n414), .ZN(new_n592));
  NOR4_X1   g406(.A1(new_n592), .A2(new_n438), .A3(G469), .A4(G902), .ZN(new_n593));
  AOI21_X1  g407(.A(KEYINPUT83), .B1(new_n440), .B2(new_n436), .ZN(new_n594));
  OAI21_X1  g408(.A(new_n450), .B1(new_n593), .B2(new_n594), .ZN(new_n595));
  INV_X1    g409(.A(new_n376), .ZN(new_n596));
  NAND3_X1  g410(.A1(new_n595), .A2(new_n596), .A3(new_n583), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n597), .A2(new_n372), .ZN(new_n598));
  OAI21_X1  g412(.A(new_n299), .B1(new_n279), .B2(new_n281), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n599), .A2(G472), .ZN(new_n600));
  NAND4_X1  g414(.A1(new_n598), .A2(new_n284), .A3(new_n292), .A4(new_n600), .ZN(new_n601));
  NAND2_X1  g415(.A1(new_n479), .A2(new_n489), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n602), .A2(new_n490), .ZN(new_n603));
  INV_X1    g417(.A(new_n454), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n479), .A2(new_n489), .A3(new_n491), .ZN(new_n605));
  NAND3_X1  g419(.A1(new_n603), .A2(new_n604), .A3(new_n605), .ZN(new_n606));
  INV_X1    g420(.A(new_n606), .ZN(new_n607));
  NOR2_X1   g421(.A1(new_n539), .A2(KEYINPUT20), .ZN(new_n608));
  AOI21_X1  g422(.A(new_n546), .B1(new_n545), .B2(new_n500), .ZN(new_n609));
  OAI21_X1  g423(.A(new_n586), .B1(new_n608), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n610), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT95), .B(KEYINPUT33), .Z(new_n612));
  INV_X1    g426(.A(new_n612), .ZN(new_n613));
  NAND3_X1  g427(.A1(new_n570), .A2(new_n571), .A3(new_n613), .ZN(new_n614));
  NAND3_X1  g428(.A1(new_n566), .A2(KEYINPUT33), .A3(new_n569), .ZN(new_n615));
  NAND4_X1  g429(.A1(new_n614), .A2(G478), .A3(new_n299), .A4(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n572), .A2(new_n573), .ZN(new_n617));
  NAND2_X1  g431(.A1(new_n616), .A2(new_n617), .ZN(new_n618));
  INV_X1    g432(.A(new_n618), .ZN(new_n619));
  NOR2_X1   g433(.A1(new_n611), .A2(new_n619), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n607), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n601), .A2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT34), .B(G104), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G6));
  INV_X1    g438(.A(new_n576), .ZN(new_n625));
  NAND2_X1  g439(.A1(new_n611), .A2(new_n625), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NAND2_X1  g441(.A1(new_n607), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n601), .A2(new_n628), .ZN(new_n629));
  XNOR2_X1  g443(.A(KEYINPUT35), .B(G107), .ZN(new_n630));
  XNOR2_X1  g444(.A(new_n630), .B(KEYINPUT96), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n629), .B(new_n631), .ZN(G9));
  INV_X1    g446(.A(new_n495), .ZN(new_n633));
  NAND3_X1  g447(.A1(new_n479), .A2(new_n489), .A3(new_n493), .ZN(new_n634));
  AOI21_X1  g448(.A(new_n454), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n358), .A2(new_n299), .ZN(new_n636));
  NAND2_X1  g450(.A1(new_n636), .A2(KEYINPUT25), .ZN(new_n637));
  NAND2_X1  g451(.A1(new_n364), .A2(new_n365), .ZN(new_n638));
  NAND3_X1  g452(.A1(new_n637), .A2(new_n638), .A3(new_n363), .ZN(new_n639));
  NOR2_X1   g453(.A1(new_n354), .A2(KEYINPUT36), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n348), .B(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n359), .ZN(new_n642));
  AOI21_X1  g456(.A(new_n587), .B1(new_n639), .B2(new_n642), .ZN(new_n643));
  AND4_X1   g457(.A1(new_n635), .A2(new_n643), .A3(new_n596), .A4(new_n595), .ZN(new_n644));
  NAND4_X1  g458(.A1(new_n644), .A2(new_n284), .A3(new_n292), .A4(new_n600), .ZN(new_n645));
  XOR2_X1   g459(.A(KEYINPUT37), .B(G110), .Z(new_n646));
  XNOR2_X1  g460(.A(new_n645), .B(new_n646), .ZN(G12));
  AOI21_X1  g461(.A(new_n452), .B1(new_n293), .B2(new_n313), .ZN(new_n648));
  INV_X1    g462(.A(G900), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n580), .A2(new_n649), .ZN(new_n650));
  NAND2_X1  g464(.A1(new_n650), .A2(new_n578), .ZN(new_n651));
  INV_X1    g465(.A(new_n651), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n626), .A2(new_n652), .ZN(new_n653));
  INV_X1    g467(.A(new_n366), .ZN(new_n654));
  AOI22_X1  g468(.A1(new_n654), .A2(new_n638), .B1(new_n359), .B2(new_n641), .ZN(new_n655));
  NOR2_X1   g469(.A1(new_n606), .A2(new_n655), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n648), .A2(new_n653), .A3(new_n656), .ZN(new_n657));
  XNOR2_X1  g471(.A(new_n657), .B(G128), .ZN(G30));
  NAND3_X1  g472(.A1(new_n291), .A2(KEYINPUT32), .A3(new_n187), .ZN(new_n659));
  INV_X1    g473(.A(new_n264), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n660), .B1(new_n272), .B2(new_n307), .ZN(new_n661));
  OAI21_X1  g475(.A(G472), .B1(new_n661), .B2(G902), .ZN(new_n662));
  AND2_X1   g476(.A1(new_n659), .A2(new_n662), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n293), .ZN(new_n664));
  INV_X1    g478(.A(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n651), .B(KEYINPUT39), .ZN(new_n666));
  NAND2_X1  g480(.A1(new_n451), .A2(new_n666), .ZN(new_n667));
  XNOR2_X1  g481(.A(new_n667), .B(KEYINPUT40), .ZN(new_n668));
  XNOR2_X1  g482(.A(new_n496), .B(KEYINPUT38), .ZN(new_n669));
  NOR3_X1   g483(.A1(new_n611), .A2(new_n454), .A3(new_n576), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n655), .ZN(new_n671));
  OR4_X1    g485(.A1(new_n665), .A2(new_n668), .A3(new_n669), .A4(new_n671), .ZN(new_n672));
  XNOR2_X1  g486(.A(new_n672), .B(G143), .ZN(G45));
  NAND4_X1  g487(.A1(new_n656), .A2(new_n451), .A3(new_n620), .A4(new_n651), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n674), .B1(new_n293), .B2(new_n313), .ZN(new_n675));
  INV_X1    g489(.A(KEYINPUT97), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n675), .B(new_n676), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G146), .ZN(G48));
  AOI21_X1  g492(.A(new_n372), .B1(new_n293), .B2(new_n313), .ZN(new_n679));
  OAI21_X1  g493(.A(G469), .B1(new_n592), .B2(G902), .ZN(new_n680));
  NAND3_X1  g494(.A1(new_n442), .A2(new_n596), .A3(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(new_n681), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n583), .ZN(new_n683));
  NOR2_X1   g497(.A1(new_n683), .A2(new_n621), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n679), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n685), .B(KEYINPUT41), .ZN(new_n686));
  XNOR2_X1  g500(.A(new_n686), .B(G113), .ZN(G15));
  NOR2_X1   g501(.A1(new_n683), .A2(new_n628), .ZN(new_n688));
  NAND3_X1  g502(.A1(new_n314), .A2(new_n373), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g503(.A(new_n689), .B(G116), .ZN(G18));
  NOR4_X1   g504(.A1(new_n681), .A2(new_n606), .A3(new_n655), .A4(new_n587), .ZN(new_n691));
  NAND2_X1  g505(.A1(new_n314), .A2(new_n691), .ZN(new_n692));
  XNOR2_X1  g506(.A(new_n692), .B(G119), .ZN(G21));
  OR2_X1    g507(.A1(new_n300), .A2(KEYINPUT98), .ZN(new_n694));
  NAND2_X1  g508(.A1(new_n300), .A2(KEYINPUT98), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n694), .A2(new_n307), .A3(new_n695), .ZN(new_n696));
  AOI21_X1  g510(.A(new_n294), .B1(new_n696), .B2(new_n269), .ZN(new_n697));
  AOI21_X1  g511(.A(G902), .B1(new_n289), .B2(new_n290), .ZN(new_n698));
  INV_X1    g512(.A(G472), .ZN(new_n699));
  OAI21_X1  g513(.A(KEYINPUT99), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  INV_X1    g514(.A(KEYINPUT99), .ZN(new_n701));
  NAND3_X1  g515(.A1(new_n599), .A2(new_n701), .A3(G472), .ZN(new_n702));
  AOI21_X1  g516(.A(new_n697), .B1(new_n700), .B2(new_n702), .ZN(new_n703));
  NAND3_X1  g517(.A1(new_n670), .A2(new_n603), .A3(new_n605), .ZN(new_n704));
  NOR2_X1   g518(.A1(new_n683), .A2(new_n704), .ZN(new_n705));
  INV_X1    g519(.A(new_n368), .ZN(new_n706));
  NAND3_X1  g520(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(new_n707));
  XNOR2_X1  g521(.A(new_n707), .B(KEYINPUT100), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NAND2_X1  g523(.A1(new_n700), .A2(new_n702), .ZN(new_n710));
  INV_X1    g524(.A(new_n655), .ZN(new_n711));
  INV_X1    g525(.A(new_n697), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n610), .A2(new_n618), .A3(new_n651), .ZN(new_n713));
  NOR3_X1   g527(.A1(new_n681), .A2(new_n606), .A3(new_n713), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n715), .B(KEYINPUT101), .ZN(new_n716));
  XNOR2_X1  g530(.A(new_n716), .B(new_n338), .ZN(G27));
  AOI21_X1  g531(.A(new_n376), .B1(new_n595), .B2(KEYINPUT102), .ZN(new_n718));
  NOR4_X1   g532(.A1(new_n713), .A2(new_n494), .A3(new_n495), .A4(new_n454), .ZN(new_n719));
  INV_X1    g533(.A(KEYINPUT102), .ZN(new_n720));
  NAND3_X1  g534(.A1(new_n442), .A2(new_n720), .A3(new_n450), .ZN(new_n721));
  NAND3_X1  g535(.A1(new_n718), .A2(new_n719), .A3(new_n721), .ZN(new_n722));
  INV_X1    g536(.A(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT42), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n312), .A2(G472), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n659), .A2(new_n725), .ZN(new_n726));
  NOR2_X1   g540(.A1(new_n295), .A2(KEYINPUT32), .ZN(new_n727));
  OAI21_X1  g541(.A(new_n706), .B1(new_n726), .B2(new_n727), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n728), .A2(KEYINPUT104), .ZN(new_n729));
  INV_X1    g543(.A(KEYINPUT104), .ZN(new_n730));
  OAI211_X1 g544(.A(new_n730), .B(new_n706), .C1(new_n726), .C2(new_n727), .ZN(new_n731));
  AOI21_X1  g545(.A(new_n724), .B1(new_n729), .B2(new_n731), .ZN(new_n732));
  INV_X1    g546(.A(new_n732), .ZN(new_n733));
  INV_X1    g547(.A(KEYINPUT103), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n679), .A2(new_n723), .ZN(new_n735));
  INV_X1    g549(.A(KEYINPUT42), .ZN(new_n736));
  AOI21_X1  g550(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  AOI211_X1 g551(.A(KEYINPUT103), .B(KEYINPUT42), .C1(new_n679), .C2(new_n723), .ZN(new_n738));
  OAI21_X1  g552(.A(new_n733), .B1(new_n737), .B2(new_n738), .ZN(new_n739));
  INV_X1    g553(.A(KEYINPUT105), .ZN(new_n740));
  NAND2_X1  g554(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  OAI211_X1 g555(.A(new_n733), .B(KEYINPUT105), .C1(new_n737), .C2(new_n738), .ZN(new_n742));
  AND2_X1   g556(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G131), .ZN(G33));
  NAND2_X1  g558(.A1(new_n496), .A2(new_n604), .ZN(new_n745));
  INV_X1    g559(.A(new_n745), .ZN(new_n746));
  AND4_X1   g560(.A1(new_n653), .A2(new_n746), .A3(new_n718), .A4(new_n721), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n679), .A2(new_n747), .ZN(new_n748));
  XNOR2_X1  g562(.A(new_n748), .B(KEYINPUT106), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(G134), .ZN(G36));
  AND2_X1   g564(.A1(new_n449), .A2(KEYINPUT45), .ZN(new_n751));
  OAI21_X1  g565(.A(G469), .B1(new_n449), .B2(KEYINPUT45), .ZN(new_n752));
  OR2_X1    g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g567(.A1(G469), .A2(G902), .ZN(new_n754));
  AOI21_X1  g568(.A(KEYINPUT46), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  AOI21_X1  g569(.A(new_n755), .B1(new_n439), .B2(new_n441), .ZN(new_n756));
  NAND3_X1  g570(.A1(new_n753), .A2(KEYINPUT46), .A3(new_n754), .ZN(new_n757));
  NAND2_X1  g571(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND3_X1  g572(.A1(new_n758), .A2(new_n596), .A3(new_n666), .ZN(new_n759));
  XNOR2_X1  g573(.A(KEYINPUT107), .B(KEYINPUT43), .ZN(new_n760));
  INV_X1    g574(.A(KEYINPUT107), .ZN(new_n761));
  NOR2_X1   g575(.A1(new_n761), .A2(KEYINPUT43), .ZN(new_n762));
  NOR2_X1   g576(.A1(new_n610), .A2(new_n619), .ZN(new_n763));
  MUX2_X1   g577(.A(new_n760), .B(new_n762), .S(new_n763), .Z(new_n764));
  XNOR2_X1  g578(.A(new_n764), .B(KEYINPUT108), .ZN(new_n765));
  NOR2_X1   g579(.A1(new_n295), .A2(KEYINPUT71), .ZN(new_n766));
  AOI211_X1 g580(.A(new_n283), .B(new_n294), .C1(new_n289), .C2(new_n290), .ZN(new_n767));
  NOR2_X1   g581(.A1(new_n766), .A2(new_n767), .ZN(new_n768));
  AOI21_X1  g582(.A(new_n655), .B1(new_n768), .B2(new_n600), .ZN(new_n769));
  INV_X1    g583(.A(KEYINPUT109), .ZN(new_n770));
  AND2_X1   g584(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n769), .A2(new_n770), .ZN(new_n772));
  OAI21_X1  g586(.A(new_n765), .B1(new_n771), .B2(new_n772), .ZN(new_n773));
  INV_X1    g587(.A(KEYINPUT44), .ZN(new_n774));
  AOI211_X1 g588(.A(new_n745), .B(new_n759), .C1(new_n773), .C2(new_n774), .ZN(new_n775));
  OR2_X1    g589(.A1(new_n773), .A2(new_n774), .ZN(new_n776));
  NAND2_X1  g590(.A1(new_n775), .A2(new_n776), .ZN(new_n777));
  XNOR2_X1  g591(.A(new_n777), .B(KEYINPUT110), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G137), .ZN(G39));
  NAND2_X1  g593(.A1(new_n758), .A2(new_n596), .ZN(new_n780));
  XNOR2_X1  g594(.A(new_n780), .B(KEYINPUT47), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n719), .A2(new_n372), .ZN(new_n782));
  NOR3_X1   g596(.A1(new_n781), .A2(new_n314), .A3(new_n782), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(new_n315), .ZN(G42));
  AND4_X1   g598(.A1(new_n706), .A2(new_n763), .A3(new_n604), .A4(new_n596), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n442), .A2(new_n680), .ZN(new_n786));
  XOR2_X1   g600(.A(new_n786), .B(KEYINPUT49), .Z(new_n787));
  NAND4_X1  g601(.A1(new_n665), .A2(new_n669), .A3(new_n785), .A4(new_n787), .ZN(new_n788));
  AOI211_X1 g602(.A(new_n368), .B(new_n697), .C1(new_n700), .C2(new_n702), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  NOR3_X1   g604(.A1(new_n790), .A2(new_n578), .A3(new_n764), .ZN(new_n791));
  NAND4_X1  g605(.A1(new_n791), .A2(new_n454), .A3(new_n669), .A4(new_n682), .ZN(new_n792));
  XOR2_X1   g606(.A(new_n792), .B(KEYINPUT50), .Z(new_n793));
  NOR4_X1   g607(.A1(new_n764), .A2(new_n578), .A3(new_n681), .A4(new_n745), .ZN(new_n794));
  NAND3_X1  g608(.A1(new_n794), .A2(new_n711), .A3(new_n703), .ZN(new_n795));
  NOR3_X1   g609(.A1(new_n745), .A2(new_n681), .A3(new_n578), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n665), .A2(new_n373), .A3(new_n796), .ZN(new_n797));
  NAND2_X1  g611(.A1(new_n611), .A2(new_n619), .ZN(new_n798));
  OAI211_X1 g612(.A(new_n793), .B(new_n795), .C1(new_n797), .C2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n799), .A2(KEYINPUT117), .ZN(new_n800));
  OAI21_X1  g614(.A(new_n781), .B1(new_n596), .B2(new_n786), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n801), .A2(new_n746), .A3(new_n791), .ZN(new_n802));
  AOI21_X1  g616(.A(KEYINPUT51), .B1(new_n800), .B2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n635), .A2(new_n627), .ZN(new_n804));
  OAI21_X1  g618(.A(new_n645), .B1(new_n601), .B2(new_n804), .ZN(new_n805));
  INV_X1    g619(.A(KEYINPUT112), .ZN(new_n806));
  NAND2_X1  g620(.A1(new_n805), .A2(new_n806), .ZN(new_n807));
  INV_X1    g621(.A(new_n804), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n768), .A2(new_n600), .A3(new_n598), .A4(new_n808), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(KEYINPUT112), .A3(new_n645), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n635), .A2(new_n620), .ZN(new_n811));
  INV_X1    g625(.A(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n768), .A2(new_n812), .A3(new_n600), .A4(new_n598), .ZN(new_n813));
  NAND4_X1  g627(.A1(new_n807), .A2(new_n589), .A3(new_n810), .A4(new_n813), .ZN(new_n814));
  NOR4_X1   g628(.A1(new_n745), .A2(new_n625), .A3(new_n610), .A4(new_n652), .ZN(new_n815));
  AOI22_X1  g629(.A1(new_n648), .A2(new_n815), .B1(new_n703), .B2(new_n723), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n748), .B1(new_n816), .B2(new_n655), .ZN(new_n817));
  OAI21_X1  g631(.A(KEYINPUT115), .B1(new_n814), .B2(new_n817), .ZN(new_n818));
  AND3_X1   g632(.A1(new_n314), .A2(new_n373), .A3(new_n747), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n314), .A2(new_n451), .A3(new_n815), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n703), .A2(new_n723), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  AOI21_X1  g636(.A(new_n819), .B1(new_n822), .B2(new_n711), .ZN(new_n823));
  NAND2_X1  g637(.A1(new_n589), .A2(new_n813), .ZN(new_n824));
  AOI21_X1  g638(.A(KEYINPUT112), .B1(new_n809), .B2(new_n645), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n824), .A2(new_n825), .ZN(new_n826));
  INV_X1    g640(.A(KEYINPUT115), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n823), .A2(new_n826), .A3(new_n827), .A4(new_n810), .ZN(new_n828));
  AND3_X1   g642(.A1(new_n818), .A2(new_n828), .A3(KEYINPUT53), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT116), .ZN(new_n830));
  AOI211_X1 g644(.A(new_n372), .B(new_n722), .C1(new_n293), .C2(new_n313), .ZN(new_n831));
  OAI21_X1  g645(.A(KEYINPUT103), .B1(new_n831), .B2(KEYINPUT42), .ZN(new_n832));
  NAND3_X1  g646(.A1(new_n735), .A2(new_n734), .A3(new_n736), .ZN(new_n833));
  AOI21_X1  g647(.A(new_n732), .B1(new_n832), .B2(new_n833), .ZN(new_n834));
  NAND4_X1  g648(.A1(new_n685), .A2(new_n689), .A3(new_n692), .A4(new_n707), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n830), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  INV_X1    g650(.A(new_n835), .ZN(new_n837));
  NAND3_X1  g651(.A1(new_n739), .A2(KEYINPUT116), .A3(new_n837), .ZN(new_n838));
  NAND2_X1  g652(.A1(new_n836), .A2(new_n838), .ZN(new_n839));
  INV_X1    g653(.A(KEYINPUT52), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n718), .A2(new_n721), .ZN(new_n841));
  XOR2_X1   g655(.A(new_n651), .B(KEYINPUT113), .Z(new_n842));
  NOR4_X1   g656(.A1(new_n841), .A2(new_n711), .A3(new_n704), .A4(new_n842), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n843), .A2(new_n664), .ZN(new_n844));
  AOI211_X1 g658(.A(KEYINPUT97), .B(new_n674), .C1(new_n293), .C2(new_n313), .ZN(new_n845));
  INV_X1    g659(.A(new_n674), .ZN(new_n846));
  AOI21_X1  g660(.A(new_n676), .B1(new_n314), .B2(new_n846), .ZN(new_n847));
  OAI211_X1 g661(.A(new_n657), .B(new_n844), .C1(new_n845), .C2(new_n847), .ZN(new_n848));
  OAI21_X1  g662(.A(new_n840), .B1(new_n848), .B2(new_n716), .ZN(new_n849));
  INV_X1    g663(.A(KEYINPUT101), .ZN(new_n850));
  XNOR2_X1  g664(.A(new_n715), .B(new_n850), .ZN(new_n851));
  AOI21_X1  g665(.A(new_n840), .B1(new_n843), .B2(new_n664), .ZN(new_n852));
  NAND4_X1  g666(.A1(new_n851), .A2(new_n677), .A3(new_n852), .A4(new_n657), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT114), .B1(new_n849), .B2(new_n853), .ZN(new_n854));
  AND3_X1   g668(.A1(new_n849), .A2(KEYINPUT114), .A3(new_n853), .ZN(new_n855));
  OAI211_X1 g669(.A(new_n829), .B(new_n839), .C1(new_n854), .C2(new_n855), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT53), .ZN(new_n857));
  INV_X1    g671(.A(KEYINPUT111), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n835), .A2(new_n858), .ZN(new_n859));
  AOI22_X1  g673(.A1(new_n789), .A2(new_n705), .B1(new_n679), .B2(new_n688), .ZN(new_n860));
  AOI22_X1  g674(.A1(new_n679), .A2(new_n684), .B1(new_n314), .B2(new_n691), .ZN(new_n861));
  AOI21_X1  g675(.A(KEYINPUT111), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  NOR2_X1   g676(.A1(new_n859), .A2(new_n862), .ZN(new_n863));
  NOR2_X1   g677(.A1(new_n814), .A2(new_n817), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n741), .A2(new_n863), .A3(new_n742), .A4(new_n864), .ZN(new_n865));
  AND2_X1   g679(.A1(new_n657), .A2(new_n844), .ZN(new_n866));
  NAND4_X1  g680(.A1(new_n866), .A2(new_n851), .A3(KEYINPUT52), .A4(new_n677), .ZN(new_n867));
  AND2_X1   g681(.A1(new_n849), .A2(new_n867), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n857), .B1(new_n865), .B2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(KEYINPUT54), .ZN(new_n870));
  NAND3_X1  g684(.A1(new_n856), .A2(new_n869), .A3(new_n870), .ZN(new_n871));
  OAI21_X1  g685(.A(KEYINPUT53), .B1(new_n865), .B2(new_n868), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n743), .A2(new_n857), .A3(new_n863), .A4(new_n864), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n855), .A2(new_n854), .ZN(new_n874));
  OAI21_X1  g688(.A(new_n872), .B1(new_n873), .B2(new_n874), .ZN(new_n875));
  OAI21_X1  g689(.A(new_n871), .B1(new_n875), .B2(new_n870), .ZN(new_n876));
  NAND2_X1  g690(.A1(new_n729), .A2(new_n731), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n877), .A2(new_n794), .ZN(new_n878));
  XOR2_X1   g692(.A(new_n878), .B(KEYINPUT48), .Z(new_n879));
  NAND3_X1  g693(.A1(new_n791), .A2(new_n607), .A3(new_n682), .ZN(new_n880));
  INV_X1    g694(.A(new_n620), .ZN(new_n881));
  OAI211_X1 g695(.A(new_n880), .B(new_n577), .C1(new_n881), .C2(new_n797), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n879), .A2(new_n882), .ZN(new_n883));
  INV_X1    g697(.A(KEYINPUT51), .ZN(new_n884));
  NAND2_X1  g698(.A1(new_n884), .A2(KEYINPUT117), .ZN(new_n885));
  OAI21_X1  g699(.A(new_n885), .B1(new_n802), .B2(new_n884), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n883), .B1(new_n799), .B2(new_n886), .ZN(new_n887));
  NOR3_X1   g701(.A1(new_n803), .A2(new_n876), .A3(new_n887), .ZN(new_n888));
  NOR2_X1   g702(.A1(G952), .A2(G953), .ZN(new_n889));
  OAI21_X1  g703(.A(new_n788), .B1(new_n888), .B2(new_n889), .ZN(G75));
  AOI21_X1  g704(.A(new_n299), .B1(new_n856), .B2(new_n869), .ZN(new_n891));
  AND2_X1   g705(.A1(new_n891), .A2(G210), .ZN(new_n892));
  NOR2_X1   g706(.A1(new_n892), .A2(KEYINPUT56), .ZN(new_n893));
  NAND2_X1  g707(.A1(new_n476), .A2(new_n478), .ZN(new_n894));
  XNOR2_X1  g708(.A(new_n894), .B(new_n461), .ZN(new_n895));
  XNOR2_X1  g709(.A(new_n895), .B(KEYINPUT55), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n893), .A2(new_n896), .ZN(new_n897));
  NOR2_X1   g711(.A1(new_n459), .A2(G952), .ZN(new_n898));
  INV_X1    g712(.A(new_n898), .ZN(new_n899));
  XOR2_X1   g713(.A(KEYINPUT118), .B(KEYINPUT56), .Z(new_n900));
  NAND2_X1  g714(.A1(new_n896), .A2(new_n900), .ZN(new_n901));
  OAI21_X1  g715(.A(new_n899), .B1(new_n892), .B2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n897), .A2(new_n902), .ZN(G51));
  AOI211_X1 g717(.A(new_n299), .B(new_n753), .C1(new_n856), .C2(new_n869), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n754), .B(KEYINPUT57), .Z(new_n905));
  AND3_X1   g719(.A1(new_n856), .A2(new_n869), .A3(new_n870), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n870), .B1(new_n856), .B2(new_n869), .ZN(new_n907));
  OAI21_X1  g721(.A(new_n905), .B1(new_n906), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n904), .B1(new_n908), .B2(new_n435), .ZN(new_n909));
  OAI21_X1  g723(.A(KEYINPUT119), .B1(new_n909), .B2(new_n898), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT119), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n856), .A2(new_n869), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n912), .A2(KEYINPUT54), .ZN(new_n913));
  NAND2_X1  g727(.A1(new_n913), .A2(new_n871), .ZN(new_n914));
  AOI21_X1  g728(.A(new_n592), .B1(new_n914), .B2(new_n905), .ZN(new_n915));
  OAI211_X1 g729(.A(new_n911), .B(new_n899), .C1(new_n915), .C2(new_n904), .ZN(new_n916));
  NAND2_X1  g730(.A1(new_n910), .A2(new_n916), .ZN(G54));
  NAND3_X1  g731(.A1(new_n891), .A2(KEYINPUT58), .A3(G475), .ZN(new_n918));
  INV_X1    g732(.A(new_n545), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n920), .A2(new_n899), .ZN(new_n921));
  NOR2_X1   g735(.A1(new_n918), .A2(new_n919), .ZN(new_n922));
  OAI21_X1  g736(.A(KEYINPUT120), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  AOI21_X1  g737(.A(new_n898), .B1(new_n918), .B2(new_n919), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT120), .ZN(new_n925));
  OAI211_X1 g739(.A(new_n924), .B(new_n925), .C1(new_n919), .C2(new_n918), .ZN(new_n926));
  NAND2_X1  g740(.A1(new_n923), .A2(new_n926), .ZN(G60));
  NAND2_X1  g741(.A1(G478), .A2(G902), .ZN(new_n928));
  XOR2_X1   g742(.A(new_n928), .B(KEYINPUT59), .Z(new_n929));
  INV_X1    g743(.A(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n876), .A2(new_n930), .ZN(new_n931));
  AND2_X1   g745(.A1(new_n614), .A2(new_n615), .ZN(new_n932));
  INV_X1    g746(.A(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g748(.A(KEYINPUT121), .ZN(new_n935));
  OAI211_X1 g749(.A(new_n932), .B(new_n930), .C1(new_n906), .C2(new_n907), .ZN(new_n936));
  NAND4_X1  g750(.A1(new_n934), .A2(new_n935), .A3(new_n899), .A4(new_n936), .ZN(new_n937));
  NAND2_X1  g751(.A1(new_n936), .A2(new_n899), .ZN(new_n938));
  AOI21_X1  g752(.A(new_n932), .B1(new_n876), .B2(new_n930), .ZN(new_n939));
  OAI21_X1  g753(.A(KEYINPUT121), .B1(new_n938), .B2(new_n939), .ZN(new_n940));
  NAND2_X1  g754(.A1(new_n937), .A2(new_n940), .ZN(G63));
  NAND2_X1  g755(.A1(G217), .A2(G902), .ZN(new_n942));
  XNOR2_X1  g756(.A(new_n942), .B(KEYINPUT60), .ZN(new_n943));
  AOI21_X1  g757(.A(new_n943), .B1(new_n856), .B2(new_n869), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n898), .B1(new_n944), .B2(new_n641), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n945), .B1(new_n358), .B2(new_n944), .ZN(new_n946));
  AOI21_X1  g760(.A(KEYINPUT122), .B1(new_n944), .B2(new_n641), .ZN(new_n947));
  NOR2_X1   g761(.A1(new_n947), .A2(KEYINPUT61), .ZN(new_n948));
  XNOR2_X1  g762(.A(new_n946), .B(new_n948), .ZN(G66));
  NAND3_X1  g763(.A1(new_n863), .A2(new_n810), .A3(new_n826), .ZN(new_n950));
  XNOR2_X1  g764(.A(new_n950), .B(KEYINPUT123), .ZN(new_n951));
  INV_X1    g765(.A(new_n951), .ZN(new_n952));
  NAND2_X1  g766(.A1(G224), .A2(G953), .ZN(new_n953));
  OAI22_X1  g767(.A1(new_n952), .A2(G953), .B1(new_n581), .B2(new_n953), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n894), .B1(G898), .B2(new_n459), .ZN(new_n955));
  XOR2_X1   g769(.A(new_n954), .B(new_n955), .Z(G69));
  NAND2_X1  g770(.A1(new_n259), .A2(new_n260), .ZN(new_n957));
  XNOR2_X1  g771(.A(new_n957), .B(KEYINPUT124), .ZN(new_n958));
  NOR2_X1   g772(.A1(new_n533), .A2(new_n534), .ZN(new_n959));
  XNOR2_X1  g773(.A(new_n958), .B(new_n959), .ZN(new_n960));
  AND3_X1   g774(.A1(new_n851), .A2(new_n657), .A3(new_n677), .ZN(new_n961));
  NAND2_X1  g775(.A1(new_n961), .A2(new_n672), .ZN(new_n962));
  OR2_X1    g776(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n963));
  NAND2_X1  g777(.A1(new_n962), .A2(KEYINPUT62), .ZN(new_n964));
  NOR2_X1   g778(.A1(new_n627), .A2(new_n620), .ZN(new_n965));
  OR2_X1    g779(.A1(new_n965), .A2(KEYINPUT125), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n746), .ZN(new_n967));
  AOI211_X1 g781(.A(new_n667), .B(new_n967), .C1(KEYINPUT125), .C2(new_n965), .ZN(new_n968));
  AND2_X1   g782(.A1(new_n968), .A2(new_n679), .ZN(new_n969));
  NOR2_X1   g783(.A1(new_n783), .A2(new_n969), .ZN(new_n970));
  NAND4_X1  g784(.A1(new_n963), .A2(new_n777), .A3(new_n964), .A4(new_n970), .ZN(new_n971));
  OR2_X1    g785(.A1(new_n971), .A2(G953), .ZN(new_n972));
  NAND3_X1  g786(.A1(G227), .A2(G900), .A3(G953), .ZN(new_n973));
  AOI21_X1  g787(.A(new_n960), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g788(.A1(new_n743), .A2(new_n748), .ZN(new_n975));
  XNOR2_X1  g789(.A(new_n975), .B(KEYINPUT126), .ZN(new_n976));
  NOR2_X1   g790(.A1(new_n759), .A2(new_n704), .ZN(new_n977));
  AOI21_X1  g791(.A(new_n783), .B1(new_n877), .B2(new_n977), .ZN(new_n978));
  AND3_X1   g792(.A1(new_n978), .A2(new_n777), .A3(new_n961), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n976), .A2(new_n459), .A3(new_n979), .ZN(new_n980));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n981));
  NAND3_X1  g795(.A1(new_n981), .A2(new_n412), .A3(G900), .ZN(new_n982));
  OAI211_X1 g796(.A(new_n982), .B(G953), .C1(new_n981), .C2(G900), .ZN(new_n983));
  AND2_X1   g797(.A1(new_n960), .A2(new_n983), .ZN(new_n984));
  AOI21_X1  g798(.A(new_n974), .B1(new_n980), .B2(new_n984), .ZN(G72));
  NAND2_X1  g799(.A1(G472), .A2(G902), .ZN(new_n986));
  XOR2_X1   g800(.A(new_n986), .B(KEYINPUT63), .Z(new_n987));
  OAI21_X1  g801(.A(new_n987), .B1(new_n952), .B2(new_n971), .ZN(new_n988));
  NAND3_X1  g802(.A1(new_n988), .A2(new_n250), .A3(new_n306), .ZN(new_n989));
  INV_X1    g803(.A(new_n308), .ZN(new_n990));
  OAI21_X1  g804(.A(new_n987), .B1(new_n990), .B2(new_n660), .ZN(new_n991));
  OAI211_X1 g805(.A(new_n989), .B(new_n899), .C1(new_n875), .C2(new_n991), .ZN(new_n992));
  NAND3_X1  g806(.A1(new_n976), .A2(new_n951), .A3(new_n979), .ZN(new_n993));
  AOI211_X1 g807(.A(new_n250), .B(new_n306), .C1(new_n993), .C2(new_n987), .ZN(new_n994));
  NOR2_X1   g808(.A1(new_n992), .A2(new_n994), .ZN(G57));
endmodule


