//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 0 1 1 0 0 1 0 1 1 1 0 1 0 1 0 1 0 1 0 0 1 1 0 1 0 1 1 0 0 1 0 1 1 0 0 0 1 1 0 0 1 0 0 0 1 0 0 0 1 0 0 1 0 1 1 1 0 0 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:22:06 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n690, new_n691, new_n692, new_n693, new_n694, new_n696, new_n697,
    new_n698, new_n699, new_n700, new_n701, new_n702, new_n703, new_n704,
    new_n705, new_n706, new_n707, new_n708, new_n709, new_n711, new_n712,
    new_n713, new_n715, new_n716, new_n717, new_n718, new_n719, new_n721,
    new_n722, new_n723, new_n724, new_n725, new_n726, new_n727, new_n728,
    new_n729, new_n730, new_n731, new_n732, new_n733, new_n735, new_n736,
    new_n737, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n776, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n906, new_n907, new_n908, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n923, new_n924, new_n925, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n970, new_n971, new_n972,
    new_n973, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982;
  XNOR2_X1  g000(.A(KEYINPUT9), .B(G234), .ZN(new_n187));
  OAI21_X1  g001(.A(G221), .B1(new_n187), .B2(G902), .ZN(new_n188));
  INV_X1    g002(.A(G107), .ZN(new_n189));
  NAND3_X1  g003(.A1(new_n189), .A2(KEYINPUT79), .A3(G104), .ZN(new_n190));
  INV_X1    g004(.A(KEYINPUT3), .ZN(new_n191));
  NAND2_X1  g005(.A1(new_n190), .A2(new_n191), .ZN(new_n192));
  NAND4_X1  g006(.A1(new_n189), .A2(KEYINPUT79), .A3(KEYINPUT3), .A4(G104), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G104), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G107), .ZN(new_n196));
  NAND2_X1  g010(.A1(new_n194), .A2(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(G101), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT4), .ZN(new_n199));
  INV_X1    g013(.A(G101), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n200), .A2(KEYINPUT80), .ZN(new_n201));
  INV_X1    g015(.A(KEYINPUT80), .ZN(new_n202));
  NAND2_X1  g016(.A1(new_n202), .A2(G101), .ZN(new_n203));
  AND3_X1   g017(.A1(new_n201), .A2(new_n203), .A3(new_n196), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n199), .B1(new_n194), .B2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n198), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(KEYINPUT0), .A2(G128), .ZN(new_n207));
  OR2_X1    g021(.A1(KEYINPUT0), .A2(G128), .ZN(new_n208));
  INV_X1    g022(.A(G143), .ZN(new_n209));
  NOR2_X1   g023(.A1(new_n209), .A2(G146), .ZN(new_n210));
  INV_X1    g024(.A(G146), .ZN(new_n211));
  NOR2_X1   g025(.A1(new_n211), .A2(G143), .ZN(new_n212));
  OAI211_X1 g026(.A(new_n207), .B(new_n208), .C1(new_n210), .C2(new_n212), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT64), .B1(new_n209), .B2(G146), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT64), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n215), .A2(new_n211), .A3(G143), .ZN(new_n216));
  NAND2_X1  g030(.A1(new_n209), .A2(G146), .ZN(new_n217));
  INV_X1    g031(.A(new_n207), .ZN(new_n218));
  NAND4_X1  g032(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n218), .ZN(new_n219));
  NAND2_X1  g033(.A1(new_n213), .A2(new_n219), .ZN(new_n220));
  NAND2_X1  g034(.A1(new_n220), .A2(KEYINPUT69), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT69), .ZN(new_n222));
  NAND3_X1  g036(.A1(new_n213), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  AOI21_X1  g037(.A(new_n200), .B1(new_n194), .B2(new_n196), .ZN(new_n224));
  XOR2_X1   g038(.A(KEYINPUT81), .B(KEYINPUT4), .Z(new_n225));
  NAND2_X1  g039(.A1(new_n224), .A2(new_n225), .ZN(new_n226));
  NAND4_X1  g040(.A1(new_n206), .A2(new_n221), .A3(new_n223), .A4(new_n226), .ZN(new_n227));
  INV_X1    g041(.A(G128), .ZN(new_n228));
  NOR2_X1   g042(.A1(new_n228), .A2(KEYINPUT1), .ZN(new_n229));
  NAND4_X1  g043(.A1(new_n214), .A2(new_n216), .A3(new_n217), .A4(new_n229), .ZN(new_n230));
  AND3_X1   g044(.A1(new_n214), .A2(new_n216), .A3(new_n217), .ZN(new_n231));
  NAND2_X1  g045(.A1(new_n211), .A2(G143), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n228), .B1(new_n232), .B2(KEYINPUT1), .ZN(new_n233));
  OAI21_X1  g047(.A(new_n230), .B1(new_n231), .B2(new_n233), .ZN(new_n234));
  NAND2_X1  g048(.A1(new_n189), .A2(G104), .ZN(new_n235));
  AOI21_X1  g049(.A(new_n200), .B1(new_n235), .B2(new_n196), .ZN(new_n236));
  AOI21_X1  g050(.A(new_n236), .B1(new_n194), .B2(new_n204), .ZN(new_n237));
  NAND2_X1  g051(.A1(new_n234), .A2(new_n237), .ZN(new_n238));
  XNOR2_X1  g052(.A(KEYINPUT82), .B(KEYINPUT10), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT10), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT1), .ZN(new_n241));
  OAI21_X1  g055(.A(G128), .B1(new_n210), .B2(new_n241), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n232), .A2(new_n217), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n242), .A2(new_n243), .ZN(new_n244));
  AOI21_X1  g058(.A(new_n240), .B1(new_n244), .B2(new_n230), .ZN(new_n245));
  AOI22_X1  g059(.A1(new_n238), .A2(new_n239), .B1(new_n237), .B2(new_n245), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n227), .A2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(KEYINPUT11), .ZN(new_n248));
  INV_X1    g062(.A(G134), .ZN(new_n249));
  OAI21_X1  g063(.A(new_n248), .B1(new_n249), .B2(G137), .ZN(new_n250));
  INV_X1    g064(.A(G137), .ZN(new_n251));
  NAND3_X1  g065(.A1(new_n251), .A2(KEYINPUT11), .A3(G134), .ZN(new_n252));
  NAND2_X1  g066(.A1(new_n249), .A2(G137), .ZN(new_n253));
  NAND3_X1  g067(.A1(new_n250), .A2(new_n252), .A3(new_n253), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n254), .A2(G131), .ZN(new_n255));
  INV_X1    g069(.A(G131), .ZN(new_n256));
  NAND4_X1  g070(.A1(new_n250), .A2(new_n252), .A3(new_n256), .A4(new_n253), .ZN(new_n257));
  NAND2_X1  g071(.A1(new_n255), .A2(new_n257), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n247), .A2(new_n258), .ZN(new_n259));
  INV_X1    g073(.A(new_n258), .ZN(new_n260));
  NAND3_X1  g074(.A1(new_n227), .A2(new_n260), .A3(new_n246), .ZN(new_n261));
  NAND2_X1  g075(.A1(new_n259), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g076(.A1(KEYINPUT70), .A2(G953), .ZN(new_n263));
  NOR2_X1   g077(.A1(KEYINPUT70), .A2(G953), .ZN(new_n264));
  NOR2_X1   g078(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(G227), .ZN(new_n266));
  XOR2_X1   g080(.A(G110), .B(G140), .Z(new_n267));
  XNOR2_X1  g081(.A(new_n266), .B(new_n267), .ZN(new_n268));
  NAND2_X1  g082(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(new_n268), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n244), .A2(new_n230), .ZN(new_n271));
  OR2_X1    g085(.A1(new_n237), .A2(new_n271), .ZN(new_n272));
  NAND2_X1  g086(.A1(new_n272), .A2(new_n238), .ZN(new_n273));
  AOI21_X1  g087(.A(KEYINPUT12), .B1(new_n273), .B2(new_n258), .ZN(new_n274));
  INV_X1    g088(.A(KEYINPUT12), .ZN(new_n275));
  AOI211_X1 g089(.A(new_n275), .B(new_n260), .C1(new_n272), .C2(new_n238), .ZN(new_n276));
  OAI211_X1 g090(.A(new_n261), .B(new_n270), .C1(new_n274), .C2(new_n276), .ZN(new_n277));
  AOI211_X1 g091(.A(G469), .B(G902), .C1(new_n269), .C2(new_n277), .ZN(new_n278));
  OAI21_X1  g092(.A(new_n261), .B1(new_n274), .B2(new_n276), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n279), .A2(new_n268), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n259), .A2(new_n261), .A3(new_n270), .ZN(new_n281));
  NAND3_X1  g095(.A1(new_n280), .A2(new_n281), .A3(G469), .ZN(new_n282));
  INV_X1    g096(.A(G469), .ZN(new_n283));
  INV_X1    g097(.A(G902), .ZN(new_n284));
  NOR2_X1   g098(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g099(.A(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n282), .A2(new_n286), .ZN(new_n287));
  OAI21_X1  g101(.A(new_n188), .B1(new_n278), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  INV_X1    g103(.A(KEYINPUT90), .ZN(new_n290));
  INV_X1    g104(.A(G475), .ZN(new_n291));
  OR2_X1    g105(.A1(KEYINPUT70), .A2(G953), .ZN(new_n292));
  INV_X1    g106(.A(G237), .ZN(new_n293));
  NAND2_X1  g107(.A1(KEYINPUT70), .A2(G953), .ZN(new_n294));
  NAND4_X1  g108(.A1(new_n292), .A2(G214), .A3(new_n293), .A4(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n209), .ZN(new_n296));
  NAND4_X1  g110(.A1(new_n265), .A2(G143), .A3(G214), .A4(new_n293), .ZN(new_n297));
  NAND2_X1  g111(.A1(new_n296), .A2(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(KEYINPUT18), .A2(G131), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n298), .A2(new_n300), .ZN(new_n301));
  INV_X1    g115(.A(G140), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n302), .A2(G125), .ZN(new_n303));
  INV_X1    g117(.A(G125), .ZN(new_n304));
  NAND2_X1  g118(.A1(new_n304), .A2(G140), .ZN(new_n305));
  NAND2_X1  g119(.A1(new_n303), .A2(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(G146), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n303), .A2(new_n305), .A3(new_n211), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g123(.A1(new_n296), .A2(new_n297), .A3(new_n299), .ZN(new_n310));
  NAND3_X1  g124(.A1(new_n301), .A2(new_n309), .A3(new_n310), .ZN(new_n311));
  XNOR2_X1  g125(.A(G113), .B(G122), .ZN(new_n312));
  XNOR2_X1  g126(.A(new_n312), .B(new_n195), .ZN(new_n313));
  XNOR2_X1  g127(.A(new_n313), .B(KEYINPUT88), .ZN(new_n314));
  AND3_X1   g128(.A1(new_n296), .A2(new_n297), .A3(new_n256), .ZN(new_n315));
  AOI21_X1  g129(.A(new_n256), .B1(new_n296), .B2(new_n297), .ZN(new_n316));
  NOR3_X1   g130(.A1(new_n315), .A2(new_n316), .A3(KEYINPUT17), .ZN(new_n317));
  NAND3_X1  g131(.A1(new_n298), .A2(KEYINPUT17), .A3(G131), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT16), .ZN(new_n319));
  OR3_X1    g133(.A1(new_n304), .A2(KEYINPUT16), .A3(G140), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g135(.A1(new_n321), .A2(new_n211), .ZN(new_n322));
  NAND3_X1  g136(.A1(new_n319), .A2(new_n320), .A3(G146), .ZN(new_n323));
  NAND3_X1  g137(.A1(new_n318), .A2(new_n322), .A3(new_n323), .ZN(new_n324));
  OAI211_X1 g138(.A(new_n311), .B(new_n314), .C1(new_n317), .C2(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n322), .A2(new_n323), .ZN(new_n326));
  AOI21_X1  g140(.A(new_n326), .B1(KEYINPUT17), .B2(new_n316), .ZN(new_n327));
  NAND2_X1  g141(.A1(new_n298), .A2(G131), .ZN(new_n328));
  INV_X1    g142(.A(KEYINPUT17), .ZN(new_n329));
  NAND3_X1  g143(.A1(new_n296), .A2(new_n297), .A3(new_n256), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n328), .A2(new_n329), .A3(new_n330), .ZN(new_n331));
  AND2_X1   g145(.A1(new_n310), .A2(new_n309), .ZN(new_n332));
  AOI22_X1  g146(.A1(new_n327), .A2(new_n331), .B1(new_n301), .B2(new_n332), .ZN(new_n333));
  OAI21_X1  g147(.A(new_n325), .B1(new_n333), .B2(new_n313), .ZN(new_n334));
  AOI21_X1  g148(.A(new_n291), .B1(new_n334), .B2(new_n284), .ZN(new_n335));
  INV_X1    g149(.A(new_n313), .ZN(new_n336));
  AND3_X1   g150(.A1(new_n301), .A2(new_n309), .A3(new_n310), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT19), .ZN(new_n338));
  AOI21_X1  g152(.A(KEYINPUT19), .B1(new_n303), .B2(new_n305), .ZN(new_n339));
  NOR2_X1   g153(.A1(new_n338), .A2(new_n339), .ZN(new_n340));
  OAI21_X1  g154(.A(new_n323), .B1(new_n340), .B2(G146), .ZN(new_n341));
  AOI21_X1  g155(.A(new_n341), .B1(new_n328), .B2(new_n330), .ZN(new_n342));
  OAI21_X1  g156(.A(new_n336), .B1(new_n337), .B2(new_n342), .ZN(new_n343));
  AOI21_X1  g157(.A(KEYINPUT89), .B1(new_n325), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(KEYINPUT19), .ZN(new_n345));
  NAND2_X1  g159(.A1(new_n306), .A2(new_n345), .ZN(new_n346));
  NAND3_X1  g160(.A1(new_n303), .A2(new_n305), .A3(KEYINPUT19), .ZN(new_n347));
  AOI21_X1  g161(.A(G146), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  INV_X1    g162(.A(new_n323), .ZN(new_n349));
  NOR2_X1   g163(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n315), .B2(new_n316), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n313), .B1(new_n351), .B2(new_n311), .ZN(new_n352));
  AOI21_X1  g166(.A(new_n352), .B1(new_n333), .B2(new_n314), .ZN(new_n353));
  NOR2_X1   g167(.A1(G475), .A2(G902), .ZN(new_n354));
  INV_X1    g168(.A(new_n354), .ZN(new_n355));
  OAI22_X1  g169(.A1(new_n344), .A2(KEYINPUT20), .B1(new_n353), .B2(new_n355), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n325), .A2(new_n343), .ZN(new_n357));
  INV_X1    g171(.A(KEYINPUT20), .ZN(new_n358));
  NAND4_X1  g172(.A1(new_n357), .A2(KEYINPUT89), .A3(new_n358), .A4(new_n354), .ZN(new_n359));
  AOI211_X1 g173(.A(new_n290), .B(new_n335), .C1(new_n356), .C2(new_n359), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n356), .A2(new_n359), .ZN(new_n361));
  INV_X1    g175(.A(new_n335), .ZN(new_n362));
  AOI21_X1  g176(.A(KEYINPUT90), .B1(new_n361), .B2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n360), .A2(new_n363), .ZN(new_n364));
  INV_X1    g178(.A(G122), .ZN(new_n365));
  NAND2_X1  g179(.A1(new_n365), .A2(G116), .ZN(new_n366));
  INV_X1    g180(.A(G116), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n367), .A2(G122), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n366), .A2(new_n368), .A3(new_n189), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n209), .A2(G128), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n228), .A2(G143), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n370), .A2(new_n371), .A3(new_n249), .ZN(new_n372));
  INV_X1    g186(.A(new_n372), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n249), .B1(new_n370), .B2(new_n371), .ZN(new_n374));
  OAI21_X1  g188(.A(new_n369), .B1(new_n373), .B2(new_n374), .ZN(new_n375));
  OR3_X1    g189(.A1(new_n365), .A2(KEYINPUT14), .A3(G116), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT93), .ZN(new_n377));
  NOR2_X1   g191(.A1(new_n377), .A2(new_n189), .ZN(new_n378));
  NAND2_X1  g192(.A1(new_n368), .A2(KEYINPUT14), .ZN(new_n379));
  NAND4_X1  g193(.A1(new_n376), .A2(new_n379), .A3(KEYINPUT93), .A4(new_n366), .ZN(new_n380));
  AOI21_X1  g194(.A(new_n375), .B1(new_n378), .B2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(new_n381), .ZN(new_n382));
  INV_X1    g196(.A(G217), .ZN(new_n383));
  NOR3_X1   g197(.A1(new_n187), .A2(new_n383), .A3(G953), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n209), .A2(KEYINPUT13), .A3(G128), .ZN(new_n385));
  NOR2_X1   g199(.A1(new_n385), .A2(KEYINPUT91), .ZN(new_n386));
  NOR2_X1   g200(.A1(new_n386), .A2(new_n249), .ZN(new_n387));
  INV_X1    g201(.A(KEYINPUT13), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n370), .A2(new_n388), .ZN(new_n389));
  NAND4_X1  g203(.A1(new_n389), .A2(new_n385), .A3(KEYINPUT91), .A4(new_n371), .ZN(new_n390));
  NAND3_X1  g204(.A1(new_n387), .A2(KEYINPUT92), .A3(new_n390), .ZN(new_n391));
  INV_X1    g205(.A(new_n391), .ZN(new_n392));
  AOI21_X1  g206(.A(KEYINPUT92), .B1(new_n387), .B2(new_n390), .ZN(new_n393));
  NOR2_X1   g207(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n366), .A2(new_n368), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n395), .A2(G107), .ZN(new_n396));
  NAND2_X1  g210(.A1(new_n396), .A2(new_n369), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n397), .A2(new_n372), .ZN(new_n398));
  OAI211_X1 g212(.A(new_n382), .B(new_n384), .C1(new_n394), .C2(new_n398), .ZN(new_n399));
  INV_X1    g213(.A(new_n384), .ZN(new_n400));
  NAND2_X1  g214(.A1(new_n387), .A2(new_n390), .ZN(new_n401));
  INV_X1    g215(.A(KEYINPUT92), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n401), .A2(new_n402), .ZN(new_n403));
  AOI21_X1  g217(.A(new_n398), .B1(new_n403), .B2(new_n391), .ZN(new_n404));
  OAI21_X1  g218(.A(new_n400), .B1(new_n404), .B2(new_n381), .ZN(new_n405));
  NAND2_X1  g219(.A1(new_n399), .A2(new_n405), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n406), .A2(new_n284), .ZN(new_n407));
  INV_X1    g221(.A(G478), .ZN(new_n408));
  NOR2_X1   g222(.A1(new_n408), .A2(KEYINPUT15), .ZN(new_n409));
  NAND2_X1  g223(.A1(new_n407), .A2(new_n409), .ZN(new_n410));
  INV_X1    g224(.A(new_n409), .ZN(new_n411));
  NAND3_X1  g225(.A1(new_n406), .A2(new_n284), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g226(.A1(new_n410), .A2(KEYINPUT94), .A3(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT94), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n411), .B1(new_n406), .B2(new_n284), .ZN(new_n415));
  AOI211_X1 g229(.A(G902), .B(new_n409), .C1(new_n399), .C2(new_n405), .ZN(new_n416));
  OAI21_X1  g230(.A(new_n414), .B1(new_n415), .B2(new_n416), .ZN(new_n417));
  AND2_X1   g231(.A1(new_n413), .A2(new_n417), .ZN(new_n418));
  INV_X1    g232(.A(G953), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI211_X1 g234(.A(G952), .B(new_n419), .C1(new_n420), .C2(new_n293), .ZN(new_n421));
  XOR2_X1   g235(.A(new_n421), .B(KEYINPUT95), .Z(new_n422));
  INV_X1    g236(.A(new_n422), .ZN(new_n423));
  INV_X1    g237(.A(new_n265), .ZN(new_n424));
  OAI211_X1 g238(.A(new_n424), .B(G902), .C1(new_n420), .C2(new_n293), .ZN(new_n425));
  XNOR2_X1  g239(.A(new_n425), .B(KEYINPUT96), .ZN(new_n426));
  XNOR2_X1  g240(.A(KEYINPUT21), .B(G898), .ZN(new_n427));
  XNOR2_X1  g241(.A(new_n427), .B(KEYINPUT97), .ZN(new_n428));
  AOI21_X1  g242(.A(new_n423), .B1(new_n426), .B2(new_n428), .ZN(new_n429));
  NOR2_X1   g243(.A1(new_n418), .A2(new_n429), .ZN(new_n430));
  AND3_X1   g244(.A1(new_n289), .A2(new_n364), .A3(new_n430), .ZN(new_n431));
  INV_X1    g245(.A(KEYINPUT87), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT6), .ZN(new_n433));
  XNOR2_X1  g247(.A(G110), .B(G122), .ZN(new_n434));
  INV_X1    g248(.A(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(new_n205), .ZN(new_n436));
  OAI21_X1  g250(.A(new_n226), .B1(new_n436), .B2(new_n224), .ZN(new_n437));
  OAI21_X1  g251(.A(KEYINPUT66), .B1(new_n367), .B2(G119), .ZN(new_n438));
  INV_X1    g252(.A(KEYINPUT66), .ZN(new_n439));
  INV_X1    g253(.A(G119), .ZN(new_n440));
  NAND3_X1  g254(.A1(new_n439), .A2(new_n440), .A3(G116), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n438), .A2(new_n441), .ZN(new_n442));
  INV_X1    g256(.A(G113), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(KEYINPUT2), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT2), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n445), .A2(G113), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n444), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(KEYINPUT67), .B1(new_n440), .B2(G116), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT67), .ZN(new_n449));
  NAND3_X1  g263(.A1(new_n449), .A2(new_n367), .A3(G119), .ZN(new_n450));
  NAND4_X1  g264(.A1(new_n442), .A2(new_n447), .A3(new_n448), .A4(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT68), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n451), .A2(new_n452), .ZN(new_n453));
  AND2_X1   g267(.A1(new_n448), .A2(new_n450), .ZN(new_n454));
  NAND4_X1  g268(.A1(new_n454), .A2(KEYINPUT68), .A3(new_n447), .A4(new_n442), .ZN(new_n455));
  INV_X1    g269(.A(new_n447), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n454), .A2(new_n442), .ZN(new_n457));
  AOI22_X1  g271(.A1(new_n453), .A2(new_n455), .B1(new_n456), .B2(new_n457), .ZN(new_n458));
  NOR2_X1   g272(.A1(new_n437), .A2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n453), .A2(new_n455), .ZN(new_n460));
  NOR2_X1   g274(.A1(new_n367), .A2(G119), .ZN(new_n461));
  INV_X1    g275(.A(KEYINPUT5), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n443), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  OAI21_X1  g277(.A(new_n463), .B1(new_n457), .B2(new_n462), .ZN(new_n464));
  AND3_X1   g278(.A1(new_n460), .A2(new_n237), .A3(new_n464), .ZN(new_n465));
  OAI211_X1 g279(.A(new_n433), .B(new_n435), .C1(new_n459), .C2(new_n465), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n460), .A2(new_n237), .A3(new_n464), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n467), .B(new_n434), .C1(new_n437), .C2(new_n458), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n468), .A2(KEYINPUT6), .ZN(new_n469));
  NAND2_X1  g283(.A1(new_n457), .A2(new_n456), .ZN(new_n470));
  NAND2_X1  g284(.A1(new_n460), .A2(new_n470), .ZN(new_n471));
  NAND3_X1  g285(.A1(new_n471), .A2(new_n206), .A3(new_n226), .ZN(new_n472));
  AOI21_X1  g286(.A(new_n434), .B1(new_n472), .B2(new_n467), .ZN(new_n473));
  OAI211_X1 g287(.A(KEYINPUT83), .B(new_n466), .C1(new_n469), .C2(new_n473), .ZN(new_n474));
  OAI21_X1  g288(.A(new_n435), .B1(new_n459), .B2(new_n465), .ZN(new_n475));
  INV_X1    g289(.A(KEYINPUT83), .ZN(new_n476));
  NAND4_X1  g290(.A1(new_n475), .A2(new_n476), .A3(KEYINPUT6), .A4(new_n468), .ZN(new_n477));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n477), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n220), .A2(G125), .ZN(new_n479));
  NAND3_X1  g293(.A1(new_n244), .A2(new_n304), .A3(new_n230), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  INV_X1    g295(.A(G224), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n482), .A2(G953), .ZN(new_n483));
  XOR2_X1   g297(.A(new_n481), .B(new_n483), .Z(new_n484));
  INV_X1    g298(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g299(.A1(new_n478), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g300(.A(new_n434), .B(KEYINPUT8), .ZN(new_n487));
  AOI21_X1  g301(.A(new_n237), .B1(new_n460), .B2(new_n464), .ZN(new_n488));
  OAI21_X1  g302(.A(new_n487), .B1(new_n465), .B2(new_n488), .ZN(new_n489));
  AOI21_X1  g303(.A(new_n304), .B1(new_n213), .B2(new_n219), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT84), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT7), .ZN(new_n492));
  OAI22_X1  g306(.A1(new_n490), .A2(new_n491), .B1(new_n492), .B2(new_n483), .ZN(new_n493));
  XNOR2_X1  g307(.A(new_n493), .B(new_n481), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n489), .A2(new_n468), .A3(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT85), .ZN(new_n496));
  AND3_X1   g310(.A1(new_n495), .A2(new_n496), .A3(new_n284), .ZN(new_n497));
  AOI21_X1  g311(.A(new_n496), .B1(new_n495), .B2(new_n284), .ZN(new_n498));
  NOR2_X1   g312(.A1(new_n497), .A2(new_n498), .ZN(new_n499));
  NAND2_X1  g313(.A1(new_n486), .A2(new_n499), .ZN(new_n500));
  OAI21_X1  g314(.A(G210), .B1(G237), .B2(G902), .ZN(new_n501));
  NOR2_X1   g315(.A1(new_n501), .A2(KEYINPUT86), .ZN(new_n502));
  NAND2_X1  g316(.A1(new_n500), .A2(new_n502), .ZN(new_n503));
  OAI211_X1 g317(.A(new_n486), .B(new_n499), .C1(KEYINPUT86), .C2(new_n501), .ZN(new_n504));
  NAND2_X1  g318(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g319(.A(G214), .B1(G237), .B2(G902), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n432), .B1(new_n505), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n506), .ZN(new_n508));
  AOI211_X1 g322(.A(KEYINPUT87), .B(new_n508), .C1(new_n503), .C2(new_n504), .ZN(new_n509));
  OAI21_X1  g323(.A(new_n431), .B1(new_n507), .B2(new_n509), .ZN(new_n510));
  INV_X1    g324(.A(KEYINPUT98), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT25), .ZN(new_n513));
  XNOR2_X1  g327(.A(KEYINPUT24), .B(G110), .ZN(new_n514));
  INV_X1    g328(.A(KEYINPUT76), .ZN(new_n515));
  XNOR2_X1  g329(.A(new_n514), .B(new_n515), .ZN(new_n516));
  XNOR2_X1  g330(.A(G119), .B(G128), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  OAI21_X1  g332(.A(KEYINPUT77), .B1(new_n440), .B2(G128), .ZN(new_n519));
  AOI22_X1  g333(.A1(new_n519), .A2(KEYINPUT23), .B1(new_n440), .B2(G128), .ZN(new_n520));
  OAI21_X1  g334(.A(new_n520), .B1(KEYINPUT23), .B2(new_n519), .ZN(new_n521));
  NOR2_X1   g335(.A1(new_n521), .A2(G110), .ZN(new_n522));
  OAI211_X1 g336(.A(new_n323), .B(new_n308), .C1(new_n518), .C2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n516), .A2(new_n517), .ZN(new_n524));
  NAND2_X1  g338(.A1(new_n521), .A2(G110), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n326), .ZN(new_n526));
  NAND2_X1  g340(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  XNOR2_X1  g341(.A(KEYINPUT22), .B(G137), .ZN(new_n528));
  XNOR2_X1  g342(.A(new_n528), .B(KEYINPUT78), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n265), .A2(G221), .A3(G234), .ZN(new_n530));
  XNOR2_X1  g344(.A(new_n529), .B(new_n530), .ZN(new_n531));
  NOR2_X1   g345(.A1(new_n527), .A2(new_n531), .ZN(new_n532));
  INV_X1    g346(.A(new_n531), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n523), .B2(new_n526), .ZN(new_n534));
  NOR2_X1   g348(.A1(new_n532), .A2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(new_n513), .B1(new_n535), .B2(G902), .ZN(new_n536));
  OAI211_X1 g350(.A(KEYINPUT25), .B(new_n284), .C1(new_n532), .C2(new_n534), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  AOI21_X1  g352(.A(new_n383), .B1(G234), .B2(new_n284), .ZN(new_n539));
  INV_X1    g353(.A(new_n535), .ZN(new_n540));
  NOR2_X1   g354(.A1(new_n539), .A2(G902), .ZN(new_n541));
  AOI22_X1  g355(.A1(new_n538), .A2(new_n539), .B1(new_n540), .B2(new_n541), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  INV_X1    g357(.A(KEYINPUT30), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n260), .A2(new_n220), .ZN(new_n545));
  NAND3_X1  g359(.A1(new_n251), .A2(KEYINPUT65), .A3(G134), .ZN(new_n546));
  INV_X1    g360(.A(new_n253), .ZN(new_n547));
  INV_X1    g361(.A(KEYINPUT65), .ZN(new_n548));
  OAI21_X1  g362(.A(new_n548), .B1(new_n249), .B2(G137), .ZN(new_n549));
  OAI211_X1 g363(.A(G131), .B(new_n546), .C1(new_n547), .C2(new_n549), .ZN(new_n550));
  AND3_X1   g364(.A1(new_n271), .A2(new_n257), .A3(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n544), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  NAND3_X1  g366(.A1(new_n221), .A2(new_n258), .A3(new_n223), .ZN(new_n553));
  NAND3_X1  g367(.A1(new_n271), .A2(new_n257), .A3(new_n550), .ZN(new_n554));
  NAND3_X1  g368(.A1(new_n553), .A2(KEYINPUT30), .A3(new_n554), .ZN(new_n555));
  NAND3_X1  g369(.A1(new_n552), .A2(new_n555), .A3(new_n471), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n265), .A2(G210), .A3(new_n293), .ZN(new_n557));
  XOR2_X1   g371(.A(KEYINPUT71), .B(KEYINPUT27), .Z(new_n558));
  XNOR2_X1  g372(.A(new_n557), .B(new_n558), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  NAND3_X1  g375(.A1(new_n458), .A2(new_n553), .A3(new_n554), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n556), .A2(new_n561), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(KEYINPUT28), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n562), .A2(new_n565), .ZN(new_n566));
  OAI21_X1  g380(.A(new_n471), .B1(new_n551), .B2(new_n545), .ZN(new_n567));
  NAND4_X1  g381(.A1(new_n458), .A2(new_n553), .A3(KEYINPUT28), .A4(new_n554), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n566), .A2(new_n567), .A3(new_n568), .ZN(new_n569));
  INV_X1    g383(.A(new_n561), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT72), .B(KEYINPUT31), .ZN(new_n572));
  NAND4_X1  g386(.A1(new_n556), .A2(new_n561), .A3(new_n562), .A4(new_n572), .ZN(new_n573));
  NAND3_X1  g387(.A1(new_n564), .A2(new_n571), .A3(new_n573), .ZN(new_n574));
  NOR2_X1   g388(.A1(G472), .A2(G902), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(KEYINPUT73), .ZN(new_n577));
  NAND2_X1  g391(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND3_X1  g392(.A1(new_n574), .A2(KEYINPUT73), .A3(new_n575), .ZN(new_n579));
  XNOR2_X1  g393(.A(KEYINPUT74), .B(KEYINPUT32), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(new_n581));
  AND2_X1   g395(.A1(new_n574), .A2(new_n575), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n556), .A2(new_n562), .ZN(new_n583));
  NAND2_X1  g397(.A1(new_n583), .A2(new_n570), .ZN(new_n584));
  NAND4_X1  g398(.A1(new_n566), .A2(new_n561), .A3(new_n567), .A4(new_n568), .ZN(new_n585));
  INV_X1    g399(.A(KEYINPUT29), .ZN(new_n586));
  NAND3_X1  g400(.A1(new_n584), .A2(new_n585), .A3(new_n586), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n553), .A2(new_n554), .ZN(new_n588));
  NAND2_X1  g402(.A1(new_n588), .A2(new_n471), .ZN(new_n589));
  NAND3_X1  g403(.A1(new_n589), .A2(KEYINPUT75), .A3(new_n562), .ZN(new_n590));
  INV_X1    g404(.A(KEYINPUT75), .ZN(new_n591));
  NAND3_X1  g405(.A1(new_n588), .A2(new_n591), .A3(new_n471), .ZN(new_n592));
  NAND3_X1  g406(.A1(new_n590), .A2(KEYINPUT28), .A3(new_n592), .ZN(new_n593));
  NAND4_X1  g407(.A1(new_n593), .A2(KEYINPUT29), .A3(new_n561), .A4(new_n566), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n587), .A2(new_n284), .A3(new_n594), .ZN(new_n595));
  AOI22_X1  g409(.A1(new_n582), .A2(KEYINPUT32), .B1(new_n595), .B2(G472), .ZN(new_n596));
  AOI21_X1  g410(.A(new_n543), .B1(new_n581), .B2(new_n596), .ZN(new_n597));
  OAI211_X1 g411(.A(KEYINPUT98), .B(new_n431), .C1(new_n507), .C2(new_n509), .ZN(new_n598));
  NAND3_X1  g412(.A1(new_n512), .A2(new_n597), .A3(new_n598), .ZN(new_n599));
  NAND2_X1  g413(.A1(new_n201), .A2(new_n203), .ZN(new_n600));
  XNOR2_X1  g414(.A(new_n599), .B(new_n600), .ZN(G3));
  AND2_X1   g415(.A1(new_n578), .A2(new_n579), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n574), .A2(new_n284), .ZN(new_n603));
  NAND2_X1  g417(.A1(new_n603), .A2(G472), .ZN(new_n604));
  NAND2_X1  g418(.A1(new_n602), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n269), .A2(new_n277), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n606), .A2(new_n283), .A3(new_n284), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n607), .A2(new_n286), .A3(new_n282), .ZN(new_n608));
  NAND3_X1  g422(.A1(new_n542), .A2(new_n608), .A3(new_n188), .ZN(new_n609));
  OAI21_X1  g423(.A(KEYINPUT99), .B1(new_n605), .B2(new_n609), .ZN(new_n610));
  INV_X1    g424(.A(new_n609), .ZN(new_n611));
  INV_X1    g425(.A(KEYINPUT99), .ZN(new_n612));
  NAND4_X1  g426(.A1(new_n611), .A2(new_n612), .A3(new_n602), .A4(new_n604), .ZN(new_n613));
  AND2_X1   g427(.A1(new_n610), .A2(new_n613), .ZN(new_n614));
  INV_X1    g428(.A(KEYINPUT100), .ZN(new_n615));
  AOI21_X1  g429(.A(new_n508), .B1(new_n500), .B2(new_n501), .ZN(new_n616));
  INV_X1    g430(.A(new_n501), .ZN(new_n617));
  NAND3_X1  g431(.A1(new_n486), .A2(new_n499), .A3(new_n617), .ZN(new_n618));
  AOI21_X1  g432(.A(new_n615), .B1(new_n616), .B2(new_n618), .ZN(new_n619));
  NAND2_X1  g433(.A1(new_n495), .A2(new_n284), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(KEYINPUT85), .ZN(new_n621));
  NAND3_X1  g435(.A1(new_n495), .A2(new_n496), .A3(new_n284), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n621), .A2(new_n622), .ZN(new_n623));
  AOI21_X1  g437(.A(new_n484), .B1(new_n474), .B2(new_n477), .ZN(new_n624));
  OAI21_X1  g438(.A(new_n501), .B1(new_n623), .B2(new_n624), .ZN(new_n625));
  NAND4_X1  g439(.A1(new_n625), .A2(new_n618), .A3(new_n615), .A4(new_n506), .ZN(new_n626));
  INV_X1    g440(.A(new_n626), .ZN(new_n627));
  NOR2_X1   g441(.A1(new_n619), .A2(new_n627), .ZN(new_n628));
  NOR2_X1   g442(.A1(new_n407), .A2(G478), .ZN(new_n629));
  NOR2_X1   g443(.A1(new_n408), .A2(new_n284), .ZN(new_n630));
  NOR2_X1   g444(.A1(new_n629), .A2(new_n630), .ZN(new_n631));
  OR2_X1    g445(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n406), .A2(KEYINPUT33), .ZN(new_n633));
  AND2_X1   g447(.A1(new_n632), .A2(new_n633), .ZN(new_n634));
  INV_X1    g448(.A(new_n634), .ZN(new_n635));
  OAI21_X1  g449(.A(new_n631), .B1(new_n635), .B2(new_n408), .ZN(new_n636));
  NOR3_X1   g450(.A1(new_n364), .A2(new_n429), .A3(new_n636), .ZN(new_n637));
  NAND3_X1  g451(.A1(new_n614), .A2(new_n628), .A3(new_n637), .ZN(new_n638));
  XOR2_X1   g452(.A(KEYINPUT34), .B(G104), .Z(new_n639));
  XNOR2_X1  g453(.A(new_n638), .B(new_n639), .ZN(G6));
  AND3_X1   g454(.A1(new_n413), .A2(new_n417), .A3(new_n362), .ZN(new_n641));
  INV_X1    g455(.A(new_n429), .ZN(new_n642));
  OAI211_X1 g456(.A(new_n357), .B(new_n354), .C1(KEYINPUT101), .C2(new_n358), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n355), .B1(new_n325), .B2(new_n343), .ZN(new_n644));
  XNOR2_X1  g458(.A(KEYINPUT101), .B(KEYINPUT20), .ZN(new_n645));
  OAI21_X1  g459(.A(new_n643), .B1(new_n644), .B2(new_n645), .ZN(new_n646));
  NAND4_X1  g460(.A1(new_n641), .A2(KEYINPUT102), .A3(new_n642), .A4(new_n646), .ZN(new_n647));
  INV_X1    g461(.A(KEYINPUT102), .ZN(new_n648));
  NAND4_X1  g462(.A1(new_n646), .A2(new_n413), .A3(new_n417), .A4(new_n362), .ZN(new_n649));
  OAI21_X1  g463(.A(new_n648), .B1(new_n649), .B2(new_n429), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n647), .A2(new_n650), .ZN(new_n651));
  NAND3_X1  g465(.A1(new_n614), .A2(new_n628), .A3(new_n651), .ZN(new_n652));
  XNOR2_X1  g466(.A(KEYINPUT104), .B(G107), .ZN(new_n653));
  XNOR2_X1  g467(.A(new_n652), .B(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT103), .B(KEYINPUT35), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(G9));
  INV_X1    g470(.A(KEYINPUT36), .ZN(new_n657));
  NAND2_X1  g471(.A1(new_n531), .A2(new_n657), .ZN(new_n658));
  XOR2_X1   g472(.A(new_n658), .B(KEYINPUT105), .Z(new_n659));
  XNOR2_X1  g473(.A(new_n659), .B(new_n527), .ZN(new_n660));
  NAND2_X1  g474(.A1(new_n660), .A2(new_n541), .ZN(new_n661));
  NAND2_X1  g475(.A1(new_n538), .A2(new_n539), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n661), .A2(new_n662), .ZN(new_n663));
  NAND3_X1  g477(.A1(new_n602), .A2(new_n604), .A3(new_n663), .ZN(new_n664));
  XNOR2_X1  g478(.A(new_n664), .B(KEYINPUT106), .ZN(new_n665));
  NAND3_X1  g479(.A1(new_n512), .A2(new_n598), .A3(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(KEYINPUT37), .B(G110), .Z(new_n667));
  XNOR2_X1  g481(.A(new_n666), .B(new_n667), .ZN(G12));
  AOI22_X1  g482(.A1(new_n660), .A2(new_n541), .B1(new_n538), .B2(new_n539), .ZN(new_n669));
  AOI211_X1 g483(.A(new_n288), .B(new_n669), .C1(new_n581), .C2(new_n596), .ZN(new_n670));
  INV_X1    g484(.A(G900), .ZN(new_n671));
  AOI21_X1  g485(.A(new_n423), .B1(new_n426), .B2(new_n671), .ZN(new_n672));
  NOR2_X1   g486(.A1(new_n649), .A2(new_n672), .ZN(new_n673));
  NAND3_X1  g487(.A1(new_n628), .A2(new_n670), .A3(new_n673), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(G128), .ZN(G30));
  NAND2_X1  g489(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n590), .A2(new_n570), .A3(new_n592), .ZN(new_n677));
  AND2_X1   g491(.A1(new_n677), .A2(new_n563), .ZN(new_n678));
  OAI21_X1  g492(.A(G472), .B1(new_n678), .B2(G902), .ZN(new_n679));
  NAND3_X1  g493(.A1(new_n581), .A2(new_n676), .A3(new_n679), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  XOR2_X1   g495(.A(new_n672), .B(KEYINPUT39), .Z(new_n682));
  NAND2_X1  g496(.A1(new_n289), .A2(new_n682), .ZN(new_n683));
  AOI211_X1 g497(.A(new_n508), .B(new_n663), .C1(new_n683), .C2(KEYINPUT40), .ZN(new_n684));
  OAI21_X1  g498(.A(new_n684), .B1(KEYINPUT40), .B2(new_n683), .ZN(new_n685));
  OAI21_X1  g499(.A(new_n418), .B1(new_n360), .B2(new_n363), .ZN(new_n686));
  XOR2_X1   g500(.A(new_n505), .B(KEYINPUT38), .Z(new_n687));
  OR4_X1    g501(.A1(new_n681), .A2(new_n685), .A3(new_n686), .A4(new_n687), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(G143), .ZN(G45));
  AOI211_X1 g503(.A(new_n629), .B(new_n630), .C1(new_n634), .C2(G478), .ZN(new_n690));
  INV_X1    g504(.A(new_n672), .ZN(new_n691));
  OAI211_X1 g505(.A(new_n690), .B(new_n691), .C1(new_n360), .C2(new_n363), .ZN(new_n692));
  INV_X1    g506(.A(new_n692), .ZN(new_n693));
  NAND3_X1  g507(.A1(new_n628), .A2(new_n670), .A3(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G146), .ZN(G48));
  NAND2_X1  g509(.A1(new_n606), .A2(new_n284), .ZN(new_n696));
  NAND2_X1  g510(.A1(new_n696), .A2(G469), .ZN(new_n697));
  NAND3_X1  g511(.A1(new_n697), .A2(new_n188), .A3(new_n607), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n597), .A2(new_n699), .ZN(new_n700));
  NAND4_X1  g514(.A1(new_n700), .A2(new_n628), .A3(KEYINPUT107), .A4(new_n637), .ZN(new_n701));
  INV_X1    g515(.A(KEYINPUT107), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n625), .A2(new_n618), .A3(new_n506), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n703), .A2(KEYINPUT100), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n637), .A2(new_n626), .A3(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n597), .A2(new_n699), .ZN(new_n706));
  OAI21_X1  g520(.A(new_n702), .B1(new_n705), .B2(new_n706), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n701), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(KEYINPUT41), .B(G113), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n708), .B(new_n709), .ZN(G15));
  NAND3_X1  g524(.A1(new_n651), .A2(new_n626), .A3(new_n704), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n706), .ZN(new_n712));
  XOR2_X1   g526(.A(KEYINPUT108), .B(G116), .Z(new_n713));
  XNOR2_X1  g527(.A(new_n712), .B(new_n713), .ZN(G18));
  AND2_X1   g528(.A1(new_n364), .A2(new_n430), .ZN(new_n715));
  NAND4_X1  g529(.A1(new_n715), .A2(new_n704), .A3(new_n626), .A4(new_n699), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n581), .A2(new_n596), .ZN(new_n717));
  NAND2_X1  g531(.A1(new_n717), .A2(new_n663), .ZN(new_n718));
  NOR2_X1   g532(.A1(new_n716), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g533(.A(new_n719), .B(new_n440), .ZN(G21));
  AND2_X1   g534(.A1(new_n593), .A2(new_n566), .ZN(new_n721));
  OAI211_X1 g535(.A(new_n564), .B(new_n573), .C1(new_n721), .C2(new_n561), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n722), .A2(new_n575), .ZN(new_n723));
  AND2_X1   g537(.A1(new_n723), .A2(new_n604), .ZN(new_n724));
  NAND2_X1  g538(.A1(new_n724), .A2(new_n542), .ZN(new_n725));
  NOR3_X1   g539(.A1(new_n725), .A2(new_n429), .A3(new_n698), .ZN(new_n726));
  INV_X1    g540(.A(KEYINPUT109), .ZN(new_n727));
  NAND2_X1  g541(.A1(new_n686), .A2(new_n727), .ZN(new_n728));
  OAI211_X1 g542(.A(KEYINPUT109), .B(new_n418), .C1(new_n360), .C2(new_n363), .ZN(new_n729));
  NAND4_X1  g543(.A1(new_n728), .A2(new_n704), .A3(new_n626), .A4(new_n729), .ZN(new_n730));
  AND2_X1   g544(.A1(new_n730), .A2(KEYINPUT110), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n730), .A2(KEYINPUT110), .ZN(new_n732));
  OAI21_X1  g546(.A(new_n726), .B1(new_n731), .B2(new_n732), .ZN(new_n733));
  XNOR2_X1  g547(.A(new_n733), .B(G122), .ZN(G24));
  NAND3_X1  g548(.A1(new_n663), .A2(new_n604), .A3(new_n723), .ZN(new_n735));
  NOR2_X1   g549(.A1(new_n735), .A2(new_n692), .ZN(new_n736));
  NAND3_X1  g550(.A1(new_n628), .A2(new_n699), .A3(new_n736), .ZN(new_n737));
  XNOR2_X1  g551(.A(new_n737), .B(G125), .ZN(G27));
  XNOR2_X1  g552(.A(new_n288), .B(KEYINPUT111), .ZN(new_n739));
  NOR2_X1   g553(.A1(new_n505), .A2(new_n508), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n739), .A2(new_n597), .A3(new_n740), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n692), .A2(KEYINPUT42), .ZN(new_n742));
  OR2_X1    g556(.A1(new_n582), .A2(KEYINPUT32), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n543), .B1(new_n743), .B2(new_n596), .ZN(new_n744));
  NAND4_X1  g558(.A1(new_n739), .A2(new_n693), .A3(new_n740), .A4(new_n744), .ZN(new_n745));
  AOI22_X1  g559(.A1(new_n741), .A2(new_n742), .B1(new_n745), .B2(KEYINPUT42), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G131), .ZN(G33));
  NAND4_X1  g561(.A1(new_n739), .A2(new_n740), .A3(new_n673), .A4(new_n597), .ZN(new_n748));
  XNOR2_X1  g562(.A(KEYINPUT112), .B(G134), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n748), .B(new_n749), .ZN(G36));
  NAND2_X1  g564(.A1(new_n280), .A2(new_n281), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT45), .ZN(new_n752));
  AOI21_X1  g566(.A(new_n283), .B1(new_n751), .B2(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n753), .B1(new_n752), .B2(new_n751), .ZN(new_n754));
  INV_X1    g568(.A(KEYINPUT113), .ZN(new_n755));
  XNOR2_X1  g569(.A(new_n754), .B(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n286), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  NAND2_X1  g572(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n756), .A2(KEYINPUT46), .A3(new_n286), .ZN(new_n760));
  NAND3_X1  g574(.A1(new_n759), .A2(new_n607), .A3(new_n760), .ZN(new_n761));
  NAND3_X1  g575(.A1(new_n761), .A2(new_n188), .A3(new_n682), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT114), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  NAND4_X1  g578(.A1(new_n761), .A2(KEYINPUT114), .A3(new_n188), .A4(new_n682), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n364), .A2(new_n690), .ZN(new_n766));
  XOR2_X1   g580(.A(new_n766), .B(KEYINPUT43), .Z(new_n767));
  AOI21_X1  g581(.A(new_n669), .B1(new_n602), .B2(new_n604), .ZN(new_n768));
  NAND3_X1  g582(.A1(new_n767), .A2(KEYINPUT44), .A3(new_n768), .ZN(new_n769));
  AOI21_X1  g583(.A(KEYINPUT44), .B1(new_n767), .B2(new_n768), .ZN(new_n770));
  INV_X1    g584(.A(new_n740), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n770), .A2(new_n771), .ZN(new_n772));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n765), .A3(new_n769), .A4(new_n772), .ZN(new_n773));
  XOR2_X1   g587(.A(KEYINPUT115), .B(G137), .Z(new_n774));
  XNOR2_X1  g588(.A(new_n773), .B(new_n774), .ZN(G39));
  NOR4_X1   g589(.A1(new_n771), .A2(new_n717), .A3(new_n542), .A4(new_n692), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n761), .A2(KEYINPUT47), .A3(new_n188), .ZN(new_n777));
  INV_X1    g591(.A(new_n777), .ZN(new_n778));
  AOI21_X1  g592(.A(KEYINPUT47), .B1(new_n761), .B2(new_n188), .ZN(new_n779));
  OAI21_X1  g593(.A(new_n776), .B1(new_n778), .B2(new_n779), .ZN(new_n780));
  NAND2_X1  g594(.A1(new_n780), .A2(KEYINPUT116), .ZN(new_n781));
  INV_X1    g595(.A(new_n779), .ZN(new_n782));
  NAND2_X1  g596(.A1(new_n782), .A2(new_n777), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT116), .ZN(new_n784));
  NAND3_X1  g598(.A1(new_n783), .A2(new_n784), .A3(new_n776), .ZN(new_n785));
  NAND2_X1  g599(.A1(new_n781), .A2(new_n785), .ZN(new_n786));
  XNOR2_X1  g600(.A(new_n786), .B(G140), .ZN(G42));
  INV_X1    g601(.A(KEYINPUT53), .ZN(new_n788));
  OAI22_X1  g602(.A1(new_n716), .A2(new_n718), .B1(new_n711), .B2(new_n706), .ZN(new_n789));
  INV_X1    g603(.A(new_n789), .ZN(new_n790));
  AND4_X1   g604(.A1(new_n708), .A2(new_n733), .A3(new_n746), .A4(new_n790), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n674), .A2(new_n694), .A3(new_n737), .ZN(new_n792));
  NAND4_X1  g606(.A1(new_n680), .A2(new_n289), .A3(new_n669), .A4(new_n691), .ZN(new_n793));
  INV_X1    g607(.A(new_n793), .ZN(new_n794));
  OAI21_X1  g608(.A(new_n794), .B1(new_n731), .B2(new_n732), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND3_X1  g610(.A1(new_n792), .A2(new_n795), .A3(new_n796), .ZN(new_n797));
  INV_X1    g611(.A(KEYINPUT110), .ZN(new_n798));
  NAND4_X1  g612(.A1(new_n628), .A2(new_n798), .A3(new_n729), .A4(new_n728), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n730), .A2(KEYINPUT110), .ZN(new_n800));
  AOI21_X1  g614(.A(new_n793), .B1(new_n799), .B2(new_n800), .ZN(new_n801));
  NAND3_X1  g615(.A1(new_n674), .A2(new_n694), .A3(new_n737), .ZN(new_n802));
  OAI21_X1  g616(.A(KEYINPUT52), .B1(new_n801), .B2(new_n802), .ZN(new_n803));
  NOR3_X1   g617(.A1(new_n415), .A2(new_n416), .A3(new_n672), .ZN(new_n804));
  NAND3_X1  g618(.A1(new_n804), .A2(new_n646), .A3(new_n362), .ZN(new_n805));
  XNOR2_X1  g619(.A(new_n805), .B(KEYINPUT118), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n670), .A2(new_n740), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g621(.A1(new_n736), .A2(new_n739), .A3(new_n740), .ZN(new_n808));
  AND3_X1   g622(.A1(new_n807), .A2(new_n748), .A3(new_n808), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n791), .A2(new_n797), .A3(new_n803), .A4(new_n809), .ZN(new_n810));
  OR2_X1    g624(.A1(new_n507), .A2(new_n509), .ZN(new_n811));
  NAND3_X1  g625(.A1(new_n614), .A2(new_n811), .A3(new_n637), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n599), .A2(new_n812), .ZN(new_n813));
  INV_X1    g627(.A(KEYINPUT117), .ZN(new_n814));
  NAND2_X1  g628(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n599), .A2(new_n812), .A3(KEYINPUT117), .ZN(new_n816));
  OAI21_X1  g630(.A(new_n364), .B1(new_n415), .B2(new_n416), .ZN(new_n817));
  NOR2_X1   g631(.A1(new_n817), .A2(new_n429), .ZN(new_n818));
  NAND3_X1  g632(.A1(new_n614), .A2(new_n811), .A3(new_n818), .ZN(new_n819));
  NAND4_X1  g633(.A1(new_n815), .A2(new_n666), .A3(new_n816), .A4(new_n819), .ZN(new_n820));
  OAI21_X1  g634(.A(new_n788), .B1(new_n810), .B2(new_n820), .ZN(new_n821));
  NAND2_X1  g635(.A1(new_n797), .A2(new_n803), .ZN(new_n822));
  NAND2_X1  g636(.A1(new_n799), .A2(new_n800), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n789), .B1(new_n823), .B2(new_n726), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n824), .A2(new_n708), .A3(new_n746), .A4(new_n809), .ZN(new_n825));
  NOR2_X1   g639(.A1(new_n822), .A2(new_n825), .ZN(new_n826));
  AND3_X1   g640(.A1(new_n599), .A2(new_n812), .A3(KEYINPUT117), .ZN(new_n827));
  AOI21_X1  g641(.A(KEYINPUT117), .B1(new_n599), .B2(new_n812), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n666), .A2(new_n819), .ZN(new_n829));
  NOR3_X1   g643(.A1(new_n827), .A2(new_n828), .A3(new_n829), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n826), .A2(new_n830), .ZN(new_n831));
  NAND2_X1  g645(.A1(new_n674), .A2(new_n737), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n832), .A2(KEYINPUT52), .ZN(new_n833));
  NAND2_X1  g647(.A1(new_n833), .A2(new_n788), .ZN(new_n834));
  INV_X1    g648(.A(new_n834), .ZN(new_n835));
  OAI21_X1  g649(.A(new_n821), .B1(new_n831), .B2(new_n835), .ZN(new_n836));
  NAND2_X1  g650(.A1(new_n836), .A2(KEYINPUT54), .ZN(new_n837));
  NAND4_X1  g651(.A1(new_n733), .A2(new_n708), .A3(new_n790), .A4(new_n746), .ZN(new_n838));
  INV_X1    g652(.A(KEYINPUT119), .ZN(new_n839));
  NAND2_X1  g653(.A1(new_n838), .A2(new_n839), .ZN(new_n840));
  NAND4_X1  g654(.A1(new_n824), .A2(KEYINPUT119), .A3(new_n708), .A4(new_n746), .ZN(new_n841));
  NAND2_X1  g655(.A1(new_n840), .A2(new_n841), .ZN(new_n842));
  NAND4_X1  g656(.A1(new_n807), .A2(new_n808), .A3(new_n748), .A4(KEYINPUT53), .ZN(new_n843));
  AOI21_X1  g657(.A(new_n843), .B1(KEYINPUT52), .B2(new_n832), .ZN(new_n844));
  AND3_X1   g658(.A1(new_n797), .A2(new_n803), .A3(new_n844), .ZN(new_n845));
  NAND3_X1  g659(.A1(new_n842), .A2(new_n830), .A3(new_n845), .ZN(new_n846));
  XNOR2_X1  g660(.A(KEYINPUT120), .B(KEYINPUT54), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n821), .A2(new_n846), .A3(new_n847), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT121), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n821), .A2(KEYINPUT121), .A3(new_n846), .A4(new_n847), .ZN(new_n851));
  NAND3_X1  g665(.A1(new_n837), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n767), .A2(new_n423), .ZN(new_n853));
  NOR2_X1   g667(.A1(new_n771), .A2(new_n698), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n853), .A2(new_n854), .ZN(new_n855));
  NAND4_X1  g669(.A1(new_n854), .A2(new_n542), .A3(new_n423), .A4(new_n681), .ZN(new_n856));
  NAND2_X1  g670(.A1(new_n364), .A2(new_n636), .ZN(new_n857));
  OAI22_X1  g671(.A1(new_n855), .A2(new_n735), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  INV_X1    g672(.A(new_n725), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n853), .A2(new_n859), .ZN(new_n860));
  INV_X1    g674(.A(KEYINPUT50), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n687), .A2(new_n508), .A3(new_n699), .ZN(new_n862));
  OR3_X1    g676(.A1(new_n860), .A2(new_n861), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n861), .B1(new_n860), .B2(new_n862), .ZN(new_n864));
  AOI21_X1  g678(.A(new_n858), .B1(new_n863), .B2(new_n864), .ZN(new_n865));
  INV_X1    g679(.A(new_n860), .ZN(new_n866));
  NAND2_X1  g680(.A1(new_n697), .A2(new_n607), .ZN(new_n867));
  NOR2_X1   g681(.A1(new_n867), .A2(new_n188), .ZN(new_n868));
  OAI211_X1 g682(.A(new_n740), .B(new_n866), .C1(new_n783), .C2(new_n868), .ZN(new_n869));
  AND3_X1   g683(.A1(new_n865), .A2(new_n869), .A3(KEYINPUT51), .ZN(new_n870));
  AOI21_X1  g684(.A(KEYINPUT51), .B1(new_n865), .B2(new_n869), .ZN(new_n871));
  NAND3_X1  g685(.A1(new_n853), .A2(new_n744), .A3(new_n854), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(KEYINPUT48), .ZN(new_n873));
  NOR2_X1   g687(.A1(new_n364), .A2(new_n636), .ZN(new_n874));
  INV_X1    g688(.A(new_n874), .ZN(new_n875));
  OAI211_X1 g689(.A(G952), .B(new_n419), .C1(new_n856), .C2(new_n875), .ZN(new_n876));
  NOR3_X1   g690(.A1(new_n619), .A2(new_n627), .A3(new_n698), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n876), .B1(new_n866), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n873), .A2(new_n878), .ZN(new_n879));
  OR3_X1    g693(.A1(new_n870), .A2(new_n871), .A3(new_n879), .ZN(new_n880));
  OAI22_X1  g694(.A1(new_n852), .A2(new_n880), .B1(G952), .B2(G953), .ZN(new_n881));
  AND2_X1   g695(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n882));
  NOR2_X1   g696(.A1(new_n867), .A2(KEYINPUT49), .ZN(new_n883));
  NAND3_X1  g697(.A1(new_n542), .A2(new_n506), .A3(new_n188), .ZN(new_n884));
  NOR3_X1   g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND4_X1  g699(.A1(new_n687), .A2(new_n364), .A3(new_n690), .A4(new_n885), .ZN(new_n886));
  OAI21_X1  g700(.A(new_n881), .B1(new_n680), .B2(new_n886), .ZN(G75));
  INV_X1    g701(.A(KEYINPUT56), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n821), .A2(new_n846), .ZN(new_n889));
  NAND2_X1  g703(.A1(new_n889), .A2(G902), .ZN(new_n890));
  INV_X1    g704(.A(G210), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n888), .B1(new_n890), .B2(new_n891), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n478), .B(new_n485), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  AND2_X1   g708(.A1(new_n892), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n892), .A2(new_n894), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n265), .A2(G952), .ZN(new_n897));
  NOR3_X1   g711(.A1(new_n895), .A2(new_n896), .A3(new_n897), .ZN(G51));
  AND3_X1   g712(.A1(new_n821), .A2(new_n846), .A3(new_n847), .ZN(new_n899));
  AOI21_X1  g713(.A(new_n847), .B1(new_n821), .B2(new_n846), .ZN(new_n900));
  NOR2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  XOR2_X1   g715(.A(new_n285), .B(KEYINPUT57), .Z(new_n902));
  OAI21_X1  g716(.A(new_n606), .B1(new_n901), .B2(new_n902), .ZN(new_n903));
  OR2_X1    g717(.A1(new_n890), .A2(new_n756), .ZN(new_n904));
  AOI21_X1  g718(.A(new_n897), .B1(new_n903), .B2(new_n904), .ZN(G54));
  NAND4_X1  g719(.A1(new_n889), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n906));
  AND2_X1   g720(.A1(new_n906), .A2(new_n353), .ZN(new_n907));
  NOR2_X1   g721(.A1(new_n906), .A2(new_n353), .ZN(new_n908));
  NOR3_X1   g722(.A1(new_n907), .A2(new_n908), .A3(new_n897), .ZN(G60));
  XOR2_X1   g723(.A(KEYINPUT122), .B(KEYINPUT59), .Z(new_n910));
  XNOR2_X1  g724(.A(new_n910), .B(new_n630), .ZN(new_n911));
  NAND2_X1  g725(.A1(new_n635), .A2(new_n911), .ZN(new_n912));
  INV_X1    g726(.A(new_n847), .ZN(new_n913));
  AND3_X1   g727(.A1(new_n842), .A2(new_n830), .A3(new_n845), .ZN(new_n914));
  AOI21_X1  g728(.A(KEYINPUT53), .B1(new_n826), .B2(new_n830), .ZN(new_n915));
  OAI21_X1  g729(.A(new_n913), .B1(new_n914), .B2(new_n915), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n912), .B1(new_n916), .B2(new_n848), .ZN(new_n917));
  OAI21_X1  g731(.A(KEYINPUT123), .B1(new_n917), .B2(new_n897), .ZN(new_n918));
  INV_X1    g732(.A(new_n912), .ZN(new_n919));
  OAI21_X1  g733(.A(new_n919), .B1(new_n899), .B2(new_n900), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT123), .ZN(new_n921));
  INV_X1    g735(.A(new_n897), .ZN(new_n922));
  NAND3_X1  g736(.A1(new_n920), .A2(new_n921), .A3(new_n922), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n918), .A2(new_n923), .ZN(new_n924));
  AOI21_X1  g738(.A(new_n635), .B1(new_n852), .B2(new_n911), .ZN(new_n925));
  NOR2_X1   g739(.A1(new_n924), .A2(new_n925), .ZN(G63));
  XNOR2_X1  g740(.A(KEYINPUT124), .B(KEYINPUT61), .ZN(new_n927));
  NAND2_X1  g741(.A1(G217), .A2(G902), .ZN(new_n928));
  XNOR2_X1  g742(.A(new_n928), .B(KEYINPUT60), .ZN(new_n929));
  AOI21_X1  g743(.A(new_n929), .B1(new_n821), .B2(new_n846), .ZN(new_n930));
  OAI21_X1  g744(.A(new_n922), .B1(new_n930), .B2(new_n540), .ZN(new_n931));
  INV_X1    g745(.A(new_n929), .ZN(new_n932));
  AND3_X1   g746(.A1(new_n889), .A2(new_n660), .A3(new_n932), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n927), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND2_X1  g748(.A1(new_n934), .A2(KEYINPUT125), .ZN(new_n935));
  NOR2_X1   g749(.A1(new_n931), .A2(new_n933), .ZN(new_n936));
  NAND2_X1  g750(.A1(new_n936), .A2(KEYINPUT61), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT125), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n927), .C1(new_n931), .C2(new_n933), .ZN(new_n939));
  NAND3_X1  g753(.A1(new_n935), .A2(new_n937), .A3(new_n939), .ZN(G66));
  OAI21_X1  g754(.A(G953), .B1(new_n428), .B2(new_n482), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n830), .A2(new_n708), .A3(new_n824), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n424), .ZN(new_n943));
  OAI211_X1 g757(.A(new_n474), .B(new_n477), .C1(G898), .C2(new_n265), .ZN(new_n944));
  XNOR2_X1  g758(.A(new_n943), .B(new_n944), .ZN(G69));
  INV_X1    g759(.A(G227), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n424), .B1(new_n946), .B2(new_n671), .ZN(new_n947));
  XNOR2_X1  g761(.A(new_n947), .B(KEYINPUT127), .ZN(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND2_X1  g763(.A1(new_n552), .A2(new_n555), .ZN(new_n950));
  XOR2_X1   g764(.A(new_n950), .B(KEYINPUT126), .Z(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(new_n340), .ZN(new_n952));
  INV_X1    g766(.A(new_n786), .ZN(new_n953));
  NAND4_X1  g767(.A1(new_n764), .A2(new_n823), .A3(new_n744), .A4(new_n765), .ZN(new_n954));
  AND2_X1   g768(.A1(new_n746), .A2(new_n748), .ZN(new_n955));
  NAND4_X1  g769(.A1(new_n954), .A2(new_n773), .A3(new_n792), .A4(new_n955), .ZN(new_n956));
  OAI21_X1  g770(.A(new_n265), .B1(new_n953), .B2(new_n956), .ZN(new_n957));
  NOR2_X1   g771(.A1(new_n265), .A2(G900), .ZN(new_n958));
  INV_X1    g772(.A(new_n958), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n952), .B1(new_n957), .B2(new_n959), .ZN(new_n960));
  INV_X1    g774(.A(new_n960), .ZN(new_n961));
  INV_X1    g775(.A(new_n952), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n688), .A2(new_n792), .ZN(new_n963));
  OR2_X1    g777(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n963), .A2(KEYINPUT62), .ZN(new_n965));
  AOI211_X1 g779(.A(new_n683), .B(new_n771), .C1(new_n875), .C2(new_n817), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n597), .ZN(new_n967));
  AND2_X1   g781(.A1(new_n773), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g782(.A1(new_n964), .A2(new_n786), .A3(new_n965), .A4(new_n968), .ZN(new_n969));
  AOI21_X1  g783(.A(new_n962), .B1(new_n969), .B2(new_n265), .ZN(new_n970));
  INV_X1    g784(.A(new_n970), .ZN(new_n971));
  AOI21_X1  g785(.A(new_n949), .B1(new_n961), .B2(new_n971), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n960), .A2(new_n948), .A3(new_n970), .ZN(new_n973));
  NOR2_X1   g787(.A1(new_n972), .A2(new_n973), .ZN(G72));
  NAND2_X1  g788(.A1(new_n584), .A2(new_n563), .ZN(new_n975));
  NAND2_X1  g789(.A1(new_n969), .A2(new_n561), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n570), .B1(new_n953), .B2(new_n956), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n976), .A2(new_n977), .A3(new_n942), .ZN(new_n978));
  NAND2_X1  g792(.A1(G472), .A2(G902), .ZN(new_n979));
  XOR2_X1   g793(.A(new_n979), .B(KEYINPUT63), .Z(new_n980));
  AOI21_X1  g794(.A(new_n975), .B1(new_n978), .B2(new_n980), .ZN(new_n981));
  AND3_X1   g795(.A1(new_n836), .A2(new_n975), .A3(new_n980), .ZN(new_n982));
  NOR3_X1   g796(.A1(new_n981), .A2(new_n897), .A3(new_n982), .ZN(G57));
endmodule


