//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 1 0 0 0 0 0 0 0 1 1 1 1 0 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 0 1 1 1 0 1 1 1 0 1 1 0 0 1 1 0 0 0 0 1 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:47 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n442, new_n443, new_n444, new_n449, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n481, new_n482, new_n483, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n532, new_n533, new_n534, new_n535, new_n536, new_n537, new_n538,
    new_n539, new_n540, new_n541, new_n542, new_n543, new_n544, new_n545,
    new_n547, new_n548, new_n549, new_n550, new_n551, new_n552, new_n553,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n562, new_n563,
    new_n564, new_n565, new_n566, new_n569, new_n570, new_n572, new_n573,
    new_n574, new_n575, new_n576, new_n577, new_n578, new_n579, new_n580,
    new_n583, new_n584, new_n585, new_n586, new_n587, new_n588, new_n589,
    new_n590, new_n592, new_n593, new_n594, new_n595, new_n597, new_n598,
    new_n599, new_n600, new_n601, new_n603, new_n604, new_n605, new_n606,
    new_n607, new_n608, new_n609, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n622, new_n625,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n675, new_n676, new_n677, new_n678, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n697, new_n698, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1155, new_n1156;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  INV_X1    g016(.A(G2072), .ZN(new_n442));
  INV_X1    g017(.A(G2078), .ZN(new_n443));
  NOR2_X1   g018(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  NAND3_X1  g019(.A1(new_n444), .A2(G2084), .A3(G2090), .ZN(G158));
  NAND3_X1  g020(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g021(.A(G452), .Z(G391));
  AND2_X1   g022(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g023(.A1(G7), .A2(G661), .ZN(new_n449));
  XOR2_X1   g024(.A(new_n449), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g025(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g026(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g027(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n453));
  XNOR2_X1  g028(.A(new_n453), .B(KEYINPUT2), .ZN(new_n454));
  NAND4_X1  g029(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT64), .Z(new_n456));
  NAND2_X1  g031(.A1(new_n454), .A2(new_n456), .ZN(G261));
  INV_X1    g032(.A(G261), .ZN(G325));
  INV_X1    g033(.A(G2106), .ZN(new_n459));
  INV_X1    g034(.A(G567), .ZN(new_n460));
  OAI22_X1  g035(.A1(new_n454), .A2(new_n459), .B1(new_n460), .B2(new_n456), .ZN(new_n461));
  XOR2_X1   g036(.A(new_n461), .B(KEYINPUT65), .Z(G319));
  INV_X1    g037(.A(G2105), .ZN(new_n463));
  NAND2_X1  g038(.A1(new_n463), .A2(G2104), .ZN(new_n464));
  XOR2_X1   g039(.A(new_n464), .B(KEYINPUT68), .Z(new_n465));
  INV_X1    g040(.A(new_n465), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(G2104), .ZN(new_n468));
  OAI21_X1  g043(.A(new_n467), .B1(new_n468), .B2(KEYINPUT67), .ZN(new_n469));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n470));
  NAND3_X1  g045(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n471));
  AOI21_X1  g046(.A(G2105), .B1(new_n469), .B2(new_n471), .ZN(new_n472));
  AOI22_X1  g047(.A1(new_n466), .A2(G101), .B1(G137), .B2(new_n472), .ZN(new_n473));
  NOR2_X1   g048(.A1(new_n467), .A2(G2104), .ZN(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n475));
  OAI21_X1  g050(.A(KEYINPUT66), .B1(new_n474), .B2(new_n475), .ZN(new_n476));
  NAND2_X1  g051(.A1(new_n468), .A2(KEYINPUT3), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n467), .A2(G2104), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT66), .ZN(new_n479));
  NAND3_X1  g054(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n476), .A2(new_n480), .ZN(new_n481));
  AOI22_X1  g056(.A1(new_n481), .A2(G125), .B1(G113), .B2(G2104), .ZN(new_n482));
  OAI21_X1  g057(.A(new_n473), .B1(new_n463), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g058(.A(new_n483), .B(KEYINPUT69), .ZN(G160));
  INV_X1    g059(.A(G100), .ZN(new_n485));
  AND3_X1   g060(.A1(new_n485), .A2(new_n463), .A3(KEYINPUT72), .ZN(new_n486));
  AOI21_X1  g061(.A(KEYINPUT72), .B1(new_n485), .B2(new_n463), .ZN(new_n487));
  OAI221_X1 g062(.A(G2104), .B1(G112), .B2(new_n463), .C1(new_n486), .C2(new_n487), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n469), .A2(new_n471), .ZN(new_n489));
  OR2_X1    g064(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n490));
  NAND2_X1  g065(.A1(new_n489), .A2(KEYINPUT70), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n490), .A2(G2105), .A3(new_n491), .ZN(new_n492));
  INV_X1    g067(.A(G124), .ZN(new_n493));
  OAI21_X1  g068(.A(new_n488), .B1(new_n492), .B2(new_n493), .ZN(new_n494));
  NAND3_X1  g069(.A1(new_n490), .A2(new_n463), .A3(new_n491), .ZN(new_n495));
  XNOR2_X1  g070(.A(new_n495), .B(KEYINPUT71), .ZN(new_n496));
  AOI21_X1  g071(.A(new_n494), .B1(new_n496), .B2(G136), .ZN(G162));
  NAND3_X1  g072(.A1(new_n489), .A2(G126), .A3(G2105), .ZN(new_n498));
  OR2_X1    g073(.A1(G102), .A2(G2105), .ZN(new_n499));
  OAI211_X1 g074(.A(new_n499), .B(G2104), .C1(G114), .C2(new_n463), .ZN(new_n500));
  NAND2_X1  g075(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  INV_X1    g076(.A(G138), .ZN(new_n502));
  NOR3_X1   g077(.A1(new_n502), .A2(KEYINPUT4), .A3(G2105), .ZN(new_n503));
  AND3_X1   g078(.A1(new_n477), .A2(new_n478), .A3(new_n479), .ZN(new_n504));
  AOI21_X1  g079(.A(new_n479), .B1(new_n477), .B2(new_n478), .ZN(new_n505));
  OAI21_X1  g080(.A(new_n503), .B1(new_n504), .B2(new_n505), .ZN(new_n506));
  NAND2_X1  g081(.A1(new_n506), .A2(KEYINPUT74), .ZN(new_n507));
  INV_X1    g082(.A(KEYINPUT74), .ZN(new_n508));
  NAND3_X1  g083(.A1(new_n481), .A2(new_n508), .A3(new_n503), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n507), .A2(new_n509), .ZN(new_n510));
  AOI211_X1 g085(.A(new_n502), .B(G2105), .C1(new_n469), .C2(new_n471), .ZN(new_n511));
  INV_X1    g086(.A(KEYINPUT4), .ZN(new_n512));
  OAI21_X1  g087(.A(KEYINPUT73), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  AND3_X1   g088(.A1(new_n470), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n514));
  AOI21_X1  g089(.A(KEYINPUT3), .B1(new_n470), .B2(G2104), .ZN(new_n515));
  OAI211_X1 g090(.A(G138), .B(new_n463), .C1(new_n514), .C2(new_n515), .ZN(new_n516));
  INV_X1    g091(.A(KEYINPUT73), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n516), .A2(new_n517), .A3(KEYINPUT4), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n513), .A2(new_n518), .ZN(new_n519));
  AOI21_X1  g094(.A(new_n501), .B1(new_n510), .B2(new_n519), .ZN(G164));
  INV_X1    g095(.A(G651), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT75), .ZN(new_n523));
  OR2_X1    g098(.A1(new_n521), .A2(KEYINPUT6), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n523), .A2(new_n524), .ZN(new_n525));
  INV_X1    g100(.A(G543), .ZN(new_n526));
  INV_X1    g101(.A(KEYINPUT5), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n527), .B2(KEYINPUT77), .ZN(new_n528));
  INV_X1    g103(.A(KEYINPUT77), .ZN(new_n529));
  NAND3_X1  g104(.A1(new_n529), .A2(KEYINPUT5), .A3(G543), .ZN(new_n530));
  NAND2_X1  g105(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  INV_X1    g106(.A(new_n531), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n525), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g108(.A1(new_n533), .A2(G88), .ZN(new_n534));
  INV_X1    g109(.A(KEYINPUT76), .ZN(new_n535));
  INV_X1    g110(.A(new_n525), .ZN(new_n536));
  INV_X1    g111(.A(G50), .ZN(new_n537));
  NOR2_X1   g112(.A1(new_n537), .A2(new_n526), .ZN(new_n538));
  AOI21_X1  g113(.A(new_n535), .B1(new_n536), .B2(new_n538), .ZN(new_n539));
  NOR4_X1   g114(.A1(new_n525), .A2(KEYINPUT76), .A3(new_n537), .A4(new_n526), .ZN(new_n540));
  OAI21_X1  g115(.A(new_n534), .B1(new_n539), .B2(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n531), .A2(G62), .ZN(new_n542));
  OR2_X1    g117(.A1(new_n542), .A2(KEYINPUT78), .ZN(new_n543));
  AOI22_X1  g118(.A1(new_n542), .A2(KEYINPUT78), .B1(G75), .B2(G543), .ZN(new_n544));
  AOI21_X1  g119(.A(new_n521), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n541), .A2(new_n545), .ZN(G166));
  XOR2_X1   g121(.A(new_n531), .B(KEYINPUT79), .Z(new_n547));
  NAND3_X1  g122(.A1(new_n547), .A2(G63), .A3(G651), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n533), .A2(G89), .ZN(new_n549));
  NOR2_X1   g124(.A1(new_n525), .A2(new_n526), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G51), .ZN(new_n551));
  NAND3_X1  g126(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT7), .ZN(new_n553));
  NAND4_X1  g128(.A1(new_n548), .A2(new_n549), .A3(new_n551), .A4(new_n553), .ZN(G286));
  INV_X1    g129(.A(G286), .ZN(G168));
  AOI22_X1  g130(.A1(G52), .A2(new_n550), .B1(new_n533), .B2(G90), .ZN(new_n556));
  INV_X1    g131(.A(new_n556), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n547), .A2(G64), .ZN(new_n558));
  NAND2_X1  g133(.A1(G77), .A2(G543), .ZN(new_n559));
  AOI21_X1  g134(.A(new_n521), .B1(new_n558), .B2(new_n559), .ZN(new_n560));
  NOR2_X1   g135(.A1(new_n557), .A2(new_n560), .ZN(G171));
  AOI22_X1  g136(.A1(new_n547), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n562));
  OR2_X1    g137(.A1(new_n562), .A2(new_n521), .ZN(new_n563));
  AOI22_X1  g138(.A1(G43), .A2(new_n550), .B1(new_n533), .B2(G81), .ZN(new_n564));
  NAND2_X1  g139(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g140(.A(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n566), .A2(G860), .ZN(G153));
  NAND4_X1  g142(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g143(.A1(G1), .A2(G3), .ZN(new_n569));
  XNOR2_X1  g144(.A(new_n569), .B(KEYINPUT8), .ZN(new_n570));
  NAND4_X1  g145(.A1(G319), .A2(G483), .A3(G661), .A4(new_n570), .ZN(G188));
  NAND2_X1  g146(.A1(new_n536), .A2(new_n531), .ZN(new_n572));
  INV_X1    g147(.A(G91), .ZN(new_n573));
  AOI22_X1  g148(.A1(new_n531), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n574));
  OAI22_X1  g149(.A1(new_n572), .A2(new_n573), .B1(new_n521), .B2(new_n574), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n536), .A2(G53), .A3(G543), .ZN(new_n576));
  NAND2_X1  g151(.A1(new_n576), .A2(KEYINPUT9), .ZN(new_n577));
  INV_X1    g152(.A(KEYINPUT9), .ZN(new_n578));
  NAND3_X1  g153(.A1(new_n550), .A2(new_n578), .A3(G53), .ZN(new_n579));
  AOI21_X1  g154(.A(new_n575), .B1(new_n577), .B2(new_n579), .ZN(new_n580));
  INV_X1    g155(.A(new_n580), .ZN(G299));
  INV_X1    g156(.A(G171), .ZN(G301));
  INV_X1    g157(.A(KEYINPUT80), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n583), .B1(new_n541), .B2(new_n545), .ZN(new_n584));
  NAND2_X1  g159(.A1(new_n536), .A2(new_n538), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(KEYINPUT76), .ZN(new_n586));
  NAND3_X1  g161(.A1(new_n536), .A2(new_n535), .A3(new_n538), .ZN(new_n587));
  NAND2_X1  g162(.A1(new_n586), .A2(new_n587), .ZN(new_n588));
  INV_X1    g163(.A(new_n545), .ZN(new_n589));
  NAND4_X1  g164(.A1(new_n588), .A2(KEYINPUT80), .A3(new_n589), .A4(new_n534), .ZN(new_n590));
  AND2_X1   g165(.A1(new_n584), .A2(new_n590), .ZN(G303));
  AOI22_X1  g166(.A1(G49), .A2(new_n550), .B1(new_n533), .B2(G87), .ZN(new_n592));
  OAI21_X1  g167(.A(G651), .B1(new_n547), .B2(G74), .ZN(new_n593));
  NAND2_X1  g168(.A1(new_n592), .A2(new_n593), .ZN(new_n594));
  INV_X1    g169(.A(KEYINPUT81), .ZN(new_n595));
  XNOR2_X1  g170(.A(new_n594), .B(new_n595), .ZN(G288));
  NAND2_X1  g171(.A1(new_n533), .A2(G86), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n550), .A2(G48), .ZN(new_n598));
  AND2_X1   g173(.A1(new_n531), .A2(G61), .ZN(new_n599));
  AND2_X1   g174(.A1(G73), .A2(G543), .ZN(new_n600));
  OAI21_X1  g175(.A(G651), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NAND3_X1  g176(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(G305));
  NAND2_X1  g177(.A1(new_n547), .A2(G60), .ZN(new_n603));
  NAND2_X1  g178(.A1(G72), .A2(G543), .ZN(new_n604));
  AOI21_X1  g179(.A(new_n521), .B1(new_n603), .B2(new_n604), .ZN(new_n605));
  NAND2_X1  g180(.A1(new_n550), .A2(G47), .ZN(new_n606));
  INV_X1    g181(.A(G85), .ZN(new_n607));
  OAI21_X1  g182(.A(new_n606), .B1(new_n607), .B2(new_n572), .ZN(new_n608));
  NOR2_X1   g183(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g184(.A(new_n609), .ZN(G290));
  INV_X1    g185(.A(G868), .ZN(new_n611));
  NOR2_X1   g186(.A1(G301), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n550), .A2(G54), .ZN(new_n613));
  AOI22_X1  g188(.A1(new_n531), .A2(G66), .B1(G79), .B2(G543), .ZN(new_n614));
  AND3_X1   g189(.A1(new_n533), .A2(KEYINPUT10), .A3(G92), .ZN(new_n615));
  AOI21_X1  g190(.A(KEYINPUT10), .B1(new_n533), .B2(G92), .ZN(new_n616));
  OAI221_X1 g191(.A(new_n613), .B1(new_n521), .B2(new_n614), .C1(new_n615), .C2(new_n616), .ZN(new_n617));
  INV_X1    g192(.A(KEYINPUT82), .ZN(new_n618));
  XNOR2_X1  g193(.A(new_n617), .B(new_n618), .ZN(new_n619));
  AOI21_X1  g194(.A(new_n612), .B1(new_n619), .B2(new_n611), .ZN(G284));
  AOI21_X1  g195(.A(new_n612), .B1(new_n619), .B2(new_n611), .ZN(G321));
  NAND2_X1  g196(.A1(G286), .A2(G868), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(new_n580), .B2(G868), .ZN(G280));
  XOR2_X1   g198(.A(G280), .B(KEYINPUT83), .Z(G297));
  INV_X1    g199(.A(G559), .ZN(new_n625));
  OAI21_X1  g200(.A(new_n619), .B1(new_n625), .B2(G860), .ZN(G148));
  NOR2_X1   g201(.A1(new_n566), .A2(G868), .ZN(new_n627));
  NAND2_X1  g202(.A1(new_n619), .A2(new_n625), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n627), .B1(new_n628), .B2(G868), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT84), .Z(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n466), .A2(new_n481), .ZN(new_n632));
  XOR2_X1   g207(.A(new_n632), .B(KEYINPUT12), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XOR2_X1   g209(.A(new_n634), .B(G2100), .Z(new_n635));
  AND2_X1   g210(.A1(new_n496), .A2(G135), .ZN(new_n636));
  OAI21_X1  g211(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n637));
  INV_X1    g212(.A(G111), .ZN(new_n638));
  AOI22_X1  g213(.A1(new_n637), .A2(KEYINPUT85), .B1(new_n638), .B2(G2105), .ZN(new_n639));
  OAI21_X1  g214(.A(new_n639), .B1(KEYINPUT85), .B2(new_n637), .ZN(new_n640));
  INV_X1    g215(.A(G123), .ZN(new_n641));
  OAI21_X1  g216(.A(new_n640), .B1(new_n492), .B2(new_n641), .ZN(new_n642));
  NOR2_X1   g217(.A1(new_n636), .A2(new_n642), .ZN(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  OR2_X1    g219(.A1(new_n644), .A2(G2096), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n644), .A2(G2096), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n635), .A2(new_n645), .A3(new_n646), .ZN(G156));
  XOR2_X1   g222(.A(G2451), .B(G2454), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT16), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT87), .ZN(new_n651));
  XOR2_X1   g226(.A(new_n649), .B(new_n651), .Z(new_n652));
  INV_X1    g227(.A(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(KEYINPUT86), .B(G2438), .ZN(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(new_n656));
  XOR2_X1   g231(.A(G2427), .B(G2430), .Z(new_n657));
  AOI21_X1  g232(.A(new_n653), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n658), .B1(new_n657), .B2(new_n656), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n652), .B(new_n659), .ZN(new_n660));
  INV_X1    g235(.A(new_n660), .ZN(new_n661));
  XNOR2_X1  g236(.A(G2443), .B(G2446), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  OAI21_X1  g238(.A(G14), .B1(new_n661), .B2(new_n663), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n664), .B1(new_n663), .B2(new_n661), .ZN(G401));
  XNOR2_X1  g240(.A(G2067), .B(G2678), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n666), .B(KEYINPUT88), .ZN(new_n667));
  XOR2_X1   g242(.A(G2072), .B(G2078), .Z(new_n668));
  XOR2_X1   g243(.A(G2084), .B(G2090), .Z(new_n669));
  INV_X1    g244(.A(new_n669), .ZN(new_n670));
  NOR3_X1   g245(.A1(new_n667), .A2(new_n668), .A3(new_n670), .ZN(new_n671));
  XNOR2_X1  g246(.A(new_n671), .B(KEYINPUT18), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n667), .A2(new_n668), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n668), .B(KEYINPUT17), .ZN(new_n674));
  OAI211_X1 g249(.A(new_n673), .B(new_n670), .C1(new_n667), .C2(new_n674), .ZN(new_n675));
  NAND3_X1  g250(.A1(new_n674), .A2(new_n667), .A3(new_n669), .ZN(new_n676));
  NAND3_X1  g251(.A1(new_n672), .A2(new_n675), .A3(new_n676), .ZN(new_n677));
  XOR2_X1   g252(.A(G2096), .B(G2100), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n677), .B(new_n678), .ZN(G227));
  XNOR2_X1  g254(.A(G1971), .B(G1976), .ZN(new_n680));
  INV_X1    g255(.A(KEYINPUT19), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n680), .B(new_n681), .ZN(new_n682));
  XOR2_X1   g257(.A(G1956), .B(G2474), .Z(new_n683));
  XOR2_X1   g258(.A(G1961), .B(G1966), .Z(new_n684));
  AND2_X1   g259(.A1(new_n683), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g260(.A1(new_n682), .A2(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n686), .B(KEYINPUT20), .ZN(new_n687));
  NOR2_X1   g262(.A1(new_n683), .A2(new_n684), .ZN(new_n688));
  NOR3_X1   g263(.A1(new_n682), .A2(new_n685), .A3(new_n688), .ZN(new_n689));
  AOI21_X1  g264(.A(new_n689), .B1(new_n682), .B2(new_n688), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n687), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT89), .ZN(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT90), .ZN(new_n693));
  XOR2_X1   g268(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n694));
  XNOR2_X1  g269(.A(new_n693), .B(new_n694), .ZN(new_n695));
  XNOR2_X1  g270(.A(G1991), .B(G1996), .ZN(new_n696));
  XNOR2_X1  g271(.A(new_n695), .B(new_n696), .ZN(new_n697));
  XNOR2_X1  g272(.A(G1981), .B(G1986), .ZN(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(G229));
  INV_X1    g274(.A(G29), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G25), .ZN(new_n701));
  OR2_X1    g276(.A1(G95), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G107), .C2(new_n463), .ZN(new_n703));
  XOR2_X1   g278(.A(new_n703), .B(KEYINPUT91), .Z(new_n704));
  INV_X1    g279(.A(G119), .ZN(new_n705));
  OAI21_X1  g280(.A(new_n704), .B1(new_n492), .B2(new_n705), .ZN(new_n706));
  AOI21_X1  g281(.A(new_n706), .B1(new_n496), .B2(G131), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT92), .ZN(new_n708));
  INV_X1    g283(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n701), .B1(new_n709), .B2(new_n700), .ZN(new_n710));
  XOR2_X1   g285(.A(KEYINPUT35), .B(G1991), .Z(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  OR2_X1    g287(.A1(new_n712), .A2(KEYINPUT93), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n712), .A2(KEYINPUT93), .ZN(new_n714));
  XOR2_X1   g289(.A(KEYINPUT94), .B(G16), .Z(new_n715));
  INV_X1    g290(.A(new_n715), .ZN(new_n716));
  NOR2_X1   g291(.A1(new_n716), .A2(G24), .ZN(new_n717));
  AOI21_X1  g292(.A(new_n717), .B1(new_n609), .B2(new_n716), .ZN(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(G1986), .ZN(new_n719));
  NOR2_X1   g294(.A1(new_n716), .A2(G22), .ZN(new_n720));
  AOI21_X1  g295(.A(new_n720), .B1(G166), .B2(new_n716), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n721), .B(G1971), .ZN(new_n722));
  INV_X1    g297(.A(G16), .ZN(new_n723));
  NAND2_X1  g298(.A1(new_n723), .A2(G23), .ZN(new_n724));
  INV_X1    g299(.A(new_n594), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n724), .B1(new_n725), .B2(new_n723), .ZN(new_n726));
  XOR2_X1   g301(.A(KEYINPUT33), .B(G1976), .Z(new_n727));
  XNOR2_X1  g302(.A(new_n726), .B(new_n727), .ZN(new_n728));
  NOR2_X1   g303(.A1(G6), .A2(G16), .ZN(new_n729));
  AND3_X1   g304(.A1(new_n597), .A2(new_n598), .A3(new_n601), .ZN(new_n730));
  AOI21_X1  g305(.A(new_n729), .B1(new_n730), .B2(G16), .ZN(new_n731));
  XNOR2_X1  g306(.A(KEYINPUT32), .B(G1981), .ZN(new_n732));
  XNOR2_X1  g307(.A(new_n731), .B(new_n732), .ZN(new_n733));
  NOR3_X1   g308(.A1(new_n722), .A2(new_n728), .A3(new_n733), .ZN(new_n734));
  INV_X1    g309(.A(KEYINPUT34), .ZN(new_n735));
  AOI21_X1  g310(.A(new_n719), .B1(new_n734), .B2(new_n735), .ZN(new_n736));
  NAND3_X1  g311(.A1(new_n713), .A2(new_n714), .A3(new_n736), .ZN(new_n737));
  OR2_X1    g312(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n738));
  NAND2_X1  g313(.A1(new_n737), .A2(KEYINPUT95), .ZN(new_n739));
  OAI211_X1 g314(.A(new_n738), .B(new_n739), .C1(new_n735), .C2(new_n734), .ZN(new_n740));
  NAND2_X1  g315(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n741));
  OR2_X1    g316(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OR2_X1    g317(.A1(KEYINPUT96), .A2(KEYINPUT36), .ZN(new_n743));
  NAND3_X1  g318(.A1(new_n740), .A2(new_n741), .A3(new_n743), .ZN(new_n744));
  NAND2_X1  g319(.A1(new_n496), .A2(G139), .ZN(new_n745));
  NAND3_X1  g320(.A1(new_n463), .A2(G103), .A3(G2104), .ZN(new_n746));
  XOR2_X1   g321(.A(new_n746), .B(KEYINPUT25), .Z(new_n747));
  AOI22_X1  g322(.A1(new_n481), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n748));
  OAI211_X1 g323(.A(new_n745), .B(new_n747), .C1(new_n463), .C2(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G33), .B(new_n749), .S(G29), .Z(new_n750));
  XNOR2_X1  g325(.A(new_n750), .B(new_n442), .ZN(new_n751));
  INV_X1    g326(.A(G2084), .ZN(new_n752));
  NAND2_X1  g327(.A1(G160), .A2(G29), .ZN(new_n753));
  INV_X1    g328(.A(G34), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n754), .A2(KEYINPUT24), .ZN(new_n755));
  AOI21_X1  g330(.A(G29), .B1(new_n754), .B2(KEYINPUT24), .ZN(new_n756));
  AOI21_X1  g331(.A(new_n755), .B1(new_n756), .B2(KEYINPUT97), .ZN(new_n757));
  OAI21_X1  g332(.A(new_n757), .B1(KEYINPUT97), .B2(new_n756), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n753), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n700), .A2(G32), .ZN(new_n760));
  NAND2_X1  g335(.A1(new_n496), .A2(G141), .ZN(new_n761));
  NAND4_X1  g336(.A1(new_n490), .A2(G129), .A3(G2105), .A4(new_n491), .ZN(new_n762));
  NAND3_X1  g337(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n763));
  INV_X1    g338(.A(KEYINPUT26), .ZN(new_n764));
  NAND2_X1  g339(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  OR2_X1    g340(.A1(new_n763), .A2(new_n764), .ZN(new_n766));
  AOI22_X1  g341(.A1(new_n466), .A2(G105), .B1(new_n765), .B2(new_n766), .ZN(new_n767));
  NAND3_X1  g342(.A1(new_n761), .A2(new_n762), .A3(new_n767), .ZN(new_n768));
  INV_X1    g343(.A(new_n768), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n760), .B1(new_n769), .B2(new_n700), .ZN(new_n770));
  XOR2_X1   g345(.A(KEYINPUT27), .B(G1996), .Z(new_n771));
  OAI221_X1 g346(.A(new_n751), .B1(new_n752), .B2(new_n759), .C1(new_n770), .C2(new_n771), .ZN(new_n772));
  OR2_X1    g347(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n772), .A2(KEYINPUT98), .ZN(new_n774));
  NOR2_X1   g349(.A1(new_n716), .A2(G19), .ZN(new_n775));
  AOI21_X1  g350(.A(new_n775), .B1(new_n566), .B2(new_n716), .ZN(new_n776));
  NOR2_X1   g351(.A1(new_n776), .A2(G1341), .ZN(new_n777));
  NOR2_X1   g352(.A1(G286), .A2(new_n723), .ZN(new_n778));
  INV_X1    g353(.A(new_n778), .ZN(new_n779));
  OAI211_X1 g354(.A(new_n779), .B(KEYINPUT99), .C1(G16), .C2(G21), .ZN(new_n780));
  OAI21_X1  g355(.A(new_n780), .B1(KEYINPUT99), .B2(new_n779), .ZN(new_n781));
  AOI21_X1  g356(.A(new_n777), .B1(new_n781), .B2(G1966), .ZN(new_n782));
  XNOR2_X1  g357(.A(KEYINPUT31), .B(G11), .ZN(new_n783));
  XNOR2_X1  g358(.A(new_n783), .B(KEYINPUT100), .ZN(new_n784));
  INV_X1    g359(.A(G28), .ZN(new_n785));
  AOI21_X1  g360(.A(G29), .B1(new_n785), .B2(KEYINPUT30), .ZN(new_n786));
  OAI21_X1  g361(.A(new_n786), .B1(KEYINPUT30), .B2(new_n785), .ZN(new_n787));
  OAI211_X1 g362(.A(new_n784), .B(new_n787), .C1(new_n644), .C2(new_n700), .ZN(new_n788));
  NOR2_X1   g363(.A1(G171), .A2(new_n723), .ZN(new_n789));
  AOI21_X1  g364(.A(new_n789), .B1(G5), .B2(new_n723), .ZN(new_n790));
  INV_X1    g365(.A(new_n790), .ZN(new_n791));
  AOI21_X1  g366(.A(new_n788), .B1(new_n791), .B2(G1961), .ZN(new_n792));
  NAND2_X1  g367(.A1(new_n715), .A2(G20), .ZN(new_n793));
  XOR2_X1   g368(.A(new_n793), .B(KEYINPUT102), .Z(new_n794));
  XNOR2_X1  g369(.A(new_n794), .B(KEYINPUT23), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n795), .B1(G299), .B2(G16), .ZN(new_n796));
  XNOR2_X1  g371(.A(new_n796), .B(G1956), .ZN(new_n797));
  NAND2_X1  g372(.A1(new_n759), .A2(new_n752), .ZN(new_n798));
  NAND4_X1  g373(.A1(new_n782), .A2(new_n792), .A3(new_n797), .A4(new_n798), .ZN(new_n799));
  NAND2_X1  g374(.A1(new_n700), .A2(G26), .ZN(new_n800));
  XNOR2_X1  g375(.A(new_n800), .B(KEYINPUT28), .ZN(new_n801));
  INV_X1    g376(.A(G128), .ZN(new_n802));
  NOR2_X1   g377(.A1(new_n463), .A2(G116), .ZN(new_n803));
  OAI21_X1  g378(.A(G2104), .B1(G104), .B2(G2105), .ZN(new_n804));
  OAI22_X1  g379(.A1(new_n492), .A2(new_n802), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  AOI21_X1  g380(.A(new_n805), .B1(new_n496), .B2(G140), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n801), .B1(new_n806), .B2(new_n700), .ZN(new_n807));
  XNOR2_X1  g382(.A(new_n807), .B(G2067), .ZN(new_n808));
  INV_X1    g383(.A(G1961), .ZN(new_n809));
  AOI22_X1  g384(.A1(new_n790), .A2(new_n809), .B1(new_n776), .B2(G1341), .ZN(new_n810));
  OAI21_X1  g385(.A(new_n810), .B1(G1966), .B2(new_n781), .ZN(new_n811));
  NOR3_X1   g386(.A1(new_n799), .A2(new_n808), .A3(new_n811), .ZN(new_n812));
  NAND3_X1  g387(.A1(new_n773), .A2(new_n774), .A3(new_n812), .ZN(new_n813));
  NAND2_X1  g388(.A1(new_n700), .A2(G35), .ZN(new_n814));
  XOR2_X1   g389(.A(new_n814), .B(KEYINPUT101), .Z(new_n815));
  OAI21_X1  g390(.A(new_n815), .B1(G162), .B2(new_n700), .ZN(new_n816));
  XOR2_X1   g391(.A(new_n816), .B(KEYINPUT29), .Z(new_n817));
  INV_X1    g392(.A(G2090), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NOR2_X1   g394(.A1(G164), .A2(new_n700), .ZN(new_n820));
  AOI21_X1  g395(.A(new_n820), .B1(G27), .B2(new_n700), .ZN(new_n821));
  AOI22_X1  g396(.A1(new_n770), .A2(new_n771), .B1(new_n821), .B2(new_n443), .ZN(new_n822));
  OAI211_X1 g397(.A(new_n819), .B(new_n822), .C1(new_n443), .C2(new_n821), .ZN(new_n823));
  NOR2_X1   g398(.A1(G4), .A2(G16), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n824), .B1(new_n619), .B2(G16), .ZN(new_n825));
  INV_X1    g400(.A(G1348), .ZN(new_n826));
  XNOR2_X1  g401(.A(new_n825), .B(new_n826), .ZN(new_n827));
  OAI21_X1  g402(.A(new_n827), .B1(new_n818), .B2(new_n817), .ZN(new_n828));
  NOR3_X1   g403(.A1(new_n813), .A2(new_n823), .A3(new_n828), .ZN(new_n829));
  AND3_X1   g404(.A1(new_n742), .A2(new_n744), .A3(new_n829), .ZN(G311));
  NAND3_X1  g405(.A1(new_n742), .A2(new_n744), .A3(new_n829), .ZN(G150));
  NAND2_X1  g406(.A1(new_n550), .A2(G55), .ZN(new_n832));
  INV_X1    g407(.A(G93), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n832), .B1(new_n833), .B2(new_n572), .ZN(new_n834));
  NAND2_X1  g409(.A1(new_n547), .A2(G67), .ZN(new_n835));
  INV_X1    g410(.A(G80), .ZN(new_n836));
  OAI21_X1  g411(.A(new_n835), .B1(new_n836), .B2(new_n526), .ZN(new_n837));
  AOI21_X1  g412(.A(new_n834), .B1(G651), .B2(new_n837), .ZN(new_n838));
  XNOR2_X1  g413(.A(new_n838), .B(KEYINPUT104), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n839), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT37), .Z(new_n841));
  NAND2_X1  g416(.A1(new_n839), .A2(new_n565), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n566), .A2(new_n838), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XNOR2_X1  g419(.A(new_n844), .B(KEYINPUT105), .ZN(new_n845));
  INV_X1    g420(.A(new_n619), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n846), .A2(new_n625), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n845), .B(new_n847), .ZN(new_n848));
  XOR2_X1   g423(.A(KEYINPUT103), .B(KEYINPUT38), .Z(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  AND2_X1   g425(.A1(new_n850), .A2(KEYINPUT39), .ZN(new_n851));
  INV_X1    g426(.A(G860), .ZN(new_n852));
  OAI21_X1  g427(.A(new_n852), .B1(new_n850), .B2(KEYINPUT39), .ZN(new_n853));
  OAI21_X1  g428(.A(new_n841), .B1(new_n851), .B2(new_n853), .ZN(G145));
  NOR2_X1   g429(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n855));
  INV_X1    g430(.A(new_n501), .ZN(new_n856));
  INV_X1    g431(.A(KEYINPUT106), .ZN(new_n857));
  AND3_X1   g432(.A1(new_n510), .A2(new_n519), .A3(new_n857), .ZN(new_n858));
  AOI21_X1  g433(.A(new_n857), .B1(new_n510), .B2(new_n519), .ZN(new_n859));
  OAI21_X1  g434(.A(new_n856), .B1(new_n858), .B2(new_n859), .ZN(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n806), .ZN(new_n861));
  AOI21_X1  g436(.A(new_n855), .B1(new_n861), .B2(new_n768), .ZN(new_n862));
  OAI21_X1  g437(.A(new_n862), .B1(new_n768), .B2(new_n861), .ZN(new_n863));
  NAND2_X1  g438(.A1(new_n749), .A2(KEYINPUT107), .ZN(new_n864));
  XOR2_X1   g439(.A(new_n863), .B(new_n864), .Z(new_n865));
  INV_X1    g440(.A(G130), .ZN(new_n866));
  NOR2_X1   g441(.A1(new_n463), .A2(G118), .ZN(new_n867));
  OAI21_X1  g442(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n868));
  OAI22_X1  g443(.A1(new_n492), .A2(new_n866), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  AOI21_X1  g444(.A(new_n869), .B1(new_n496), .B2(G142), .ZN(new_n870));
  XOR2_X1   g445(.A(new_n870), .B(new_n633), .Z(new_n871));
  XNOR2_X1  g446(.A(new_n871), .B(new_n708), .ZN(new_n872));
  INV_X1    g447(.A(new_n872), .ZN(new_n873));
  AND2_X1   g448(.A1(new_n865), .A2(new_n873), .ZN(new_n874));
  NOR2_X1   g449(.A1(new_n865), .A2(new_n873), .ZN(new_n875));
  XOR2_X1   g450(.A(new_n643), .B(G160), .Z(new_n876));
  XNOR2_X1  g451(.A(new_n876), .B(G162), .ZN(new_n877));
  INV_X1    g452(.A(new_n877), .ZN(new_n878));
  OR3_X1    g453(.A1(new_n874), .A2(new_n875), .A3(new_n878), .ZN(new_n879));
  INV_X1    g454(.A(G37), .ZN(new_n880));
  OAI21_X1  g455(.A(new_n878), .B1(new_n874), .B2(new_n875), .ZN(new_n881));
  NAND3_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n881), .ZN(new_n882));
  XNOR2_X1  g457(.A(new_n882), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g458(.A1(new_n839), .A2(new_n611), .ZN(new_n884));
  XOR2_X1   g459(.A(new_n844), .B(new_n628), .Z(new_n885));
  XNOR2_X1  g460(.A(G299), .B(new_n617), .ZN(new_n886));
  XOR2_X1   g461(.A(new_n886), .B(KEYINPUT41), .Z(new_n887));
  NAND2_X1  g462(.A1(new_n885), .A2(new_n887), .ZN(new_n888));
  INV_X1    g463(.A(new_n886), .ZN(new_n889));
  OAI21_X1  g464(.A(new_n888), .B1(new_n889), .B2(new_n885), .ZN(new_n890));
  XNOR2_X1  g465(.A(new_n890), .B(KEYINPUT42), .ZN(new_n891));
  XNOR2_X1  g466(.A(G166), .B(new_n609), .ZN(new_n892));
  XNOR2_X1  g467(.A(new_n594), .B(new_n730), .ZN(new_n893));
  XNOR2_X1  g468(.A(new_n892), .B(new_n893), .ZN(new_n894));
  XNOR2_X1  g469(.A(new_n891), .B(new_n894), .ZN(new_n895));
  OAI21_X1  g470(.A(new_n884), .B1(new_n895), .B2(new_n611), .ZN(G295));
  OAI21_X1  g471(.A(new_n884), .B1(new_n895), .B2(new_n611), .ZN(G331));
  XNOR2_X1  g472(.A(G171), .B(G286), .ZN(new_n898));
  XNOR2_X1  g473(.A(new_n844), .B(new_n898), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n899), .A2(new_n889), .ZN(new_n900));
  NOR2_X1   g475(.A1(new_n899), .A2(new_n887), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n900), .A2(new_n901), .A3(new_n894), .ZN(new_n902));
  OAI21_X1  g477(.A(new_n894), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n902), .A2(new_n880), .A3(new_n903), .ZN(new_n904));
  NAND2_X1  g479(.A1(new_n904), .A2(KEYINPUT43), .ZN(new_n905));
  INV_X1    g480(.A(KEYINPUT43), .ZN(new_n906));
  NAND4_X1  g481(.A1(new_n902), .A2(new_n906), .A3(new_n880), .A4(new_n903), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n905), .A2(KEYINPUT44), .A3(new_n907), .ZN(new_n908));
  INV_X1    g483(.A(KEYINPUT108), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n905), .A2(new_n909), .A3(new_n907), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n904), .A2(KEYINPUT108), .A3(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n910), .A2(new_n911), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n908), .B1(new_n912), .B2(KEYINPUT44), .ZN(G397));
  NAND2_X1  g488(.A1(G286), .A2(G8), .ZN(new_n914));
  XOR2_X1   g489(.A(new_n914), .B(KEYINPUT123), .Z(new_n915));
  INV_X1    g490(.A(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT112), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n508), .B1(new_n481), .B2(new_n503), .ZN(new_n918));
  INV_X1    g493(.A(new_n503), .ZN(new_n919));
  AOI211_X1 g494(.A(KEYINPUT74), .B(new_n919), .C1(new_n476), .C2(new_n480), .ZN(new_n920));
  AOI211_X1 g495(.A(KEYINPUT73), .B(new_n512), .C1(new_n472), .C2(G138), .ZN(new_n921));
  AOI21_X1  g496(.A(new_n517), .B1(new_n516), .B2(KEYINPUT4), .ZN(new_n922));
  OAI22_X1  g497(.A1(new_n918), .A2(new_n920), .B1(new_n921), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n923), .A2(KEYINPUT106), .ZN(new_n924));
  NAND3_X1  g499(.A1(new_n510), .A2(new_n519), .A3(new_n857), .ZN(new_n925));
  AOI21_X1  g500(.A(new_n501), .B1(new_n924), .B2(new_n925), .ZN(new_n926));
  OAI21_X1  g501(.A(new_n917), .B1(new_n926), .B2(G1384), .ZN(new_n927));
  INV_X1    g502(.A(G1384), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n860), .A2(KEYINPUT112), .A3(new_n928), .ZN(new_n929));
  INV_X1    g504(.A(KEYINPUT50), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n927), .A2(new_n929), .A3(new_n930), .ZN(new_n931));
  NOR2_X1   g506(.A1(G164), .A2(G1384), .ZN(new_n932));
  NAND2_X1  g507(.A1(new_n932), .A2(KEYINPUT50), .ZN(new_n933));
  NAND2_X1  g508(.A1(new_n931), .A2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(G40), .ZN(new_n935));
  NOR2_X1   g510(.A1(new_n483), .A2(new_n935), .ZN(new_n936));
  INV_X1    g511(.A(new_n936), .ZN(new_n937));
  NOR2_X1   g512(.A1(new_n937), .A2(G2084), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n934), .A2(KEYINPUT114), .A3(new_n938), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT45), .ZN(new_n940));
  NAND3_X1  g515(.A1(new_n927), .A2(new_n929), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n937), .B1(new_n932), .B2(KEYINPUT45), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(G1966), .ZN(new_n944));
  NAND2_X1  g519(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n939), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(new_n938), .ZN(new_n947));
  AOI21_X1  g522(.A(new_n947), .B1(new_n931), .B2(new_n933), .ZN(new_n948));
  NOR2_X1   g523(.A1(new_n948), .A2(KEYINPUT114), .ZN(new_n949));
  OAI21_X1  g524(.A(new_n916), .B1(new_n946), .B2(new_n949), .ZN(new_n950));
  INV_X1    g525(.A(G8), .ZN(new_n951));
  AOI22_X1  g526(.A1(new_n948), .A2(KEYINPUT114), .B1(new_n943), .B2(new_n944), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n934), .A2(new_n938), .ZN(new_n953));
  INV_X1    g528(.A(KEYINPUT114), .ZN(new_n954));
  NAND2_X1  g529(.A1(new_n953), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n951), .B1(new_n952), .B2(new_n955), .ZN(new_n956));
  OAI211_X1 g531(.A(new_n950), .B(KEYINPUT51), .C1(new_n956), .C2(new_n916), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT124), .ZN(new_n958));
  OAI21_X1  g533(.A(G8), .B1(new_n946), .B2(new_n949), .ZN(new_n959));
  INV_X1    g534(.A(KEYINPUT51), .ZN(new_n960));
  NAND3_X1  g535(.A1(new_n959), .A2(new_n960), .A3(new_n915), .ZN(new_n961));
  AND3_X1   g536(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n962));
  AOI21_X1  g537(.A(new_n958), .B1(new_n957), .B2(new_n961), .ZN(new_n963));
  OAI21_X1  g538(.A(KEYINPUT62), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  NAND2_X1  g539(.A1(new_n950), .A2(KEYINPUT51), .ZN(new_n965));
  NAND2_X1  g540(.A1(new_n952), .A2(new_n955), .ZN(new_n966));
  AOI21_X1  g541(.A(new_n916), .B1(new_n966), .B2(G8), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n961), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND2_X1  g543(.A1(new_n968), .A2(KEYINPUT124), .ZN(new_n969));
  INV_X1    g544(.A(KEYINPUT62), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n957), .A2(new_n958), .A3(new_n961), .ZN(new_n971));
  NAND3_X1  g546(.A1(new_n969), .A2(new_n970), .A3(new_n971), .ZN(new_n972));
  INV_X1    g547(.A(KEYINPUT53), .ZN(new_n973));
  NOR2_X1   g548(.A1(new_n973), .A2(G2078), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n941), .A2(new_n942), .A3(new_n974), .ZN(new_n975));
  AOI21_X1  g550(.A(new_n937), .B1(new_n931), .B2(new_n933), .ZN(new_n976));
  OAI21_X1  g551(.A(new_n975), .B1(new_n976), .B2(G1961), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n977), .A2(KEYINPUT125), .ZN(new_n978));
  INV_X1    g553(.A(KEYINPUT125), .ZN(new_n979));
  OAI211_X1 g554(.A(new_n979), .B(new_n975), .C1(new_n976), .C2(G1961), .ZN(new_n980));
  NAND2_X1  g555(.A1(new_n978), .A2(new_n980), .ZN(new_n981));
  XOR2_X1   g556(.A(KEYINPUT109), .B(G1384), .Z(new_n982));
  NAND2_X1  g557(.A1(new_n924), .A2(new_n925), .ZN(new_n983));
  AOI21_X1  g558(.A(new_n982), .B1(new_n983), .B2(new_n856), .ZN(new_n984));
  AOI21_X1  g559(.A(new_n937), .B1(new_n984), .B2(KEYINPUT45), .ZN(new_n985));
  OAI21_X1  g560(.A(new_n940), .B1(G164), .B2(G1384), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n985), .A2(new_n986), .ZN(new_n987));
  OAI21_X1  g562(.A(new_n973), .B1(new_n987), .B2(G2078), .ZN(new_n988));
  AOI21_X1  g563(.A(G301), .B1(new_n981), .B2(new_n988), .ZN(new_n989));
  NAND3_X1  g564(.A1(new_n927), .A2(new_n929), .A3(KEYINPUT50), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n937), .B1(new_n932), .B2(new_n930), .ZN(new_n991));
  NAND3_X1  g566(.A1(new_n990), .A2(new_n818), .A3(new_n991), .ZN(new_n992));
  AND2_X1   g567(.A1(new_n985), .A2(new_n986), .ZN(new_n993));
  OAI21_X1  g568(.A(new_n992), .B1(new_n993), .B2(G1971), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(G8), .ZN(new_n995));
  NAND3_X1  g570(.A1(new_n584), .A2(new_n590), .A3(G8), .ZN(new_n996));
  INV_X1    g571(.A(KEYINPUT55), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  NAND4_X1  g573(.A1(new_n584), .A2(new_n590), .A3(KEYINPUT55), .A4(G8), .ZN(new_n999));
  AND2_X1   g574(.A1(new_n998), .A2(new_n999), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n995), .A2(new_n1000), .ZN(new_n1001));
  NAND2_X1  g576(.A1(new_n927), .A2(new_n929), .ZN(new_n1002));
  AOI21_X1  g577(.A(new_n951), .B1(new_n1002), .B2(new_n936), .ZN(new_n1003));
  NAND2_X1  g578(.A1(new_n725), .A2(G1976), .ZN(new_n1004));
  INV_X1    g579(.A(G1976), .ZN(new_n1005));
  AOI21_X1  g580(.A(KEYINPUT52), .B1(G288), .B2(new_n1005), .ZN(new_n1006));
  NAND3_X1  g581(.A1(new_n1003), .A2(new_n1004), .A3(new_n1006), .ZN(new_n1007));
  NAND2_X1  g582(.A1(new_n1002), .A2(new_n936), .ZN(new_n1008));
  INV_X1    g583(.A(G1981), .ZN(new_n1009));
  NAND2_X1  g584(.A1(new_n730), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(G305), .A2(G1981), .ZN(new_n1011));
  AND2_X1   g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  OR2_X1    g587(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1012), .A2(KEYINPUT49), .ZN(new_n1014));
  NAND4_X1  g589(.A1(new_n1008), .A2(new_n1013), .A3(G8), .A4(new_n1014), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1007), .A2(new_n1015), .ZN(new_n1016));
  INV_X1    g591(.A(KEYINPUT52), .ZN(new_n1017));
  AOI21_X1  g592(.A(new_n1017), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1018));
  NOR2_X1   g593(.A1(new_n1016), .A2(new_n1018), .ZN(new_n1019));
  INV_X1    g594(.A(KEYINPUT113), .ZN(new_n1020));
  AND3_X1   g595(.A1(new_n998), .A2(new_n1020), .A3(new_n999), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n1020), .B1(new_n998), .B2(new_n999), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1021), .A2(new_n1022), .ZN(new_n1023));
  NOR2_X1   g598(.A1(new_n993), .A2(G1971), .ZN(new_n1024));
  AOI211_X1 g599(.A(G2090), .B(new_n937), .C1(new_n931), .C2(new_n933), .ZN(new_n1025));
  OAI211_X1 g600(.A(new_n1023), .B(G8), .C1(new_n1024), .C2(new_n1025), .ZN(new_n1026));
  AND2_X1   g601(.A1(new_n1019), .A2(new_n1026), .ZN(new_n1027));
  AND3_X1   g602(.A1(new_n989), .A2(new_n1001), .A3(new_n1027), .ZN(new_n1028));
  NAND3_X1  g603(.A1(new_n964), .A2(new_n972), .A3(new_n1028), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n1030));
  NAND2_X1  g605(.A1(new_n934), .A2(new_n936), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(new_n809), .ZN(new_n1032));
  OAI211_X1 g607(.A(new_n985), .B(new_n974), .C1(KEYINPUT45), .C2(new_n984), .ZN(new_n1033));
  AND2_X1   g608(.A1(new_n1033), .A2(KEYINPUT126), .ZN(new_n1034));
  NOR2_X1   g609(.A1(new_n1033), .A2(KEYINPUT126), .ZN(new_n1035));
  OAI211_X1 g610(.A(new_n1032), .B(new_n988), .C1(new_n1034), .C2(new_n1035), .ZN(new_n1036));
  NOR2_X1   g611(.A1(new_n1036), .A2(G171), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1030), .B1(new_n989), .B2(new_n1037), .ZN(new_n1038));
  NAND3_X1  g613(.A1(new_n1001), .A2(new_n1019), .A3(new_n1026), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n981), .A2(G301), .A3(new_n988), .ZN(new_n1040));
  AOI21_X1  g615(.A(new_n1030), .B1(new_n1036), .B2(G171), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1039), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  AND2_X1   g617(.A1(new_n1038), .A2(new_n1042), .ZN(new_n1043));
  INV_X1    g618(.A(KEYINPUT122), .ZN(new_n1044));
  INV_X1    g619(.A(KEYINPUT57), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1045), .B1(new_n580), .B2(KEYINPUT117), .ZN(new_n1046));
  INV_X1    g621(.A(KEYINPUT120), .ZN(new_n1047));
  INV_X1    g622(.A(KEYINPUT117), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n577), .A2(new_n579), .ZN(new_n1049));
  OAI211_X1 g624(.A(new_n1048), .B(KEYINPUT57), .C1(new_n1049), .C2(new_n575), .ZN(new_n1050));
  AND3_X1   g625(.A1(new_n1046), .A2(new_n1047), .A3(new_n1050), .ZN(new_n1051));
  AOI21_X1  g626(.A(new_n1047), .B1(new_n1046), .B2(new_n1050), .ZN(new_n1052));
  NOR2_X1   g627(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1053));
  AOI21_X1  g628(.A(G1956), .B1(new_n990), .B2(new_n991), .ZN(new_n1054));
  INV_X1    g629(.A(new_n982), .ZN(new_n1055));
  NAND3_X1  g630(.A1(new_n860), .A2(KEYINPUT45), .A3(new_n1055), .ZN(new_n1056));
  XNOR2_X1  g631(.A(KEYINPUT118), .B(KEYINPUT56), .ZN(new_n1057));
  XNOR2_X1  g632(.A(new_n1057), .B(new_n442), .ZN(new_n1058));
  AND4_X1   g633(.A1(new_n936), .A2(new_n1056), .A3(new_n986), .A4(new_n1058), .ZN(new_n1059));
  OAI21_X1  g634(.A(new_n1053), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1060));
  NAND2_X1  g635(.A1(new_n1060), .A2(KEYINPUT61), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1046), .A2(new_n1050), .ZN(new_n1062));
  NOR3_X1   g637(.A1(new_n1054), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1063));
  OAI21_X1  g638(.A(new_n1044), .B1(new_n1061), .B2(new_n1063), .ZN(new_n1064));
  OR3_X1    g639(.A1(new_n1054), .A2(new_n1059), .A3(new_n1062), .ZN(new_n1065));
  NAND4_X1  g640(.A1(new_n1065), .A2(KEYINPUT122), .A3(KEYINPUT61), .A4(new_n1060), .ZN(new_n1066));
  AND2_X1   g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1062), .B1(new_n1054), .B2(new_n1059), .ZN(new_n1068));
  AOI21_X1  g643(.A(KEYINPUT61), .B1(new_n1065), .B2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(G1996), .ZN(new_n1070));
  NAND4_X1  g645(.A1(new_n985), .A2(KEYINPUT121), .A3(new_n1070), .A4(new_n986), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n1056), .A2(new_n1070), .A3(new_n986), .A4(new_n936), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1072), .A2(new_n1073), .ZN(new_n1074));
  NAND2_X1  g649(.A1(new_n1071), .A2(new_n1074), .ZN(new_n1075));
  AOI21_X1  g650(.A(KEYINPUT119), .B1(new_n1002), .B2(new_n936), .ZN(new_n1076));
  INV_X1    g651(.A(KEYINPUT119), .ZN(new_n1077));
  AOI211_X1 g652(.A(new_n1077), .B(new_n937), .C1(new_n927), .C2(new_n929), .ZN(new_n1078));
  NOR2_X1   g653(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1079));
  XOR2_X1   g654(.A(KEYINPUT58), .B(G1341), .Z(new_n1080));
  AOI21_X1  g655(.A(new_n1075), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  OAI21_X1  g656(.A(KEYINPUT59), .B1(new_n1081), .B2(new_n565), .ZN(new_n1082));
  INV_X1    g657(.A(KEYINPUT59), .ZN(new_n1083));
  INV_X1    g658(.A(new_n1080), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1076), .A2(new_n1078), .A3(new_n1084), .ZN(new_n1085));
  OAI211_X1 g660(.A(new_n1083), .B(new_n566), .C1(new_n1085), .C2(new_n1075), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1069), .B1(new_n1082), .B2(new_n1086), .ZN(new_n1087));
  NAND2_X1  g662(.A1(new_n1031), .A2(new_n826), .ZN(new_n1088));
  INV_X1    g663(.A(G2067), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1089), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1090));
  NAND2_X1  g665(.A1(new_n1088), .A2(new_n1090), .ZN(new_n1091));
  INV_X1    g666(.A(KEYINPUT60), .ZN(new_n1092));
  OAI21_X1  g667(.A(new_n846), .B1(new_n1091), .B2(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n1091), .A2(new_n1092), .ZN(new_n1094));
  NAND4_X1  g669(.A1(new_n1088), .A2(new_n1090), .A3(KEYINPUT60), .A4(new_n619), .ZN(new_n1095));
  NAND3_X1  g670(.A1(new_n1093), .A2(new_n1094), .A3(new_n1095), .ZN(new_n1096));
  NAND3_X1  g671(.A1(new_n1067), .A2(new_n1087), .A3(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(new_n1060), .ZN(new_n1098));
  AOI21_X1  g673(.A(new_n846), .B1(new_n1088), .B2(new_n1090), .ZN(new_n1099));
  AOI21_X1  g674(.A(new_n1098), .B1(new_n1099), .B2(new_n1065), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1097), .A2(new_n1100), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n969), .A2(new_n971), .ZN(new_n1102));
  NAND3_X1  g677(.A1(new_n1043), .A2(new_n1101), .A3(new_n1102), .ZN(new_n1103));
  NAND2_X1  g678(.A1(new_n956), .A2(G168), .ZN(new_n1104));
  INV_X1    g679(.A(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(KEYINPUT63), .ZN(new_n1106));
  OAI21_X1  g681(.A(G8), .B1(new_n1024), .B2(new_n1025), .ZN(new_n1107));
  AOI21_X1  g682(.A(new_n1106), .B1(new_n1107), .B2(new_n1000), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1105), .A2(new_n1027), .A3(new_n1108), .ZN(new_n1109));
  INV_X1    g684(.A(KEYINPUT116), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  OAI21_X1  g686(.A(new_n1106), .B1(new_n1039), .B2(new_n1104), .ZN(new_n1112));
  NAND2_X1  g687(.A1(new_n1112), .A2(KEYINPUT115), .ZN(new_n1113));
  INV_X1    g688(.A(KEYINPUT115), .ZN(new_n1114));
  OAI211_X1 g689(.A(new_n1114), .B(new_n1106), .C1(new_n1039), .C2(new_n1104), .ZN(new_n1115));
  NAND4_X1  g690(.A1(new_n1105), .A2(new_n1027), .A3(KEYINPUT116), .A4(new_n1108), .ZN(new_n1116));
  NAND4_X1  g691(.A1(new_n1111), .A2(new_n1113), .A3(new_n1115), .A4(new_n1116), .ZN(new_n1117));
  NOR3_X1   g692(.A1(new_n1026), .A2(new_n1018), .A3(new_n1016), .ZN(new_n1118));
  INV_X1    g693(.A(G288), .ZN(new_n1119));
  NAND3_X1  g694(.A1(new_n1015), .A2(new_n1005), .A3(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1120), .A2(new_n1010), .ZN(new_n1121));
  AOI21_X1  g696(.A(new_n1118), .B1(new_n1003), .B2(new_n1121), .ZN(new_n1122));
  NAND4_X1  g697(.A1(new_n1029), .A2(new_n1103), .A3(new_n1117), .A4(new_n1122), .ZN(new_n1123));
  INV_X1    g698(.A(new_n984), .ZN(new_n1124));
  NAND3_X1  g699(.A1(new_n1124), .A2(new_n940), .A3(new_n936), .ZN(new_n1125));
  INV_X1    g700(.A(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n708), .B(new_n711), .ZN(new_n1127));
  XOR2_X1   g702(.A(new_n1127), .B(KEYINPUT111), .Z(new_n1128));
  XNOR2_X1  g703(.A(new_n768), .B(new_n1070), .ZN(new_n1129));
  XNOR2_X1  g704(.A(new_n806), .B(G2067), .ZN(new_n1130));
  AND2_X1   g705(.A1(new_n1129), .A2(new_n1130), .ZN(new_n1131));
  NAND2_X1  g706(.A1(new_n1128), .A2(new_n1131), .ZN(new_n1132));
  OR2_X1    g707(.A1(G290), .A2(G1986), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT110), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  NAND2_X1  g710(.A1(G290), .A2(G1986), .ZN(new_n1136));
  XNOR2_X1  g711(.A(new_n1135), .B(new_n1136), .ZN(new_n1137));
  OAI21_X1  g712(.A(new_n1126), .B1(new_n1132), .B2(new_n1137), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1123), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1125), .B1(new_n1130), .B2(new_n769), .ZN(new_n1140));
  OR3_X1    g715(.A1(new_n1125), .A2(KEYINPUT46), .A3(G1996), .ZN(new_n1141));
  OAI21_X1  g716(.A(KEYINPUT46), .B1(new_n1125), .B2(G1996), .ZN(new_n1142));
  AOI21_X1  g717(.A(new_n1140), .B1(new_n1141), .B2(new_n1142), .ZN(new_n1143));
  XNOR2_X1  g718(.A(new_n1143), .B(KEYINPUT47), .ZN(new_n1144));
  NAND3_X1  g719(.A1(new_n1131), .A2(new_n711), .A3(new_n709), .ZN(new_n1145));
  NAND2_X1  g720(.A1(new_n806), .A2(new_n1089), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1125), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1132), .A2(new_n1126), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1125), .A2(new_n1133), .ZN(new_n1149));
  XOR2_X1   g724(.A(new_n1149), .B(KEYINPUT48), .Z(new_n1150));
  AOI211_X1 g725(.A(new_n1144), .B(new_n1147), .C1(new_n1148), .C2(new_n1150), .ZN(new_n1151));
  XNOR2_X1  g726(.A(new_n1151), .B(KEYINPUT127), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n1139), .A2(new_n1152), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g728(.A(G319), .ZN(new_n1155));
  NOR4_X1   g729(.A1(G229), .A2(new_n1155), .A3(G401), .A4(G227), .ZN(new_n1156));
  NAND4_X1  g730(.A1(new_n910), .A2(new_n1156), .A3(new_n882), .A4(new_n911), .ZN(G225));
  INV_X1    g731(.A(G225), .ZN(G308));
endmodule


