

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584;

  XNOR2_X1 U319 ( .A(n342), .B(n341), .ZN(n346) );
  XOR2_X1 U320 ( .A(G78GAT), .B(KEYINPUT13), .Z(n287) );
  XOR2_X1 U321 ( .A(G43GAT), .B(KEYINPUT83), .Z(n288) );
  XNOR2_X1 U322 ( .A(KEYINPUT48), .B(KEYINPUT112), .ZN(n389) );
  XNOR2_X1 U323 ( .A(n340), .B(n406), .ZN(n341) );
  XNOR2_X1 U324 ( .A(n436), .B(n288), .ZN(n437) );
  AND2_X1 U325 ( .A1(n512), .A2(n411), .ZN(n567) );
  XNOR2_X1 U326 ( .A(n390), .B(n389), .ZN(n522) );
  XNOR2_X1 U327 ( .A(n438), .B(n437), .ZN(n439) );
  INV_X1 U328 ( .A(G169GAT), .ZN(n444) );
  XOR2_X1 U329 ( .A(n442), .B(n441), .Z(n516) );
  XNOR2_X1 U330 ( .A(n466), .B(n465), .ZN(n493) );
  XNOR2_X1 U331 ( .A(n444), .B(KEYINPUT122), .ZN(n445) );
  XNOR2_X1 U332 ( .A(G43GAT), .B(KEYINPUT40), .ZN(n471) );
  XNOR2_X1 U333 ( .A(n446), .B(n445), .ZN(G1348GAT) );
  XNOR2_X1 U334 ( .A(n472), .B(n471), .ZN(G1330GAT) );
  XOR2_X1 U335 ( .A(G141GAT), .B(G113GAT), .Z(n290) );
  XNOR2_X1 U336 ( .A(G36GAT), .B(G50GAT), .ZN(n289) );
  XNOR2_X1 U337 ( .A(n290), .B(n289), .ZN(n294) );
  XOR2_X1 U338 ( .A(KEYINPUT72), .B(KEYINPUT70), .Z(n292) );
  XNOR2_X1 U339 ( .A(KEYINPUT69), .B(KEYINPUT68), .ZN(n291) );
  XNOR2_X1 U340 ( .A(n292), .B(n291), .ZN(n293) );
  XOR2_X1 U341 ( .A(n294), .B(n293), .Z(n299) );
  XOR2_X1 U342 ( .A(KEYINPUT29), .B(KEYINPUT30), .Z(n296) );
  NAND2_X1 U343 ( .A1(G229GAT), .A2(G233GAT), .ZN(n295) );
  XNOR2_X1 U344 ( .A(n296), .B(n295), .ZN(n297) );
  XNOR2_X1 U345 ( .A(KEYINPUT67), .B(n297), .ZN(n298) );
  XNOR2_X1 U346 ( .A(n299), .B(n298), .ZN(n303) );
  XOR2_X1 U347 ( .A(G22GAT), .B(G8GAT), .Z(n301) );
  XNOR2_X1 U348 ( .A(G169GAT), .B(G197GAT), .ZN(n300) );
  XNOR2_X1 U349 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U350 ( .A(n303), .B(n302), .Z(n308) );
  XOR2_X1 U351 ( .A(G29GAT), .B(G43GAT), .Z(n305) );
  XNOR2_X1 U352 ( .A(KEYINPUT7), .B(KEYINPUT8), .ZN(n304) );
  XNOR2_X1 U353 ( .A(n305), .B(n304), .ZN(n379) );
  XNOR2_X1 U354 ( .A(G1GAT), .B(KEYINPUT71), .ZN(n306) );
  XNOR2_X1 U355 ( .A(n306), .B(G15GAT), .ZN(n351) );
  XNOR2_X1 U356 ( .A(n379), .B(n351), .ZN(n307) );
  XOR2_X1 U357 ( .A(n308), .B(n307), .Z(n495) );
  INV_X1 U358 ( .A(n495), .ZN(n568) );
  XOR2_X1 U359 ( .A(G120GAT), .B(G148GAT), .Z(n344) );
  XOR2_X1 U360 ( .A(G57GAT), .B(G162GAT), .Z(n310) );
  XNOR2_X1 U361 ( .A(G29GAT), .B(G85GAT), .ZN(n309) );
  XNOR2_X1 U362 ( .A(n310), .B(n309), .ZN(n311) );
  XOR2_X1 U363 ( .A(n344), .B(n311), .Z(n313) );
  NAND2_X1 U364 ( .A1(G225GAT), .A2(G233GAT), .ZN(n312) );
  XNOR2_X1 U365 ( .A(n313), .B(n312), .ZN(n316) );
  XOR2_X1 U366 ( .A(KEYINPUT3), .B(KEYINPUT2), .Z(n315) );
  XNOR2_X1 U367 ( .A(G141GAT), .B(KEYINPUT86), .ZN(n314) );
  XNOR2_X1 U368 ( .A(n315), .B(n314), .ZN(n417) );
  XOR2_X1 U369 ( .A(n316), .B(n417), .Z(n318) );
  XNOR2_X1 U370 ( .A(G1GAT), .B(KEYINPUT4), .ZN(n317) );
  XNOR2_X1 U371 ( .A(n318), .B(n317), .ZN(n322) );
  XOR2_X1 U372 ( .A(KEYINPUT88), .B(G155GAT), .Z(n320) );
  XNOR2_X1 U373 ( .A(KEYINPUT87), .B(KEYINPUT1), .ZN(n319) );
  XNOR2_X1 U374 ( .A(n320), .B(n319), .ZN(n321) );
  XOR2_X1 U375 ( .A(n322), .B(n321), .Z(n330) );
  XOR2_X1 U376 ( .A(KEYINPUT82), .B(G134GAT), .Z(n324) );
  XNOR2_X1 U377 ( .A(KEYINPUT0), .B(G127GAT), .ZN(n323) );
  XNOR2_X1 U378 ( .A(n324), .B(n323), .ZN(n325) );
  XNOR2_X1 U379 ( .A(G113GAT), .B(n325), .ZN(n441) );
  XOR2_X1 U380 ( .A(KEYINPUT6), .B(KEYINPUT90), .Z(n327) );
  XNOR2_X1 U381 ( .A(KEYINPUT89), .B(KEYINPUT5), .ZN(n326) );
  XNOR2_X1 U382 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U383 ( .A(n441), .B(n328), .Z(n329) );
  XOR2_X1 U384 ( .A(n330), .B(n329), .Z(n512) );
  INV_X1 U385 ( .A(KEYINPUT47), .ZN(n382) );
  INV_X1 U386 ( .A(G71GAT), .ZN(n333) );
  XNOR2_X1 U387 ( .A(G57GAT), .B(KEYINPUT73), .ZN(n331) );
  XNOR2_X1 U388 ( .A(n287), .B(n331), .ZN(n332) );
  XNOR2_X1 U389 ( .A(n333), .B(n332), .ZN(n361) );
  XOR2_X1 U390 ( .A(KEYINPUT32), .B(KEYINPUT31), .Z(n335) );
  XNOR2_X1 U391 ( .A(G92GAT), .B(G204GAT), .ZN(n334) );
  XNOR2_X1 U392 ( .A(n335), .B(n334), .ZN(n336) );
  XNOR2_X1 U393 ( .A(n361), .B(n336), .ZN(n342) );
  XOR2_X1 U394 ( .A(KEYINPUT75), .B(KEYINPUT33), .Z(n338) );
  NAND2_X1 U395 ( .A1(G230GAT), .A2(G233GAT), .ZN(n337) );
  XNOR2_X1 U396 ( .A(n338), .B(n337), .ZN(n339) );
  XNOR2_X1 U397 ( .A(n339), .B(KEYINPUT74), .ZN(n340) );
  XOR2_X1 U398 ( .A(G176GAT), .B(G64GAT), .Z(n406) );
  XNOR2_X1 U399 ( .A(G99GAT), .B(G85GAT), .ZN(n343) );
  XNOR2_X1 U400 ( .A(n343), .B(G106GAT), .ZN(n372) );
  XNOR2_X1 U401 ( .A(n344), .B(n372), .ZN(n345) );
  XNOR2_X1 U402 ( .A(n346), .B(n345), .ZN(n572) );
  XNOR2_X1 U403 ( .A(n572), .B(KEYINPUT41), .ZN(n553) );
  NOR2_X1 U404 ( .A1(n568), .A2(n553), .ZN(n348) );
  INV_X1 U405 ( .A(KEYINPUT111), .ZN(n347) );
  XNOR2_X1 U406 ( .A(n348), .B(n347), .ZN(n349) );
  XNOR2_X1 U407 ( .A(n349), .B(KEYINPUT46), .ZN(n366) );
  XNOR2_X1 U408 ( .A(G8GAT), .B(G183GAT), .ZN(n350) );
  XNOR2_X1 U409 ( .A(n350), .B(G211GAT), .ZN(n393) );
  XNOR2_X1 U410 ( .A(n351), .B(n393), .ZN(n365) );
  XOR2_X1 U411 ( .A(KEYINPUT14), .B(KEYINPUT79), .Z(n353) );
  XNOR2_X1 U412 ( .A(KEYINPUT78), .B(KEYINPUT15), .ZN(n352) );
  XNOR2_X1 U413 ( .A(n353), .B(n352), .ZN(n354) );
  XOR2_X1 U414 ( .A(G22GAT), .B(G155GAT), .Z(n420) );
  XOR2_X1 U415 ( .A(n354), .B(n420), .Z(n356) );
  XNOR2_X1 U416 ( .A(G127GAT), .B(G64GAT), .ZN(n355) );
  XNOR2_X1 U417 ( .A(n356), .B(n355), .ZN(n360) );
  XOR2_X1 U418 ( .A(KEYINPUT12), .B(KEYINPUT80), .Z(n358) );
  NAND2_X1 U419 ( .A1(G231GAT), .A2(G233GAT), .ZN(n357) );
  XNOR2_X1 U420 ( .A(n358), .B(n357), .ZN(n359) );
  XOR2_X1 U421 ( .A(n360), .B(n359), .Z(n363) );
  XNOR2_X1 U422 ( .A(n361), .B(KEYINPUT77), .ZN(n362) );
  XNOR2_X1 U423 ( .A(n363), .B(n362), .ZN(n364) );
  XOR2_X1 U424 ( .A(n365), .B(n364), .Z(n547) );
  XOR2_X1 U425 ( .A(n547), .B(KEYINPUT110), .Z(n557) );
  NOR2_X1 U426 ( .A1(n366), .A2(n557), .ZN(n380) );
  XOR2_X1 U427 ( .A(KEYINPUT10), .B(KEYINPUT9), .Z(n368) );
  NAND2_X1 U428 ( .A1(G232GAT), .A2(G233GAT), .ZN(n367) );
  XNOR2_X1 U429 ( .A(n368), .B(n367), .ZN(n371) );
  XOR2_X1 U430 ( .A(G218GAT), .B(G92GAT), .Z(n370) );
  XNOR2_X1 U431 ( .A(G36GAT), .B(G190GAT), .ZN(n369) );
  XNOR2_X1 U432 ( .A(n370), .B(n369), .ZN(n400) );
  XOR2_X1 U433 ( .A(n371), .B(n400), .Z(n374) );
  XNOR2_X1 U434 ( .A(G134GAT), .B(n372), .ZN(n373) );
  XNOR2_X1 U435 ( .A(n374), .B(n373), .ZN(n375) );
  XOR2_X1 U436 ( .A(G50GAT), .B(G162GAT), .Z(n412) );
  XOR2_X1 U437 ( .A(n375), .B(n412), .Z(n377) );
  XNOR2_X1 U438 ( .A(KEYINPUT11), .B(KEYINPUT65), .ZN(n376) );
  XNOR2_X1 U439 ( .A(n377), .B(n376), .ZN(n378) );
  XNOR2_X1 U440 ( .A(n379), .B(n378), .ZN(n550) );
  AND2_X1 U441 ( .A1(n380), .A2(n550), .ZN(n381) );
  XNOR2_X1 U442 ( .A(n382), .B(n381), .ZN(n388) );
  XNOR2_X1 U443 ( .A(KEYINPUT76), .B(n550), .ZN(n562) );
  XNOR2_X1 U444 ( .A(KEYINPUT36), .B(n562), .ZN(n582) );
  NOR2_X1 U445 ( .A1(n582), .A2(n547), .ZN(n384) );
  XNOR2_X1 U446 ( .A(KEYINPUT64), .B(KEYINPUT45), .ZN(n383) );
  XNOR2_X1 U447 ( .A(n384), .B(n383), .ZN(n385) );
  NAND2_X1 U448 ( .A1(n385), .A2(n568), .ZN(n386) );
  NOR2_X1 U449 ( .A1(n572), .A2(n386), .ZN(n387) );
  NOR2_X1 U450 ( .A1(n388), .A2(n387), .ZN(n390) );
  XOR2_X1 U451 ( .A(KEYINPUT85), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U452 ( .A(G197GAT), .B(G204GAT), .ZN(n391) );
  XNOR2_X1 U453 ( .A(n392), .B(n391), .ZN(n413) );
  XNOR2_X1 U454 ( .A(n393), .B(n413), .ZN(n404) );
  XOR2_X1 U455 ( .A(KEYINPUT92), .B(KEYINPUT91), .Z(n402) );
  INV_X1 U456 ( .A(KEYINPUT18), .ZN(n394) );
  NAND2_X1 U457 ( .A1(KEYINPUT19), .A2(n394), .ZN(n397) );
  INV_X1 U458 ( .A(KEYINPUT19), .ZN(n395) );
  NAND2_X1 U459 ( .A1(n395), .A2(KEYINPUT18), .ZN(n396) );
  NAND2_X1 U460 ( .A1(n397), .A2(n396), .ZN(n399) );
  XNOR2_X1 U461 ( .A(G169GAT), .B(KEYINPUT17), .ZN(n398) );
  XNOR2_X1 U462 ( .A(n399), .B(n398), .ZN(n431) );
  XNOR2_X1 U463 ( .A(n431), .B(n400), .ZN(n401) );
  XNOR2_X1 U464 ( .A(n402), .B(n401), .ZN(n403) );
  XNOR2_X1 U465 ( .A(n404), .B(n403), .ZN(n405) );
  XOR2_X1 U466 ( .A(n406), .B(n405), .Z(n408) );
  NAND2_X1 U467 ( .A1(G226GAT), .A2(G233GAT), .ZN(n407) );
  XOR2_X1 U468 ( .A(n408), .B(n407), .Z(n514) );
  XOR2_X1 U469 ( .A(n514), .B(KEYINPUT121), .Z(n409) );
  NOR2_X1 U470 ( .A1(n522), .A2(n409), .ZN(n410) );
  XNOR2_X1 U471 ( .A(KEYINPUT54), .B(n410), .ZN(n411) );
  XOR2_X1 U472 ( .A(n413), .B(n412), .Z(n415) );
  NAND2_X1 U473 ( .A1(G228GAT), .A2(G233GAT), .ZN(n414) );
  XNOR2_X1 U474 ( .A(n415), .B(n414), .ZN(n416) );
  XOR2_X1 U475 ( .A(n416), .B(KEYINPUT24), .Z(n419) );
  XNOR2_X1 U476 ( .A(n417), .B(KEYINPUT23), .ZN(n418) );
  XNOR2_X1 U477 ( .A(n419), .B(n418), .ZN(n421) );
  XNOR2_X1 U478 ( .A(n421), .B(n420), .ZN(n423) );
  XOR2_X1 U479 ( .A(G106GAT), .B(G218GAT), .Z(n422) );
  XNOR2_X1 U480 ( .A(n423), .B(n422), .ZN(n427) );
  XOR2_X1 U481 ( .A(KEYINPUT22), .B(G211GAT), .Z(n425) );
  XNOR2_X1 U482 ( .A(G148GAT), .B(G78GAT), .ZN(n424) );
  XNOR2_X1 U483 ( .A(n425), .B(n424), .ZN(n426) );
  XNOR2_X1 U484 ( .A(n427), .B(n426), .ZN(n455) );
  NAND2_X1 U485 ( .A1(n567), .A2(n455), .ZN(n428) );
  XNOR2_X1 U486 ( .A(n428), .B(KEYINPUT55), .ZN(n443) );
  XOR2_X1 U487 ( .A(G183GAT), .B(G71GAT), .Z(n430) );
  XNOR2_X1 U488 ( .A(G15GAT), .B(G176GAT), .ZN(n429) );
  XNOR2_X1 U489 ( .A(n430), .B(n429), .ZN(n440) );
  XOR2_X1 U490 ( .A(G190GAT), .B(G99GAT), .Z(n433) );
  XNOR2_X1 U491 ( .A(G120GAT), .B(n431), .ZN(n432) );
  XNOR2_X1 U492 ( .A(n433), .B(n432), .ZN(n438) );
  XOR2_X1 U493 ( .A(KEYINPUT20), .B(KEYINPUT84), .Z(n435) );
  NAND2_X1 U494 ( .A1(G227GAT), .A2(G233GAT), .ZN(n434) );
  XNOR2_X1 U495 ( .A(n435), .B(n434), .ZN(n436) );
  XNOR2_X1 U496 ( .A(n440), .B(n439), .ZN(n442) );
  INV_X1 U497 ( .A(n516), .ZN(n523) );
  NAND2_X1 U498 ( .A1(n443), .A2(n523), .ZN(n561) );
  NOR2_X1 U499 ( .A1(n568), .A2(n561), .ZN(n446) );
  XOR2_X1 U500 ( .A(n514), .B(KEYINPUT27), .Z(n457) );
  NOR2_X1 U501 ( .A1(n523), .A2(n455), .ZN(n448) );
  XNOR2_X1 U502 ( .A(KEYINPUT95), .B(KEYINPUT26), .ZN(n447) );
  XNOR2_X1 U503 ( .A(n448), .B(n447), .ZN(n449) );
  XOR2_X1 U504 ( .A(KEYINPUT94), .B(n449), .Z(n566) );
  NAND2_X1 U505 ( .A1(n457), .A2(n566), .ZN(n453) );
  INV_X1 U506 ( .A(n514), .ZN(n467) );
  NAND2_X1 U507 ( .A1(n467), .A2(n523), .ZN(n450) );
  NAND2_X1 U508 ( .A1(n455), .A2(n450), .ZN(n451) );
  XOR2_X1 U509 ( .A(KEYINPUT25), .B(n451), .Z(n452) );
  NAND2_X1 U510 ( .A1(n453), .A2(n452), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n454), .A2(n512), .ZN(n461) );
  XNOR2_X1 U512 ( .A(KEYINPUT28), .B(KEYINPUT66), .ZN(n456) );
  XOR2_X1 U513 ( .A(n456), .B(n455), .Z(n492) );
  INV_X1 U514 ( .A(n512), .ZN(n489) );
  NAND2_X1 U515 ( .A1(n489), .A2(n457), .ZN(n521) );
  NOR2_X1 U516 ( .A1(n492), .A2(n521), .ZN(n458) );
  XOR2_X1 U517 ( .A(KEYINPUT93), .B(n458), .Z(n459) );
  NAND2_X1 U518 ( .A1(n516), .A2(n459), .ZN(n460) );
  NAND2_X1 U519 ( .A1(n461), .A2(n460), .ZN(n476) );
  NAND2_X1 U520 ( .A1(n476), .A2(n547), .ZN(n462) );
  XOR2_X1 U521 ( .A(n462), .B(KEYINPUT99), .Z(n463) );
  NOR2_X1 U522 ( .A1(n582), .A2(n463), .ZN(n464) );
  XOR2_X1 U523 ( .A(KEYINPUT37), .B(n464), .Z(n511) );
  NOR2_X1 U524 ( .A1(n568), .A2(n572), .ZN(n477) );
  NAND2_X1 U525 ( .A1(n511), .A2(n477), .ZN(n466) );
  XOR2_X1 U526 ( .A(KEYINPUT100), .B(KEYINPUT38), .Z(n465) );
  NAND2_X1 U527 ( .A1(n493), .A2(n467), .ZN(n470) );
  XOR2_X1 U528 ( .A(KEYINPUT102), .B(KEYINPUT103), .Z(n468) );
  XNOR2_X1 U529 ( .A(n468), .B(G36GAT), .ZN(n469) );
  XNOR2_X1 U530 ( .A(n470), .B(n469), .ZN(G1329GAT) );
  NAND2_X1 U531 ( .A1(n523), .A2(n493), .ZN(n472) );
  INV_X1 U532 ( .A(n547), .ZN(n576) );
  NAND2_X1 U533 ( .A1(n576), .A2(n562), .ZN(n473) );
  XOR2_X1 U534 ( .A(KEYINPUT16), .B(n473), .Z(n474) );
  XOR2_X1 U535 ( .A(KEYINPUT81), .B(n474), .Z(n475) );
  AND2_X1 U536 ( .A1(n476), .A2(n475), .ZN(n496) );
  NAND2_X1 U537 ( .A1(n477), .A2(n496), .ZN(n485) );
  NOR2_X1 U538 ( .A1(n512), .A2(n485), .ZN(n479) );
  XNOR2_X1 U539 ( .A(KEYINPUT96), .B(KEYINPUT34), .ZN(n478) );
  XNOR2_X1 U540 ( .A(n479), .B(n478), .ZN(n480) );
  XOR2_X1 U541 ( .A(G1GAT), .B(n480), .Z(G1324GAT) );
  NOR2_X1 U542 ( .A1(n514), .A2(n485), .ZN(n481) );
  XOR2_X1 U543 ( .A(G8GAT), .B(n481), .Z(G1325GAT) );
  NOR2_X1 U544 ( .A1(n516), .A2(n485), .ZN(n483) );
  XNOR2_X1 U545 ( .A(KEYINPUT97), .B(KEYINPUT35), .ZN(n482) );
  XNOR2_X1 U546 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U547 ( .A(G15GAT), .B(n484), .Z(G1326GAT) );
  INV_X1 U548 ( .A(n492), .ZN(n525) );
  NOR2_X1 U549 ( .A1(n525), .A2(n485), .ZN(n486) );
  XOR2_X1 U550 ( .A(G22GAT), .B(n486), .Z(G1327GAT) );
  XOR2_X1 U551 ( .A(KEYINPUT98), .B(KEYINPUT101), .Z(n488) );
  XNOR2_X1 U552 ( .A(G29GAT), .B(KEYINPUT39), .ZN(n487) );
  XNOR2_X1 U553 ( .A(n488), .B(n487), .ZN(n491) );
  NAND2_X1 U554 ( .A1(n493), .A2(n489), .ZN(n490) );
  XOR2_X1 U555 ( .A(n491), .B(n490), .Z(G1328GAT) );
  NAND2_X1 U556 ( .A1(n493), .A2(n492), .ZN(n494) );
  XNOR2_X1 U557 ( .A(n494), .B(G50GAT), .ZN(G1331GAT) );
  NOR2_X1 U558 ( .A1(n495), .A2(n553), .ZN(n510) );
  NAND2_X1 U559 ( .A1(n510), .A2(n496), .ZN(n497) );
  XOR2_X1 U560 ( .A(KEYINPUT105), .B(n497), .Z(n506) );
  NOR2_X1 U561 ( .A1(n512), .A2(n506), .ZN(n499) );
  XNOR2_X1 U562 ( .A(G57GAT), .B(KEYINPUT104), .ZN(n498) );
  XNOR2_X1 U563 ( .A(n499), .B(n498), .ZN(n501) );
  XOR2_X1 U564 ( .A(KEYINPUT42), .B(KEYINPUT106), .Z(n500) );
  XNOR2_X1 U565 ( .A(n501), .B(n500), .ZN(G1332GAT) );
  NOR2_X1 U566 ( .A1(n514), .A2(n506), .ZN(n503) );
  XNOR2_X1 U567 ( .A(KEYINPUT107), .B(KEYINPUT108), .ZN(n502) );
  XNOR2_X1 U568 ( .A(n503), .B(n502), .ZN(n504) );
  XNOR2_X1 U569 ( .A(G64GAT), .B(n504), .ZN(G1333GAT) );
  NOR2_X1 U570 ( .A1(n516), .A2(n506), .ZN(n505) );
  XOR2_X1 U571 ( .A(G71GAT), .B(n505), .Z(G1334GAT) );
  NOR2_X1 U572 ( .A1(n525), .A2(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(KEYINPUT109), .B(KEYINPUT43), .ZN(n507) );
  XNOR2_X1 U574 ( .A(n508), .B(n507), .ZN(n509) );
  XOR2_X1 U575 ( .A(G78GAT), .B(n509), .Z(G1335GAT) );
  NAND2_X1 U576 ( .A1(n511), .A2(n510), .ZN(n518) );
  NOR2_X1 U577 ( .A1(n512), .A2(n518), .ZN(n513) );
  XOR2_X1 U578 ( .A(G85GAT), .B(n513), .Z(G1336GAT) );
  NOR2_X1 U579 ( .A1(n514), .A2(n518), .ZN(n515) );
  XOR2_X1 U580 ( .A(G92GAT), .B(n515), .Z(G1337GAT) );
  NOR2_X1 U581 ( .A1(n516), .A2(n518), .ZN(n517) );
  XOR2_X1 U582 ( .A(G99GAT), .B(n517), .Z(G1338GAT) );
  NOR2_X1 U583 ( .A1(n525), .A2(n518), .ZN(n519) );
  XOR2_X1 U584 ( .A(KEYINPUT44), .B(n519), .Z(n520) );
  XNOR2_X1 U585 ( .A(G106GAT), .B(n520), .ZN(G1339GAT) );
  NOR2_X1 U586 ( .A1(n522), .A2(n521), .ZN(n540) );
  NAND2_X1 U587 ( .A1(n540), .A2(n523), .ZN(n524) );
  XNOR2_X1 U588 ( .A(n524), .B(KEYINPUT113), .ZN(n526) );
  NAND2_X1 U589 ( .A1(n526), .A2(n525), .ZN(n527) );
  XOR2_X1 U590 ( .A(KEYINPUT114), .B(n527), .Z(n533) );
  INV_X1 U591 ( .A(n533), .ZN(n537) );
  NOR2_X1 U592 ( .A1(n568), .A2(n537), .ZN(n528) );
  XOR2_X1 U593 ( .A(G113GAT), .B(n528), .Z(G1340GAT) );
  NOR2_X1 U594 ( .A1(n553), .A2(n537), .ZN(n532) );
  XOR2_X1 U595 ( .A(KEYINPUT116), .B(KEYINPUT49), .Z(n530) );
  XNOR2_X1 U596 ( .A(G120GAT), .B(KEYINPUT115), .ZN(n529) );
  XNOR2_X1 U597 ( .A(n530), .B(n529), .ZN(n531) );
  XNOR2_X1 U598 ( .A(n532), .B(n531), .ZN(G1341GAT) );
  XOR2_X1 U599 ( .A(KEYINPUT117), .B(KEYINPUT50), .Z(n535) );
  NAND2_X1 U600 ( .A1(n533), .A2(n557), .ZN(n534) );
  XNOR2_X1 U601 ( .A(n535), .B(n534), .ZN(n536) );
  XNOR2_X1 U602 ( .A(G127GAT), .B(n536), .ZN(G1342GAT) );
  XNOR2_X1 U603 ( .A(G134GAT), .B(KEYINPUT51), .ZN(n539) );
  NOR2_X1 U604 ( .A1(n562), .A2(n537), .ZN(n538) );
  XNOR2_X1 U605 ( .A(n539), .B(n538), .ZN(G1343GAT) );
  NAND2_X1 U606 ( .A1(n540), .A2(n566), .ZN(n549) );
  NOR2_X1 U607 ( .A1(n568), .A2(n549), .ZN(n541) );
  XOR2_X1 U608 ( .A(G141GAT), .B(n541), .Z(n542) );
  XNOR2_X1 U609 ( .A(KEYINPUT118), .B(n542), .ZN(G1344GAT) );
  NOR2_X1 U610 ( .A1(n549), .A2(n553), .ZN(n546) );
  XOR2_X1 U611 ( .A(KEYINPUT119), .B(KEYINPUT52), .Z(n544) );
  XNOR2_X1 U612 ( .A(G148GAT), .B(KEYINPUT53), .ZN(n543) );
  XNOR2_X1 U613 ( .A(n544), .B(n543), .ZN(n545) );
  XNOR2_X1 U614 ( .A(n546), .B(n545), .ZN(G1345GAT) );
  NOR2_X1 U615 ( .A1(n547), .A2(n549), .ZN(n548) );
  XOR2_X1 U616 ( .A(G155GAT), .B(n548), .Z(G1346GAT) );
  NOR2_X1 U617 ( .A1(n550), .A2(n549), .ZN(n551) );
  XOR2_X1 U618 ( .A(KEYINPUT120), .B(n551), .Z(n552) );
  XNOR2_X1 U619 ( .A(G162GAT), .B(n552), .ZN(G1347GAT) );
  NOR2_X1 U620 ( .A1(n553), .A2(n561), .ZN(n555) );
  XNOR2_X1 U621 ( .A(KEYINPUT56), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(G176GAT), .B(n556), .ZN(G1349GAT) );
  XOR2_X1 U624 ( .A(G183GAT), .B(KEYINPUT123), .Z(n560) );
  INV_X1 U625 ( .A(n561), .ZN(n558) );
  NAND2_X1 U626 ( .A1(n558), .A2(n557), .ZN(n559) );
  XNOR2_X1 U627 ( .A(n560), .B(n559), .ZN(G1350GAT) );
  INV_X1 U628 ( .A(KEYINPUT58), .ZN(n564) );
  NOR2_X1 U629 ( .A1(n562), .A2(n561), .ZN(n563) );
  XNOR2_X1 U630 ( .A(n564), .B(n563), .ZN(n565) );
  XNOR2_X1 U631 ( .A(G190GAT), .B(n565), .ZN(G1351GAT) );
  NAND2_X1 U632 ( .A1(n567), .A2(n566), .ZN(n581) );
  NOR2_X1 U633 ( .A1(n568), .A2(n581), .ZN(n570) );
  XNOR2_X1 U634 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n569) );
  XNOR2_X1 U635 ( .A(n570), .B(n569), .ZN(n571) );
  XNOR2_X1 U636 ( .A(G197GAT), .B(n571), .ZN(G1352GAT) );
  XOR2_X1 U637 ( .A(KEYINPUT124), .B(KEYINPUT61), .Z(n574) );
  INV_X1 U638 ( .A(n581), .ZN(n577) );
  NAND2_X1 U639 ( .A1(n577), .A2(n572), .ZN(n573) );
  XNOR2_X1 U640 ( .A(n574), .B(n573), .ZN(n575) );
  XNOR2_X1 U641 ( .A(G204GAT), .B(n575), .ZN(G1353GAT) );
  XOR2_X1 U642 ( .A(KEYINPUT125), .B(KEYINPUT126), .Z(n579) );
  NAND2_X1 U643 ( .A1(n577), .A2(n576), .ZN(n578) );
  XNOR2_X1 U644 ( .A(n579), .B(n578), .ZN(n580) );
  XNOR2_X1 U645 ( .A(G211GAT), .B(n580), .ZN(G1354GAT) );
  NOR2_X1 U646 ( .A1(n582), .A2(n581), .ZN(n583) );
  XOR2_X1 U647 ( .A(KEYINPUT62), .B(n583), .Z(n584) );
  XNOR2_X1 U648 ( .A(G218GAT), .B(n584), .ZN(G1355GAT) );
endmodule

