//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 1 0 1 1 0 1 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 0 1 1 1 1 1 0 1 1 1 1 0 1 1 1 1 1 0 1 0 1 1 1 0 0 0 1 1 1 0 1 0 1 1 0 0 1 1 0' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:41:46 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n201, new_n202, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n226, new_n227, new_n228, new_n229, new_n230, new_n231,
    new_n232, new_n233, new_n235, new_n236, new_n237, new_n238, new_n239,
    new_n240, new_n241, new_n242, new_n244, new_n245, new_n246, new_n247,
    new_n248, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n604, new_n605,
    new_n606, new_n607, new_n608, new_n609, new_n610, new_n611, new_n612,
    new_n613, new_n614, new_n615, new_n616, new_n617, new_n618, new_n619,
    new_n620, new_n621, new_n622, new_n623, new_n624, new_n625, new_n626,
    new_n628, new_n629, new_n630, new_n631, new_n632, new_n633, new_n634,
    new_n635, new_n636, new_n637, new_n638, new_n639, new_n640, new_n641,
    new_n642, new_n643, new_n644, new_n645, new_n646, new_n647, new_n648,
    new_n649, new_n650, new_n651, new_n652, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n703, new_n704, new_n705, new_n706,
    new_n707, new_n708, new_n709, new_n710, new_n711, new_n712, new_n713,
    new_n714, new_n715, new_n716, new_n717, new_n718, new_n719, new_n720,
    new_n721, new_n722, new_n723, new_n724, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n830, new_n831, new_n832, new_n833, new_n834,
    new_n835, new_n836, new_n837, new_n838, new_n839, new_n840, new_n841,
    new_n842, new_n843, new_n844, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n900, new_n901, new_n902, new_n903, new_n904, new_n905,
    new_n906, new_n907, new_n908, new_n909, new_n910, new_n911, new_n912,
    new_n913, new_n914, new_n915, new_n916, new_n917, new_n918, new_n919,
    new_n920, new_n921, new_n922, new_n923, new_n924, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1018, new_n1019, new_n1020, new_n1021, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1047,
    new_n1048, new_n1049, new_n1050, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1109, new_n1110, new_n1111, new_n1112, new_n1113, new_n1114,
    new_n1115, new_n1116, new_n1117, new_n1118, new_n1119, new_n1120,
    new_n1121, new_n1122, new_n1123, new_n1124, new_n1125, new_n1126,
    new_n1127, new_n1128, new_n1129, new_n1130, new_n1131, new_n1132,
    new_n1133, new_n1134, new_n1135, new_n1136, new_n1137, new_n1138,
    new_n1139, new_n1140, new_n1141, new_n1142, new_n1143, new_n1144,
    new_n1145, new_n1146, new_n1147, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1177, new_n1178, new_n1179, new_n1180, new_n1181,
    new_n1182, new_n1183, new_n1184, new_n1185, new_n1186, new_n1187,
    new_n1188, new_n1189, new_n1190, new_n1191, new_n1192, new_n1193,
    new_n1194, new_n1195, new_n1196, new_n1197, new_n1198, new_n1199,
    new_n1200, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1210, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219, new_n1220,
    new_n1221, new_n1222, new_n1223, new_n1224, new_n1225, new_n1226,
    new_n1227, new_n1228, new_n1229, new_n1230, new_n1231, new_n1232,
    new_n1233, new_n1234, new_n1235, new_n1236, new_n1237, new_n1238,
    new_n1239, new_n1240, new_n1241, new_n1242, new_n1243, new_n1244,
    new_n1245, new_n1246, new_n1247, new_n1248, new_n1249, new_n1250,
    new_n1251, new_n1252, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1269,
    new_n1270, new_n1271, new_n1272, new_n1273, new_n1274, new_n1275,
    new_n1276, new_n1277, new_n1278, new_n1279, new_n1280;
  NOR2_X1   g0000(.A1(G58), .A2(G68), .ZN(new_n201));
  INV_X1    g0001(.A(new_n201), .ZN(new_n202));
  NOR3_X1   g0002(.A1(new_n202), .A2(G50), .A3(G77), .ZN(G353));
  OAI21_X1  g0003(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  INV_X1    g0004(.A(G1), .ZN(new_n205));
  INV_X1    g0005(.A(G20), .ZN(new_n206));
  NOR2_X1   g0006(.A1(new_n205), .A2(new_n206), .ZN(new_n207));
  INV_X1    g0007(.A(new_n207), .ZN(new_n208));
  NOR2_X1   g0008(.A1(new_n208), .A2(G13), .ZN(new_n209));
  OAI211_X1 g0009(.A(new_n209), .B(G250), .C1(G257), .C2(G264), .ZN(new_n210));
  XNOR2_X1  g0010(.A(new_n210), .B(KEYINPUT0), .ZN(new_n211));
  NAND2_X1  g0011(.A1(new_n202), .A2(G50), .ZN(new_n212));
  INV_X1    g0012(.A(new_n212), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G1), .A2(G13), .ZN(new_n214));
  NOR2_X1   g0014(.A1(new_n214), .A2(new_n206), .ZN(new_n215));
  NAND2_X1  g0015(.A1(new_n213), .A2(new_n215), .ZN(new_n216));
  AOI22_X1  g0016(.A1(G50), .A2(G226), .B1(G68), .B2(G238), .ZN(new_n217));
  AOI22_X1  g0017(.A1(G77), .A2(G244), .B1(G107), .B2(G264), .ZN(new_n218));
  NAND2_X1  g0018(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  AOI22_X1  g0019(.A1(G87), .A2(G250), .B1(G116), .B2(G270), .ZN(new_n220));
  AOI22_X1  g0020(.A1(G58), .A2(G232), .B1(G97), .B2(G257), .ZN(new_n221));
  NAND2_X1  g0021(.A1(new_n220), .A2(new_n221), .ZN(new_n222));
  OAI21_X1  g0022(.A(new_n208), .B1(new_n219), .B2(new_n222), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n211), .B(new_n216), .C1(KEYINPUT1), .C2(new_n223), .ZN(new_n224));
  AOI21_X1  g0024(.A(new_n224), .B1(KEYINPUT1), .B2(new_n223), .ZN(G361));
  XOR2_X1   g0025(.A(G238), .B(G244), .Z(new_n226));
  XNOR2_X1  g0026(.A(KEYINPUT64), .B(KEYINPUT2), .ZN(new_n227));
  XNOR2_X1  g0027(.A(new_n226), .B(new_n227), .ZN(new_n228));
  XNOR2_X1  g0028(.A(G226), .B(G232), .ZN(new_n229));
  XNOR2_X1  g0029(.A(new_n228), .B(new_n229), .ZN(new_n230));
  XNOR2_X1  g0030(.A(G250), .B(G257), .ZN(new_n231));
  XNOR2_X1  g0031(.A(G264), .B(G270), .ZN(new_n232));
  XNOR2_X1  g0032(.A(new_n231), .B(new_n232), .ZN(new_n233));
  XOR2_X1   g0033(.A(new_n230), .B(new_n233), .Z(G358));
  XNOR2_X1  g0034(.A(G68), .B(G77), .ZN(new_n235));
  INV_X1    g0035(.A(G58), .ZN(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XOR2_X1   g0037(.A(KEYINPUT65), .B(G50), .Z(new_n238));
  XNOR2_X1  g0038(.A(new_n237), .B(new_n238), .ZN(new_n239));
  XOR2_X1   g0039(.A(G107), .B(G116), .Z(new_n240));
  XNOR2_X1  g0040(.A(G87), .B(G97), .ZN(new_n241));
  XNOR2_X1  g0041(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XOR2_X1   g0042(.A(new_n239), .B(new_n242), .Z(G351));
  XNOR2_X1  g0043(.A(KEYINPUT3), .B(G33), .ZN(new_n244));
  INV_X1    g0044(.A(G1698), .ZN(new_n245));
  NAND3_X1  g0045(.A1(new_n244), .A2(G222), .A3(new_n245), .ZN(new_n246));
  INV_X1    g0046(.A(G77), .ZN(new_n247));
  NAND2_X1  g0047(.A1(new_n244), .A2(G1698), .ZN(new_n248));
  INV_X1    g0048(.A(G223), .ZN(new_n249));
  OAI221_X1 g0049(.A(new_n246), .B1(new_n247), .B2(new_n244), .C1(new_n248), .C2(new_n249), .ZN(new_n250));
  INV_X1    g0050(.A(new_n214), .ZN(new_n251));
  NAND2_X1  g0051(.A1(G33), .A2(G41), .ZN(new_n252));
  AND3_X1   g0052(.A1(new_n251), .A2(KEYINPUT67), .A3(new_n252), .ZN(new_n253));
  AOI21_X1  g0053(.A(KEYINPUT67), .B1(new_n251), .B2(new_n252), .ZN(new_n254));
  NOR2_X1   g0054(.A1(new_n253), .A2(new_n254), .ZN(new_n255));
  NAND2_X1  g0055(.A1(new_n250), .A2(new_n255), .ZN(new_n256));
  INV_X1    g0056(.A(G274), .ZN(new_n257));
  AOI21_X1  g0057(.A(new_n257), .B1(new_n251), .B2(new_n252), .ZN(new_n258));
  NOR2_X1   g0058(.A1(G41), .A2(G45), .ZN(new_n259));
  NOR2_X1   g0059(.A1(new_n259), .A2(G1), .ZN(new_n260));
  NAND2_X1  g0060(.A1(new_n258), .A2(new_n260), .ZN(new_n261));
  INV_X1    g0061(.A(KEYINPUT66), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n262), .B1(new_n259), .B2(G1), .ZN(new_n263));
  NAND2_X1  g0063(.A1(new_n251), .A2(new_n252), .ZN(new_n264));
  OAI211_X1 g0064(.A(new_n205), .B(KEYINPUT66), .C1(G41), .C2(G45), .ZN(new_n265));
  AND3_X1   g0065(.A1(new_n263), .A2(new_n264), .A3(new_n265), .ZN(new_n266));
  NAND2_X1  g0066(.A1(new_n266), .A2(G226), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n256), .A2(new_n261), .A3(new_n267), .ZN(new_n268));
  INV_X1    g0068(.A(G190), .ZN(new_n269));
  NOR2_X1   g0069(.A1(new_n268), .A2(new_n269), .ZN(new_n270));
  AOI21_X1  g0070(.A(new_n270), .B1(G200), .B2(new_n268), .ZN(new_n271));
  INV_X1    g0071(.A(KEYINPUT9), .ZN(new_n272));
  INV_X1    g0072(.A(G50), .ZN(new_n273));
  AOI21_X1  g0073(.A(new_n206), .B1(new_n201), .B2(new_n273), .ZN(new_n274));
  INV_X1    g0074(.A(KEYINPUT69), .ZN(new_n275));
  XNOR2_X1  g0075(.A(new_n274), .B(new_n275), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n206), .A2(G33), .ZN(new_n277));
  INV_X1    g0077(.A(new_n277), .ZN(new_n278));
  XOR2_X1   g0078(.A(KEYINPUT8), .B(G58), .Z(new_n279));
  INV_X1    g0079(.A(G33), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n206), .A2(new_n280), .A3(KEYINPUT68), .ZN(new_n281));
  INV_X1    g0081(.A(KEYINPUT68), .ZN(new_n282));
  OAI21_X1  g0082(.A(new_n282), .B1(G20), .B2(G33), .ZN(new_n283));
  NAND2_X1  g0083(.A1(new_n281), .A2(new_n283), .ZN(new_n284));
  AOI22_X1  g0084(.A1(new_n278), .A2(new_n279), .B1(new_n284), .B2(G150), .ZN(new_n285));
  NAND2_X1  g0085(.A1(new_n276), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g0086(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n287));
  NAND2_X1  g0087(.A1(new_n287), .A2(new_n214), .ZN(new_n288));
  NAND3_X1  g0088(.A1(new_n205), .A2(G13), .A3(G20), .ZN(new_n289));
  INV_X1    g0089(.A(new_n289), .ZN(new_n290));
  AOI22_X1  g0090(.A1(new_n286), .A2(new_n288), .B1(new_n273), .B2(new_n290), .ZN(new_n291));
  INV_X1    g0091(.A(new_n288), .ZN(new_n292));
  NAND2_X1  g0092(.A1(new_n292), .A2(new_n289), .ZN(new_n293));
  XNOR2_X1  g0093(.A(new_n293), .B(KEYINPUT70), .ZN(new_n294));
  NAND2_X1  g0094(.A1(new_n205), .A2(G20), .ZN(new_n295));
  NAND3_X1  g0095(.A1(new_n294), .A2(G50), .A3(new_n295), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT73), .ZN(new_n297));
  AND3_X1   g0097(.A1(new_n291), .A2(new_n296), .A3(new_n297), .ZN(new_n298));
  AOI21_X1  g0098(.A(new_n297), .B1(new_n291), .B2(new_n296), .ZN(new_n299));
  OAI21_X1  g0099(.A(new_n272), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g0100(.A1(new_n291), .A2(new_n296), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n301), .A2(KEYINPUT73), .ZN(new_n302));
  NAND3_X1  g0102(.A1(new_n291), .A2(new_n296), .A3(new_n297), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n302), .A2(KEYINPUT9), .A3(new_n303), .ZN(new_n304));
  NAND3_X1  g0104(.A1(new_n271), .A2(new_n300), .A3(new_n304), .ZN(new_n305));
  NAND2_X1  g0105(.A1(new_n305), .A2(KEYINPUT10), .ZN(new_n306));
  INV_X1    g0106(.A(KEYINPUT10), .ZN(new_n307));
  NAND4_X1  g0107(.A1(new_n271), .A2(new_n300), .A3(new_n304), .A4(new_n307), .ZN(new_n308));
  NAND2_X1  g0108(.A1(new_n306), .A2(new_n308), .ZN(new_n309));
  NAND3_X1  g0109(.A1(new_n244), .A2(G232), .A3(new_n245), .ZN(new_n310));
  XNOR2_X1  g0110(.A(KEYINPUT72), .B(G107), .ZN(new_n311));
  INV_X1    g0111(.A(G238), .ZN(new_n312));
  OAI221_X1 g0112(.A(new_n310), .B1(new_n244), .B2(new_n311), .C1(new_n248), .C2(new_n312), .ZN(new_n313));
  NAND2_X1  g0113(.A1(new_n313), .A2(new_n255), .ZN(new_n314));
  INV_X1    g0114(.A(new_n261), .ZN(new_n315));
  AOI21_X1  g0115(.A(new_n315), .B1(new_n266), .B2(G244), .ZN(new_n316));
  NAND2_X1  g0116(.A1(new_n314), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(G169), .ZN(new_n318));
  NAND2_X1  g0118(.A1(new_n317), .A2(new_n318), .ZN(new_n319));
  NAND4_X1  g0119(.A1(new_n292), .A2(G77), .A3(new_n289), .A4(new_n295), .ZN(new_n320));
  XNOR2_X1  g0120(.A(KEYINPUT15), .B(G87), .ZN(new_n321));
  OAI22_X1  g0121(.A1(new_n321), .A2(new_n277), .B1(new_n206), .B2(new_n247), .ZN(new_n322));
  AOI21_X1  g0122(.A(new_n322), .B1(new_n284), .B2(new_n279), .ZN(new_n323));
  OAI221_X1 g0123(.A(new_n320), .B1(G77), .B2(new_n289), .C1(new_n323), .C2(new_n292), .ZN(new_n324));
  AND2_X1   g0124(.A1(new_n319), .A2(new_n324), .ZN(new_n325));
  INV_X1    g0125(.A(new_n317), .ZN(new_n326));
  INV_X1    g0126(.A(G179), .ZN(new_n327));
  NAND2_X1  g0127(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  AOI21_X1  g0128(.A(new_n324), .B1(new_n317), .B2(G200), .ZN(new_n329));
  NAND2_X1  g0129(.A1(new_n326), .A2(G190), .ZN(new_n330));
  AOI22_X1  g0130(.A1(new_n325), .A2(new_n328), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OR2_X1    g0131(.A1(new_n268), .A2(G179), .ZN(new_n332));
  NAND2_X1  g0132(.A1(new_n268), .A2(new_n318), .ZN(new_n333));
  NAND3_X1  g0133(.A1(new_n332), .A2(new_n301), .A3(new_n333), .ZN(new_n334));
  XNOR2_X1  g0134(.A(new_n334), .B(KEYINPUT71), .ZN(new_n335));
  NAND3_X1  g0135(.A1(new_n309), .A2(new_n331), .A3(new_n335), .ZN(new_n336));
  INV_X1    g0136(.A(G68), .ZN(new_n337));
  NAND2_X1  g0137(.A1(new_n290), .A2(new_n337), .ZN(new_n338));
  XNOR2_X1  g0138(.A(new_n338), .B(KEYINPUT12), .ZN(new_n339));
  NAND2_X1  g0139(.A1(new_n295), .A2(G68), .ZN(new_n340));
  INV_X1    g0140(.A(new_n284), .ZN(new_n341));
  NOR2_X1   g0141(.A1(new_n341), .A2(new_n273), .ZN(new_n342));
  OAI22_X1  g0142(.A1(new_n277), .A2(new_n247), .B1(new_n206), .B2(G68), .ZN(new_n343));
  OAI21_X1  g0143(.A(new_n288), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  INV_X1    g0144(.A(KEYINPUT11), .ZN(new_n345));
  OAI221_X1 g0145(.A(new_n339), .B1(new_n293), .B2(new_n340), .C1(new_n344), .C2(new_n345), .ZN(new_n346));
  AND2_X1   g0146(.A1(new_n344), .A2(new_n345), .ZN(new_n347));
  NOR2_X1   g0147(.A1(new_n346), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n348), .ZN(new_n349));
  INV_X1    g0149(.A(KEYINPUT14), .ZN(new_n350));
  NAND3_X1  g0150(.A1(new_n244), .A2(G226), .A3(new_n245), .ZN(new_n351));
  NAND3_X1  g0151(.A1(new_n244), .A2(G232), .A3(G1698), .ZN(new_n352));
  NAND2_X1  g0152(.A1(G33), .A2(G97), .ZN(new_n353));
  NAND3_X1  g0153(.A1(new_n351), .A2(new_n352), .A3(new_n353), .ZN(new_n354));
  INV_X1    g0154(.A(KEYINPUT74), .ZN(new_n355));
  NAND2_X1  g0155(.A1(new_n354), .A2(new_n355), .ZN(new_n356));
  NAND4_X1  g0156(.A1(new_n351), .A2(new_n352), .A3(KEYINPUT74), .A4(new_n353), .ZN(new_n357));
  NAND3_X1  g0157(.A1(new_n356), .A2(new_n357), .A3(new_n255), .ZN(new_n358));
  NAND4_X1  g0158(.A1(new_n263), .A2(new_n264), .A3(G238), .A4(new_n265), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT75), .ZN(new_n360));
  AND3_X1   g0160(.A1(new_n359), .A2(new_n360), .A3(new_n261), .ZN(new_n361));
  AOI21_X1  g0161(.A(new_n360), .B1(new_n359), .B2(new_n261), .ZN(new_n362));
  NOR2_X1   g0162(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  INV_X1    g0163(.A(KEYINPUT13), .ZN(new_n364));
  NAND3_X1  g0164(.A1(new_n358), .A2(new_n363), .A3(new_n364), .ZN(new_n365));
  INV_X1    g0165(.A(new_n365), .ZN(new_n366));
  AOI21_X1  g0166(.A(new_n364), .B1(new_n358), .B2(new_n363), .ZN(new_n367));
  OAI211_X1 g0167(.A(new_n350), .B(G169), .C1(new_n366), .C2(new_n367), .ZN(new_n368));
  NAND2_X1  g0168(.A1(new_n358), .A2(new_n363), .ZN(new_n369));
  NAND2_X1  g0169(.A1(new_n369), .A2(KEYINPUT13), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n370), .A2(G179), .A3(new_n365), .ZN(new_n371));
  NAND2_X1  g0171(.A1(new_n368), .A2(new_n371), .ZN(new_n372));
  NAND2_X1  g0172(.A1(new_n370), .A2(new_n365), .ZN(new_n373));
  AOI21_X1  g0173(.A(new_n350), .B1(new_n373), .B2(G169), .ZN(new_n374));
  OAI21_X1  g0174(.A(new_n349), .B1(new_n372), .B2(new_n374), .ZN(new_n375));
  NAND2_X1  g0175(.A1(new_n373), .A2(G200), .ZN(new_n376));
  OAI211_X1 g0176(.A(new_n376), .B(new_n348), .C1(new_n269), .C2(new_n373), .ZN(new_n377));
  NAND2_X1  g0177(.A1(new_n375), .A2(new_n377), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT7), .ZN(new_n379));
  OAI21_X1  g0179(.A(new_n379), .B1(new_n244), .B2(G20), .ZN(new_n380));
  AND2_X1   g0180(.A1(KEYINPUT3), .A2(G33), .ZN(new_n381));
  NOR2_X1   g0181(.A1(KEYINPUT3), .A2(G33), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n381), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g0183(.A1(new_n383), .A2(KEYINPUT7), .A3(new_n206), .ZN(new_n384));
  AOI21_X1  g0184(.A(new_n337), .B1(new_n380), .B2(new_n384), .ZN(new_n385));
  XNOR2_X1  g0185(.A(G58), .B(G68), .ZN(new_n386));
  AOI22_X1  g0186(.A1(new_n284), .A2(G159), .B1(new_n386), .B2(G20), .ZN(new_n387));
  INV_X1    g0187(.A(new_n387), .ZN(new_n388));
  NOR2_X1   g0188(.A1(new_n385), .A2(new_n388), .ZN(new_n389));
  AOI21_X1  g0189(.A(new_n292), .B1(new_n389), .B2(KEYINPUT16), .ZN(new_n390));
  INV_X1    g0190(.A(KEYINPUT16), .ZN(new_n391));
  OAI21_X1  g0191(.A(new_n391), .B1(new_n385), .B2(new_n388), .ZN(new_n392));
  NAND3_X1  g0192(.A1(new_n390), .A2(KEYINPUT76), .A3(new_n392), .ZN(new_n393));
  NOR3_X1   g0193(.A1(new_n244), .A2(new_n379), .A3(G20), .ZN(new_n394));
  AOI21_X1  g0194(.A(KEYINPUT7), .B1(new_n383), .B2(new_n206), .ZN(new_n395));
  OAI21_X1  g0195(.A(G68), .B1(new_n394), .B2(new_n395), .ZN(new_n396));
  NAND3_X1  g0196(.A1(new_n396), .A2(KEYINPUT16), .A3(new_n387), .ZN(new_n397));
  NAND3_X1  g0197(.A1(new_n397), .A2(new_n392), .A3(new_n288), .ZN(new_n398));
  INV_X1    g0198(.A(KEYINPUT76), .ZN(new_n399));
  NAND2_X1  g0199(.A1(new_n398), .A2(new_n399), .ZN(new_n400));
  NAND2_X1  g0200(.A1(new_n393), .A2(new_n400), .ZN(new_n401));
  AND2_X1   g0201(.A1(new_n279), .A2(new_n295), .ZN(new_n402));
  INV_X1    g0202(.A(new_n279), .ZN(new_n403));
  AOI22_X1  g0203(.A1(new_n294), .A2(new_n402), .B1(new_n290), .B2(new_n403), .ZN(new_n404));
  NAND2_X1  g0204(.A1(new_n401), .A2(new_n404), .ZN(new_n405));
  INV_X1    g0205(.A(KEYINPUT18), .ZN(new_n406));
  AOI21_X1  g0206(.A(new_n315), .B1(new_n266), .B2(G232), .ZN(new_n407));
  NAND3_X1  g0207(.A1(new_n244), .A2(G223), .A3(new_n245), .ZN(new_n408));
  NAND2_X1  g0208(.A1(G33), .A2(G87), .ZN(new_n409));
  INV_X1    g0209(.A(G226), .ZN(new_n410));
  OAI211_X1 g0210(.A(new_n408), .B(new_n409), .C1(new_n248), .C2(new_n410), .ZN(new_n411));
  NAND2_X1  g0211(.A1(new_n411), .A2(new_n255), .ZN(new_n412));
  NAND2_X1  g0212(.A1(new_n407), .A2(new_n412), .ZN(new_n413));
  NOR2_X1   g0213(.A1(new_n413), .A2(new_n327), .ZN(new_n414));
  AOI21_X1  g0214(.A(new_n414), .B1(G169), .B2(new_n413), .ZN(new_n415));
  INV_X1    g0215(.A(new_n415), .ZN(new_n416));
  NAND3_X1  g0216(.A1(new_n405), .A2(new_n406), .A3(new_n416), .ZN(new_n417));
  NOR2_X1   g0217(.A1(new_n413), .A2(new_n269), .ZN(new_n418));
  INV_X1    g0218(.A(G200), .ZN(new_n419));
  AOI21_X1  g0219(.A(new_n419), .B1(new_n412), .B2(new_n407), .ZN(new_n420));
  NOR2_X1   g0220(.A1(new_n418), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g0221(.A1(new_n401), .A2(new_n404), .A3(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(KEYINPUT17), .ZN(new_n423));
  NAND2_X1  g0223(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  INV_X1    g0224(.A(new_n404), .ZN(new_n425));
  AOI21_X1  g0225(.A(new_n425), .B1(new_n393), .B2(new_n400), .ZN(new_n426));
  OAI21_X1  g0226(.A(KEYINPUT18), .B1(new_n426), .B2(new_n415), .ZN(new_n427));
  NAND3_X1  g0227(.A1(new_n426), .A2(KEYINPUT17), .A3(new_n421), .ZN(new_n428));
  NAND4_X1  g0228(.A1(new_n417), .A2(new_n424), .A3(new_n427), .A4(new_n428), .ZN(new_n429));
  NOR3_X1   g0229(.A1(new_n336), .A2(new_n378), .A3(new_n429), .ZN(new_n430));
  OAI211_X1 g0230(.A(G264), .B(G1698), .C1(new_n381), .C2(new_n382), .ZN(new_n431));
  INV_X1    g0231(.A(KEYINPUT80), .ZN(new_n432));
  NAND2_X1  g0232(.A1(new_n431), .A2(new_n432), .ZN(new_n433));
  NAND4_X1  g0233(.A1(new_n244), .A2(KEYINPUT80), .A3(G264), .A4(G1698), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n383), .A2(G303), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n244), .A2(G257), .A3(new_n245), .ZN(new_n436));
  NAND4_X1  g0236(.A1(new_n433), .A2(new_n434), .A3(new_n435), .A4(new_n436), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n437), .A2(new_n255), .ZN(new_n438));
  INV_X1    g0238(.A(G45), .ZN(new_n439));
  NOR2_X1   g0239(.A1(new_n439), .A2(G1), .ZN(new_n440));
  INV_X1    g0240(.A(KEYINPUT77), .ZN(new_n441));
  INV_X1    g0241(.A(G41), .ZN(new_n442));
  OAI211_X1 g0242(.A(new_n440), .B(new_n441), .C1(KEYINPUT5), .C2(new_n442), .ZN(new_n443));
  OAI211_X1 g0243(.A(new_n205), .B(G45), .C1(new_n442), .C2(KEYINPUT5), .ZN(new_n444));
  NAND2_X1  g0244(.A1(new_n444), .A2(KEYINPUT77), .ZN(new_n445));
  NAND2_X1  g0245(.A1(new_n442), .A2(KEYINPUT5), .ZN(new_n446));
  NAND4_X1  g0246(.A1(new_n443), .A2(new_n445), .A3(new_n258), .A4(new_n446), .ZN(new_n447));
  INV_X1    g0247(.A(new_n446), .ZN(new_n448));
  OAI211_X1 g0248(.A(new_n264), .B(G270), .C1(new_n444), .C2(new_n448), .ZN(new_n449));
  AND2_X1   g0249(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  NAND2_X1  g0250(.A1(new_n438), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g0251(.A1(G33), .A2(G283), .ZN(new_n452));
  INV_X1    g0252(.A(G97), .ZN(new_n453));
  OAI211_X1 g0253(.A(new_n452), .B(new_n206), .C1(G33), .C2(new_n453), .ZN(new_n454));
  INV_X1    g0254(.A(G116), .ZN(new_n455));
  NAND2_X1  g0255(.A1(new_n455), .A2(G20), .ZN(new_n456));
  NAND3_X1  g0256(.A1(new_n454), .A2(new_n288), .A3(new_n456), .ZN(new_n457));
  INV_X1    g0257(.A(KEYINPUT20), .ZN(new_n458));
  NAND2_X1  g0258(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND4_X1  g0259(.A1(new_n454), .A2(KEYINPUT20), .A3(new_n288), .A4(new_n456), .ZN(new_n460));
  NAND2_X1  g0260(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  NOR2_X1   g0261(.A1(new_n289), .A2(G116), .ZN(new_n462));
  NOR2_X1   g0262(.A1(new_n280), .A2(G1), .ZN(new_n463));
  NOR3_X1   g0263(.A1(new_n290), .A2(new_n288), .A3(new_n463), .ZN(new_n464));
  AOI21_X1  g0264(.A(new_n462), .B1(new_n464), .B2(G116), .ZN(new_n465));
  AOI21_X1  g0265(.A(new_n318), .B1(new_n461), .B2(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n451), .A2(new_n466), .A3(KEYINPUT21), .ZN(new_n467));
  NAND2_X1  g0267(.A1(new_n467), .A2(KEYINPUT81), .ZN(new_n468));
  NAND3_X1  g0268(.A1(new_n438), .A2(new_n450), .A3(G179), .ZN(new_n469));
  INV_X1    g0269(.A(new_n469), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n461), .A2(new_n465), .ZN(new_n471));
  NAND2_X1  g0271(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  INV_X1    g0272(.A(KEYINPUT81), .ZN(new_n473));
  NAND4_X1  g0273(.A1(new_n451), .A2(new_n466), .A3(new_n473), .A4(KEYINPUT21), .ZN(new_n474));
  NAND3_X1  g0274(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n475));
  NAND2_X1  g0275(.A1(new_n475), .A2(KEYINPUT82), .ZN(new_n476));
  INV_X1    g0276(.A(KEYINPUT82), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n468), .A2(new_n472), .A3(new_n477), .A4(new_n474), .ZN(new_n478));
  AND2_X1   g0278(.A1(new_n451), .A2(new_n466), .ZN(new_n479));
  NOR2_X1   g0279(.A1(new_n479), .A2(KEYINPUT21), .ZN(new_n480));
  INV_X1    g0280(.A(new_n480), .ZN(new_n481));
  AOI21_X1  g0281(.A(new_n471), .B1(new_n451), .B2(G200), .ZN(new_n482));
  OAI21_X1  g0282(.A(new_n482), .B1(new_n269), .B2(new_n451), .ZN(new_n483));
  NAND4_X1  g0283(.A1(new_n476), .A2(new_n478), .A3(new_n481), .A4(new_n483), .ZN(new_n484));
  INV_X1    g0284(.A(new_n484), .ZN(new_n485));
  OAI211_X1 g0285(.A(G257), .B(G1698), .C1(new_n381), .C2(new_n382), .ZN(new_n486));
  OAI211_X1 g0286(.A(G250), .B(new_n245), .C1(new_n381), .C2(new_n382), .ZN(new_n487));
  AND2_X1   g0287(.A1(KEYINPUT85), .A2(G294), .ZN(new_n488));
  NOR2_X1   g0288(.A1(KEYINPUT85), .A2(G294), .ZN(new_n489));
  OAI21_X1  g0289(.A(G33), .B1(new_n488), .B2(new_n489), .ZN(new_n490));
  NAND3_X1  g0290(.A1(new_n486), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND2_X1  g0291(.A1(new_n255), .A2(new_n491), .ZN(new_n492));
  OAI211_X1 g0292(.A(new_n264), .B(G264), .C1(new_n444), .C2(new_n448), .ZN(new_n493));
  NAND3_X1  g0293(.A1(new_n492), .A2(new_n447), .A3(new_n493), .ZN(new_n494));
  NAND2_X1  g0294(.A1(new_n494), .A2(new_n318), .ZN(new_n495));
  OAI21_X1  g0295(.A(new_n495), .B1(G179), .B2(new_n494), .ZN(new_n496));
  OAI211_X1 g0296(.A(new_n206), .B(G87), .C1(new_n381), .C2(new_n382), .ZN(new_n497));
  NAND2_X1  g0297(.A1(new_n497), .A2(KEYINPUT22), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT83), .ZN(new_n499));
  NOR2_X1   g0299(.A1(KEYINPUT22), .A2(G20), .ZN(new_n500));
  NAND2_X1  g0300(.A1(new_n500), .A2(G87), .ZN(new_n501));
  OAI21_X1  g0301(.A(new_n499), .B1(new_n383), .B2(new_n501), .ZN(new_n502));
  NAND4_X1  g0302(.A1(new_n244), .A2(KEYINPUT83), .A3(G87), .A4(new_n500), .ZN(new_n503));
  NAND3_X1  g0303(.A1(new_n498), .A2(new_n502), .A3(new_n503), .ZN(new_n504));
  INV_X1    g0304(.A(KEYINPUT23), .ZN(new_n505));
  INV_X1    g0305(.A(G107), .ZN(new_n506));
  NAND3_X1  g0306(.A1(new_n505), .A2(new_n506), .A3(G20), .ZN(new_n507));
  OAI21_X1  g0307(.A(new_n507), .B1(new_n455), .B2(new_n277), .ZN(new_n508));
  NAND2_X1  g0308(.A1(new_n311), .A2(G20), .ZN(new_n509));
  AOI21_X1  g0309(.A(new_n508), .B1(new_n509), .B2(KEYINPUT23), .ZN(new_n510));
  NAND2_X1  g0310(.A1(new_n504), .A2(new_n510), .ZN(new_n511));
  INV_X1    g0311(.A(KEYINPUT84), .ZN(new_n512));
  INV_X1    g0312(.A(KEYINPUT24), .ZN(new_n513));
  NAND3_X1  g0313(.A1(new_n511), .A2(new_n512), .A3(new_n513), .ZN(new_n514));
  NAND3_X1  g0314(.A1(new_n504), .A2(KEYINPUT84), .A3(new_n510), .ZN(new_n515));
  NAND2_X1  g0315(.A1(new_n515), .A2(KEYINPUT24), .ZN(new_n516));
  AOI21_X1  g0316(.A(KEYINPUT84), .B1(new_n504), .B2(new_n510), .ZN(new_n517));
  OAI211_X1 g0317(.A(new_n288), .B(new_n514), .C1(new_n516), .C2(new_n517), .ZN(new_n518));
  INV_X1    g0318(.A(KEYINPUT25), .ZN(new_n519));
  NOR3_X1   g0319(.A1(new_n289), .A2(new_n519), .A3(G107), .ZN(new_n520));
  INV_X1    g0320(.A(new_n520), .ZN(new_n521));
  OAI21_X1  g0321(.A(new_n519), .B1(new_n289), .B2(G107), .ZN(new_n522));
  AOI22_X1  g0322(.A1(new_n464), .A2(G107), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI21_X1  g0323(.A(new_n496), .B1(new_n518), .B2(new_n523), .ZN(new_n524));
  NAND2_X1  g0324(.A1(new_n494), .A2(new_n419), .ZN(new_n525));
  NAND4_X1  g0325(.A1(new_n492), .A2(new_n269), .A3(new_n447), .A4(new_n493), .ZN(new_n526));
  NAND2_X1  g0326(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  NOR2_X1   g0327(.A1(new_n516), .A2(new_n517), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n514), .A2(new_n288), .ZN(new_n529));
  OAI211_X1 g0329(.A(new_n523), .B(new_n527), .C1(new_n528), .C2(new_n529), .ZN(new_n530));
  NAND2_X1  g0330(.A1(new_n530), .A2(KEYINPUT86), .ZN(new_n531));
  INV_X1    g0331(.A(KEYINPUT86), .ZN(new_n532));
  NAND4_X1  g0332(.A1(new_n518), .A2(new_n532), .A3(new_n523), .A4(new_n527), .ZN(new_n533));
  AOI21_X1  g0333(.A(new_n524), .B1(new_n531), .B2(new_n533), .ZN(new_n534));
  INV_X1    g0334(.A(KEYINPUT87), .ZN(new_n535));
  XNOR2_X1  g0335(.A(new_n534), .B(new_n535), .ZN(new_n536));
  NAND4_X1  g0336(.A1(new_n244), .A2(KEYINPUT4), .A3(G244), .A4(new_n245), .ZN(new_n537));
  AND2_X1   g0337(.A1(new_n244), .A2(G244), .ZN(new_n538));
  OAI211_X1 g0338(.A(new_n452), .B(new_n537), .C1(new_n538), .C2(KEYINPUT4), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n244), .A2(G250), .ZN(new_n540));
  AOI21_X1  g0340(.A(new_n245), .B1(new_n540), .B2(KEYINPUT4), .ZN(new_n541));
  OAI21_X1  g0341(.A(new_n255), .B1(new_n539), .B2(new_n541), .ZN(new_n542));
  OAI211_X1 g0342(.A(new_n264), .B(G257), .C1(new_n444), .C2(new_n448), .ZN(new_n543));
  AND2_X1   g0343(.A1(new_n447), .A2(new_n543), .ZN(new_n544));
  NAND2_X1  g0344(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  NAND2_X1  g0345(.A1(new_n545), .A2(new_n318), .ZN(new_n546));
  NAND3_X1  g0346(.A1(new_n506), .A2(KEYINPUT6), .A3(G97), .ZN(new_n547));
  NOR2_X1   g0347(.A1(new_n453), .A2(new_n506), .ZN(new_n548));
  NOR2_X1   g0348(.A1(G97), .A2(G107), .ZN(new_n549));
  NOR2_X1   g0349(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  OAI21_X1  g0350(.A(new_n547), .B1(new_n550), .B2(KEYINPUT6), .ZN(new_n551));
  AOI22_X1  g0351(.A1(new_n551), .A2(G20), .B1(G77), .B2(new_n284), .ZN(new_n552));
  INV_X1    g0352(.A(new_n311), .ZN(new_n553));
  OAI21_X1  g0353(.A(new_n553), .B1(new_n394), .B2(new_n395), .ZN(new_n554));
  NAND2_X1  g0354(.A1(new_n552), .A2(new_n554), .ZN(new_n555));
  NAND2_X1  g0355(.A1(new_n555), .A2(new_n288), .ZN(new_n556));
  NOR2_X1   g0356(.A1(new_n289), .A2(G97), .ZN(new_n557));
  AOI21_X1  g0357(.A(new_n557), .B1(new_n464), .B2(G97), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND3_X1  g0359(.A1(new_n542), .A2(new_n327), .A3(new_n544), .ZN(new_n560));
  NAND3_X1  g0360(.A1(new_n546), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  INV_X1    g0361(.A(new_n558), .ZN(new_n562));
  AOI21_X1  g0362(.A(new_n562), .B1(new_n555), .B2(new_n288), .ZN(new_n563));
  NAND3_X1  g0363(.A1(new_n542), .A2(G190), .A3(new_n544), .ZN(new_n564));
  AND2_X1   g0364(.A1(new_n542), .A2(new_n544), .ZN(new_n565));
  OAI211_X1 g0365(.A(new_n563), .B(new_n564), .C1(new_n565), .C2(new_n419), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n244), .A2(G238), .A3(new_n245), .ZN(new_n567));
  NAND3_X1  g0367(.A1(new_n244), .A2(G244), .A3(G1698), .ZN(new_n568));
  OAI211_X1 g0368(.A(new_n567), .B(new_n568), .C1(new_n280), .C2(new_n455), .ZN(new_n569));
  NAND2_X1  g0369(.A1(new_n569), .A2(new_n255), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n440), .A2(new_n257), .ZN(new_n571));
  INV_X1    g0371(.A(G250), .ZN(new_n572));
  OAI21_X1  g0372(.A(new_n572), .B1(new_n439), .B2(G1), .ZN(new_n573));
  NAND3_X1  g0373(.A1(new_n571), .A2(new_n264), .A3(new_n573), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n570), .A2(new_n574), .ZN(new_n575));
  NAND2_X1  g0375(.A1(new_n575), .A2(new_n318), .ZN(new_n576));
  XNOR2_X1  g0376(.A(KEYINPUT78), .B(G87), .ZN(new_n577));
  NAND3_X1  g0377(.A1(new_n311), .A2(new_n577), .A3(new_n453), .ZN(new_n578));
  INV_X1    g0378(.A(KEYINPUT19), .ZN(new_n579));
  OAI21_X1  g0379(.A(new_n206), .B1(new_n353), .B2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  INV_X1    g0381(.A(new_n581), .ZN(new_n582));
  OAI21_X1  g0382(.A(new_n579), .B1(new_n277), .B2(new_n453), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n244), .A2(new_n206), .ZN(new_n584));
  OAI21_X1  g0384(.A(new_n583), .B1(new_n584), .B2(new_n337), .ZN(new_n585));
  OAI21_X1  g0385(.A(new_n288), .B1(new_n582), .B2(new_n585), .ZN(new_n586));
  NAND2_X1  g0386(.A1(new_n321), .A2(new_n290), .ZN(new_n587));
  INV_X1    g0387(.A(new_n321), .ZN(new_n588));
  NAND2_X1  g0388(.A1(new_n464), .A2(new_n588), .ZN(new_n589));
  NAND3_X1  g0389(.A1(new_n586), .A2(new_n587), .A3(new_n589), .ZN(new_n590));
  INV_X1    g0390(.A(new_n574), .ZN(new_n591));
  AOI21_X1  g0391(.A(new_n591), .B1(new_n569), .B2(new_n255), .ZN(new_n592));
  NAND2_X1  g0392(.A1(new_n592), .A2(new_n327), .ZN(new_n593));
  NAND3_X1  g0393(.A1(new_n576), .A2(new_n590), .A3(new_n593), .ZN(new_n594));
  NAND2_X1  g0394(.A1(new_n575), .A2(G200), .ZN(new_n595));
  OAI211_X1 g0395(.A(new_n581), .B(new_n583), .C1(new_n337), .C2(new_n584), .ZN(new_n596));
  AOI22_X1  g0396(.A1(new_n596), .A2(new_n288), .B1(new_n290), .B2(new_n321), .ZN(new_n597));
  NAND2_X1  g0397(.A1(new_n592), .A2(G190), .ZN(new_n598));
  NAND2_X1  g0398(.A1(new_n464), .A2(G87), .ZN(new_n599));
  NAND4_X1  g0399(.A1(new_n595), .A2(new_n597), .A3(new_n598), .A4(new_n599), .ZN(new_n600));
  AND4_X1   g0400(.A1(new_n561), .A2(new_n566), .A3(new_n594), .A4(new_n600), .ZN(new_n601));
  XNOR2_X1  g0401(.A(new_n601), .B(KEYINPUT79), .ZN(new_n602));
  AND4_X1   g0402(.A1(new_n430), .A2(new_n485), .A3(new_n536), .A4(new_n602), .ZN(G372));
  NAND2_X1  g0403(.A1(new_n424), .A2(new_n428), .ZN(new_n604));
  AND2_X1   g0404(.A1(new_n325), .A2(new_n328), .ZN(new_n605));
  NAND2_X1  g0405(.A1(new_n377), .A2(new_n605), .ZN(new_n606));
  AOI21_X1  g0406(.A(new_n604), .B1(new_n606), .B2(new_n375), .ZN(new_n607));
  NAND2_X1  g0407(.A1(new_n417), .A2(new_n427), .ZN(new_n608));
  OAI21_X1  g0408(.A(new_n309), .B1(new_n607), .B2(new_n608), .ZN(new_n609));
  AND2_X1   g0409(.A1(new_n609), .A2(new_n335), .ZN(new_n610));
  AND3_X1   g0410(.A1(new_n468), .A2(new_n472), .A3(new_n474), .ZN(new_n611));
  NAND2_X1  g0411(.A1(new_n518), .A2(new_n523), .ZN(new_n612));
  INV_X1    g0412(.A(new_n496), .ZN(new_n613));
  NAND2_X1  g0413(.A1(new_n612), .A2(new_n613), .ZN(new_n614));
  NAND3_X1  g0414(.A1(new_n611), .A2(new_n481), .A3(new_n614), .ZN(new_n615));
  NAND2_X1  g0415(.A1(new_n531), .A2(new_n533), .ZN(new_n616));
  NAND3_X1  g0416(.A1(new_n615), .A2(new_n601), .A3(new_n616), .ZN(new_n617));
  INV_X1    g0417(.A(new_n594), .ZN(new_n618));
  AND3_X1   g0418(.A1(new_n546), .A2(new_n559), .A3(new_n560), .ZN(new_n619));
  NAND4_X1  g0419(.A1(new_n619), .A2(KEYINPUT26), .A3(new_n594), .A4(new_n600), .ZN(new_n620));
  INV_X1    g0420(.A(KEYINPUT26), .ZN(new_n621));
  NAND2_X1  g0421(.A1(new_n600), .A2(new_n594), .ZN(new_n622));
  OAI21_X1  g0422(.A(new_n621), .B1(new_n622), .B2(new_n561), .ZN(new_n623));
  AOI21_X1  g0423(.A(new_n618), .B1(new_n620), .B2(new_n623), .ZN(new_n624));
  NAND2_X1  g0424(.A1(new_n617), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g0425(.A1(new_n430), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n610), .A2(new_n626), .ZN(G369));
  INV_X1    g0427(.A(KEYINPUT88), .ZN(new_n628));
  NAND2_X1  g0428(.A1(new_n484), .A2(new_n628), .ZN(new_n629));
  AOI21_X1  g0429(.A(new_n480), .B1(new_n475), .B2(KEYINPUT82), .ZN(new_n630));
  NAND4_X1  g0430(.A1(new_n630), .A2(KEYINPUT88), .A3(new_n478), .A4(new_n483), .ZN(new_n631));
  NAND3_X1  g0431(.A1(new_n205), .A2(new_n206), .A3(G13), .ZN(new_n632));
  OR2_X1    g0432(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n633));
  NAND2_X1  g0433(.A1(new_n632), .A2(KEYINPUT27), .ZN(new_n634));
  NAND3_X1  g0434(.A1(new_n633), .A2(G213), .A3(new_n634), .ZN(new_n635));
  INV_X1    g0435(.A(G343), .ZN(new_n636));
  NOR2_X1   g0436(.A1(new_n635), .A2(new_n636), .ZN(new_n637));
  AOI22_X1  g0437(.A1(new_n629), .A2(new_n631), .B1(new_n471), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n471), .A2(new_n637), .ZN(new_n639));
  AOI21_X1  g0439(.A(new_n639), .B1(new_n611), .B2(new_n481), .ZN(new_n640));
  OAI21_X1  g0440(.A(G330), .B1(new_n638), .B2(new_n640), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n612), .A2(new_n637), .ZN(new_n642));
  AOI21_X1  g0442(.A(new_n535), .B1(new_n616), .B2(new_n614), .ZN(new_n643));
  AOI211_X1 g0443(.A(KEYINPUT87), .B(new_n524), .C1(new_n531), .C2(new_n533), .ZN(new_n644));
  OAI21_X1  g0444(.A(new_n642), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  NAND2_X1  g0445(.A1(new_n524), .A2(new_n637), .ZN(new_n646));
  AND2_X1   g0446(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NOR2_X1   g0447(.A1(new_n641), .A2(new_n647), .ZN(new_n648));
  INV_X1    g0448(.A(new_n648), .ZN(new_n649));
  NOR2_X1   g0449(.A1(new_n614), .A2(new_n637), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n637), .B1(new_n630), .B2(new_n478), .ZN(new_n651));
  AOI21_X1  g0451(.A(new_n650), .B1(new_n536), .B2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n649), .A2(new_n652), .ZN(G399));
  INV_X1    g0453(.A(new_n209), .ZN(new_n654));
  NOR2_X1   g0454(.A1(new_n654), .A2(G41), .ZN(new_n655));
  INV_X1    g0455(.A(new_n655), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(G1), .ZN(new_n657));
  OR2_X1    g0457(.A1(new_n578), .A2(G116), .ZN(new_n658));
  OAI22_X1  g0458(.A1(new_n657), .A2(new_n658), .B1(new_n212), .B2(new_n656), .ZN(new_n659));
  XOR2_X1   g0459(.A(KEYINPUT89), .B(KEYINPUT28), .Z(new_n660));
  XNOR2_X1  g0460(.A(new_n659), .B(new_n660), .ZN(new_n661));
  INV_X1    g0461(.A(G330), .ZN(new_n662));
  INV_X1    g0462(.A(new_n637), .ZN(new_n663));
  NAND4_X1  g0463(.A1(new_n536), .A2(new_n485), .A3(new_n602), .A4(new_n663), .ZN(new_n664));
  INV_X1    g0464(.A(KEYINPUT91), .ZN(new_n665));
  NOR2_X1   g0465(.A1(new_n592), .A2(G179), .ZN(new_n666));
  NAND4_X1  g0466(.A1(new_n545), .A2(new_n666), .A3(new_n451), .A4(new_n494), .ZN(new_n667));
  INV_X1    g0467(.A(KEYINPUT90), .ZN(new_n668));
  NAND2_X1  g0468(.A1(new_n667), .A2(new_n668), .ZN(new_n669));
  AND3_X1   g0469(.A1(new_n575), .A2(new_n327), .A3(new_n494), .ZN(new_n670));
  NAND4_X1  g0470(.A1(new_n670), .A2(KEYINPUT90), .A3(new_n451), .A4(new_n545), .ZN(new_n671));
  AND2_X1   g0471(.A1(new_n492), .A2(new_n493), .ZN(new_n672));
  AND2_X1   g0472(.A1(new_n672), .A2(new_n592), .ZN(new_n673));
  NAND4_X1  g0473(.A1(new_n565), .A2(new_n673), .A3(new_n470), .A4(KEYINPUT30), .ZN(new_n674));
  INV_X1    g0474(.A(KEYINPUT30), .ZN(new_n675));
  NAND4_X1  g0475(.A1(new_n542), .A2(new_n672), .A3(new_n544), .A4(new_n592), .ZN(new_n676));
  OAI21_X1  g0476(.A(new_n675), .B1(new_n676), .B2(new_n469), .ZN(new_n677));
  NAND4_X1  g0477(.A1(new_n669), .A2(new_n671), .A3(new_n674), .A4(new_n677), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n678), .A2(new_n637), .ZN(new_n679));
  INV_X1    g0479(.A(KEYINPUT31), .ZN(new_n680));
  NAND2_X1  g0480(.A1(new_n679), .A2(new_n680), .ZN(new_n681));
  NAND3_X1  g0481(.A1(new_n674), .A2(new_n677), .A3(new_n667), .ZN(new_n682));
  NAND3_X1  g0482(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n665), .B1(new_n681), .B2(new_n683), .ZN(new_n684));
  AOI21_X1  g0484(.A(KEYINPUT31), .B1(new_n678), .B2(new_n637), .ZN(new_n685));
  AND3_X1   g0485(.A1(new_n682), .A2(KEYINPUT31), .A3(new_n637), .ZN(new_n686));
  NOR3_X1   g0486(.A1(new_n685), .A2(new_n686), .A3(KEYINPUT91), .ZN(new_n687));
  NOR2_X1   g0487(.A1(new_n684), .A2(new_n687), .ZN(new_n688));
  AOI21_X1  g0488(.A(new_n662), .B1(new_n664), .B2(new_n688), .ZN(new_n689));
  NAND2_X1  g0489(.A1(new_n625), .A2(new_n663), .ZN(new_n690));
  INV_X1    g0490(.A(KEYINPUT29), .ZN(new_n691));
  NAND3_X1  g0491(.A1(new_n690), .A2(KEYINPUT92), .A3(new_n691), .ZN(new_n692));
  INV_X1    g0492(.A(KEYINPUT92), .ZN(new_n693));
  AOI21_X1  g0493(.A(new_n637), .B1(new_n617), .B2(new_n624), .ZN(new_n694));
  OAI21_X1  g0494(.A(new_n693), .B1(new_n694), .B2(KEYINPUT29), .ZN(new_n695));
  AND2_X1   g0495(.A1(new_n692), .A2(new_n695), .ZN(new_n696));
  NAND3_X1  g0496(.A1(new_n630), .A2(new_n478), .A3(new_n614), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n697), .A2(new_n616), .A3(new_n601), .ZN(new_n698));
  AOI21_X1  g0498(.A(new_n637), .B1(new_n698), .B2(new_n624), .ZN(new_n699));
  NAND2_X1  g0499(.A1(new_n699), .A2(KEYINPUT29), .ZN(new_n700));
  AOI21_X1  g0500(.A(new_n689), .B1(new_n696), .B2(new_n700), .ZN(new_n701));
  OAI21_X1  g0501(.A(new_n661), .B1(new_n701), .B2(G1), .ZN(G364));
  AND2_X1   g0502(.A1(new_n206), .A2(G13), .ZN(new_n703));
  NAND2_X1  g0503(.A1(new_n703), .A2(G45), .ZN(new_n704));
  NAND2_X1  g0504(.A1(new_n704), .A2(G1), .ZN(new_n705));
  OR3_X1    g0505(.A1(new_n655), .A2(KEYINPUT93), .A3(new_n705), .ZN(new_n706));
  OAI21_X1  g0506(.A(KEYINPUT93), .B1(new_n655), .B2(new_n705), .ZN(new_n707));
  NAND2_X1  g0507(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g0508(.A(new_n708), .ZN(new_n709));
  NOR2_X1   g0509(.A1(new_n654), .A2(new_n383), .ZN(new_n710));
  INV_X1    g0510(.A(KEYINPUT94), .ZN(new_n711));
  NAND2_X1  g0511(.A1(G355), .A2(new_n711), .ZN(new_n712));
  OR2_X1    g0512(.A1(G355), .A2(new_n711), .ZN(new_n713));
  NAND3_X1  g0513(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  OAI21_X1  g0514(.A(new_n714), .B1(G116), .B2(new_n209), .ZN(new_n715));
  NAND2_X1  g0515(.A1(new_n239), .A2(G45), .ZN(new_n716));
  NOR2_X1   g0516(.A1(new_n654), .A2(new_n244), .ZN(new_n717));
  INV_X1    g0517(.A(new_n717), .ZN(new_n718));
  AOI21_X1  g0518(.A(new_n718), .B1(new_n439), .B2(new_n213), .ZN(new_n719));
  AOI21_X1  g0519(.A(new_n715), .B1(new_n716), .B2(new_n719), .ZN(new_n720));
  NOR2_X1   g0520(.A1(G13), .A2(G33), .ZN(new_n721));
  INV_X1    g0521(.A(new_n721), .ZN(new_n722));
  NOR2_X1   g0522(.A1(new_n722), .A2(G20), .ZN(new_n723));
  AOI21_X1  g0523(.A(new_n214), .B1(G20), .B2(new_n318), .ZN(new_n724));
  NOR2_X1   g0524(.A1(new_n723), .A2(new_n724), .ZN(new_n725));
  INV_X1    g0525(.A(new_n725), .ZN(new_n726));
  OAI21_X1  g0526(.A(new_n709), .B1(new_n720), .B2(new_n726), .ZN(new_n727));
  NOR2_X1   g0527(.A1(new_n419), .A2(G179), .ZN(new_n728));
  XNOR2_X1  g0528(.A(new_n728), .B(KEYINPUT97), .ZN(new_n729));
  NOR2_X1   g0529(.A1(new_n206), .A2(new_n269), .ZN(new_n730));
  NAND2_X1  g0530(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  XOR2_X1   g0531(.A(new_n731), .B(KEYINPUT99), .Z(new_n732));
  NAND2_X1  g0532(.A1(new_n732), .A2(G303), .ZN(new_n733));
  OR3_X1    g0533(.A1(new_n206), .A2(KEYINPUT96), .A3(G190), .ZN(new_n734));
  NOR2_X1   g0534(.A1(G179), .A2(G200), .ZN(new_n735));
  OAI21_X1  g0535(.A(KEYINPUT96), .B1(new_n206), .B2(G190), .ZN(new_n736));
  NAND3_X1  g0536(.A1(new_n734), .A2(new_n735), .A3(new_n736), .ZN(new_n737));
  INV_X1    g0537(.A(new_n737), .ZN(new_n738));
  OR2_X1    g0538(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n739));
  NAND2_X1  g0539(.A1(new_n738), .A2(KEYINPUT100), .ZN(new_n740));
  NAND2_X1  g0540(.A1(new_n739), .A2(new_n740), .ZN(new_n741));
  INV_X1    g0541(.A(new_n741), .ZN(new_n742));
  NAND2_X1  g0542(.A1(new_n742), .A2(G329), .ZN(new_n743));
  NAND3_X1  g0543(.A1(new_n729), .A2(new_n736), .A3(new_n734), .ZN(new_n744));
  INV_X1    g0544(.A(new_n744), .ZN(new_n745));
  NAND2_X1  g0545(.A1(new_n745), .A2(G283), .ZN(new_n746));
  INV_X1    g0546(.A(G311), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n206), .A2(new_n327), .ZN(new_n748));
  NAND3_X1  g0548(.A1(new_n748), .A2(new_n269), .A3(new_n419), .ZN(new_n749));
  NAND2_X1  g0549(.A1(new_n748), .A2(G200), .ZN(new_n750));
  NOR2_X1   g0550(.A1(new_n750), .A2(new_n269), .ZN(new_n751));
  INV_X1    g0551(.A(new_n751), .ZN(new_n752));
  INV_X1    g0552(.A(G326), .ZN(new_n753));
  OAI221_X1 g0553(.A(new_n383), .B1(new_n747), .B2(new_n749), .C1(new_n752), .C2(new_n753), .ZN(new_n754));
  NOR2_X1   g0554(.A1(new_n488), .A2(new_n489), .ZN(new_n755));
  INV_X1    g0555(.A(new_n755), .ZN(new_n756));
  AOI21_X1  g0556(.A(new_n206), .B1(new_n735), .B2(G190), .ZN(new_n757));
  INV_X1    g0557(.A(new_n757), .ZN(new_n758));
  AOI21_X1  g0558(.A(new_n754), .B1(new_n756), .B2(new_n758), .ZN(new_n759));
  NAND4_X1  g0559(.A1(new_n733), .A2(new_n743), .A3(new_n746), .A4(new_n759), .ZN(new_n760));
  NAND3_X1  g0560(.A1(new_n730), .A2(G179), .A3(new_n419), .ZN(new_n761));
  NAND2_X1  g0561(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n762));
  INV_X1    g0562(.A(new_n762), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n761), .A2(KEYINPUT95), .ZN(new_n764));
  NOR2_X1   g0564(.A1(new_n763), .A2(new_n764), .ZN(new_n765));
  INV_X1    g0565(.A(G322), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n750), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  XOR2_X1   g0568(.A(KEYINPUT33), .B(G317), .Z(new_n769));
  OAI22_X1  g0569(.A1(new_n765), .A2(new_n766), .B1(new_n768), .B2(new_n769), .ZN(new_n770));
  XNOR2_X1  g0570(.A(new_n770), .B(KEYINPUT101), .ZN(new_n771));
  NAND2_X1  g0571(.A1(new_n738), .A2(G159), .ZN(new_n772));
  XOR2_X1   g0572(.A(new_n772), .B(KEYINPUT32), .Z(new_n773));
  INV_X1    g0573(.A(new_n749), .ZN(new_n774));
  AOI22_X1  g0574(.A1(new_n774), .A2(G77), .B1(new_n758), .B2(G97), .ZN(new_n775));
  INV_X1    g0575(.A(new_n765), .ZN(new_n776));
  AOI22_X1  g0576(.A1(new_n776), .A2(G58), .B1(G107), .B2(new_n745), .ZN(new_n777));
  AOI22_X1  g0577(.A1(new_n767), .A2(G68), .B1(new_n751), .B2(G50), .ZN(new_n778));
  NAND4_X1  g0578(.A1(new_n773), .A2(new_n775), .A3(new_n777), .A4(new_n778), .ZN(new_n779));
  OAI21_X1  g0579(.A(new_n244), .B1(new_n731), .B2(new_n577), .ZN(new_n780));
  XNOR2_X1  g0580(.A(new_n780), .B(KEYINPUT98), .ZN(new_n781));
  OAI22_X1  g0581(.A1(new_n760), .A2(new_n771), .B1(new_n779), .B2(new_n781), .ZN(new_n782));
  AOI21_X1  g0582(.A(new_n727), .B1(new_n782), .B2(new_n724), .ZN(new_n783));
  OR2_X1    g0583(.A1(new_n638), .A2(new_n640), .ZN(new_n784));
  INV_X1    g0584(.A(new_n723), .ZN(new_n785));
  OAI21_X1  g0585(.A(new_n783), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  NOR2_X1   g0586(.A1(new_n784), .A2(G330), .ZN(new_n787));
  NAND2_X1  g0587(.A1(new_n641), .A2(new_n708), .ZN(new_n788));
  OAI21_X1  g0588(.A(new_n786), .B1(new_n787), .B2(new_n788), .ZN(new_n789));
  XNOR2_X1  g0589(.A(new_n789), .B(KEYINPUT102), .ZN(G396));
  OAI21_X1  g0590(.A(new_n383), .B1(new_n749), .B2(new_n455), .ZN(new_n791));
  XOR2_X1   g0591(.A(KEYINPUT103), .B(G283), .Z(new_n792));
  INV_X1    g0592(.A(G303), .ZN(new_n793));
  OAI22_X1  g0593(.A1(new_n768), .A2(new_n792), .B1(new_n752), .B2(new_n793), .ZN(new_n794));
  AOI211_X1 g0594(.A(new_n791), .B(new_n794), .C1(G97), .C2(new_n758), .ZN(new_n795));
  AOI22_X1  g0595(.A1(new_n776), .A2(G294), .B1(G87), .B2(new_n745), .ZN(new_n796));
  AND2_X1   g0596(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  INV_X1    g0597(.A(new_n732), .ZN(new_n798));
  OAI221_X1 g0598(.A(new_n797), .B1(new_n506), .B2(new_n798), .C1(new_n747), .C2(new_n741), .ZN(new_n799));
  NAND2_X1  g0599(.A1(new_n742), .A2(G132), .ZN(new_n800));
  OAI21_X1  g0600(.A(new_n244), .B1(new_n757), .B2(new_n236), .ZN(new_n801));
  AOI21_X1  g0601(.A(new_n801), .B1(new_n745), .B2(G68), .ZN(new_n802));
  OAI211_X1 g0602(.A(new_n800), .B(new_n802), .C1(new_n798), .C2(new_n273), .ZN(new_n803));
  AOI22_X1  g0603(.A1(G137), .A2(new_n751), .B1(new_n774), .B2(G159), .ZN(new_n804));
  INV_X1    g0604(.A(G150), .ZN(new_n805));
  OAI21_X1  g0605(.A(new_n804), .B1(new_n805), .B2(new_n768), .ZN(new_n806));
  AOI21_X1  g0606(.A(new_n806), .B1(G143), .B2(new_n776), .ZN(new_n807));
  XNOR2_X1  g0607(.A(new_n807), .B(KEYINPUT34), .ZN(new_n808));
  OAI21_X1  g0608(.A(new_n799), .B1(new_n803), .B2(new_n808), .ZN(new_n809));
  NAND2_X1  g0609(.A1(new_n809), .A2(new_n724), .ZN(new_n810));
  NOR2_X1   g0610(.A1(new_n724), .A2(new_n721), .ZN(new_n811));
  AOI21_X1  g0611(.A(new_n708), .B1(new_n247), .B2(new_n811), .ZN(new_n812));
  NAND4_X1  g0612(.A1(new_n328), .A2(new_n324), .A3(new_n319), .A4(new_n637), .ZN(new_n813));
  XNOR2_X1  g0613(.A(new_n813), .B(KEYINPUT104), .ZN(new_n814));
  NAND2_X1  g0614(.A1(new_n324), .A2(new_n637), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n331), .A2(new_n815), .ZN(new_n816));
  NAND2_X1  g0616(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  OAI211_X1 g0617(.A(new_n810), .B(new_n812), .C1(new_n817), .C2(new_n722), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n664), .A2(new_n688), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n819), .A2(G330), .ZN(new_n820));
  INV_X1    g0620(.A(new_n817), .ZN(new_n821));
  XNOR2_X1  g0621(.A(new_n694), .B(new_n821), .ZN(new_n822));
  INV_X1    g0622(.A(new_n822), .ZN(new_n823));
  AOI21_X1  g0623(.A(new_n709), .B1(new_n820), .B2(new_n823), .ZN(new_n824));
  INV_X1    g0624(.A(new_n824), .ZN(new_n825));
  NOR2_X1   g0625(.A1(new_n820), .A2(new_n823), .ZN(new_n826));
  OAI21_X1  g0626(.A(new_n818), .B1(new_n825), .B2(new_n826), .ZN(G384));
  NOR2_X1   g0627(.A1(new_n679), .A2(new_n680), .ZN(new_n828));
  NOR2_X1   g0628(.A1(new_n828), .A2(new_n685), .ZN(new_n829));
  NAND2_X1  g0629(.A1(new_n664), .A2(new_n829), .ZN(new_n830));
  NAND3_X1  g0630(.A1(new_n375), .A2(KEYINPUT105), .A3(new_n377), .ZN(new_n831));
  NAND2_X1  g0631(.A1(new_n349), .A2(new_n637), .ZN(new_n832));
  NAND2_X1  g0632(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  INV_X1    g0633(.A(KEYINPUT105), .ZN(new_n834));
  NAND3_X1  g0634(.A1(new_n375), .A2(new_n834), .A3(new_n377), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n372), .A2(new_n374), .A3(new_n832), .ZN(new_n836));
  NAND2_X1  g0636(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g0637(.A1(new_n833), .A2(new_n837), .A3(new_n817), .ZN(new_n838));
  INV_X1    g0638(.A(new_n838), .ZN(new_n839));
  INV_X1    g0639(.A(KEYINPUT106), .ZN(new_n840));
  OAI21_X1  g0640(.A(new_n391), .B1(new_n389), .B2(new_n840), .ZN(new_n841));
  NOR3_X1   g0641(.A1(new_n385), .A2(new_n388), .A3(KEYINPUT106), .ZN(new_n842));
  OAI21_X1  g0642(.A(new_n390), .B1(new_n841), .B2(new_n842), .ZN(new_n843));
  AOI21_X1  g0643(.A(new_n635), .B1(new_n843), .B2(new_n404), .ZN(new_n844));
  NAND2_X1  g0644(.A1(new_n429), .A2(new_n844), .ZN(new_n845));
  NAND2_X1  g0645(.A1(new_n405), .A2(new_n416), .ZN(new_n846));
  INV_X1    g0646(.A(new_n635), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n405), .A2(new_n847), .ZN(new_n848));
  INV_X1    g0648(.A(KEYINPUT37), .ZN(new_n849));
  NAND4_X1  g0649(.A1(new_n846), .A2(new_n848), .A3(new_n849), .A4(new_n422), .ZN(new_n850));
  INV_X1    g0650(.A(new_n422), .ZN(new_n851));
  AOI22_X1  g0651(.A1(new_n415), .A2(new_n635), .B1(new_n404), .B2(new_n843), .ZN(new_n852));
  OAI21_X1  g0652(.A(KEYINPUT37), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  NAND2_X1  g0653(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NAND3_X1  g0654(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n855));
  OAI21_X1  g0655(.A(new_n422), .B1(new_n426), .B2(new_n415), .ZN(new_n856));
  NOR2_X1   g0656(.A1(new_n426), .A2(new_n635), .ZN(new_n857));
  OAI21_X1  g0657(.A(KEYINPUT37), .B1(new_n856), .B2(new_n857), .ZN(new_n858));
  AOI22_X1  g0658(.A1(new_n850), .A2(new_n858), .B1(new_n429), .B2(new_n857), .ZN(new_n859));
  OAI21_X1  g0659(.A(new_n855), .B1(new_n859), .B2(KEYINPUT38), .ZN(new_n860));
  NAND3_X1  g0660(.A1(new_n830), .A2(new_n839), .A3(new_n860), .ZN(new_n861));
  AOI21_X1  g0661(.A(new_n838), .B1(new_n664), .B2(new_n829), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n845), .A2(new_n854), .ZN(new_n863));
  INV_X1    g0663(.A(KEYINPUT38), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  AOI21_X1  g0665(.A(KEYINPUT40), .B1(new_n865), .B2(new_n855), .ZN(new_n866));
  AOI22_X1  g0666(.A1(new_n861), .A2(KEYINPUT40), .B1(new_n862), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(new_n867), .ZN(new_n868));
  AND2_X1   g0668(.A1(new_n830), .A2(new_n430), .ZN(new_n869));
  AND2_X1   g0669(.A1(new_n868), .A2(new_n869), .ZN(new_n870));
  NOR2_X1   g0670(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NOR3_X1   g0671(.A1(new_n870), .A2(new_n871), .A3(new_n662), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT39), .ZN(new_n873));
  NAND2_X1  g0673(.A1(new_n860), .A2(new_n873), .ZN(new_n874));
  OR2_X1    g0674(.A1(new_n375), .A2(new_n637), .ZN(new_n875));
  INV_X1    g0675(.A(new_n875), .ZN(new_n876));
  NAND3_X1  g0676(.A1(new_n865), .A2(KEYINPUT39), .A3(new_n855), .ZN(new_n877));
  NAND3_X1  g0677(.A1(new_n874), .A2(new_n876), .A3(new_n877), .ZN(new_n878));
  NAND2_X1  g0678(.A1(new_n605), .A2(new_n663), .ZN(new_n879));
  INV_X1    g0679(.A(new_n879), .ZN(new_n880));
  AOI21_X1  g0680(.A(new_n880), .B1(new_n694), .B2(new_n817), .ZN(new_n881));
  NAND2_X1  g0681(.A1(new_n833), .A2(new_n837), .ZN(new_n882));
  NOR2_X1   g0682(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g0683(.A1(new_n865), .A2(new_n855), .ZN(new_n884));
  AOI22_X1  g0684(.A1(new_n883), .A2(new_n884), .B1(new_n608), .B2(new_n635), .ZN(new_n885));
  NAND2_X1  g0685(.A1(new_n878), .A2(new_n885), .ZN(new_n886));
  NAND4_X1  g0686(.A1(new_n700), .A2(new_n430), .A3(new_n692), .A4(new_n695), .ZN(new_n887));
  NAND2_X1  g0687(.A1(new_n887), .A2(new_n610), .ZN(new_n888));
  XOR2_X1   g0688(.A(new_n886), .B(new_n888), .Z(new_n889));
  OAI22_X1  g0689(.A1(new_n872), .A2(new_n889), .B1(new_n205), .B2(new_n703), .ZN(new_n890));
  AOI21_X1  g0690(.A(new_n890), .B1(new_n889), .B2(new_n872), .ZN(new_n891));
  OR2_X1    g0691(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n551), .A2(KEYINPUT35), .ZN(new_n893));
  NAND4_X1  g0693(.A1(new_n892), .A2(G116), .A3(new_n215), .A4(new_n893), .ZN(new_n894));
  XOR2_X1   g0694(.A(new_n894), .B(KEYINPUT36), .Z(new_n895));
  OAI211_X1 g0695(.A(new_n213), .B(G77), .C1(new_n236), .C2(new_n337), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n273), .A2(G68), .ZN(new_n897));
  AOI211_X1 g0697(.A(new_n205), .B(G13), .C1(new_n896), .C2(new_n897), .ZN(new_n898));
  OR3_X1    g0698(.A1(new_n891), .A2(new_n895), .A3(new_n898), .ZN(G367));
  OAI211_X1 g0699(.A(new_n561), .B(new_n566), .C1(new_n563), .C2(new_n663), .ZN(new_n900));
  NAND2_X1  g0700(.A1(new_n619), .A2(new_n637), .ZN(new_n901));
  NAND2_X1  g0701(.A1(new_n900), .A2(new_n901), .ZN(new_n902));
  NAND3_X1  g0702(.A1(new_n536), .A2(new_n651), .A3(new_n902), .ZN(new_n903));
  OR2_X1    g0703(.A1(new_n903), .A2(KEYINPUT42), .ZN(new_n904));
  OAI21_X1  g0704(.A(new_n561), .B1(new_n900), .B2(new_n614), .ZN(new_n905));
  AOI22_X1  g0705(.A1(new_n903), .A2(KEYINPUT42), .B1(new_n663), .B2(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n597), .A2(new_n599), .ZN(new_n907));
  NAND2_X1  g0707(.A1(new_n907), .A2(new_n637), .ZN(new_n908));
  NAND3_X1  g0708(.A1(new_n908), .A2(new_n594), .A3(new_n600), .ZN(new_n909));
  OAI21_X1  g0709(.A(new_n909), .B1(new_n594), .B2(new_n908), .ZN(new_n910));
  AOI22_X1  g0710(.A1(new_n904), .A2(new_n906), .B1(KEYINPUT43), .B2(new_n910), .ZN(new_n911));
  OR2_X1    g0711(.A1(new_n910), .A2(KEYINPUT43), .ZN(new_n912));
  XNOR2_X1  g0712(.A(new_n911), .B(new_n912), .ZN(new_n913));
  INV_X1    g0713(.A(new_n902), .ZN(new_n914));
  NOR2_X1   g0714(.A1(new_n649), .A2(new_n914), .ZN(new_n915));
  XNOR2_X1  g0715(.A(new_n913), .B(new_n915), .ZN(new_n916));
  XOR2_X1   g0716(.A(new_n705), .B(KEYINPUT110), .Z(new_n917));
  XOR2_X1   g0717(.A(new_n655), .B(KEYINPUT41), .Z(new_n918));
  INV_X1    g0718(.A(KEYINPUT108), .ZN(new_n919));
  INV_X1    g0719(.A(new_n651), .ZN(new_n920));
  NAND3_X1  g0720(.A1(new_n645), .A2(new_n646), .A3(new_n920), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n651), .B1(new_n643), .B2(new_n644), .ZN(new_n922));
  NAND2_X1  g0722(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  XNOR2_X1  g0723(.A(new_n923), .B(new_n641), .ZN(new_n924));
  NAND3_X1  g0724(.A1(new_n700), .A2(new_n692), .A3(new_n695), .ZN(new_n925));
  NAND2_X1  g0725(.A1(new_n820), .A2(new_n925), .ZN(new_n926));
  OAI21_X1  g0726(.A(new_n919), .B1(new_n924), .B2(new_n926), .ZN(new_n927));
  NAND3_X1  g0727(.A1(new_n923), .A2(new_n784), .A3(G330), .ZN(new_n928));
  NAND3_X1  g0728(.A1(new_n641), .A2(new_n922), .A3(new_n921), .ZN(new_n929));
  NAND2_X1  g0729(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  NAND3_X1  g0730(.A1(new_n701), .A2(new_n930), .A3(KEYINPUT108), .ZN(new_n931));
  NAND3_X1  g0731(.A1(new_n652), .A2(KEYINPUT45), .A3(new_n902), .ZN(new_n932));
  INV_X1    g0732(.A(KEYINPUT45), .ZN(new_n933));
  INV_X1    g0733(.A(new_n650), .ZN(new_n934));
  NAND2_X1  g0734(.A1(new_n922), .A2(new_n934), .ZN(new_n935));
  OAI21_X1  g0735(.A(new_n933), .B1(new_n935), .B2(new_n914), .ZN(new_n936));
  NAND2_X1  g0736(.A1(new_n932), .A2(new_n936), .ZN(new_n937));
  XOR2_X1   g0737(.A(KEYINPUT107), .B(KEYINPUT44), .Z(new_n938));
  NAND3_X1  g0738(.A1(new_n935), .A2(new_n914), .A3(new_n938), .ZN(new_n939));
  INV_X1    g0739(.A(new_n938), .ZN(new_n940));
  OAI21_X1  g0740(.A(new_n940), .B1(new_n652), .B2(new_n902), .ZN(new_n941));
  NAND4_X1  g0741(.A1(new_n649), .A2(new_n937), .A3(new_n939), .A4(new_n941), .ZN(new_n942));
  AND2_X1   g0742(.A1(new_n932), .A2(new_n936), .ZN(new_n943));
  NAND2_X1  g0743(.A1(new_n941), .A2(new_n939), .ZN(new_n944));
  OAI21_X1  g0744(.A(new_n648), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND4_X1  g0745(.A1(new_n927), .A2(new_n931), .A3(new_n942), .A4(new_n945), .ZN(new_n946));
  AOI21_X1  g0746(.A(new_n918), .B1(new_n946), .B2(new_n701), .ZN(new_n947));
  OAI21_X1  g0747(.A(new_n917), .B1(new_n947), .B2(KEYINPUT109), .ZN(new_n948));
  INV_X1    g0748(.A(KEYINPUT109), .ZN(new_n949));
  AOI211_X1 g0749(.A(new_n949), .B(new_n918), .C1(new_n946), .C2(new_n701), .ZN(new_n950));
  OAI21_X1  g0750(.A(new_n916), .B1(new_n948), .B2(new_n950), .ZN(new_n951));
  AOI21_X1  g0751(.A(new_n726), .B1(new_n654), .B2(new_n588), .ZN(new_n952));
  NAND2_X1  g0752(.A1(new_n717), .A2(new_n233), .ZN(new_n953));
  AND2_X1   g0753(.A1(new_n952), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g0754(.A(new_n244), .B1(new_n749), .B2(new_n273), .ZN(new_n955));
  INV_X1    g0755(.A(G159), .ZN(new_n956));
  OAI22_X1  g0756(.A1(new_n768), .A2(new_n956), .B1(new_n757), .B2(new_n337), .ZN(new_n957));
  AOI211_X1 g0757(.A(new_n955), .B(new_n957), .C1(G143), .C2(new_n751), .ZN(new_n958));
  INV_X1    g0758(.A(new_n731), .ZN(new_n959));
  AOI22_X1  g0759(.A1(new_n959), .A2(G58), .B1(G137), .B2(new_n738), .ZN(new_n960));
  NAND2_X1  g0760(.A1(new_n745), .A2(G77), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n776), .A2(G150), .ZN(new_n962));
  NAND4_X1  g0762(.A1(new_n958), .A2(new_n960), .A3(new_n961), .A4(new_n962), .ZN(new_n963));
  OAI21_X1  g0763(.A(new_n383), .B1(new_n749), .B2(new_n792), .ZN(new_n964));
  OAI22_X1  g0764(.A1(new_n755), .A2(new_n768), .B1(new_n752), .B2(new_n747), .ZN(new_n965));
  AOI211_X1 g0765(.A(new_n964), .B(new_n965), .C1(new_n553), .C2(new_n758), .ZN(new_n966));
  NAND3_X1  g0766(.A1(new_n732), .A2(KEYINPUT46), .A3(G116), .ZN(new_n967));
  NAND2_X1  g0767(.A1(new_n738), .A2(G317), .ZN(new_n968));
  NOR2_X1   g0768(.A1(new_n744), .A2(new_n453), .ZN(new_n969));
  AOI21_X1  g0769(.A(new_n969), .B1(new_n776), .B2(G303), .ZN(new_n970));
  NAND4_X1  g0770(.A1(new_n966), .A2(new_n967), .A3(new_n968), .A4(new_n970), .ZN(new_n971));
  AOI21_X1  g0771(.A(KEYINPUT46), .B1(new_n959), .B2(G116), .ZN(new_n972));
  XNOR2_X1  g0772(.A(new_n972), .B(KEYINPUT111), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n963), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  XNOR2_X1  g0774(.A(KEYINPUT112), .B(KEYINPUT47), .ZN(new_n975));
  XOR2_X1   g0775(.A(new_n974), .B(new_n975), .Z(new_n976));
  AOI211_X1 g0776(.A(new_n708), .B(new_n954), .C1(new_n976), .C2(new_n724), .ZN(new_n977));
  OR2_X1    g0777(.A1(new_n977), .A2(KEYINPUT113), .ZN(new_n978));
  NAND2_X1  g0778(.A1(new_n977), .A2(KEYINPUT113), .ZN(new_n979));
  OAI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n785), .C2(new_n910), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n951), .A2(new_n980), .ZN(G387));
  NAND2_X1  g0781(.A1(new_n924), .A2(new_n926), .ZN(new_n982));
  NAND2_X1  g0782(.A1(new_n701), .A2(new_n930), .ZN(new_n983));
  NAND3_X1  g0783(.A1(new_n982), .A2(new_n983), .A3(new_n655), .ZN(new_n984));
  AND2_X1   g0784(.A1(new_n647), .A2(new_n723), .ZN(new_n985));
  OR2_X1    g0785(.A1(new_n230), .A2(new_n439), .ZN(new_n986));
  AOI22_X1  g0786(.A1(new_n986), .A2(new_n717), .B1(new_n658), .B2(new_n710), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n279), .A2(new_n273), .ZN(new_n988));
  XNOR2_X1  g0788(.A(new_n988), .B(KEYINPUT50), .ZN(new_n989));
  OAI21_X1  g0789(.A(new_n439), .B1(new_n337), .B2(new_n247), .ZN(new_n990));
  NOR3_X1   g0790(.A1(new_n989), .A2(new_n658), .A3(new_n990), .ZN(new_n991));
  OAI22_X1  g0791(.A1(new_n987), .A2(new_n991), .B1(G107), .B2(new_n209), .ZN(new_n992));
  AOI21_X1  g0792(.A(new_n708), .B1(new_n992), .B2(new_n725), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n765), .A2(new_n273), .B1(new_n805), .B2(new_n737), .ZN(new_n994));
  NOR2_X1   g0794(.A1(new_n757), .A2(new_n321), .ZN(new_n995));
  AOI21_X1  g0795(.A(new_n995), .B1(new_n767), .B2(new_n279), .ZN(new_n996));
  AOI21_X1  g0796(.A(new_n383), .B1(new_n774), .B2(G68), .ZN(new_n997));
  OAI211_X1 g0797(.A(new_n996), .B(new_n997), .C1(new_n956), .C2(new_n752), .ZN(new_n998));
  NOR2_X1   g0798(.A1(new_n731), .A2(new_n247), .ZN(new_n999));
  NOR4_X1   g0799(.A1(new_n994), .A2(new_n998), .A3(new_n969), .A4(new_n999), .ZN(new_n1000));
  AOI22_X1  g0800(.A1(G311), .A2(new_n767), .B1(new_n774), .B2(G303), .ZN(new_n1001));
  INV_X1    g0801(.A(G317), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1001), .B1(new_n766), .B2(new_n752), .C1(new_n765), .C2(new_n1002), .ZN(new_n1003));
  INV_X1    g0803(.A(KEYINPUT48), .ZN(new_n1004));
  AND2_X1   g0804(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1005));
  NOR2_X1   g0805(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1006));
  OAI22_X1  g0806(.A1(new_n731), .A2(new_n755), .B1(new_n757), .B2(new_n792), .ZN(new_n1007));
  OR3_X1    g0807(.A1(new_n1005), .A2(new_n1006), .A3(new_n1007), .ZN(new_n1008));
  INV_X1    g0808(.A(new_n1008), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n1009), .A2(KEYINPUT49), .ZN(new_n1010));
  OAI221_X1 g0810(.A(new_n383), .B1(new_n753), .B2(new_n737), .C1(new_n744), .C2(new_n455), .ZN(new_n1011));
  XOR2_X1   g0811(.A(new_n1011), .B(KEYINPUT114), .Z(new_n1012));
  AOI21_X1  g0812(.A(new_n1012), .B1(new_n1009), .B2(KEYINPUT49), .ZN(new_n1013));
  AOI21_X1  g0813(.A(new_n1000), .B1(new_n1010), .B2(new_n1013), .ZN(new_n1014));
  INV_X1    g0814(.A(new_n724), .ZN(new_n1015));
  OAI21_X1  g0815(.A(new_n993), .B1(new_n1014), .B2(new_n1015), .ZN(new_n1016));
  OAI221_X1 g0816(.A(new_n984), .B1(new_n924), .B2(new_n917), .C1(new_n985), .C2(new_n1016), .ZN(G393));
  NAND3_X1  g0817(.A1(new_n945), .A2(KEYINPUT115), .A3(new_n942), .ZN(new_n1018));
  OAI21_X1  g0818(.A(new_n1018), .B1(KEYINPUT115), .B2(new_n942), .ZN(new_n1019));
  INV_X1    g0819(.A(new_n983), .ZN(new_n1020));
  OAI211_X1 g0820(.A(new_n655), .B(new_n946), .C1(new_n1019), .C2(new_n1020), .ZN(new_n1021));
  INV_X1    g0821(.A(new_n917), .ZN(new_n1022));
  NAND2_X1  g0822(.A1(new_n914), .A2(new_n723), .ZN(new_n1023));
  OAI221_X1 g0823(.A(new_n725), .B1(new_n453), .B2(new_n209), .C1(new_n718), .C2(new_n242), .ZN(new_n1024));
  NAND2_X1  g0824(.A1(new_n709), .A2(new_n1024), .ZN(new_n1025));
  OAI221_X1 g0825(.A(new_n244), .B1(new_n403), .B2(new_n749), .C1(new_n768), .C2(new_n273), .ZN(new_n1026));
  AOI22_X1  g0826(.A1(new_n745), .A2(G87), .B1(G143), .B2(new_n738), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n1027), .B1(new_n337), .B2(new_n731), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1026), .B(new_n1028), .C1(G77), .C2(new_n758), .ZN(new_n1029));
  OAI22_X1  g0829(.A1(new_n765), .A2(new_n956), .B1(new_n805), .B2(new_n752), .ZN(new_n1030));
  XOR2_X1   g0830(.A(new_n1030), .B(KEYINPUT116), .Z(new_n1031));
  NAND2_X1  g0831(.A1(new_n1031), .A2(KEYINPUT51), .ZN(new_n1032));
  NAND2_X1  g0832(.A1(new_n1029), .A2(new_n1032), .ZN(new_n1033));
  NOR2_X1   g0833(.A1(new_n1031), .A2(KEYINPUT51), .ZN(new_n1034));
  OAI22_X1  g0834(.A1(new_n731), .A2(new_n792), .B1(new_n766), .B2(new_n737), .ZN(new_n1035));
  AOI211_X1 g0835(.A(new_n244), .B(new_n1035), .C1(G107), .C2(new_n745), .ZN(new_n1036));
  XOR2_X1   g0836(.A(new_n1036), .B(KEYINPUT117), .Z(new_n1037));
  OAI22_X1  g0837(.A1(new_n765), .A2(new_n747), .B1(new_n1002), .B2(new_n752), .ZN(new_n1038));
  XNOR2_X1  g0838(.A(new_n1038), .B(KEYINPUT52), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n767), .A2(G303), .ZN(new_n1040));
  AOI22_X1  g0840(.A1(new_n774), .A2(G294), .B1(new_n758), .B2(G116), .ZN(new_n1041));
  NAND3_X1  g0841(.A1(new_n1039), .A2(new_n1040), .A3(new_n1041), .ZN(new_n1042));
  OAI22_X1  g0842(.A1(new_n1033), .A2(new_n1034), .B1(new_n1037), .B2(new_n1042), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1025), .B1(new_n1043), .B2(new_n724), .ZN(new_n1044));
  AOI22_X1  g0844(.A1(new_n1019), .A2(new_n1022), .B1(new_n1023), .B2(new_n1044), .ZN(new_n1045));
  NAND2_X1  g0845(.A1(new_n1021), .A2(new_n1045), .ZN(G390));
  INV_X1    g0846(.A(new_n881), .ZN(new_n1047));
  AOI22_X1  g0847(.A1(new_n832), .A2(new_n831), .B1(new_n835), .B2(new_n836), .ZN(new_n1048));
  AOI21_X1  g0848(.A(new_n1048), .B1(new_n689), .B2(new_n817), .ZN(new_n1049));
  AND3_X1   g0849(.A1(new_n830), .A2(new_n839), .A3(G330), .ZN(new_n1050));
  OAI21_X1  g0850(.A(new_n1047), .B1(new_n1049), .B2(new_n1050), .ZN(new_n1051));
  NAND4_X1  g0851(.A1(new_n819), .A2(G330), .A3(new_n817), .A4(new_n1048), .ZN(new_n1052));
  AOI21_X1  g0852(.A(new_n880), .B1(new_n699), .B2(new_n817), .ZN(new_n1053));
  AOI211_X1 g0853(.A(new_n662), .B(new_n821), .C1(new_n664), .C2(new_n829), .ZN(new_n1054));
  OAI211_X1 g0854(.A(new_n1052), .B(new_n1053), .C1(new_n1054), .C2(new_n1048), .ZN(new_n1055));
  NAND2_X1  g0855(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n662), .B1(new_n664), .B2(new_n829), .ZN(new_n1057));
  NAND2_X1  g0857(.A1(new_n1057), .A2(new_n430), .ZN(new_n1058));
  NAND3_X1  g0858(.A1(new_n1058), .A2(new_n610), .A3(new_n887), .ZN(new_n1059));
  INV_X1    g0859(.A(new_n1059), .ZN(new_n1060));
  NAND2_X1  g0860(.A1(new_n1056), .A2(new_n1060), .ZN(new_n1061));
  AND3_X1   g0861(.A1(new_n625), .A2(new_n663), .A3(new_n817), .ZN(new_n1062));
  OAI21_X1  g0862(.A(new_n1048), .B1(new_n1062), .B2(new_n880), .ZN(new_n1063));
  AOI22_X1  g0863(.A1(new_n874), .A2(new_n877), .B1(new_n1063), .B2(new_n875), .ZN(new_n1064));
  NAND2_X1  g0864(.A1(new_n699), .A2(new_n817), .ZN(new_n1065));
  AOI21_X1  g0865(.A(new_n882), .B1(new_n1065), .B2(new_n879), .ZN(new_n1066));
  NAND2_X1  g0866(.A1(new_n860), .A2(new_n875), .ZN(new_n1067));
  NOR2_X1   g0867(.A1(new_n1066), .A2(new_n1067), .ZN(new_n1068));
  OAI21_X1  g0868(.A(new_n1050), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1069));
  NAND2_X1  g0869(.A1(new_n858), .A2(new_n850), .ZN(new_n1070));
  NAND2_X1  g0870(.A1(new_n429), .A2(new_n857), .ZN(new_n1071));
  NAND2_X1  g0871(.A1(new_n1070), .A2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g0872(.A1(new_n1072), .A2(new_n864), .ZN(new_n1073));
  AOI21_X1  g0873(.A(KEYINPUT39), .B1(new_n1073), .B2(new_n855), .ZN(new_n1074));
  AND3_X1   g0874(.A1(new_n845), .A2(KEYINPUT38), .A3(new_n854), .ZN(new_n1075));
  AOI21_X1  g0875(.A(KEYINPUT38), .B1(new_n845), .B2(new_n854), .ZN(new_n1076));
  NOR3_X1   g0876(.A1(new_n1075), .A2(new_n1076), .A3(new_n873), .ZN(new_n1077));
  OAI22_X1  g0877(.A1(new_n1074), .A2(new_n1077), .B1(new_n876), .B2(new_n883), .ZN(new_n1078));
  OAI211_X1 g0878(.A(new_n875), .B(new_n860), .C1(new_n1053), .C2(new_n882), .ZN(new_n1079));
  NAND3_X1  g0879(.A1(new_n1078), .A2(new_n1079), .A3(new_n1052), .ZN(new_n1080));
  NAND2_X1  g0880(.A1(new_n1069), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g0881(.A(new_n656), .B1(new_n1061), .B2(new_n1081), .ZN(new_n1082));
  OAI21_X1  g0882(.A(new_n1082), .B1(new_n1081), .B2(new_n1061), .ZN(new_n1083));
  INV_X1    g0883(.A(new_n1081), .ZN(new_n1084));
  OAI21_X1  g0884(.A(new_n721), .B1(new_n1074), .B2(new_n1077), .ZN(new_n1085));
  OAI21_X1  g0885(.A(new_n383), .B1(new_n749), .B2(new_n453), .ZN(new_n1086));
  INV_X1    g0886(.A(G283), .ZN(new_n1087));
  OAI22_X1  g0887(.A1(new_n1087), .A2(new_n752), .B1(new_n768), .B2(new_n311), .ZN(new_n1088));
  AOI211_X1 g0888(.A(new_n1086), .B(new_n1088), .C1(G77), .C2(new_n758), .ZN(new_n1089));
  NAND2_X1  g0889(.A1(new_n742), .A2(G294), .ZN(new_n1090));
  NAND2_X1  g0890(.A1(new_n732), .A2(G87), .ZN(new_n1091));
  AOI22_X1  g0891(.A1(new_n776), .A2(G116), .B1(G68), .B2(new_n745), .ZN(new_n1092));
  NAND4_X1  g0892(.A1(new_n1089), .A2(new_n1090), .A3(new_n1091), .A4(new_n1092), .ZN(new_n1093));
  XNOR2_X1  g0893(.A(KEYINPUT54), .B(G143), .ZN(new_n1094));
  OAI21_X1  g0894(.A(new_n244), .B1(new_n749), .B2(new_n1094), .ZN(new_n1095));
  INV_X1    g0895(.A(G128), .ZN(new_n1096));
  OAI22_X1  g0896(.A1(new_n752), .A2(new_n1096), .B1(new_n757), .B2(new_n956), .ZN(new_n1097));
  AOI211_X1 g0897(.A(new_n1095), .B(new_n1097), .C1(G137), .C2(new_n767), .ZN(new_n1098));
  NAND2_X1  g0898(.A1(new_n742), .A2(G125), .ZN(new_n1099));
  NOR2_X1   g0899(.A1(new_n731), .A2(new_n805), .ZN(new_n1100));
  XNOR2_X1  g0900(.A(new_n1100), .B(KEYINPUT53), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n776), .A2(G132), .B1(G50), .B2(new_n745), .ZN(new_n1102));
  NAND4_X1  g0902(.A1(new_n1098), .A2(new_n1099), .A3(new_n1101), .A4(new_n1102), .ZN(new_n1103));
  AOI21_X1  g0903(.A(new_n1015), .B1(new_n1093), .B2(new_n1103), .ZN(new_n1104));
  AOI211_X1 g0904(.A(new_n708), .B(new_n1104), .C1(new_n403), .C2(new_n811), .ZN(new_n1105));
  XOR2_X1   g0905(.A(new_n1105), .B(KEYINPUT118), .Z(new_n1106));
  AOI22_X1  g0906(.A1(new_n1084), .A2(new_n1022), .B1(new_n1085), .B2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g0907(.A1(new_n1083), .A2(new_n1107), .ZN(G378));
  AND2_X1   g0908(.A1(new_n1051), .A2(new_n1055), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1060), .B1(new_n1109), .B2(new_n1081), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1110), .A2(KEYINPUT57), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n309), .A2(new_n334), .ZN(new_n1112));
  AOI21_X1  g0912(.A(new_n635), .B1(new_n302), .B2(new_n303), .ZN(new_n1113));
  NAND2_X1  g0913(.A1(new_n1112), .A2(new_n1113), .ZN(new_n1114));
  INV_X1    g0914(.A(new_n1113), .ZN(new_n1115));
  NAND3_X1  g0915(.A1(new_n309), .A2(new_n334), .A3(new_n1115), .ZN(new_n1116));
  XNOR2_X1  g0916(.A(KEYINPUT55), .B(KEYINPUT56), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n1114), .A2(new_n1116), .A3(new_n1117), .ZN(new_n1118));
  INV_X1    g0918(.A(new_n1117), .ZN(new_n1119));
  AOI21_X1  g0919(.A(new_n1115), .B1(new_n309), .B2(new_n334), .ZN(new_n1120));
  INV_X1    g0920(.A(new_n334), .ZN(new_n1121));
  AOI211_X1 g0921(.A(new_n1121), .B(new_n1113), .C1(new_n306), .C2(new_n308), .ZN(new_n1122));
  OAI21_X1  g0922(.A(new_n1119), .B1(new_n1120), .B2(new_n1122), .ZN(new_n1123));
  NAND2_X1  g0923(.A1(new_n1118), .A2(new_n1123), .ZN(new_n1124));
  OAI21_X1  g0924(.A(new_n1124), .B1(new_n867), .B2(new_n662), .ZN(new_n1125));
  INV_X1    g0925(.A(KEYINPUT119), .ZN(new_n1126));
  NAND2_X1  g0926(.A1(new_n1124), .A2(new_n1126), .ZN(new_n1127));
  NAND3_X1  g0927(.A1(new_n1118), .A2(new_n1123), .A3(KEYINPUT119), .ZN(new_n1128));
  NAND2_X1  g0928(.A1(new_n1127), .A2(new_n1128), .ZN(new_n1129));
  INV_X1    g0929(.A(KEYINPUT40), .ZN(new_n1130));
  AOI21_X1  g0930(.A(new_n1130), .B1(new_n862), .B2(new_n860), .ZN(new_n1131));
  NAND2_X1  g0931(.A1(new_n830), .A2(new_n839), .ZN(new_n1132));
  OAI21_X1  g0932(.A(new_n1130), .B1(new_n1075), .B2(new_n1076), .ZN(new_n1133));
  NOR2_X1   g0933(.A1(new_n1132), .A2(new_n1133), .ZN(new_n1134));
  OAI211_X1 g0934(.A(new_n1129), .B(G330), .C1(new_n1131), .C2(new_n1134), .ZN(new_n1135));
  AND3_X1   g0935(.A1(new_n1125), .A2(new_n1135), .A3(new_n886), .ZN(new_n1136));
  AOI21_X1  g0936(.A(new_n886), .B1(new_n1125), .B2(new_n1135), .ZN(new_n1137));
  NOR2_X1   g0937(.A1(new_n1136), .A2(new_n1137), .ZN(new_n1138));
  OAI21_X1  g0938(.A(new_n655), .B1(new_n1111), .B2(new_n1138), .ZN(new_n1139));
  INV_X1    g0939(.A(KEYINPUT57), .ZN(new_n1140));
  INV_X1    g0940(.A(new_n1137), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1125), .A2(new_n1135), .A3(new_n886), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1141), .A2(KEYINPUT121), .A3(new_n1142), .ZN(new_n1143));
  INV_X1    g0943(.A(KEYINPUT121), .ZN(new_n1144));
  OAI21_X1  g0944(.A(new_n1144), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1145));
  NAND3_X1  g0945(.A1(new_n1143), .A2(new_n1145), .A3(new_n1110), .ZN(new_n1146));
  AOI21_X1  g0946(.A(new_n1139), .B1(new_n1140), .B2(new_n1146), .ZN(new_n1147));
  NAND3_X1  g0947(.A1(new_n1143), .A2(new_n1145), .A3(new_n1022), .ZN(new_n1148));
  AOI21_X1  g0948(.A(new_n708), .B1(new_n273), .B2(new_n811), .ZN(new_n1149));
  OAI211_X1 g0949(.A(new_n442), .B(new_n383), .C1(new_n749), .C2(new_n321), .ZN(new_n1150));
  OAI22_X1  g0950(.A1(new_n768), .A2(new_n453), .B1(new_n752), .B2(new_n455), .ZN(new_n1151));
  AOI211_X1 g0951(.A(new_n1150), .B(new_n1151), .C1(G68), .C2(new_n758), .ZN(new_n1152));
  NOR2_X1   g0952(.A1(new_n744), .A2(new_n236), .ZN(new_n1153));
  AOI211_X1 g0953(.A(new_n999), .B(new_n1153), .C1(G107), .C2(new_n776), .ZN(new_n1154));
  OAI211_X1 g0954(.A(new_n1152), .B(new_n1154), .C1(new_n1087), .C2(new_n741), .ZN(new_n1155));
  INV_X1    g0955(.A(KEYINPUT58), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1157));
  OR2_X1    g0957(.A1(new_n1155), .A2(new_n1156), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1094), .ZN(new_n1159));
  AOI22_X1  g0959(.A1(new_n776), .A2(G128), .B1(new_n959), .B2(new_n1159), .ZN(new_n1160));
  AOI22_X1  g0960(.A1(new_n774), .A2(G137), .B1(new_n758), .B2(G150), .ZN(new_n1161));
  AOI22_X1  g0961(.A1(new_n767), .A2(G132), .B1(new_n751), .B2(G125), .ZN(new_n1162));
  NAND3_X1  g0962(.A1(new_n1160), .A2(new_n1161), .A3(new_n1162), .ZN(new_n1163));
  OR2_X1    g0963(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1164));
  NAND2_X1  g0964(.A1(new_n1163), .A2(KEYINPUT59), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n745), .A2(G159), .ZN(new_n1166));
  AOI211_X1 g0966(.A(G33), .B(G41), .C1(new_n738), .C2(G124), .ZN(new_n1167));
  NAND4_X1  g0967(.A1(new_n1164), .A2(new_n1165), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI21_X1  g0968(.A(G50), .B1(new_n280), .B2(new_n442), .ZN(new_n1169));
  OAI21_X1  g0969(.A(new_n1169), .B1(new_n244), .B2(G41), .ZN(new_n1170));
  AND4_X1   g0970(.A1(new_n1157), .A2(new_n1158), .A3(new_n1168), .A4(new_n1170), .ZN(new_n1171));
  OAI21_X1  g0971(.A(new_n1149), .B1(new_n1171), .B2(new_n1015), .ZN(new_n1172));
  AOI21_X1  g0972(.A(new_n1172), .B1(new_n1129), .B2(new_n721), .ZN(new_n1173));
  XNOR2_X1  g0973(.A(new_n1173), .B(KEYINPUT120), .ZN(new_n1174));
  NAND2_X1  g0974(.A1(new_n1148), .A2(new_n1174), .ZN(new_n1175));
  OR2_X1    g0975(.A1(new_n1147), .A2(new_n1175), .ZN(G375));
  AOI22_X1  g0976(.A1(new_n732), .A2(G159), .B1(new_n742), .B2(G128), .ZN(new_n1177));
  XOR2_X1   g0977(.A(new_n1177), .B(KEYINPUT123), .Z(new_n1178));
  AOI22_X1  g0978(.A1(G132), .A2(new_n751), .B1(new_n767), .B2(new_n1159), .ZN(new_n1179));
  AOI21_X1  g0979(.A(new_n383), .B1(new_n774), .B2(G150), .ZN(new_n1180));
  OAI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(new_n273), .C2(new_n757), .ZN(new_n1181));
  AOI211_X1 g0981(.A(new_n1153), .B(new_n1181), .C1(G137), .C2(new_n776), .ZN(new_n1182));
  NAND2_X1  g0982(.A1(new_n1178), .A2(new_n1182), .ZN(new_n1183));
  OAI21_X1  g0983(.A(new_n961), .B1(new_n1087), .B2(new_n765), .ZN(new_n1184));
  OAI21_X1  g0984(.A(new_n383), .B1(new_n749), .B2(new_n311), .ZN(new_n1185));
  NAND2_X1  g0985(.A1(new_n751), .A2(G294), .ZN(new_n1186));
  OAI21_X1  g0986(.A(new_n1186), .B1(new_n768), .B2(new_n455), .ZN(new_n1187));
  NOR4_X1   g0987(.A1(new_n1184), .A2(new_n995), .A3(new_n1185), .A4(new_n1187), .ZN(new_n1188));
  OAI221_X1 g0988(.A(new_n1188), .B1(new_n453), .B2(new_n798), .C1(new_n793), .C2(new_n741), .ZN(new_n1189));
  AOI21_X1  g0989(.A(new_n1015), .B1(new_n1183), .B2(new_n1189), .ZN(new_n1190));
  AOI211_X1 g0990(.A(new_n708), .B(new_n1190), .C1(new_n337), .C2(new_n811), .ZN(new_n1191));
  OAI21_X1  g0991(.A(new_n1191), .B1(new_n1048), .B2(new_n722), .ZN(new_n1192));
  AOI21_X1  g0992(.A(new_n917), .B1(new_n1051), .B2(new_n1055), .ZN(new_n1193));
  OAI21_X1  g0993(.A(new_n1192), .B1(new_n1193), .B2(KEYINPUT122), .ZN(new_n1194));
  INV_X1    g0994(.A(KEYINPUT122), .ZN(new_n1195));
  AOI211_X1 g0995(.A(new_n1195), .B(new_n917), .C1(new_n1051), .C2(new_n1055), .ZN(new_n1196));
  NOR2_X1   g0996(.A1(new_n1194), .A2(new_n1196), .ZN(new_n1197));
  INV_X1    g0997(.A(new_n918), .ZN(new_n1198));
  NAND3_X1  g0998(.A1(new_n1051), .A2(new_n1059), .A3(new_n1055), .ZN(new_n1199));
  NAND3_X1  g0999(.A1(new_n1061), .A2(new_n1198), .A3(new_n1199), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1197), .A2(new_n1200), .ZN(G381));
  OR3_X1    g1001(.A1(new_n1147), .A2(G378), .A3(new_n1175), .ZN(new_n1202));
  INV_X1    g1002(.A(KEYINPUT124), .ZN(new_n1203));
  OR2_X1    g1003(.A1(G393), .A2(G396), .ZN(new_n1204));
  NOR4_X1   g1004(.A1(G390), .A2(G381), .A3(new_n1204), .A4(G384), .ZN(new_n1205));
  NAND3_X1  g1005(.A1(new_n1205), .A2(new_n951), .A3(new_n980), .ZN(new_n1206));
  AOI21_X1  g1006(.A(new_n1202), .B1(new_n1203), .B2(new_n1206), .ZN(new_n1207));
  OAI21_X1  g1007(.A(new_n1207), .B1(new_n1203), .B2(new_n1206), .ZN(G407));
  OAI211_X1 g1008(.A(G407), .B(G213), .C1(G343), .C2(new_n1202), .ZN(G409));
  OAI21_X1  g1009(.A(G378), .B1(new_n1147), .B2(new_n1175), .ZN(new_n1210));
  OAI21_X1  g1010(.A(new_n1022), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1211));
  AND4_X1   g1011(.A1(new_n1083), .A2(new_n1211), .A3(new_n1107), .A4(new_n1174), .ZN(new_n1212));
  NAND4_X1  g1012(.A1(new_n1143), .A2(new_n1145), .A3(new_n1198), .A4(new_n1110), .ZN(new_n1213));
  AOI22_X1  g1013(.A1(new_n1212), .A2(new_n1213), .B1(G213), .B2(new_n636), .ZN(new_n1214));
  NAND2_X1  g1014(.A1(new_n1199), .A2(KEYINPUT60), .ZN(new_n1215));
  INV_X1    g1015(.A(KEYINPUT60), .ZN(new_n1216));
  NAND4_X1  g1016(.A1(new_n1051), .A2(new_n1216), .A3(new_n1059), .A4(new_n1055), .ZN(new_n1217));
  NAND2_X1  g1017(.A1(new_n1215), .A2(new_n1217), .ZN(new_n1218));
  AOI21_X1  g1018(.A(new_n656), .B1(new_n1056), .B2(new_n1060), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1218), .A2(new_n1219), .ZN(new_n1220));
  AND3_X1   g1020(.A1(new_n1220), .A2(new_n1197), .A3(G384), .ZN(new_n1221));
  AOI21_X1  g1021(.A(G384), .B1(new_n1220), .B2(new_n1197), .ZN(new_n1222));
  NOR2_X1   g1022(.A1(new_n1221), .A2(new_n1222), .ZN(new_n1223));
  NAND3_X1  g1023(.A1(new_n1210), .A2(new_n1214), .A3(new_n1223), .ZN(new_n1224));
  NAND2_X1  g1024(.A1(new_n1224), .A2(KEYINPUT62), .ZN(new_n1225));
  NAND2_X1  g1025(.A1(new_n1210), .A2(new_n1214), .ZN(new_n1226));
  NAND3_X1  g1026(.A1(new_n636), .A2(G213), .A3(G2897), .ZN(new_n1227));
  INV_X1    g1027(.A(new_n1227), .ZN(new_n1228));
  OAI21_X1  g1028(.A(new_n1228), .B1(new_n1221), .B2(new_n1222), .ZN(new_n1229));
  INV_X1    g1029(.A(G384), .ZN(new_n1230));
  NAND2_X1  g1030(.A1(new_n1061), .A2(new_n655), .ZN(new_n1231));
  AOI21_X1  g1031(.A(new_n1231), .B1(new_n1215), .B2(new_n1217), .ZN(new_n1232));
  INV_X1    g1032(.A(new_n1196), .ZN(new_n1233));
  OAI21_X1  g1033(.A(new_n1195), .B1(new_n1109), .B2(new_n917), .ZN(new_n1234));
  NAND3_X1  g1034(.A1(new_n1233), .A2(new_n1234), .A3(new_n1192), .ZN(new_n1235));
  OAI21_X1  g1035(.A(new_n1230), .B1(new_n1232), .B2(new_n1235), .ZN(new_n1236));
  NAND3_X1  g1036(.A1(new_n1220), .A2(new_n1197), .A3(G384), .ZN(new_n1237));
  NAND3_X1  g1037(.A1(new_n1236), .A2(new_n1237), .A3(new_n1227), .ZN(new_n1238));
  NAND2_X1  g1038(.A1(new_n1229), .A2(new_n1238), .ZN(new_n1239));
  INV_X1    g1039(.A(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1226), .A2(new_n1240), .ZN(new_n1241));
  INV_X1    g1041(.A(KEYINPUT61), .ZN(new_n1242));
  INV_X1    g1042(.A(KEYINPUT62), .ZN(new_n1243));
  NAND4_X1  g1043(.A1(new_n1210), .A2(new_n1243), .A3(new_n1214), .A4(new_n1223), .ZN(new_n1244));
  NAND4_X1  g1044(.A1(new_n1225), .A2(new_n1241), .A3(new_n1242), .A4(new_n1244), .ZN(new_n1245));
  INV_X1    g1045(.A(G390), .ZN(new_n1246));
  AOI21_X1  g1046(.A(KEYINPUT125), .B1(G387), .B2(new_n1246), .ZN(new_n1247));
  XOR2_X1   g1047(.A(G393), .B(G396), .Z(new_n1248));
  NAND3_X1  g1048(.A1(new_n951), .A2(G390), .A3(new_n980), .ZN(new_n1249));
  INV_X1    g1049(.A(new_n1249), .ZN(new_n1250));
  AOI21_X1  g1050(.A(G390), .B1(new_n951), .B2(new_n980), .ZN(new_n1251));
  OAI22_X1  g1051(.A1(new_n1247), .A2(new_n1248), .B1(new_n1250), .B2(new_n1251), .ZN(new_n1252));
  INV_X1    g1052(.A(new_n1252), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1251), .ZN(new_n1254));
  INV_X1    g1054(.A(new_n1248), .ZN(new_n1255));
  NAND4_X1  g1055(.A1(new_n1254), .A2(KEYINPUT125), .A3(new_n1249), .A4(new_n1255), .ZN(new_n1256));
  INV_X1    g1056(.A(new_n1256), .ZN(new_n1257));
  NOR2_X1   g1057(.A1(new_n1253), .A2(new_n1257), .ZN(new_n1258));
  NAND2_X1  g1058(.A1(new_n1245), .A2(new_n1258), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT63), .ZN(new_n1260));
  OR2_X1    g1060(.A1(new_n1224), .A2(new_n1260), .ZN(new_n1261));
  AOI21_X1  g1061(.A(new_n1239), .B1(new_n1210), .B2(new_n1214), .ZN(new_n1262));
  OAI21_X1  g1062(.A(new_n1224), .B1(new_n1262), .B2(new_n1260), .ZN(new_n1263));
  AOI21_X1  g1063(.A(KEYINPUT61), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1264));
  INV_X1    g1064(.A(KEYINPUT126), .ZN(new_n1265));
  OAI211_X1 g1065(.A(new_n1261), .B(new_n1263), .C1(new_n1264), .C2(new_n1265), .ZN(new_n1266));
  AOI211_X1 g1066(.A(KEYINPUT126), .B(KEYINPUT61), .C1(new_n1252), .C2(new_n1256), .ZN(new_n1267));
  OAI21_X1  g1067(.A(new_n1259), .B1(new_n1266), .B2(new_n1267), .ZN(G405));
  INV_X1    g1068(.A(new_n1223), .ZN(new_n1269));
  NAND2_X1  g1069(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1270));
  NAND3_X1  g1070(.A1(new_n1202), .A2(new_n1210), .A3(new_n1270), .ZN(new_n1271));
  NOR2_X1   g1071(.A1(new_n1269), .A2(KEYINPUT127), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1272), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1252), .A2(new_n1256), .A3(new_n1273), .ZN(new_n1274));
  INV_X1    g1074(.A(new_n1274), .ZN(new_n1275));
  AOI21_X1  g1075(.A(new_n1273), .B1(new_n1252), .B2(new_n1256), .ZN(new_n1276));
  OAI21_X1  g1076(.A(new_n1271), .B1(new_n1275), .B2(new_n1276), .ZN(new_n1277));
  INV_X1    g1077(.A(new_n1276), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n1271), .ZN(new_n1279));
  NAND3_X1  g1079(.A1(new_n1278), .A2(new_n1279), .A3(new_n1274), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1277), .A2(new_n1280), .ZN(G402));
endmodule


