//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 1 1 0 1 1 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 0 1 1 0 0 0 0 1 0 1 0 0 1 0 0 1 1 1 0 1 1 0 0 1 1 0 1 0 0 1 1 1 1 0 1 0 0 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:31:55 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n447, new_n449, new_n452, new_n453, new_n454, new_n455,
    new_n458, new_n459, new_n460, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n562, new_n564, new_n565, new_n566,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n573, new_n574,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n592, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n623, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n667, new_n668, new_n669, new_n670, new_n671, new_n672,
    new_n673, new_n674, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n687,
    new_n688, new_n689, new_n690, new_n691, new_n692, new_n693, new_n694,
    new_n695, new_n696, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1168, new_n1169, new_n1170;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT64), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  XNOR2_X1  g020(.A(KEYINPUT65), .B(KEYINPUT1), .ZN(new_n446));
  AND2_X1   g021(.A1(G7), .A2(G661), .ZN(new_n447));
  XNOR2_X1  g022(.A(new_n446), .B(new_n447), .ZN(G223));
  NAND2_X1  g023(.A1(new_n447), .A2(G567), .ZN(new_n449));
  XNOR2_X1  g024(.A(new_n449), .B(KEYINPUT66), .ZN(G234));
  NAND2_X1  g025(.A1(new_n447), .A2(G2106), .ZN(G217));
  NOR4_X1   g026(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NOR4_X1   g028(.A1(G237), .A2(G235), .A3(G238), .A4(G236), .ZN(new_n454));
  NAND2_X1  g029(.A1(new_n453), .A2(new_n454), .ZN(new_n455));
  XOR2_X1   g030(.A(new_n455), .B(KEYINPUT67), .Z(G261));
  INV_X1    g031(.A(G261), .ZN(G325));
  INV_X1    g032(.A(G2106), .ZN(new_n458));
  INV_X1    g033(.A(G567), .ZN(new_n459));
  OAI22_X1  g034(.A1(new_n453), .A2(new_n458), .B1(new_n459), .B2(new_n454), .ZN(new_n460));
  XOR2_X1   g035(.A(new_n460), .B(KEYINPUT68), .Z(G319));
  XNOR2_X1  g036(.A(KEYINPUT3), .B(G2104), .ZN(new_n462));
  NAND2_X1  g037(.A1(new_n462), .A2(G137), .ZN(new_n463));
  NAND2_X1  g038(.A1(G101), .A2(G2104), .ZN(new_n464));
  AOI21_X1  g039(.A(G2105), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  INV_X1    g040(.A(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(KEYINPUT3), .ZN(new_n467));
  INV_X1    g042(.A(KEYINPUT3), .ZN(new_n468));
  NAND2_X1  g043(.A1(new_n468), .A2(G2104), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n467), .A2(new_n469), .A3(G125), .ZN(new_n470));
  INV_X1    g045(.A(KEYINPUT69), .ZN(new_n471));
  AOI22_X1  g046(.A1(new_n470), .A2(new_n471), .B1(G113), .B2(G2104), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n462), .A2(KEYINPUT69), .A3(G125), .ZN(new_n473));
  NAND2_X1  g048(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n465), .B1(new_n474), .B2(G2105), .ZN(new_n475));
  XNOR2_X1  g050(.A(new_n475), .B(KEYINPUT70), .ZN(G160));
  NAND2_X1  g051(.A1(new_n467), .A2(new_n469), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(KEYINPUT71), .ZN(new_n478));
  INV_X1    g053(.A(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n462), .A2(new_n479), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n478), .A2(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(G2105), .ZN(new_n482));
  NOR2_X1   g057(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  AOI21_X1  g058(.A(KEYINPUT72), .B1(new_n483), .B2(G124), .ZN(new_n484));
  OR2_X1    g059(.A1(G100), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G112), .C2(new_n482), .ZN(new_n486));
  XNOR2_X1  g061(.A(new_n486), .B(KEYINPUT73), .ZN(new_n487));
  NAND3_X1  g062(.A1(new_n478), .A2(new_n480), .A3(new_n482), .ZN(new_n488));
  INV_X1    g063(.A(G136), .ZN(new_n489));
  NOR2_X1   g064(.A1(new_n488), .A2(new_n489), .ZN(new_n490));
  NOR3_X1   g065(.A1(new_n484), .A2(new_n487), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n483), .A2(KEYINPUT72), .A3(G124), .ZN(new_n492));
  NAND2_X1  g067(.A1(new_n491), .A2(new_n492), .ZN(new_n493));
  INV_X1    g068(.A(new_n493), .ZN(G162));
  NOR2_X1   g069(.A1(new_n466), .A2(G2105), .ZN(new_n495));
  NAND2_X1  g070(.A1(new_n495), .A2(G102), .ZN(new_n496));
  AOI22_X1  g071(.A1(new_n462), .A2(G126), .B1(G114), .B2(G2104), .ZN(new_n497));
  OAI21_X1  g072(.A(new_n496), .B1(new_n497), .B2(new_n482), .ZN(new_n498));
  INV_X1    g073(.A(KEYINPUT4), .ZN(new_n499));
  INV_X1    g074(.A(G138), .ZN(new_n500));
  NOR2_X1   g075(.A1(new_n500), .A2(G2105), .ZN(new_n501));
  AOI21_X1  g076(.A(new_n499), .B1(new_n462), .B2(new_n501), .ZN(new_n502));
  AND4_X1   g077(.A1(new_n499), .A2(new_n501), .A3(new_n467), .A4(new_n469), .ZN(new_n503));
  NOR2_X1   g078(.A1(new_n502), .A2(new_n503), .ZN(new_n504));
  OAI21_X1  g079(.A(KEYINPUT74), .B1(new_n498), .B2(new_n504), .ZN(new_n505));
  NAND3_X1  g080(.A1(new_n467), .A2(new_n469), .A3(G126), .ZN(new_n506));
  NAND2_X1  g081(.A1(G114), .A2(G2104), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(new_n507), .ZN(new_n508));
  AOI22_X1  g083(.A1(new_n508), .A2(G2105), .B1(G102), .B2(new_n495), .ZN(new_n509));
  INV_X1    g084(.A(KEYINPUT74), .ZN(new_n510));
  NAND3_X1  g085(.A1(new_n501), .A2(new_n467), .A3(new_n469), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT4), .ZN(new_n512));
  NAND3_X1  g087(.A1(new_n462), .A2(new_n499), .A3(new_n501), .ZN(new_n513));
  NAND2_X1  g088(.A1(new_n512), .A2(new_n513), .ZN(new_n514));
  NAND3_X1  g089(.A1(new_n509), .A2(new_n510), .A3(new_n514), .ZN(new_n515));
  NAND2_X1  g090(.A1(new_n505), .A2(new_n515), .ZN(G164));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  XNOR2_X1  g092(.A(KEYINPUT6), .B(G651), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g094(.A(G88), .ZN(new_n520));
  NAND2_X1  g095(.A1(new_n518), .A2(G543), .ZN(new_n521));
  INV_X1    g096(.A(G50), .ZN(new_n522));
  OAI22_X1  g097(.A1(new_n519), .A2(new_n520), .B1(new_n521), .B2(new_n522), .ZN(new_n523));
  AOI22_X1  g098(.A1(new_n517), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n524));
  INV_X1    g099(.A(G651), .ZN(new_n525));
  NOR2_X1   g100(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  OR2_X1    g101(.A1(new_n523), .A2(new_n526), .ZN(G303));
  INV_X1    g102(.A(G303), .ZN(G166));
  NAND3_X1  g103(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n529));
  XNOR2_X1  g104(.A(new_n529), .B(KEYINPUT75), .ZN(new_n530));
  XOR2_X1   g105(.A(new_n530), .B(KEYINPUT7), .Z(new_n531));
  NAND3_X1  g106(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n532));
  INV_X1    g107(.A(G51), .ZN(new_n533));
  INV_X1    g108(.A(G89), .ZN(new_n534));
  OAI221_X1 g109(.A(new_n532), .B1(new_n521), .B2(new_n533), .C1(new_n534), .C2(new_n519), .ZN(new_n535));
  NOR2_X1   g110(.A1(new_n531), .A2(new_n535), .ZN(G168));
  INV_X1    g111(.A(new_n519), .ZN(new_n537));
  INV_X1    g112(.A(new_n521), .ZN(new_n538));
  AOI22_X1  g113(.A1(G90), .A2(new_n537), .B1(new_n538), .B2(G52), .ZN(new_n539));
  NAND2_X1  g114(.A1(G77), .A2(G543), .ZN(new_n540));
  INV_X1    g115(.A(G543), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n541), .A2(KEYINPUT5), .ZN(new_n542));
  INV_X1    g117(.A(KEYINPUT5), .ZN(new_n543));
  NAND2_X1  g118(.A1(new_n543), .A2(G543), .ZN(new_n544));
  NAND2_X1  g119(.A1(new_n542), .A2(new_n544), .ZN(new_n545));
  INV_X1    g120(.A(G64), .ZN(new_n546));
  OAI21_X1  g121(.A(new_n540), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  NAND2_X1  g122(.A1(new_n547), .A2(G651), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT76), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n548), .A2(new_n549), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n547), .A2(KEYINPUT76), .A3(G651), .ZN(new_n551));
  NAND3_X1  g126(.A1(new_n539), .A2(new_n550), .A3(new_n551), .ZN(G301));
  INV_X1    g127(.A(G301), .ZN(G171));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  INV_X1    g129(.A(G43), .ZN(new_n555));
  OAI22_X1  g130(.A1(new_n519), .A2(new_n554), .B1(new_n521), .B2(new_n555), .ZN(new_n556));
  AOI22_X1  g131(.A1(new_n517), .A2(G56), .B1(G68), .B2(G543), .ZN(new_n557));
  NOR2_X1   g132(.A1(new_n557), .A2(new_n525), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n556), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT77), .Z(G153));
  AND3_X1   g136(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n562));
  NAND2_X1  g137(.A1(new_n562), .A2(G36), .ZN(G176));
  XOR2_X1   g138(.A(KEYINPUT78), .B(KEYINPUT8), .Z(new_n564));
  NAND2_X1  g139(.A1(G1), .A2(G3), .ZN(new_n565));
  XNOR2_X1  g140(.A(new_n564), .B(new_n565), .ZN(new_n566));
  NAND2_X1  g141(.A1(new_n562), .A2(new_n566), .ZN(G188));
  NAND3_X1  g142(.A1(new_n518), .A2(G53), .A3(G543), .ZN(new_n568));
  XNOR2_X1  g143(.A(new_n568), .B(KEYINPUT9), .ZN(new_n569));
  AOI22_X1  g144(.A1(new_n517), .A2(G65), .B1(G78), .B2(G543), .ZN(new_n570));
  OR2_X1    g145(.A1(new_n570), .A2(new_n525), .ZN(new_n571));
  AND3_X1   g146(.A1(new_n517), .A2(new_n518), .A3(KEYINPUT79), .ZN(new_n572));
  AOI21_X1  g147(.A(KEYINPUT79), .B1(new_n517), .B2(new_n518), .ZN(new_n573));
  OAI21_X1  g148(.A(G91), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(G299));
  INV_X1    g150(.A(G168), .ZN(G286));
  OAI21_X1  g151(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n577));
  INV_X1    g152(.A(G49), .ZN(new_n578));
  OAI21_X1  g153(.A(new_n577), .B1(new_n578), .B2(new_n521), .ZN(new_n579));
  OR2_X1    g154(.A1(new_n572), .A2(new_n573), .ZN(new_n580));
  AOI21_X1  g155(.A(new_n579), .B1(new_n580), .B2(G87), .ZN(new_n581));
  INV_X1    g156(.A(new_n581), .ZN(G288));
  NAND4_X1  g157(.A1(new_n518), .A2(KEYINPUT80), .A3(G48), .A4(G543), .ZN(new_n583));
  NAND2_X1  g158(.A1(new_n525), .A2(KEYINPUT6), .ZN(new_n584));
  INV_X1    g159(.A(KEYINPUT6), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n585), .A2(G651), .ZN(new_n586));
  NAND4_X1  g161(.A1(new_n584), .A2(new_n586), .A3(G48), .A4(G543), .ZN(new_n587));
  INV_X1    g162(.A(KEYINPUT80), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n587), .A2(new_n588), .ZN(new_n589));
  AOI22_X1  g164(.A1(new_n517), .A2(G61), .B1(G73), .B2(G543), .ZN(new_n590));
  OAI211_X1 g165(.A(new_n583), .B(new_n589), .C1(new_n590), .C2(new_n525), .ZN(new_n591));
  AOI21_X1  g166(.A(new_n591), .B1(new_n580), .B2(G86), .ZN(new_n592));
  INV_X1    g167(.A(new_n592), .ZN(G305));
  INV_X1    g168(.A(G85), .ZN(new_n594));
  INV_X1    g169(.A(G47), .ZN(new_n595));
  OAI22_X1  g170(.A1(new_n519), .A2(new_n594), .B1(new_n521), .B2(new_n595), .ZN(new_n596));
  AOI22_X1  g171(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n597), .A2(new_n525), .ZN(new_n598));
  INV_X1    g173(.A(KEYINPUT81), .ZN(new_n599));
  OR3_X1    g174(.A1(new_n596), .A2(new_n598), .A3(new_n599), .ZN(new_n600));
  OAI21_X1  g175(.A(new_n599), .B1(new_n596), .B2(new_n598), .ZN(new_n601));
  NAND2_X1  g176(.A1(new_n600), .A2(new_n601), .ZN(G290));
  NAND2_X1  g177(.A1(G301), .A2(G868), .ZN(new_n603));
  NAND2_X1  g178(.A1(G79), .A2(G543), .ZN(new_n604));
  INV_X1    g179(.A(G66), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n604), .B1(new_n545), .B2(new_n605), .ZN(new_n606));
  AOI22_X1  g181(.A1(G54), .A2(new_n538), .B1(new_n606), .B2(G651), .ZN(new_n607));
  OAI21_X1  g182(.A(G92), .B1(new_n572), .B2(new_n573), .ZN(new_n608));
  INV_X1    g183(.A(KEYINPUT10), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n608), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n608), .A2(new_n609), .ZN(new_n611));
  OAI21_X1  g186(.A(new_n607), .B1(new_n610), .B2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n603), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  INV_X1    g191(.A(G299), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(G868), .B2(new_n617), .ZN(G280));
  XOR2_X1   g194(.A(KEYINPUT82), .B(G559), .Z(new_n620));
  OAI21_X1  g195(.A(new_n613), .B1(G860), .B2(new_n620), .ZN(G148));
  NAND2_X1  g196(.A1(new_n613), .A2(new_n620), .ZN(new_n622));
  NAND2_X1  g197(.A1(new_n622), .A2(G868), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n623), .B1(G868), .B2(new_n559), .ZN(G323));
  XNOR2_X1  g199(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g200(.A1(new_n462), .A2(new_n495), .ZN(new_n626));
  XNOR2_X1  g201(.A(new_n626), .B(KEYINPUT12), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT13), .ZN(new_n628));
  XNOR2_X1  g203(.A(new_n628), .B(G2100), .ZN(new_n629));
  NAND2_X1  g204(.A1(new_n483), .A2(G123), .ZN(new_n630));
  INV_X1    g205(.A(new_n488), .ZN(new_n631));
  NAND2_X1  g206(.A1(new_n631), .A2(G135), .ZN(new_n632));
  OR2_X1    g207(.A1(G99), .A2(G2105), .ZN(new_n633));
  OAI211_X1 g208(.A(new_n633), .B(G2104), .C1(G111), .C2(new_n482), .ZN(new_n634));
  NAND3_X1  g209(.A1(new_n630), .A2(new_n632), .A3(new_n634), .ZN(new_n635));
  INV_X1    g210(.A(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(KEYINPUT83), .B(G2096), .ZN(new_n637));
  OR2_X1    g212(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  NAND2_X1  g213(.A1(new_n636), .A2(new_n637), .ZN(new_n639));
  NAND3_X1  g214(.A1(new_n629), .A2(new_n638), .A3(new_n639), .ZN(G156));
  XOR2_X1   g215(.A(G2427), .B(G2430), .Z(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT85), .B(G2438), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  XOR2_X1   g218(.A(KEYINPUT15), .B(G2435), .Z(new_n644));
  OR2_X1    g219(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  NAND2_X1  g220(.A1(new_n643), .A2(new_n644), .ZN(new_n646));
  NAND3_X1  g221(.A1(new_n645), .A2(KEYINPUT14), .A3(new_n646), .ZN(new_n647));
  XOR2_X1   g222(.A(KEYINPUT84), .B(KEYINPUT16), .Z(new_n648));
  XNOR2_X1  g223(.A(new_n647), .B(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G2443), .B(G2446), .ZN(new_n650));
  XNOR2_X1  g225(.A(G2451), .B(G2454), .ZN(new_n651));
  XNOR2_X1  g226(.A(new_n650), .B(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(new_n649), .B(new_n652), .ZN(new_n653));
  XNOR2_X1  g228(.A(G1341), .B(G1348), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(KEYINPUT86), .ZN(new_n655));
  NOR2_X1   g230(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(new_n656), .B(KEYINPUT87), .ZN(new_n657));
  INV_X1    g232(.A(G14), .ZN(new_n658));
  AOI21_X1  g233(.A(new_n658), .B1(new_n653), .B2(new_n655), .ZN(new_n659));
  AND2_X1   g234(.A1(new_n657), .A2(new_n659), .ZN(G401));
  XNOR2_X1  g235(.A(G2067), .B(G2678), .ZN(new_n661));
  XNOR2_X1  g236(.A(new_n661), .B(KEYINPUT88), .ZN(new_n662));
  XOR2_X1   g237(.A(G2072), .B(G2078), .Z(new_n663));
  XNOR2_X1  g238(.A(G2084), .B(G2090), .ZN(new_n664));
  NOR3_X1   g239(.A1(new_n662), .A2(new_n663), .A3(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(new_n665), .B(KEYINPUT18), .ZN(new_n666));
  NAND2_X1  g241(.A1(new_n662), .A2(new_n664), .ZN(new_n667));
  INV_X1    g242(.A(new_n663), .ZN(new_n668));
  NAND3_X1  g243(.A1(new_n667), .A2(KEYINPUT17), .A3(new_n668), .ZN(new_n669));
  OAI21_X1  g244(.A(new_n669), .B1(new_n662), .B2(new_n664), .ZN(new_n670));
  AOI21_X1  g245(.A(new_n668), .B1(new_n667), .B2(KEYINPUT17), .ZN(new_n671));
  OAI21_X1  g246(.A(new_n666), .B1(new_n670), .B2(new_n671), .ZN(new_n672));
  XNOR2_X1  g247(.A(new_n672), .B(G2100), .ZN(new_n673));
  XNOR2_X1  g248(.A(KEYINPUT89), .B(G2096), .ZN(new_n674));
  XNOR2_X1  g249(.A(new_n673), .B(new_n674), .ZN(G227));
  XNOR2_X1  g250(.A(G1971), .B(G1976), .ZN(new_n676));
  INV_X1    g251(.A(KEYINPUT19), .ZN(new_n677));
  XNOR2_X1  g252(.A(new_n676), .B(new_n677), .ZN(new_n678));
  XOR2_X1   g253(.A(G1956), .B(G2474), .Z(new_n679));
  XOR2_X1   g254(.A(G1961), .B(G1966), .Z(new_n680));
  NAND3_X1  g255(.A1(new_n678), .A2(new_n679), .A3(new_n680), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT20), .ZN(new_n682));
  OR2_X1    g257(.A1(new_n678), .A2(KEYINPUT90), .ZN(new_n683));
  OR2_X1    g258(.A1(new_n679), .A2(new_n680), .ZN(new_n684));
  NAND2_X1  g259(.A1(new_n679), .A2(new_n680), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n684), .B1(new_n678), .B2(new_n685), .ZN(new_n686));
  OR2_X1    g261(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n683), .A2(new_n686), .ZN(new_n688));
  NAND3_X1  g263(.A1(new_n682), .A2(new_n687), .A3(new_n688), .ZN(new_n689));
  XNOR2_X1  g264(.A(new_n689), .B(KEYINPUT21), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(KEYINPUT22), .ZN(new_n691));
  XOR2_X1   g266(.A(G1991), .B(G1996), .Z(new_n692));
  XNOR2_X1  g267(.A(new_n692), .B(KEYINPUT91), .ZN(new_n693));
  XNOR2_X1  g268(.A(new_n691), .B(new_n693), .ZN(new_n694));
  XNOR2_X1  g269(.A(G1981), .B(G1986), .ZN(new_n695));
  XNOR2_X1  g270(.A(new_n694), .B(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n696), .ZN(G229));
  NAND2_X1  g272(.A1(new_n483), .A2(G128), .ZN(new_n698));
  OR2_X1    g273(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n699));
  NAND2_X1  g274(.A1(new_n698), .A2(KEYINPUT98), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n631), .A2(G140), .ZN(new_n701));
  OR2_X1    g276(.A1(G104), .A2(G2105), .ZN(new_n702));
  OAI211_X1 g277(.A(new_n702), .B(G2104), .C1(G116), .C2(new_n482), .ZN(new_n703));
  NAND4_X1  g278(.A1(new_n699), .A2(new_n700), .A3(new_n701), .A4(new_n703), .ZN(new_n704));
  NAND2_X1  g279(.A1(new_n704), .A2(G29), .ZN(new_n705));
  XNOR2_X1  g280(.A(new_n705), .B(KEYINPUT99), .ZN(new_n706));
  INV_X1    g281(.A(G29), .ZN(new_n707));
  NAND2_X1  g282(.A1(new_n707), .A2(G26), .ZN(new_n708));
  XNOR2_X1  g283(.A(new_n708), .B(KEYINPUT28), .ZN(new_n709));
  NAND2_X1  g284(.A1(new_n706), .A2(new_n709), .ZN(new_n710));
  INV_X1    g285(.A(G2067), .ZN(new_n711));
  XNOR2_X1  g286(.A(new_n710), .B(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G16), .ZN(new_n713));
  NAND2_X1  g288(.A1(new_n713), .A2(G4), .ZN(new_n714));
  OAI21_X1  g289(.A(new_n714), .B1(new_n613), .B2(new_n713), .ZN(new_n715));
  INV_X1    g290(.A(G1348), .ZN(new_n716));
  XNOR2_X1  g291(.A(new_n715), .B(new_n716), .ZN(new_n717));
  NAND2_X1  g292(.A1(new_n713), .A2(G19), .ZN(new_n718));
  OAI21_X1  g293(.A(new_n718), .B1(new_n559), .B2(new_n713), .ZN(new_n719));
  XOR2_X1   g294(.A(KEYINPUT97), .B(G1341), .Z(new_n720));
  XNOR2_X1  g295(.A(new_n719), .B(new_n720), .ZN(new_n721));
  NAND3_X1  g296(.A1(new_n712), .A2(new_n717), .A3(new_n721), .ZN(new_n722));
  XNOR2_X1  g297(.A(new_n722), .B(KEYINPUT100), .ZN(new_n723));
  NOR2_X1   g298(.A1(G16), .A2(G22), .ZN(new_n724));
  AOI21_X1  g299(.A(new_n724), .B1(G166), .B2(G16), .ZN(new_n725));
  XNOR2_X1  g300(.A(KEYINPUT95), .B(G1971), .ZN(new_n726));
  XNOR2_X1  g301(.A(new_n725), .B(new_n726), .ZN(new_n727));
  NOR2_X1   g302(.A1(G16), .A2(G23), .ZN(new_n728));
  AOI21_X1  g303(.A(new_n728), .B1(new_n581), .B2(G16), .ZN(new_n729));
  XOR2_X1   g304(.A(KEYINPUT33), .B(G1976), .Z(new_n730));
  OR2_X1    g305(.A1(new_n729), .A2(new_n730), .ZN(new_n731));
  NAND2_X1  g306(.A1(new_n713), .A2(G6), .ZN(new_n732));
  OAI21_X1  g307(.A(new_n732), .B1(new_n592), .B2(new_n713), .ZN(new_n733));
  XOR2_X1   g308(.A(KEYINPUT94), .B(KEYINPUT32), .Z(new_n734));
  XOR2_X1   g309(.A(new_n734), .B(G1981), .Z(new_n735));
  XNOR2_X1  g310(.A(new_n733), .B(new_n735), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n729), .A2(new_n730), .ZN(new_n737));
  NAND4_X1  g312(.A1(new_n727), .A2(new_n731), .A3(new_n736), .A4(new_n737), .ZN(new_n738));
  XOR2_X1   g313(.A(new_n738), .B(KEYINPUT34), .Z(new_n739));
  NAND2_X1  g314(.A1(new_n483), .A2(G119), .ZN(new_n740));
  NAND2_X1  g315(.A1(new_n631), .A2(G131), .ZN(new_n741));
  NOR2_X1   g316(.A1(new_n482), .A2(G107), .ZN(new_n742));
  OAI21_X1  g317(.A(G2104), .B1(G95), .B2(G2105), .ZN(new_n743));
  OAI211_X1 g318(.A(new_n740), .B(new_n741), .C1(new_n742), .C2(new_n743), .ZN(new_n744));
  MUX2_X1   g319(.A(G25), .B(new_n744), .S(G29), .Z(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT35), .B(G1991), .ZN(new_n746));
  XNOR2_X1  g321(.A(new_n745), .B(new_n746), .ZN(new_n747));
  XNOR2_X1  g322(.A(KEYINPUT92), .B(KEYINPUT93), .ZN(new_n748));
  XNOR2_X1  g323(.A(new_n747), .B(new_n748), .ZN(new_n749));
  MUX2_X1   g324(.A(G24), .B(G290), .S(G16), .Z(new_n750));
  XOR2_X1   g325(.A(new_n750), .B(G1986), .Z(new_n751));
  NAND3_X1  g326(.A1(new_n739), .A2(new_n749), .A3(new_n751), .ZN(new_n752));
  XOR2_X1   g327(.A(KEYINPUT96), .B(KEYINPUT36), .Z(new_n753));
  XNOR2_X1  g328(.A(new_n752), .B(new_n753), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n483), .A2(G129), .ZN(new_n755));
  NAND2_X1  g330(.A1(new_n631), .A2(G141), .ZN(new_n756));
  NAND3_X1  g331(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n757));
  INV_X1    g332(.A(KEYINPUT26), .ZN(new_n758));
  OR2_X1    g333(.A1(new_n757), .A2(new_n758), .ZN(new_n759));
  NAND2_X1  g334(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  AOI22_X1  g335(.A1(new_n759), .A2(new_n760), .B1(G105), .B2(new_n495), .ZN(new_n761));
  NAND3_X1  g336(.A1(new_n755), .A2(new_n756), .A3(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n707), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT103), .ZN(new_n764));
  OAI21_X1  g339(.A(new_n764), .B1(G29), .B2(G32), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n765), .B(KEYINPUT27), .ZN(new_n766));
  INV_X1    g341(.A(G1996), .ZN(new_n767));
  XNOR2_X1  g342(.A(new_n766), .B(new_n767), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n707), .A2(G35), .ZN(new_n769));
  OAI21_X1  g344(.A(new_n769), .B1(G162), .B2(new_n707), .ZN(new_n770));
  XNOR2_X1  g345(.A(new_n770), .B(KEYINPUT29), .ZN(new_n771));
  XNOR2_X1  g346(.A(new_n771), .B(G2090), .ZN(new_n772));
  OAI21_X1  g347(.A(KEYINPUT23), .B1(new_n617), .B2(new_n713), .ZN(new_n773));
  NAND2_X1  g348(.A1(new_n713), .A2(G20), .ZN(new_n774));
  MUX2_X1   g349(.A(KEYINPUT23), .B(new_n773), .S(new_n774), .Z(new_n775));
  XOR2_X1   g350(.A(new_n775), .B(G1956), .Z(new_n776));
  INV_X1    g351(.A(G2084), .ZN(new_n777));
  XNOR2_X1  g352(.A(KEYINPUT102), .B(KEYINPUT24), .ZN(new_n778));
  AND2_X1   g353(.A1(new_n778), .A2(G34), .ZN(new_n779));
  OAI21_X1  g354(.A(new_n707), .B1(new_n778), .B2(G34), .ZN(new_n780));
  OAI22_X1  g355(.A1(G160), .A2(new_n707), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  INV_X1    g356(.A(new_n781), .ZN(new_n782));
  OAI21_X1  g357(.A(new_n776), .B1(new_n777), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g358(.A1(new_n707), .A2(G33), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n631), .A2(G139), .ZN(new_n785));
  XOR2_X1   g360(.A(new_n785), .B(KEYINPUT101), .Z(new_n786));
  AND2_X1   g361(.A1(new_n495), .A2(G103), .ZN(new_n787));
  OR2_X1    g362(.A1(new_n787), .A2(KEYINPUT25), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n787), .A2(KEYINPUT25), .ZN(new_n789));
  NAND2_X1  g364(.A1(G115), .A2(G2104), .ZN(new_n790));
  INV_X1    g365(.A(G127), .ZN(new_n791));
  OAI21_X1  g366(.A(new_n790), .B1(new_n477), .B2(new_n791), .ZN(new_n792));
  AOI22_X1  g367(.A1(new_n788), .A2(new_n789), .B1(G2105), .B2(new_n792), .ZN(new_n793));
  AND2_X1   g368(.A1(new_n786), .A2(new_n793), .ZN(new_n794));
  OAI21_X1  g369(.A(new_n784), .B1(new_n794), .B2(new_n707), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n707), .A2(G27), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n796), .B1(G164), .B2(new_n707), .ZN(new_n797));
  AOI22_X1  g372(.A1(new_n795), .A2(G2072), .B1(G2078), .B2(new_n797), .ZN(new_n798));
  OR2_X1    g373(.A1(new_n797), .A2(G2078), .ZN(new_n799));
  OAI211_X1 g374(.A(new_n798), .B(new_n799), .C1(G2072), .C2(new_n795), .ZN(new_n800));
  XOR2_X1   g375(.A(KEYINPUT31), .B(G11), .Z(new_n801));
  INV_X1    g376(.A(G28), .ZN(new_n802));
  OR2_X1    g377(.A1(new_n802), .A2(KEYINPUT30), .ZN(new_n803));
  AOI21_X1  g378(.A(G29), .B1(new_n802), .B2(KEYINPUT30), .ZN(new_n804));
  AOI21_X1  g379(.A(new_n801), .B1(new_n803), .B2(new_n804), .ZN(new_n805));
  NOR2_X1   g380(.A1(G16), .A2(G21), .ZN(new_n806));
  AOI21_X1  g381(.A(new_n806), .B1(G168), .B2(G16), .ZN(new_n807));
  OAI221_X1 g382(.A(new_n805), .B1(new_n707), .B2(new_n635), .C1(new_n807), .C2(G1966), .ZN(new_n808));
  AOI21_X1  g383(.A(new_n808), .B1(G1966), .B2(new_n807), .ZN(new_n809));
  NOR2_X1   g384(.A1(G5), .A2(G16), .ZN(new_n810));
  AOI21_X1  g385(.A(new_n810), .B1(G171), .B2(G16), .ZN(new_n811));
  INV_X1    g386(.A(G1961), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  OAI211_X1 g388(.A(new_n809), .B(new_n813), .C1(G2084), .C2(new_n781), .ZN(new_n814));
  NOR4_X1   g389(.A1(new_n772), .A2(new_n783), .A3(new_n800), .A4(new_n814), .ZN(new_n815));
  NAND4_X1  g390(.A1(new_n723), .A2(new_n754), .A3(new_n768), .A4(new_n815), .ZN(G150));
  INV_X1    g391(.A(G150), .ZN(G311));
  NAND2_X1  g392(.A1(new_n613), .A2(G559), .ZN(new_n818));
  AOI22_X1  g393(.A1(new_n517), .A2(G67), .B1(G80), .B2(G543), .ZN(new_n819));
  OR2_X1    g394(.A1(new_n819), .A2(new_n525), .ZN(new_n820));
  NAND3_X1  g395(.A1(new_n517), .A2(new_n518), .A3(G93), .ZN(new_n821));
  INV_X1    g396(.A(KEYINPUT104), .ZN(new_n822));
  NAND4_X1  g397(.A1(new_n584), .A2(new_n586), .A3(G55), .A4(G543), .ZN(new_n823));
  AND3_X1   g398(.A1(new_n821), .A2(new_n822), .A3(new_n823), .ZN(new_n824));
  AOI21_X1  g399(.A(new_n822), .B1(new_n821), .B2(new_n823), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n820), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  INV_X1    g401(.A(KEYINPUT105), .ZN(new_n827));
  NAND2_X1  g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  INV_X1    g403(.A(new_n559), .ZN(new_n829));
  OAI211_X1 g404(.A(new_n820), .B(KEYINPUT105), .C1(new_n824), .C2(new_n825), .ZN(new_n830));
  NAND3_X1  g405(.A1(new_n828), .A2(new_n829), .A3(new_n830), .ZN(new_n831));
  INV_X1    g406(.A(new_n826), .ZN(new_n832));
  NAND3_X1  g407(.A1(new_n832), .A2(KEYINPUT105), .A3(new_n559), .ZN(new_n833));
  NAND2_X1  g408(.A1(new_n831), .A2(new_n833), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n818), .B(new_n834), .ZN(new_n835));
  INV_X1    g410(.A(new_n835), .ZN(new_n836));
  XNOR2_X1  g411(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n837));
  AOI21_X1  g412(.A(G860), .B1(new_n836), .B2(new_n837), .ZN(new_n838));
  OAI21_X1  g413(.A(new_n838), .B1(new_n837), .B2(new_n836), .ZN(new_n839));
  NAND2_X1  g414(.A1(new_n826), .A2(G860), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT106), .B(KEYINPUT37), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  NAND2_X1  g417(.A1(new_n839), .A2(new_n842), .ZN(G145));
  XNOR2_X1  g418(.A(new_n704), .B(new_n493), .ZN(new_n844));
  XNOR2_X1  g419(.A(G160), .B(new_n635), .ZN(new_n845));
  XNOR2_X1  g420(.A(new_n844), .B(new_n845), .ZN(new_n846));
  NAND2_X1  g421(.A1(new_n509), .A2(new_n514), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n744), .B(new_n847), .ZN(new_n848));
  XNOR2_X1  g423(.A(new_n762), .B(new_n627), .ZN(new_n849));
  XNOR2_X1  g424(.A(new_n848), .B(new_n849), .ZN(new_n850));
  OR2_X1    g425(.A1(new_n846), .A2(new_n850), .ZN(new_n851));
  NAND2_X1  g426(.A1(new_n846), .A2(new_n850), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g428(.A1(new_n483), .A2(G130), .ZN(new_n854));
  NAND2_X1  g429(.A1(new_n631), .A2(G142), .ZN(new_n855));
  NOR2_X1   g430(.A1(new_n482), .A2(G118), .ZN(new_n856));
  OAI21_X1  g431(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n857));
  OAI211_X1 g432(.A(new_n854), .B(new_n855), .C1(new_n856), .C2(new_n857), .ZN(new_n858));
  XOR2_X1   g433(.A(new_n794), .B(new_n858), .Z(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND2_X1  g435(.A1(new_n853), .A2(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(G37), .ZN(new_n862));
  NAND3_X1  g437(.A1(new_n851), .A2(new_n859), .A3(new_n852), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n861), .A2(new_n862), .A3(new_n863), .ZN(new_n864));
  XNOR2_X1  g439(.A(new_n864), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g440(.A(new_n592), .B(G303), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(G290), .A2(new_n581), .ZN(new_n868));
  NAND3_X1  g443(.A1(G288), .A2(new_n601), .A3(new_n600), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n867), .A2(new_n868), .A3(new_n869), .ZN(new_n870));
  NAND2_X1  g445(.A1(new_n868), .A2(new_n869), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n866), .ZN(new_n872));
  AND2_X1   g447(.A1(new_n870), .A2(new_n872), .ZN(new_n873));
  NAND2_X1  g448(.A1(new_n873), .A2(KEYINPUT107), .ZN(new_n874));
  XOR2_X1   g449(.A(new_n874), .B(KEYINPUT42), .Z(new_n875));
  XNOR2_X1  g450(.A(new_n622), .B(new_n834), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT41), .ZN(new_n877));
  OAI211_X1 g452(.A(G299), .B(new_n607), .C1(new_n610), .C2(new_n611), .ZN(new_n878));
  INV_X1    g453(.A(new_n878), .ZN(new_n879));
  XNOR2_X1  g454(.A(new_n608), .B(new_n609), .ZN(new_n880));
  AOI21_X1  g455(.A(G299), .B1(new_n880), .B2(new_n607), .ZN(new_n881));
  OAI21_X1  g456(.A(new_n877), .B1(new_n879), .B2(new_n881), .ZN(new_n882));
  NAND2_X1  g457(.A1(new_n612), .A2(new_n617), .ZN(new_n883));
  NAND3_X1  g458(.A1(new_n883), .A2(KEYINPUT41), .A3(new_n878), .ZN(new_n884));
  AOI21_X1  g459(.A(new_n876), .B1(new_n882), .B2(new_n884), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n879), .A2(new_n881), .ZN(new_n886));
  INV_X1    g461(.A(new_n886), .ZN(new_n887));
  AOI21_X1  g462(.A(new_n885), .B1(new_n887), .B2(new_n876), .ZN(new_n888));
  OR2_X1    g463(.A1(new_n875), .A2(new_n888), .ZN(new_n889));
  NAND2_X1  g464(.A1(new_n875), .A2(new_n888), .ZN(new_n890));
  NAND3_X1  g465(.A1(new_n889), .A2(G868), .A3(new_n890), .ZN(new_n891));
  NOR2_X1   g466(.A1(new_n832), .A2(G868), .ZN(new_n892));
  OAI21_X1  g467(.A(new_n891), .B1(KEYINPUT108), .B2(new_n892), .ZN(new_n893));
  OAI21_X1  g468(.A(new_n893), .B1(KEYINPUT108), .B2(new_n891), .ZN(G295));
  OAI21_X1  g469(.A(new_n893), .B1(KEYINPUT108), .B2(new_n891), .ZN(G331));
  AND3_X1   g470(.A1(new_n831), .A2(G286), .A3(new_n833), .ZN(new_n896));
  AOI21_X1  g471(.A(G286), .B1(new_n831), .B2(new_n833), .ZN(new_n897));
  OAI21_X1  g472(.A(G301), .B1(new_n896), .B2(new_n897), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n834), .A2(G168), .ZN(new_n899));
  NAND3_X1  g474(.A1(new_n831), .A2(G286), .A3(new_n833), .ZN(new_n900));
  NAND3_X1  g475(.A1(new_n899), .A2(G171), .A3(new_n900), .ZN(new_n901));
  AOI21_X1  g476(.A(new_n886), .B1(new_n898), .B2(new_n901), .ZN(new_n902));
  INV_X1    g477(.A(KEYINPUT109), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n870), .A2(new_n903), .A3(new_n872), .ZN(new_n904));
  NOR2_X1   g479(.A1(new_n902), .A2(new_n904), .ZN(new_n905));
  INV_X1    g480(.A(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n882), .A2(new_n884), .ZN(new_n907));
  AND3_X1   g482(.A1(new_n898), .A2(new_n901), .A3(new_n907), .ZN(new_n908));
  NOR3_X1   g483(.A1(new_n908), .A2(new_n902), .A3(new_n873), .ZN(new_n909));
  NAND2_X1  g484(.A1(new_n870), .A2(new_n872), .ZN(new_n910));
  NOR3_X1   g485(.A1(new_n896), .A2(new_n897), .A3(G301), .ZN(new_n911));
  AOI21_X1  g486(.A(G171), .B1(new_n899), .B2(new_n900), .ZN(new_n912));
  OAI21_X1  g487(.A(new_n887), .B1(new_n911), .B2(new_n912), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n901), .A2(new_n898), .A3(new_n907), .ZN(new_n914));
  AOI21_X1  g489(.A(new_n910), .B1(new_n913), .B2(new_n914), .ZN(new_n915));
  OAI21_X1  g490(.A(new_n906), .B1(new_n909), .B2(new_n915), .ZN(new_n916));
  OAI21_X1  g491(.A(new_n873), .B1(new_n908), .B2(new_n902), .ZN(new_n917));
  NAND3_X1  g492(.A1(new_n913), .A2(new_n910), .A3(new_n914), .ZN(new_n918));
  NAND3_X1  g493(.A1(new_n917), .A2(new_n918), .A3(new_n905), .ZN(new_n919));
  NAND4_X1  g494(.A1(new_n916), .A2(KEYINPUT43), .A3(new_n862), .A4(new_n919), .ZN(new_n920));
  NAND3_X1  g495(.A1(new_n917), .A2(new_n862), .A3(new_n918), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT43), .ZN(new_n922));
  NAND2_X1  g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  NAND2_X1  g498(.A1(new_n920), .A2(new_n923), .ZN(new_n924));
  NAND2_X1  g499(.A1(new_n924), .A2(KEYINPUT44), .ZN(new_n925));
  INV_X1    g500(.A(KEYINPUT44), .ZN(new_n926));
  AOI21_X1  g501(.A(new_n905), .B1(new_n917), .B2(new_n918), .ZN(new_n927));
  NOR4_X1   g502(.A1(new_n908), .A2(new_n902), .A3(KEYINPUT109), .A4(new_n910), .ZN(new_n928));
  NOR4_X1   g503(.A1(new_n927), .A2(new_n928), .A3(KEYINPUT43), .A4(G37), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n921), .A2(KEYINPUT43), .ZN(new_n930));
  INV_X1    g505(.A(new_n930), .ZN(new_n931));
  OAI21_X1  g506(.A(new_n926), .B1(new_n929), .B2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(KEYINPUT110), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n925), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  AOI21_X1  g509(.A(new_n926), .B1(new_n920), .B2(new_n923), .ZN(new_n935));
  NAND4_X1  g510(.A1(new_n916), .A2(new_n922), .A3(new_n862), .A4(new_n919), .ZN(new_n936));
  AOI21_X1  g511(.A(KEYINPUT44), .B1(new_n936), .B2(new_n930), .ZN(new_n937));
  OAI21_X1  g512(.A(KEYINPUT110), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n934), .A2(new_n938), .ZN(G397));
  XOR2_X1   g514(.A(KEYINPUT111), .B(G1384), .Z(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n847), .A2(new_n941), .ZN(new_n942));
  AOI21_X1  g517(.A(KEYINPUT45), .B1(new_n942), .B2(KEYINPUT112), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT112), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n847), .A2(new_n944), .A3(new_n941), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n943), .A2(new_n945), .ZN(new_n946));
  INV_X1    g521(.A(G40), .ZN(new_n947));
  AOI211_X1 g522(.A(new_n947), .B(new_n465), .C1(new_n474), .C2(G2105), .ZN(new_n948));
  INV_X1    g523(.A(new_n948), .ZN(new_n949));
  NOR2_X1   g524(.A1(new_n946), .A2(new_n949), .ZN(new_n950));
  XNOR2_X1  g525(.A(new_n950), .B(KEYINPUT113), .ZN(new_n951));
  NAND3_X1  g526(.A1(new_n951), .A2(G1996), .A3(new_n762), .ZN(new_n952));
  NAND2_X1  g527(.A1(new_n950), .A2(new_n767), .ZN(new_n953));
  OR2_X1    g528(.A1(new_n953), .A2(new_n762), .ZN(new_n954));
  XNOR2_X1  g529(.A(new_n704), .B(G2067), .ZN(new_n955));
  NAND2_X1  g530(.A1(new_n951), .A2(new_n955), .ZN(new_n956));
  AND3_X1   g531(.A1(new_n952), .A2(new_n954), .A3(new_n956), .ZN(new_n957));
  XOR2_X1   g532(.A(new_n744), .B(new_n746), .Z(new_n958));
  INV_X1    g533(.A(new_n951), .ZN(new_n959));
  OAI21_X1  g534(.A(new_n957), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  XNOR2_X1  g535(.A(G290), .B(G1986), .ZN(new_n961));
  AOI21_X1  g536(.A(new_n960), .B1(new_n950), .B2(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT50), .ZN(new_n963));
  INV_X1    g538(.A(G1384), .ZN(new_n964));
  AOI21_X1  g539(.A(KEYINPUT114), .B1(new_n847), .B2(new_n964), .ZN(new_n965));
  INV_X1    g540(.A(KEYINPUT114), .ZN(new_n966));
  AOI211_X1 g541(.A(new_n966), .B(G1384), .C1(new_n509), .C2(new_n514), .ZN(new_n967));
  OAI21_X1  g542(.A(new_n963), .B1(new_n965), .B2(new_n967), .ZN(new_n968));
  NAND3_X1  g543(.A1(new_n505), .A2(new_n964), .A3(new_n515), .ZN(new_n969));
  NAND2_X1  g544(.A1(new_n969), .A2(KEYINPUT50), .ZN(new_n970));
  NAND3_X1  g545(.A1(new_n968), .A2(new_n970), .A3(new_n948), .ZN(new_n971));
  NAND2_X1  g546(.A1(new_n971), .A2(new_n812), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n972), .A2(KEYINPUT126), .ZN(new_n973));
  INV_X1    g548(.A(G2078), .ZN(new_n974));
  NAND3_X1  g549(.A1(new_n847), .A2(KEYINPUT45), .A3(new_n941), .ZN(new_n975));
  AND3_X1   g550(.A1(new_n948), .A2(new_n974), .A3(new_n975), .ZN(new_n976));
  INV_X1    g551(.A(KEYINPUT45), .ZN(new_n977));
  NAND2_X1  g552(.A1(new_n969), .A2(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(new_n976), .A2(new_n978), .ZN(new_n979));
  INV_X1    g554(.A(KEYINPUT53), .ZN(new_n980));
  AOI21_X1  g555(.A(new_n980), .B1(new_n943), .B2(new_n945), .ZN(new_n981));
  AOI22_X1  g556(.A1(new_n979), .A2(new_n980), .B1(new_n981), .B2(new_n976), .ZN(new_n982));
  INV_X1    g557(.A(KEYINPUT126), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n971), .A2(new_n983), .A3(new_n812), .ZN(new_n984));
  NAND4_X1  g559(.A1(new_n973), .A2(G301), .A3(new_n982), .A4(new_n984), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n985), .A2(KEYINPUT127), .ZN(new_n986));
  NAND3_X1  g561(.A1(new_n946), .A2(new_n976), .A3(KEYINPUT53), .ZN(new_n987));
  NAND3_X1  g562(.A1(new_n948), .A2(new_n975), .A3(new_n974), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n988), .B1(new_n977), .B2(new_n969), .ZN(new_n989));
  OAI21_X1  g564(.A(new_n987), .B1(new_n989), .B2(KEYINPUT53), .ZN(new_n990));
  AOI21_X1  g565(.A(new_n983), .B1(new_n971), .B2(new_n812), .ZN(new_n991));
  NOR2_X1   g566(.A1(new_n990), .A2(new_n991), .ZN(new_n992));
  INV_X1    g567(.A(KEYINPUT127), .ZN(new_n993));
  NAND4_X1  g568(.A1(new_n992), .A2(new_n993), .A3(G301), .A4(new_n984), .ZN(new_n994));
  OAI21_X1  g569(.A(new_n964), .B1(new_n498), .B2(new_n504), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n995), .A2(new_n966), .ZN(new_n996));
  NAND3_X1  g571(.A1(new_n847), .A2(KEYINPUT114), .A3(new_n964), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n996), .A2(new_n997), .ZN(new_n998));
  AOI21_X1  g573(.A(new_n949), .B1(new_n998), .B2(new_n963), .ZN(new_n999));
  AOI21_X1  g574(.A(G1961), .B1(new_n999), .B2(new_n970), .ZN(new_n1000));
  NAND3_X1  g575(.A1(new_n996), .A2(new_n977), .A3(new_n997), .ZN(new_n1001));
  NAND4_X1  g576(.A1(new_n505), .A2(KEYINPUT45), .A3(new_n964), .A4(new_n515), .ZN(new_n1002));
  NOR2_X1   g577(.A1(new_n980), .A2(G2078), .ZN(new_n1003));
  NAND4_X1  g578(.A1(new_n1001), .A2(new_n948), .A3(new_n1002), .A4(new_n1003), .ZN(new_n1004));
  INV_X1    g579(.A(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(KEYINPUT125), .B1(new_n1000), .B2(new_n1005), .ZN(new_n1006));
  INV_X1    g581(.A(KEYINPUT125), .ZN(new_n1007));
  NAND3_X1  g582(.A1(new_n972), .A2(new_n1007), .A3(new_n1004), .ZN(new_n1008));
  AOI22_X1  g583(.A1(new_n1006), .A2(new_n1008), .B1(new_n980), .B2(new_n979), .ZN(new_n1009));
  OAI211_X1 g584(.A(new_n986), .B(new_n994), .C1(new_n1009), .C2(G301), .ZN(new_n1010));
  INV_X1    g585(.A(KEYINPUT54), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1010), .A2(new_n1011), .ZN(new_n1012));
  AND2_X1   g587(.A1(new_n948), .A2(new_n975), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1013), .A2(new_n978), .ZN(new_n1014));
  INV_X1    g589(.A(G1971), .ZN(new_n1015));
  NAND2_X1  g590(.A1(new_n1014), .A2(new_n1015), .ZN(new_n1016));
  OAI21_X1  g591(.A(new_n1016), .B1(G2090), .B2(new_n971), .ZN(new_n1017));
  NAND2_X1  g592(.A1(G303), .A2(G8), .ZN(new_n1018));
  XNOR2_X1  g593(.A(new_n1018), .B(KEYINPUT55), .ZN(new_n1019));
  INV_X1    g594(.A(new_n1019), .ZN(new_n1020));
  NAND3_X1  g595(.A1(new_n1017), .A2(G8), .A3(new_n1020), .ZN(new_n1021));
  INV_X1    g596(.A(KEYINPUT120), .ZN(new_n1022));
  OAI21_X1  g597(.A(new_n948), .B1(new_n965), .B2(new_n967), .ZN(new_n1023));
  AND2_X1   g598(.A1(new_n537), .A2(G86), .ZN(new_n1024));
  OAI21_X1  g599(.A(G1981), .B1(new_n1024), .B2(new_n591), .ZN(new_n1025));
  OAI21_X1  g600(.A(G86), .B1(new_n572), .B2(new_n573), .ZN(new_n1026));
  NAND2_X1  g601(.A1(G73), .A2(G543), .ZN(new_n1027));
  INV_X1    g602(.A(G61), .ZN(new_n1028));
  OAI21_X1  g603(.A(new_n1027), .B1(new_n545), .B2(new_n1028), .ZN(new_n1029));
  AOI22_X1  g604(.A1(new_n1029), .A2(G651), .B1(new_n588), .B2(new_n587), .ZN(new_n1030));
  XNOR2_X1  g605(.A(KEYINPUT117), .B(G1981), .ZN(new_n1031));
  NAND4_X1  g606(.A1(new_n1026), .A2(new_n1030), .A3(new_n583), .A4(new_n1031), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n1025), .A2(new_n1032), .A3(KEYINPUT49), .ZN(new_n1033));
  AND3_X1   g608(.A1(new_n1023), .A2(G8), .A3(new_n1033), .ZN(new_n1034));
  INV_X1    g609(.A(KEYINPUT118), .ZN(new_n1035));
  NAND2_X1  g610(.A1(new_n1025), .A2(new_n1032), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT49), .ZN(new_n1037));
  AOI21_X1  g612(.A(new_n1035), .B1(new_n1036), .B2(new_n1037), .ZN(new_n1038));
  AOI211_X1 g613(.A(KEYINPUT118), .B(KEYINPUT49), .C1(new_n1025), .C2(new_n1032), .ZN(new_n1039));
  NOR2_X1   g614(.A1(new_n1038), .A2(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G8), .ZN(new_n1041));
  AOI21_X1  g616(.A(new_n1041), .B1(new_n998), .B2(new_n948), .ZN(new_n1042));
  INV_X1    g617(.A(KEYINPUT116), .ZN(new_n1043));
  AOI21_X1  g618(.A(new_n1043), .B1(new_n581), .B2(G1976), .ZN(new_n1044));
  XOR2_X1   g619(.A(KEYINPUT115), .B(G1976), .Z(new_n1045));
  NOR2_X1   g620(.A1(new_n581), .A2(new_n1045), .ZN(new_n1046));
  OAI211_X1 g621(.A(new_n1042), .B(new_n1044), .C1(KEYINPUT52), .C2(new_n1046), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1023), .A2(G8), .A3(new_n1046), .ZN(new_n1048));
  NAND3_X1  g623(.A1(new_n1023), .A2(G8), .A3(new_n1044), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT52), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1048), .A2(new_n1049), .A3(new_n1050), .ZN(new_n1051));
  AOI221_X4 g626(.A(new_n1022), .B1(new_n1034), .B2(new_n1040), .C1(new_n1047), .C2(new_n1051), .ZN(new_n1052));
  NAND2_X1  g627(.A1(new_n1047), .A2(new_n1051), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1040), .A2(new_n1034), .ZN(new_n1054));
  AOI21_X1  g629(.A(KEYINPUT120), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  OAI21_X1  g630(.A(new_n1021), .B1(new_n1052), .B2(new_n1055), .ZN(new_n1056));
  INV_X1    g631(.A(KEYINPUT119), .ZN(new_n1057));
  NAND3_X1  g632(.A1(new_n996), .A2(KEYINPUT50), .A3(new_n997), .ZN(new_n1058));
  INV_X1    g633(.A(G2090), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n505), .A2(new_n963), .A3(new_n964), .A4(new_n515), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1058), .A2(new_n1059), .A3(new_n948), .A4(new_n1060), .ZN(new_n1061));
  NAND2_X1  g636(.A1(new_n1016), .A2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(new_n1062), .A2(G8), .ZN(new_n1063));
  AOI21_X1  g638(.A(new_n1057), .B1(new_n1063), .B2(new_n1019), .ZN(new_n1064));
  AOI211_X1 g639(.A(KEYINPUT119), .B(new_n1020), .C1(new_n1062), .C2(G8), .ZN(new_n1065));
  NOR2_X1   g640(.A1(new_n1064), .A2(new_n1065), .ZN(new_n1066));
  NOR2_X1   g641(.A1(new_n1056), .A2(new_n1066), .ZN(new_n1067));
  INV_X1    g642(.A(KEYINPUT124), .ZN(new_n1068));
  NAND3_X1  g643(.A1(new_n1001), .A2(new_n948), .A3(new_n1002), .ZN(new_n1069));
  INV_X1    g644(.A(G1966), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1069), .A2(new_n1070), .ZN(new_n1071));
  NAND4_X1  g646(.A1(new_n968), .A2(new_n970), .A3(new_n777), .A4(new_n948), .ZN(new_n1072));
  NAND3_X1  g647(.A1(new_n1071), .A2(G168), .A3(new_n1072), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1073), .A2(G8), .ZN(new_n1074));
  INV_X1    g649(.A(KEYINPUT51), .ZN(new_n1075));
  OAI21_X1  g650(.A(new_n1068), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n1074), .A2(new_n1075), .ZN(new_n1077));
  NAND4_X1  g652(.A1(new_n1073), .A2(KEYINPUT124), .A3(KEYINPUT51), .A4(G8), .ZN(new_n1078));
  NAND3_X1  g653(.A1(new_n1076), .A2(new_n1077), .A3(new_n1078), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1071), .A2(new_n1072), .ZN(new_n1080));
  NAND3_X1  g655(.A1(new_n1080), .A2(G8), .A3(G286), .ZN(new_n1081));
  NAND2_X1  g656(.A1(new_n1079), .A2(new_n1081), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n992), .A2(new_n984), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1011), .B1(new_n1083), .B2(G171), .ZN(new_n1084));
  NOR3_X1   g659(.A1(new_n1000), .A2(new_n1005), .A3(KEYINPUT125), .ZN(new_n1085));
  AOI21_X1  g660(.A(new_n1007), .B1(new_n972), .B2(new_n1004), .ZN(new_n1086));
  OAI22_X1  g661(.A1(new_n1085), .A2(new_n1086), .B1(KEYINPUT53), .B2(new_n989), .ZN(new_n1087));
  OAI21_X1  g662(.A(new_n1084), .B1(G171), .B2(new_n1087), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1012), .A2(new_n1067), .A3(new_n1082), .A4(new_n1088), .ZN(new_n1089));
  AOI21_X1  g664(.A(G1348), .B1(new_n999), .B2(new_n970), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT122), .ZN(new_n1091));
  NOR2_X1   g666(.A1(new_n1023), .A2(G2067), .ZN(new_n1092));
  NOR3_X1   g667(.A1(new_n1090), .A2(new_n1091), .A3(new_n1092), .ZN(new_n1093));
  NAND2_X1  g668(.A1(new_n971), .A2(new_n716), .ZN(new_n1094));
  INV_X1    g669(.A(new_n1092), .ZN(new_n1095));
  AOI21_X1  g670(.A(KEYINPUT122), .B1(new_n1094), .B2(new_n1095), .ZN(new_n1096));
  OAI211_X1 g671(.A(KEYINPUT60), .B(new_n612), .C1(new_n1093), .C2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1097), .A2(KEYINPUT123), .ZN(new_n1098));
  OAI21_X1  g673(.A(KEYINPUT60), .B1(new_n1093), .B2(new_n1096), .ZN(new_n1099));
  NAND2_X1  g674(.A1(new_n1099), .A2(new_n613), .ZN(new_n1100));
  OAI21_X1  g675(.A(new_n1091), .B1(new_n1090), .B2(new_n1092), .ZN(new_n1101));
  NAND3_X1  g676(.A1(new_n1094), .A2(KEYINPUT122), .A3(new_n1095), .ZN(new_n1102));
  NAND2_X1  g677(.A1(new_n1101), .A2(new_n1102), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT123), .ZN(new_n1104));
  NAND4_X1  g679(.A1(new_n1103), .A2(new_n1104), .A3(KEYINPUT60), .A4(new_n612), .ZN(new_n1105));
  NAND3_X1  g680(.A1(new_n1098), .A2(new_n1100), .A3(new_n1105), .ZN(new_n1106));
  OR2_X1    g681(.A1(new_n1103), .A2(KEYINPUT60), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1106), .A2(new_n1107), .ZN(new_n1108));
  NAND3_X1  g683(.A1(new_n1058), .A2(new_n948), .A3(new_n1060), .ZN(new_n1109));
  XOR2_X1   g684(.A(KEYINPUT121), .B(G1956), .Z(new_n1110));
  AND2_X1   g685(.A1(new_n1013), .A2(new_n978), .ZN(new_n1111));
  XNOR2_X1  g686(.A(KEYINPUT56), .B(G2072), .ZN(new_n1112));
  AOI22_X1  g687(.A1(new_n1109), .A2(new_n1110), .B1(new_n1111), .B2(new_n1112), .ZN(new_n1113));
  XNOR2_X1  g688(.A(G299), .B(KEYINPUT57), .ZN(new_n1114));
  INV_X1    g689(.A(new_n1114), .ZN(new_n1115));
  NOR2_X1   g690(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1116));
  INV_X1    g691(.A(new_n1116), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1113), .A2(new_n1115), .ZN(new_n1118));
  AOI21_X1  g693(.A(KEYINPUT61), .B1(new_n1117), .B2(new_n1118), .ZN(new_n1119));
  INV_X1    g694(.A(new_n1118), .ZN(new_n1120));
  INV_X1    g695(.A(KEYINPUT61), .ZN(new_n1121));
  NOR3_X1   g696(.A1(new_n1120), .A2(new_n1116), .A3(new_n1121), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1111), .A2(new_n767), .ZN(new_n1123));
  XOR2_X1   g698(.A(KEYINPUT58), .B(G1341), .Z(new_n1124));
  NAND2_X1  g699(.A1(new_n1023), .A2(new_n1124), .ZN(new_n1125));
  AOI21_X1  g700(.A(new_n829), .B1(new_n1123), .B2(new_n1125), .ZN(new_n1126));
  XNOR2_X1  g701(.A(new_n1126), .B(KEYINPUT59), .ZN(new_n1127));
  NOR3_X1   g702(.A1(new_n1119), .A2(new_n1122), .A3(new_n1127), .ZN(new_n1128));
  NAND2_X1  g703(.A1(new_n1108), .A2(new_n1128), .ZN(new_n1129));
  NOR2_X1   g704(.A1(new_n1103), .A2(new_n612), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1118), .B1(new_n1130), .B2(new_n1116), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1089), .B1(new_n1129), .B2(new_n1131), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1082), .A2(KEYINPUT62), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1087), .A2(G171), .ZN(new_n1134));
  NOR3_X1   g709(.A1(new_n1056), .A2(new_n1134), .A3(new_n1066), .ZN(new_n1135));
  INV_X1    g710(.A(KEYINPUT62), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1079), .A2(new_n1136), .A3(new_n1081), .ZN(new_n1137));
  NAND3_X1  g712(.A1(new_n1133), .A2(new_n1135), .A3(new_n1137), .ZN(new_n1138));
  AND2_X1   g713(.A1(new_n1053), .A2(new_n1054), .ZN(new_n1139));
  INV_X1    g714(.A(new_n1021), .ZN(new_n1140));
  INV_X1    g715(.A(G1976), .ZN(new_n1141));
  NAND3_X1  g716(.A1(new_n1054), .A2(new_n1141), .A3(new_n581), .ZN(new_n1142));
  NAND2_X1  g717(.A1(new_n1142), .A2(new_n1032), .ZN(new_n1143));
  AOI22_X1  g718(.A1(new_n1139), .A2(new_n1140), .B1(new_n1143), .B2(new_n1042), .ZN(new_n1144));
  OAI211_X1 g719(.A(new_n1053), .B(new_n1054), .C1(new_n1020), .C2(new_n1017), .ZN(new_n1145));
  NAND3_X1  g720(.A1(new_n1080), .A2(G8), .A3(G168), .ZN(new_n1146));
  OAI21_X1  g721(.A(KEYINPUT63), .B1(new_n1145), .B2(new_n1146), .ZN(new_n1147));
  NAND2_X1  g722(.A1(new_n1144), .A2(new_n1147), .ZN(new_n1148));
  NOR2_X1   g723(.A1(new_n1146), .A2(KEYINPUT63), .ZN(new_n1149));
  AOI21_X1  g724(.A(new_n1148), .B1(new_n1067), .B2(new_n1149), .ZN(new_n1150));
  NAND2_X1  g725(.A1(new_n1138), .A2(new_n1150), .ZN(new_n1151));
  OAI21_X1  g726(.A(new_n962), .B1(new_n1132), .B2(new_n1151), .ZN(new_n1152));
  XNOR2_X1  g727(.A(new_n953), .B(KEYINPUT46), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n951), .A2(new_n762), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1153), .A2(new_n1154), .A3(new_n956), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT47), .ZN(new_n1156));
  NOR2_X1   g731(.A1(G290), .A2(G1986), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n950), .A2(new_n1157), .ZN(new_n1158));
  XOR2_X1   g733(.A(new_n1158), .B(KEYINPUT48), .Z(new_n1159));
  OAI21_X1  g734(.A(new_n1156), .B1(new_n960), .B2(new_n1159), .ZN(new_n1160));
  NOR2_X1   g735(.A1(new_n744), .A2(new_n746), .ZN(new_n1161));
  NAND2_X1  g736(.A1(new_n957), .A2(new_n1161), .ZN(new_n1162));
  OR2_X1    g737(.A1(new_n704), .A2(G2067), .ZN(new_n1163));
  AOI21_X1  g738(.A(new_n959), .B1(new_n1162), .B2(new_n1163), .ZN(new_n1164));
  NOR2_X1   g739(.A1(new_n1160), .A2(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1152), .A2(new_n1165), .ZN(G329));
  assign    G231 = 1'b0;
  AOI211_X1 g741(.A(new_n460), .B(G227), .C1(new_n657), .C2(new_n659), .ZN(new_n1168));
  NAND3_X1  g742(.A1(new_n696), .A2(new_n864), .A3(new_n1168), .ZN(new_n1169));
  NOR2_X1   g743(.A1(new_n929), .A2(new_n931), .ZN(new_n1170));
  NOR2_X1   g744(.A1(new_n1169), .A2(new_n1170), .ZN(G308));
  OR2_X1    g745(.A1(new_n1169), .A2(new_n1170), .ZN(G225));
endmodule


