//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 0 0 1 0 1 1 0 0 0 1 1 0 1 1 0 0 0 0 1 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 1 0 0 1 1 1 0 0 1 0 0 1 1 0 1 1 0 0 0 0 0 0 0' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:23:47 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n615,
    new_n616, new_n617, new_n618, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n663, new_n664, new_n665, new_n666, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n677,
    new_n679, new_n680, new_n681, new_n682, new_n683, new_n684, new_n685,
    new_n686, new_n687, new_n688, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n729, new_n730, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n747, new_n748, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n891,
    new_n892, new_n893, new_n894, new_n895, new_n897, new_n898, new_n899,
    new_n900, new_n901, new_n902, new_n903, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n914,
    new_n916, new_n917, new_n918, new_n919, new_n921, new_n922, new_n923,
    new_n924, new_n925, new_n926, new_n927, new_n928, new_n929, new_n930,
    new_n931, new_n932, new_n933, new_n934, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n967, new_n968, new_n969, new_n970, new_n971, new_n972;
  INV_X1    g000(.A(G469), .ZN(new_n187));
  INV_X1    g001(.A(G902), .ZN(new_n188));
  AND2_X1   g002(.A1(KEYINPUT0), .A2(G128), .ZN(new_n189));
  XNOR2_X1  g003(.A(G143), .B(G146), .ZN(new_n190));
  OAI21_X1  g004(.A(new_n189), .B1(new_n190), .B2(KEYINPUT64), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NAND2_X1  g006(.A1(new_n192), .A2(G143), .ZN(new_n193));
  INV_X1    g007(.A(G143), .ZN(new_n194));
  NAND2_X1  g008(.A1(new_n194), .A2(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n193), .A2(new_n195), .ZN(new_n196));
  NOR2_X1   g010(.A1(KEYINPUT0), .A2(G128), .ZN(new_n197));
  NOR2_X1   g011(.A1(new_n189), .A2(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT64), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT68), .ZN(new_n201));
  NAND3_X1  g015(.A1(new_n191), .A2(new_n200), .A3(new_n201), .ZN(new_n202));
  AND3_X1   g016(.A1(new_n196), .A2(new_n198), .A3(new_n199), .ZN(new_n203));
  INV_X1    g017(.A(new_n189), .ZN(new_n204));
  AOI21_X1  g018(.A(new_n204), .B1(new_n196), .B2(new_n199), .ZN(new_n205));
  OAI21_X1  g019(.A(KEYINPUT68), .B1(new_n203), .B2(new_n205), .ZN(new_n206));
  INV_X1    g020(.A(G101), .ZN(new_n207));
  INV_X1    g021(.A(G104), .ZN(new_n208));
  OAI21_X1  g022(.A(KEYINPUT3), .B1(new_n208), .B2(G107), .ZN(new_n209));
  INV_X1    g023(.A(G107), .ZN(new_n210));
  NOR2_X1   g024(.A1(new_n210), .A2(G104), .ZN(new_n211));
  AND2_X1   g025(.A1(KEYINPUT79), .A2(G107), .ZN(new_n212));
  NOR2_X1   g026(.A1(KEYINPUT79), .A2(G107), .ZN(new_n213));
  NOR2_X1   g027(.A1(new_n212), .A2(new_n213), .ZN(new_n214));
  AOI21_X1  g028(.A(new_n211), .B1(new_n214), .B2(G104), .ZN(new_n215));
  OAI211_X1 g029(.A(new_n207), .B(new_n209), .C1(new_n215), .C2(KEYINPUT3), .ZN(new_n216));
  OAI21_X1  g030(.A(new_n209), .B1(new_n215), .B2(KEYINPUT3), .ZN(new_n217));
  NOR2_X1   g031(.A1(new_n207), .A2(KEYINPUT80), .ZN(new_n218));
  AOI22_X1  g032(.A1(new_n216), .A2(KEYINPUT4), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OR2_X1    g033(.A1(KEYINPUT79), .A2(G107), .ZN(new_n220));
  NAND2_X1  g034(.A1(KEYINPUT79), .A2(G107), .ZN(new_n221));
  NAND3_X1  g035(.A1(new_n220), .A2(G104), .A3(new_n221), .ZN(new_n222));
  INV_X1    g036(.A(new_n211), .ZN(new_n223));
  AOI21_X1  g037(.A(KEYINPUT3), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(new_n209), .ZN(new_n225));
  OAI211_X1 g039(.A(KEYINPUT4), .B(new_n218), .C1(new_n224), .C2(new_n225), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  OAI211_X1 g041(.A(new_n202), .B(new_n206), .C1(new_n219), .C2(new_n227), .ZN(new_n228));
  INV_X1    g042(.A(KEYINPUT11), .ZN(new_n229));
  INV_X1    g043(.A(G134), .ZN(new_n230));
  OAI21_X1  g044(.A(new_n229), .B1(new_n230), .B2(G137), .ZN(new_n231));
  INV_X1    g045(.A(G137), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n232), .A2(KEYINPUT11), .A3(G134), .ZN(new_n233));
  NAND2_X1  g047(.A1(new_n230), .A2(G137), .ZN(new_n234));
  NAND3_X1  g048(.A1(new_n231), .A2(new_n233), .A3(new_n234), .ZN(new_n235));
  NAND2_X1  g049(.A1(new_n235), .A2(G131), .ZN(new_n236));
  INV_X1    g050(.A(G131), .ZN(new_n237));
  NAND4_X1  g051(.A1(new_n231), .A2(new_n233), .A3(new_n237), .A4(new_n234), .ZN(new_n238));
  AND2_X1   g052(.A1(new_n236), .A2(new_n238), .ZN(new_n239));
  INV_X1    g053(.A(KEYINPUT82), .ZN(new_n240));
  INV_X1    g054(.A(KEYINPUT81), .ZN(new_n241));
  OAI211_X1 g055(.A(new_n241), .B(new_n208), .C1(new_n212), .C2(new_n213), .ZN(new_n242));
  NAND2_X1  g056(.A1(new_n242), .A2(G101), .ZN(new_n243));
  OAI21_X1  g057(.A(KEYINPUT81), .B1(new_n208), .B2(G107), .ZN(new_n244));
  XNOR2_X1  g058(.A(KEYINPUT79), .B(G107), .ZN(new_n245));
  AOI21_X1  g059(.A(new_n244), .B1(new_n245), .B2(new_n208), .ZN(new_n246));
  OAI21_X1  g060(.A(new_n240), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(new_n244), .ZN(new_n248));
  OAI21_X1  g062(.A(new_n248), .B1(new_n214), .B2(G104), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(KEYINPUT82), .A3(G101), .A4(new_n242), .ZN(new_n250));
  AND3_X1   g064(.A1(new_n216), .A2(new_n247), .A3(new_n250), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n193), .A2(KEYINPUT1), .ZN(new_n252));
  NAND3_X1  g066(.A1(new_n196), .A2(new_n252), .A3(G128), .ZN(new_n253));
  INV_X1    g067(.A(G128), .ZN(new_n254));
  OAI211_X1 g068(.A(new_n193), .B(new_n195), .C1(KEYINPUT1), .C2(new_n254), .ZN(new_n255));
  AND2_X1   g069(.A1(new_n253), .A2(new_n255), .ZN(new_n256));
  NAND3_X1  g070(.A1(new_n251), .A2(KEYINPUT10), .A3(new_n256), .ZN(new_n257));
  NAND4_X1  g071(.A1(new_n216), .A2(new_n247), .A3(new_n250), .A4(new_n256), .ZN(new_n258));
  INV_X1    g072(.A(KEYINPUT10), .ZN(new_n259));
  NAND2_X1  g073(.A1(new_n258), .A2(new_n259), .ZN(new_n260));
  NAND4_X1  g074(.A1(new_n228), .A2(new_n239), .A3(new_n257), .A4(new_n260), .ZN(new_n261));
  INV_X1    g075(.A(G953), .ZN(new_n262));
  NAND2_X1  g076(.A1(new_n262), .A2(G227), .ZN(new_n263));
  XNOR2_X1  g077(.A(new_n263), .B(KEYINPUT78), .ZN(new_n264));
  XNOR2_X1  g078(.A(G110), .B(G140), .ZN(new_n265));
  XNOR2_X1  g079(.A(new_n264), .B(new_n265), .ZN(new_n266));
  NAND2_X1  g080(.A1(new_n261), .A2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT83), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n216), .A2(new_n247), .A3(new_n250), .ZN(new_n269));
  INV_X1    g083(.A(new_n256), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n269), .A2(new_n270), .ZN(new_n271));
  AOI21_X1  g085(.A(new_n239), .B1(new_n271), .B2(new_n258), .ZN(new_n272));
  AOI21_X1  g086(.A(new_n268), .B1(new_n272), .B2(KEYINPUT12), .ZN(new_n273));
  NOR2_X1   g087(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n274));
  NOR2_X1   g088(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n272), .A2(new_n268), .A3(KEYINPUT12), .ZN(new_n276));
  AOI21_X1  g090(.A(new_n267), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  NAND3_X1  g091(.A1(new_n228), .A2(new_n257), .A3(new_n260), .ZN(new_n278));
  NAND2_X1  g092(.A1(new_n236), .A2(new_n238), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  AOI21_X1  g094(.A(new_n266), .B1(new_n280), .B2(new_n261), .ZN(new_n281));
  OAI211_X1 g095(.A(new_n187), .B(new_n188), .C1(new_n277), .C2(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(new_n267), .ZN(new_n283));
  NAND2_X1  g097(.A1(new_n283), .A2(new_n280), .ZN(new_n284));
  INV_X1    g098(.A(new_n261), .ZN(new_n285));
  AOI21_X1  g099(.A(new_n285), .B1(new_n275), .B2(new_n276), .ZN(new_n286));
  OAI211_X1 g100(.A(G469), .B(new_n284), .C1(new_n286), .C2(new_n266), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n187), .A2(new_n188), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND3_X1  g103(.A1(new_n282), .A2(new_n287), .A3(new_n289), .ZN(new_n290));
  XNOR2_X1  g104(.A(KEYINPUT9), .B(G234), .ZN(new_n291));
  OAI21_X1  g105(.A(G221), .B1(new_n291), .B2(G902), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n292), .B(KEYINPUT76), .ZN(new_n293));
  XOR2_X1   g107(.A(new_n293), .B(KEYINPUT77), .Z(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n290), .A2(new_n295), .ZN(new_n296));
  OAI21_X1  g110(.A(G210), .B1(G237), .B2(G902), .ZN(new_n297));
  INV_X1    g111(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g112(.A1(new_n191), .A2(new_n200), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  NAND2_X1  g114(.A1(new_n300), .A2(G125), .ZN(new_n301));
  INV_X1    g115(.A(G125), .ZN(new_n302));
  NAND2_X1  g116(.A1(new_n256), .A2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  INV_X1    g118(.A(G224), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n305), .A2(G953), .ZN(new_n306));
  XNOR2_X1  g120(.A(new_n306), .B(KEYINPUT86), .ZN(new_n307));
  XNOR2_X1  g121(.A(new_n304), .B(new_n307), .ZN(new_n308));
  INV_X1    g122(.A(new_n308), .ZN(new_n309));
  XNOR2_X1  g123(.A(G110), .B(G122), .ZN(new_n310));
  NOR2_X1   g124(.A1(new_n310), .A2(KEYINPUT85), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT67), .ZN(new_n312));
  NAND3_X1  g126(.A1(KEYINPUT65), .A2(KEYINPUT2), .A3(G113), .ZN(new_n313));
  INV_X1    g127(.A(new_n313), .ZN(new_n314));
  AOI21_X1  g128(.A(KEYINPUT65), .B1(KEYINPUT2), .B2(G113), .ZN(new_n315));
  OAI22_X1  g129(.A1(new_n314), .A2(new_n315), .B1(KEYINPUT2), .B2(G113), .ZN(new_n316));
  INV_X1    g130(.A(G119), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n317), .A2(G116), .ZN(new_n318));
  INV_X1    g132(.A(G116), .ZN(new_n319));
  NAND2_X1  g133(.A1(new_n319), .A2(G119), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n318), .A2(new_n320), .ZN(new_n321));
  OAI21_X1  g135(.A(new_n312), .B1(new_n316), .B2(new_n321), .ZN(new_n322));
  NOR2_X1   g136(.A1(KEYINPUT2), .A2(G113), .ZN(new_n323));
  INV_X1    g137(.A(new_n315), .ZN(new_n324));
  AOI21_X1  g138(.A(new_n323), .B1(new_n324), .B2(new_n313), .ZN(new_n325));
  INV_X1    g139(.A(new_n321), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n325), .A2(KEYINPUT67), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(KEYINPUT66), .ZN(new_n328));
  AOI21_X1  g142(.A(new_n326), .B1(new_n316), .B2(new_n328), .ZN(new_n329));
  NAND2_X1  g143(.A1(new_n325), .A2(KEYINPUT66), .ZN(new_n330));
  AOI22_X1  g144(.A1(new_n322), .A2(new_n327), .B1(new_n329), .B2(new_n330), .ZN(new_n331));
  OAI21_X1  g145(.A(new_n218), .B1(new_n224), .B2(new_n225), .ZN(new_n332));
  NOR3_X1   g146(.A1(new_n224), .A2(G101), .A3(new_n225), .ZN(new_n333));
  INV_X1    g147(.A(KEYINPUT4), .ZN(new_n334));
  OAI21_X1  g148(.A(new_n332), .B1(new_n333), .B2(new_n334), .ZN(new_n335));
  AOI21_X1  g149(.A(new_n331), .B1(new_n335), .B2(new_n226), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n322), .A2(new_n327), .ZN(new_n337));
  AND3_X1   g151(.A1(new_n318), .A2(new_n320), .A3(KEYINPUT5), .ZN(new_n338));
  OAI21_X1  g152(.A(G113), .B1(new_n318), .B2(KEYINPUT5), .ZN(new_n339));
  OR3_X1    g153(.A1(new_n338), .A2(new_n339), .A3(KEYINPUT84), .ZN(new_n340));
  OAI21_X1  g154(.A(KEYINPUT84), .B1(new_n338), .B2(new_n339), .ZN(new_n341));
  NAND3_X1  g155(.A1(new_n337), .A2(new_n340), .A3(new_n341), .ZN(new_n342));
  NOR2_X1   g156(.A1(new_n342), .A2(new_n269), .ZN(new_n343));
  OAI21_X1  g157(.A(new_n311), .B1(new_n336), .B2(new_n343), .ZN(new_n344));
  INV_X1    g158(.A(new_n310), .ZN(new_n345));
  NOR3_X1   g159(.A1(new_n336), .A2(new_n343), .A3(new_n345), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT6), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n344), .B1(new_n346), .B2(new_n347), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n329), .A2(new_n330), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n349), .A2(new_n337), .ZN(new_n350));
  OAI21_X1  g164(.A(new_n350), .B1(new_n219), .B2(new_n227), .ZN(new_n351));
  OR2_X1    g165(.A1(new_n342), .A2(new_n269), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  NAND3_X1  g167(.A1(new_n353), .A2(KEYINPUT6), .A3(new_n311), .ZN(new_n354));
  AOI21_X1  g168(.A(new_n309), .B1(new_n348), .B2(new_n354), .ZN(new_n355));
  OAI21_X1  g169(.A(KEYINPUT7), .B1(new_n305), .B2(G953), .ZN(new_n356));
  NAND3_X1  g170(.A1(new_n301), .A2(new_n303), .A3(new_n356), .ZN(new_n357));
  INV_X1    g171(.A(new_n356), .ZN(new_n358));
  NAND2_X1  g172(.A1(new_n304), .A2(new_n358), .ZN(new_n359));
  OAI21_X1  g173(.A(new_n337), .B1(new_n338), .B2(new_n339), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n251), .A2(new_n360), .ZN(new_n361));
  XNOR2_X1  g175(.A(new_n310), .B(KEYINPUT8), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NOR2_X1   g177(.A1(new_n251), .A2(new_n342), .ZN(new_n364));
  OAI211_X1 g178(.A(new_n357), .B(new_n359), .C1(new_n363), .C2(new_n364), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n188), .B1(new_n365), .B2(new_n346), .ZN(new_n366));
  OAI21_X1  g180(.A(new_n298), .B1(new_n355), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n351), .A2(new_n352), .A3(new_n310), .ZN(new_n368));
  AOI22_X1  g182(.A1(new_n368), .A2(KEYINPUT6), .B1(new_n353), .B2(new_n311), .ZN(new_n369));
  NOR2_X1   g183(.A1(new_n344), .A2(new_n347), .ZN(new_n370));
  OAI21_X1  g184(.A(new_n308), .B1(new_n369), .B2(new_n370), .ZN(new_n371));
  INV_X1    g185(.A(new_n366), .ZN(new_n372));
  NAND3_X1  g186(.A1(new_n371), .A2(new_n372), .A3(new_n297), .ZN(new_n373));
  NAND3_X1  g187(.A1(new_n367), .A2(new_n373), .A3(KEYINPUT87), .ZN(new_n374));
  NAND2_X1  g188(.A1(G234), .A2(G237), .ZN(new_n375));
  AND3_X1   g189(.A1(new_n375), .A2(G952), .A3(new_n262), .ZN(new_n376));
  AND3_X1   g190(.A1(new_n375), .A2(G902), .A3(G953), .ZN(new_n377));
  XNOR2_X1  g191(.A(KEYINPUT21), .B(G898), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n376), .B1(new_n377), .B2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n379), .ZN(new_n380));
  NOR2_X1   g194(.A1(G475), .A2(G902), .ZN(new_n381));
  AND2_X1   g195(.A1(KEYINPUT69), .A2(G237), .ZN(new_n382));
  NOR2_X1   g196(.A1(KEYINPUT69), .A2(G237), .ZN(new_n383));
  OAI211_X1 g197(.A(G214), .B(new_n262), .C1(new_n382), .C2(new_n383), .ZN(new_n384));
  XOR2_X1   g198(.A(KEYINPUT88), .B(G143), .Z(new_n385));
  NAND2_X1  g199(.A1(new_n384), .A2(new_n385), .ZN(new_n386));
  XNOR2_X1  g200(.A(KEYINPUT69), .B(G237), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n194), .A2(KEYINPUT88), .ZN(new_n388));
  NAND4_X1  g202(.A1(new_n387), .A2(G214), .A3(new_n262), .A4(new_n388), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n386), .A2(new_n389), .ZN(new_n390));
  NAND4_X1  g204(.A1(new_n390), .A2(KEYINPUT89), .A3(KEYINPUT18), .A4(G131), .ZN(new_n391));
  INV_X1    g205(.A(G140), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G125), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n302), .A2(G140), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT75), .ZN(new_n396));
  NOR3_X1   g210(.A1(new_n395), .A2(new_n396), .A3(G146), .ZN(new_n397));
  XNOR2_X1  g211(.A(G125), .B(G140), .ZN(new_n398));
  AOI21_X1  g212(.A(KEYINPUT75), .B1(new_n398), .B2(new_n192), .ZN(new_n399));
  OAI22_X1  g213(.A1(new_n397), .A2(new_n399), .B1(new_n192), .B2(new_n398), .ZN(new_n400));
  NAND2_X1  g214(.A1(KEYINPUT89), .A2(KEYINPUT18), .ZN(new_n401));
  NAND3_X1  g215(.A1(new_n386), .A2(new_n389), .A3(new_n401), .ZN(new_n402));
  NAND3_X1  g216(.A1(new_n386), .A2(new_n389), .A3(new_n237), .ZN(new_n403));
  NAND4_X1  g217(.A1(new_n391), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  XNOR2_X1  g218(.A(G113), .B(G122), .ZN(new_n405));
  XNOR2_X1  g219(.A(KEYINPUT91), .B(G104), .ZN(new_n406));
  XNOR2_X1  g220(.A(new_n405), .B(new_n406), .ZN(new_n407));
  INV_X1    g221(.A(KEYINPUT16), .ZN(new_n408));
  NAND3_X1  g222(.A1(new_n408), .A2(new_n392), .A3(G125), .ZN(new_n409));
  OAI21_X1  g223(.A(new_n409), .B1(new_n395), .B2(new_n408), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n410), .A2(new_n192), .ZN(new_n411));
  OAI211_X1 g225(.A(G146), .B(new_n409), .C1(new_n395), .C2(new_n408), .ZN(new_n412));
  NAND2_X1  g226(.A1(new_n411), .A2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(new_n413), .ZN(new_n414));
  AOI21_X1  g228(.A(new_n237), .B1(new_n386), .B2(new_n389), .ZN(new_n415));
  NAND2_X1  g229(.A1(new_n415), .A2(KEYINPUT17), .ZN(new_n416));
  NAND2_X1  g230(.A1(new_n414), .A2(new_n416), .ZN(new_n417));
  AND3_X1   g231(.A1(new_n386), .A2(new_n389), .A3(new_n237), .ZN(new_n418));
  NOR3_X1   g232(.A1(new_n418), .A2(new_n415), .A3(KEYINPUT17), .ZN(new_n419));
  OAI211_X1 g233(.A(new_n404), .B(new_n407), .C1(new_n417), .C2(new_n419), .ZN(new_n420));
  INV_X1    g234(.A(new_n420), .ZN(new_n421));
  OAI21_X1  g235(.A(KEYINPUT90), .B1(new_n418), .B2(new_n415), .ZN(new_n422));
  NAND2_X1  g236(.A1(new_n390), .A2(G131), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT90), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n423), .A2(new_n424), .A3(new_n403), .ZN(new_n425));
  INV_X1    g239(.A(new_n412), .ZN(new_n426));
  XNOR2_X1  g240(.A(new_n398), .B(KEYINPUT19), .ZN(new_n427));
  AOI21_X1  g241(.A(new_n426), .B1(new_n192), .B2(new_n427), .ZN(new_n428));
  NAND3_X1  g242(.A1(new_n422), .A2(new_n425), .A3(new_n428), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n407), .B1(new_n429), .B2(new_n404), .ZN(new_n430));
  OAI21_X1  g244(.A(new_n381), .B1(new_n421), .B2(new_n430), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n431), .A2(KEYINPUT20), .ZN(new_n432));
  INV_X1    g246(.A(KEYINPUT20), .ZN(new_n433));
  OAI211_X1 g247(.A(new_n433), .B(new_n381), .C1(new_n421), .C2(new_n430), .ZN(new_n434));
  NAND2_X1  g248(.A1(new_n432), .A2(new_n434), .ZN(new_n435));
  INV_X1    g249(.A(G478), .ZN(new_n436));
  NOR2_X1   g250(.A1(new_n436), .A2(KEYINPUT15), .ZN(new_n437));
  INV_X1    g251(.A(new_n437), .ZN(new_n438));
  INV_X1    g252(.A(G217), .ZN(new_n439));
  NOR3_X1   g253(.A1(new_n291), .A2(new_n439), .A3(G953), .ZN(new_n440));
  INV_X1    g254(.A(new_n440), .ZN(new_n441));
  XNOR2_X1  g255(.A(G116), .B(G122), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n214), .A2(new_n442), .ZN(new_n443));
  INV_X1    g257(.A(G122), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n444), .A2(G116), .ZN(new_n445));
  NAND2_X1  g259(.A1(new_n319), .A2(G122), .ZN(new_n446));
  NAND2_X1  g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NOR2_X1   g261(.A1(new_n447), .A2(KEYINPUT14), .ZN(new_n448));
  INV_X1    g262(.A(KEYINPUT14), .ZN(new_n449));
  OAI21_X1  g263(.A(G107), .B1(new_n446), .B2(new_n449), .ZN(new_n450));
  OAI21_X1  g264(.A(new_n443), .B1(new_n448), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g265(.A1(new_n194), .A2(G128), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n254), .A2(G143), .ZN(new_n453));
  NAND2_X1  g267(.A1(new_n452), .A2(new_n453), .ZN(new_n454));
  INV_X1    g268(.A(KEYINPUT92), .ZN(new_n455));
  NOR2_X1   g269(.A1(new_n454), .A2(new_n455), .ZN(new_n456));
  XNOR2_X1  g270(.A(G128), .B(G143), .ZN(new_n457));
  NOR2_X1   g271(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n458));
  OAI21_X1  g272(.A(new_n230), .B1(new_n456), .B2(new_n458), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n454), .A2(new_n455), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(KEYINPUT92), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(new_n461), .A3(G134), .ZN(new_n462));
  AOI21_X1  g276(.A(new_n451), .B1(new_n459), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n447), .A2(new_n245), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n464), .A2(new_n443), .ZN(new_n465));
  INV_X1    g279(.A(KEYINPUT13), .ZN(new_n466));
  NAND3_X1  g280(.A1(new_n466), .A2(new_n194), .A3(G128), .ZN(new_n467));
  OAI211_X1 g281(.A(G134), .B(new_n467), .C1(new_n454), .C2(new_n466), .ZN(new_n468));
  NAND2_X1  g282(.A1(new_n465), .A2(new_n468), .ZN(new_n469));
  AOI21_X1  g283(.A(G134), .B1(new_n460), .B2(new_n461), .ZN(new_n470));
  NOR2_X1   g284(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  OAI21_X1  g285(.A(new_n441), .B1(new_n463), .B2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(new_n450), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n442), .A2(new_n449), .ZN(new_n474));
  AOI22_X1  g288(.A1(new_n473), .A2(new_n474), .B1(new_n214), .B2(new_n442), .ZN(new_n475));
  INV_X1    g289(.A(new_n462), .ZN(new_n476));
  OAI21_X1  g290(.A(new_n475), .B1(new_n476), .B2(new_n470), .ZN(new_n477));
  NAND3_X1  g291(.A1(new_n459), .A2(new_n465), .A3(new_n468), .ZN(new_n478));
  NAND3_X1  g292(.A1(new_n477), .A2(new_n478), .A3(new_n440), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n472), .A2(new_n479), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n438), .B1(new_n480), .B2(new_n188), .ZN(new_n481));
  AOI211_X1 g295(.A(G902), .B(new_n437), .C1(new_n472), .C2(new_n479), .ZN(new_n482));
  NOR2_X1   g296(.A1(new_n481), .A2(new_n482), .ZN(new_n483));
  INV_X1    g297(.A(KEYINPUT17), .ZN(new_n484));
  NAND3_X1  g298(.A1(new_n423), .A2(new_n484), .A3(new_n403), .ZN(new_n485));
  NAND3_X1  g299(.A1(new_n485), .A2(new_n414), .A3(new_n416), .ZN(new_n486));
  AOI21_X1  g300(.A(new_n407), .B1(new_n486), .B2(new_n404), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n188), .B1(new_n421), .B2(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(G475), .ZN(new_n489));
  AND4_X1   g303(.A1(new_n380), .A2(new_n435), .A3(new_n483), .A4(new_n489), .ZN(new_n490));
  OAI21_X1  g304(.A(G214), .B1(G237), .B2(G902), .ZN(new_n491));
  INV_X1    g305(.A(KEYINPUT87), .ZN(new_n492));
  NAND4_X1  g306(.A1(new_n371), .A2(new_n372), .A3(new_n492), .A4(new_n297), .ZN(new_n493));
  NAND4_X1  g307(.A1(new_n374), .A2(new_n490), .A3(new_n491), .A4(new_n493), .ZN(new_n494));
  NOR2_X1   g308(.A1(new_n296), .A2(new_n494), .ZN(new_n495));
  INV_X1    g309(.A(KEYINPUT72), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n387), .A2(G210), .A3(new_n262), .ZN(new_n497));
  XNOR2_X1  g311(.A(new_n497), .B(KEYINPUT27), .ZN(new_n498));
  XNOR2_X1  g312(.A(KEYINPUT26), .B(G101), .ZN(new_n499));
  XNOR2_X1  g313(.A(new_n498), .B(new_n499), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  INV_X1    g315(.A(KEYINPUT71), .ZN(new_n502));
  NOR2_X1   g316(.A1(new_n230), .A2(G137), .ZN(new_n503));
  NOR2_X1   g317(.A1(new_n232), .A2(G134), .ZN(new_n504));
  OAI21_X1  g318(.A(G131), .B1(new_n503), .B2(new_n504), .ZN(new_n505));
  AND2_X1   g319(.A1(new_n238), .A2(new_n505), .ZN(new_n506));
  AOI22_X1  g320(.A1(new_n300), .A2(new_n279), .B1(new_n256), .B2(new_n506), .ZN(new_n507));
  OAI21_X1  g321(.A(new_n502), .B1(new_n507), .B2(new_n331), .ZN(new_n508));
  NAND3_X1  g322(.A1(new_n206), .A2(new_n279), .A3(new_n202), .ZN(new_n509));
  NAND4_X1  g323(.A1(new_n253), .A2(new_n238), .A3(new_n255), .A4(new_n505), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n509), .A2(new_n331), .A3(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n510), .B1(new_n239), .B2(new_n299), .ZN(new_n512));
  NAND3_X1  g326(.A1(new_n512), .A2(new_n350), .A3(KEYINPUT71), .ZN(new_n513));
  NAND3_X1  g327(.A1(new_n508), .A2(new_n511), .A3(new_n513), .ZN(new_n514));
  AND2_X1   g328(.A1(new_n514), .A2(KEYINPUT28), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT28), .ZN(new_n516));
  AND2_X1   g330(.A1(new_n511), .A2(new_n516), .ZN(new_n517));
  OAI211_X1 g331(.A(new_n496), .B(new_n501), .C1(new_n515), .C2(new_n517), .ZN(new_n518));
  AOI21_X1  g332(.A(new_n517), .B1(new_n514), .B2(KEYINPUT28), .ZN(new_n519));
  OAI21_X1  g333(.A(KEYINPUT72), .B1(new_n519), .B2(new_n500), .ZN(new_n520));
  NAND3_X1  g334(.A1(new_n509), .A2(KEYINPUT30), .A3(new_n510), .ZN(new_n521));
  INV_X1    g335(.A(KEYINPUT30), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n512), .A2(new_n522), .ZN(new_n523));
  NAND3_X1  g337(.A1(new_n521), .A2(new_n350), .A3(new_n523), .ZN(new_n524));
  NAND3_X1  g338(.A1(new_n524), .A2(new_n500), .A3(new_n511), .ZN(new_n525));
  NAND2_X1  g339(.A1(new_n525), .A2(KEYINPUT70), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT70), .ZN(new_n527));
  NAND4_X1  g341(.A1(new_n524), .A2(new_n527), .A3(new_n500), .A4(new_n511), .ZN(new_n528));
  NAND3_X1  g342(.A1(new_n526), .A2(KEYINPUT31), .A3(new_n528), .ZN(new_n529));
  OR2_X1    g343(.A1(new_n525), .A2(KEYINPUT31), .ZN(new_n530));
  NAND4_X1  g344(.A1(new_n518), .A2(new_n520), .A3(new_n529), .A4(new_n530), .ZN(new_n531));
  INV_X1    g345(.A(G472), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n531), .A2(new_n532), .A3(new_n188), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n533), .A2(KEYINPUT32), .ZN(new_n534));
  INV_X1    g348(.A(KEYINPUT32), .ZN(new_n535));
  NAND4_X1  g349(.A1(new_n531), .A2(new_n535), .A3(new_n532), .A4(new_n188), .ZN(new_n536));
  NAND2_X1  g350(.A1(new_n534), .A2(new_n536), .ZN(new_n537));
  NAND2_X1  g351(.A1(new_n519), .A2(new_n500), .ZN(new_n538));
  NAND2_X1  g352(.A1(new_n524), .A2(new_n511), .ZN(new_n539));
  AOI21_X1  g353(.A(KEYINPUT29), .B1(new_n539), .B2(new_n501), .ZN(new_n540));
  NAND3_X1  g354(.A1(new_n538), .A2(KEYINPUT73), .A3(new_n540), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n509), .A2(new_n510), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n542), .A2(new_n350), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n516), .B1(new_n543), .B2(new_n511), .ZN(new_n544));
  NOR2_X1   g358(.A1(new_n544), .A2(new_n517), .ZN(new_n545));
  AND2_X1   g359(.A1(new_n500), .A2(KEYINPUT29), .ZN(new_n546));
  AOI21_X1  g360(.A(G902), .B1(new_n545), .B2(new_n546), .ZN(new_n547));
  AND2_X1   g361(.A1(new_n541), .A2(new_n547), .ZN(new_n548));
  NAND2_X1  g362(.A1(new_n538), .A2(new_n540), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT73), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  AOI21_X1  g365(.A(new_n532), .B1(new_n548), .B2(new_n551), .ZN(new_n552));
  INV_X1    g366(.A(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n537), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n254), .A2(G119), .ZN(new_n555));
  NAND2_X1  g369(.A1(new_n555), .A2(KEYINPUT74), .ZN(new_n556));
  NAND2_X1  g370(.A1(new_n556), .A2(KEYINPUT23), .ZN(new_n557));
  INV_X1    g371(.A(KEYINPUT23), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n555), .A2(KEYINPUT74), .A3(new_n558), .ZN(new_n559));
  NAND2_X1  g373(.A1(new_n317), .A2(G128), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n557), .A2(new_n559), .A3(new_n560), .ZN(new_n561));
  AND2_X1   g375(.A1(new_n555), .A2(new_n560), .ZN(new_n562));
  XOR2_X1   g376(.A(KEYINPUT24), .B(G110), .Z(new_n563));
  OAI22_X1  g377(.A1(new_n561), .A2(G110), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  OAI211_X1 g378(.A(new_n564), .B(new_n412), .C1(new_n399), .C2(new_n397), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n561), .A2(G110), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n562), .A2(new_n563), .ZN(new_n567));
  NAND3_X1  g381(.A1(new_n413), .A2(new_n566), .A3(new_n567), .ZN(new_n568));
  NAND2_X1  g382(.A1(new_n565), .A2(new_n568), .ZN(new_n569));
  XNOR2_X1  g383(.A(KEYINPUT22), .B(G137), .ZN(new_n570));
  NAND3_X1  g384(.A1(new_n262), .A2(G221), .A3(G234), .ZN(new_n571));
  XNOR2_X1  g385(.A(new_n570), .B(new_n571), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n569), .A2(new_n573), .ZN(new_n574));
  NAND3_X1  g388(.A1(new_n565), .A2(new_n568), .A3(new_n572), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  INV_X1    g390(.A(new_n576), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n577), .A2(KEYINPUT25), .A3(new_n188), .ZN(new_n578));
  INV_X1    g392(.A(KEYINPUT25), .ZN(new_n579));
  OAI21_X1  g393(.A(new_n579), .B1(new_n576), .B2(G902), .ZN(new_n580));
  NAND2_X1  g394(.A1(new_n578), .A2(new_n580), .ZN(new_n581));
  AOI21_X1  g395(.A(new_n439), .B1(G234), .B2(new_n188), .ZN(new_n582));
  NAND2_X1  g396(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR2_X1   g397(.A1(new_n582), .A2(G902), .ZN(new_n584));
  INV_X1    g398(.A(new_n584), .ZN(new_n585));
  OAI21_X1  g399(.A(new_n583), .B1(new_n576), .B2(new_n585), .ZN(new_n586));
  INV_X1    g400(.A(new_n586), .ZN(new_n587));
  NAND3_X1  g401(.A1(new_n495), .A2(new_n554), .A3(new_n587), .ZN(new_n588));
  XNOR2_X1  g402(.A(new_n588), .B(G101), .ZN(G3));
  AOI21_X1  g403(.A(new_n532), .B1(new_n531), .B2(new_n188), .ZN(new_n590));
  INV_X1    g404(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n591), .A2(new_n533), .ZN(new_n592));
  NOR3_X1   g406(.A1(new_n592), .A2(new_n296), .A3(new_n586), .ZN(new_n593));
  INV_X1    g407(.A(new_n491), .ZN(new_n594));
  AOI21_X1  g408(.A(new_n594), .B1(new_n367), .B2(new_n373), .ZN(new_n595));
  NAND2_X1  g409(.A1(new_n595), .A2(new_n380), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n429), .A2(new_n404), .ZN(new_n597));
  OAI21_X1  g411(.A(new_n420), .B1(new_n597), .B2(new_n407), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n433), .B1(new_n598), .B2(new_n381), .ZN(new_n599));
  INV_X1    g413(.A(new_n434), .ZN(new_n600));
  OAI21_X1  g414(.A(new_n489), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  NOR2_X1   g415(.A1(new_n436), .A2(new_n188), .ZN(new_n602));
  INV_X1    g416(.A(new_n480), .ZN(new_n603));
  NOR2_X1   g417(.A1(new_n603), .A2(G902), .ZN(new_n604));
  AOI21_X1  g418(.A(new_n602), .B1(new_n604), .B2(new_n436), .ZN(new_n605));
  OR2_X1    g419(.A1(new_n480), .A2(KEYINPUT33), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n480), .A2(KEYINPUT33), .ZN(new_n607));
  NAND3_X1  g421(.A1(new_n606), .A2(G478), .A3(new_n607), .ZN(new_n608));
  AND2_X1   g422(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n601), .A2(new_n609), .ZN(new_n610));
  NOR2_X1   g424(.A1(new_n596), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g425(.A1(new_n593), .A2(new_n611), .ZN(new_n612));
  XOR2_X1   g426(.A(KEYINPUT34), .B(G104), .Z(new_n613));
  XNOR2_X1  g427(.A(new_n612), .B(new_n613), .ZN(G6));
  NOR3_X1   g428(.A1(new_n596), .A2(new_n483), .A3(new_n601), .ZN(new_n615));
  NAND2_X1  g429(.A1(new_n593), .A2(new_n615), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(new_n210), .ZN(new_n617));
  XNOR2_X1  g431(.A(KEYINPUT93), .B(KEYINPUT35), .ZN(new_n618));
  XNOR2_X1  g432(.A(new_n617), .B(new_n618), .ZN(G9));
  INV_X1    g433(.A(new_n582), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n620), .B1(new_n578), .B2(new_n580), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n573), .A2(KEYINPUT36), .ZN(new_n622));
  XNOR2_X1  g436(.A(new_n569), .B(new_n622), .ZN(new_n623));
  NAND2_X1  g437(.A1(new_n623), .A2(new_n584), .ZN(new_n624));
  INV_X1    g438(.A(new_n624), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n621), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g440(.A1(new_n626), .A2(KEYINPUT94), .ZN(new_n627));
  INV_X1    g441(.A(KEYINPUT94), .ZN(new_n628));
  OAI21_X1  g442(.A(new_n628), .B1(new_n621), .B2(new_n625), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n627), .A2(new_n629), .ZN(new_n630));
  AND3_X1   g444(.A1(new_n531), .A2(new_n532), .A3(new_n188), .ZN(new_n631));
  NOR3_X1   g445(.A1(new_n630), .A2(new_n631), .A3(new_n590), .ZN(new_n632));
  NAND2_X1  g446(.A1(new_n495), .A2(new_n632), .ZN(new_n633));
  XOR2_X1   g447(.A(KEYINPUT37), .B(G110), .Z(new_n634));
  XNOR2_X1  g448(.A(new_n633), .B(new_n634), .ZN(G12));
  AOI221_X4 g449(.A(new_n483), .B1(G475), .B2(new_n488), .C1(new_n432), .C2(new_n434), .ZN(new_n636));
  INV_X1    g450(.A(G900), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n376), .B1(new_n377), .B2(new_n637), .ZN(new_n638));
  INV_X1    g452(.A(new_n638), .ZN(new_n639));
  AND4_X1   g453(.A1(new_n295), .A2(new_n290), .A3(new_n636), .A4(new_n639), .ZN(new_n640));
  INV_X1    g454(.A(new_n630), .ZN(new_n641));
  NAND4_X1  g455(.A1(new_n554), .A2(new_n640), .A3(new_n595), .A4(new_n641), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(G128), .ZN(G30));
  INV_X1    g457(.A(new_n296), .ZN(new_n644));
  XOR2_X1   g458(.A(new_n638), .B(KEYINPUT39), .Z(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT40), .Z(new_n647));
  AND2_X1   g461(.A1(new_n526), .A2(new_n528), .ZN(new_n648));
  INV_X1    g462(.A(new_n648), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n543), .A2(new_n511), .ZN(new_n650));
  AOI21_X1  g464(.A(new_n649), .B1(new_n501), .B2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n651), .B2(G902), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n537), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g467(.A1(new_n374), .A2(new_n493), .ZN(new_n654));
  XNOR2_X1  g468(.A(KEYINPUT95), .B(KEYINPUT38), .ZN(new_n655));
  XNOR2_X1  g469(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g470(.A(new_n626), .ZN(new_n657));
  INV_X1    g471(.A(new_n483), .ZN(new_n658));
  NAND2_X1  g472(.A1(new_n601), .A2(new_n658), .ZN(new_n659));
  NOR4_X1   g473(.A1(new_n656), .A2(new_n594), .A3(new_n657), .A4(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n647), .A2(new_n653), .A3(new_n660), .ZN(new_n661));
  XNOR2_X1  g475(.A(new_n661), .B(G143), .ZN(G45));
  INV_X1    g476(.A(new_n610), .ZN(new_n663));
  NAND2_X1  g477(.A1(new_n663), .A2(new_n639), .ZN(new_n664));
  NOR2_X1   g478(.A1(new_n296), .A2(new_n664), .ZN(new_n665));
  NAND4_X1  g479(.A1(new_n554), .A2(new_n665), .A3(new_n595), .A4(new_n641), .ZN(new_n666));
  XNOR2_X1  g480(.A(new_n666), .B(G146), .ZN(G48));
  AOI21_X1  g481(.A(new_n586), .B1(new_n537), .B2(new_n553), .ZN(new_n668));
  NOR2_X1   g482(.A1(new_n277), .A2(new_n281), .ZN(new_n669));
  OAI21_X1  g483(.A(G469), .B1(new_n669), .B2(G902), .ZN(new_n670));
  NAND2_X1  g484(.A1(new_n670), .A2(new_n282), .ZN(new_n671));
  NOR2_X1   g485(.A1(new_n671), .A2(new_n293), .ZN(new_n672));
  NAND3_X1  g486(.A1(new_n668), .A2(new_n611), .A3(new_n672), .ZN(new_n673));
  XNOR2_X1  g487(.A(KEYINPUT41), .B(G113), .ZN(new_n674));
  XNOR2_X1  g488(.A(new_n674), .B(KEYINPUT96), .ZN(new_n675));
  XNOR2_X1  g489(.A(new_n673), .B(new_n675), .ZN(G15));
  NAND3_X1  g490(.A1(new_n668), .A2(new_n615), .A3(new_n672), .ZN(new_n677));
  XNOR2_X1  g491(.A(new_n677), .B(G116), .ZN(G18));
  INV_X1    g492(.A(new_n293), .ZN(new_n679));
  AND4_X1   g493(.A1(new_n679), .A2(new_n670), .A3(new_n490), .A4(new_n282), .ZN(new_n680));
  NAND4_X1  g494(.A1(new_n554), .A2(new_n595), .A3(new_n641), .A4(new_n680), .ZN(new_n681));
  INV_X1    g495(.A(KEYINPUT97), .ZN(new_n682));
  NAND2_X1  g496(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AOI21_X1  g497(.A(new_n552), .B1(new_n534), .B2(new_n536), .ZN(new_n684));
  NOR2_X1   g498(.A1(new_n684), .A2(new_n630), .ZN(new_n685));
  NAND4_X1  g499(.A1(new_n685), .A2(KEYINPUT97), .A3(new_n595), .A4(new_n680), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n683), .A2(new_n686), .ZN(new_n687));
  XNOR2_X1  g501(.A(KEYINPUT98), .B(G119), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n687), .B(new_n688), .ZN(G21));
  NOR2_X1   g503(.A1(G472), .A2(G902), .ZN(new_n690));
  INV_X1    g504(.A(KEYINPUT99), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n501), .B1(new_n544), .B2(new_n517), .ZN(new_n692));
  NAND3_X1  g506(.A1(new_n529), .A2(new_n691), .A3(new_n692), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n693), .A2(new_n530), .ZN(new_n694));
  AOI21_X1  g508(.A(new_n691), .B1(new_n529), .B2(new_n692), .ZN(new_n695));
  OAI21_X1  g509(.A(new_n690), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  AND3_X1   g510(.A1(new_n591), .A2(new_n696), .A3(new_n587), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n595), .A2(new_n670), .A3(new_n679), .A4(new_n282), .ZN(new_n698));
  INV_X1    g512(.A(new_n698), .ZN(new_n699));
  INV_X1    g513(.A(KEYINPUT100), .ZN(new_n700));
  AOI22_X1  g514(.A1(new_n432), .A2(new_n434), .B1(G475), .B2(new_n488), .ZN(new_n701));
  OAI21_X1  g515(.A(new_n700), .B1(new_n701), .B2(new_n483), .ZN(new_n702));
  NAND3_X1  g516(.A1(new_n601), .A2(KEYINPUT100), .A3(new_n658), .ZN(new_n703));
  AND3_X1   g517(.A1(new_n702), .A2(new_n703), .A3(new_n380), .ZN(new_n704));
  NAND3_X1  g518(.A1(new_n697), .A2(new_n699), .A3(new_n704), .ZN(new_n705));
  XNOR2_X1  g519(.A(new_n705), .B(G122), .ZN(G24));
  NOR2_X1   g520(.A1(new_n610), .A2(new_n638), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n591), .A2(new_n707), .A3(new_n696), .A4(new_n657), .ZN(new_n708));
  NOR2_X1   g522(.A1(new_n708), .A2(new_n698), .ZN(new_n709));
  XNOR2_X1  g523(.A(new_n709), .B(new_n302), .ZN(G27));
  NAND2_X1  g524(.A1(new_n654), .A2(new_n491), .ZN(new_n711));
  NOR2_X1   g525(.A1(new_n711), .A2(new_n293), .ZN(new_n712));
  NAND2_X1  g526(.A1(new_n290), .A2(KEYINPUT101), .ZN(new_n713));
  INV_X1    g527(.A(KEYINPUT101), .ZN(new_n714));
  NAND4_X1  g528(.A1(new_n282), .A2(new_n287), .A3(new_n714), .A4(new_n289), .ZN(new_n715));
  AND2_X1   g529(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g530(.A(KEYINPUT102), .ZN(new_n717));
  INV_X1    g531(.A(KEYINPUT42), .ZN(new_n718));
  AOI21_X1  g532(.A(new_n664), .B1(new_n717), .B2(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n668), .A2(new_n712), .A3(new_n716), .A4(new_n719), .ZN(new_n720));
  NOR2_X1   g534(.A1(new_n717), .A2(new_n718), .ZN(new_n721));
  NAND2_X1  g535(.A1(new_n720), .A2(new_n721), .ZN(new_n722));
  AOI21_X1  g536(.A(new_n594), .B1(new_n374), .B2(new_n493), .ZN(new_n723));
  AND4_X1   g537(.A1(new_n679), .A2(new_n713), .A3(new_n723), .A4(new_n715), .ZN(new_n724));
  INV_X1    g538(.A(new_n721), .ZN(new_n725));
  NAND4_X1  g539(.A1(new_n724), .A2(new_n668), .A3(new_n725), .A4(new_n719), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n722), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(new_n237), .ZN(G33));
  NAND4_X1  g542(.A1(new_n724), .A2(new_n668), .A3(new_n636), .A4(new_n639), .ZN(new_n729));
  XOR2_X1   g543(.A(KEYINPUT103), .B(G134), .Z(new_n730));
  XNOR2_X1  g544(.A(new_n729), .B(new_n730), .ZN(G36));
  INV_X1    g545(.A(KEYINPUT106), .ZN(new_n732));
  NAND2_X1  g546(.A1(new_n601), .A2(new_n732), .ZN(new_n733));
  NAND2_X1  g547(.A1(new_n701), .A2(KEYINPUT106), .ZN(new_n734));
  NAND4_X1  g548(.A1(new_n733), .A2(new_n734), .A3(KEYINPUT43), .A4(new_n609), .ZN(new_n735));
  XOR2_X1   g549(.A(KEYINPUT105), .B(KEYINPUT43), .Z(new_n736));
  NAND2_X1  g550(.A1(new_n605), .A2(new_n608), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n736), .B1(new_n601), .B2(new_n737), .ZN(new_n738));
  NAND2_X1  g552(.A1(new_n735), .A2(new_n738), .ZN(new_n739));
  OAI211_X1 g553(.A(new_n592), .B(new_n657), .C1(new_n739), .C2(KEYINPUT107), .ZN(new_n740));
  AND2_X1   g554(.A1(new_n739), .A2(KEYINPUT107), .ZN(new_n741));
  NOR2_X1   g555(.A1(new_n740), .A2(new_n741), .ZN(new_n742));
  OAI21_X1  g556(.A(KEYINPUT108), .B1(new_n742), .B2(KEYINPUT44), .ZN(new_n743));
  INV_X1    g557(.A(KEYINPUT108), .ZN(new_n744));
  INV_X1    g558(.A(KEYINPUT44), .ZN(new_n745));
  OAI211_X1 g559(.A(new_n744), .B(new_n745), .C1(new_n740), .C2(new_n741), .ZN(new_n746));
  NAND2_X1  g560(.A1(new_n743), .A2(new_n746), .ZN(new_n747));
  NAND2_X1  g561(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n748));
  NAND2_X1  g562(.A1(new_n748), .A2(KEYINPUT83), .ZN(new_n749));
  OR2_X1    g563(.A1(new_n272), .A2(KEYINPUT12), .ZN(new_n750));
  NAND3_X1  g564(.A1(new_n749), .A2(new_n276), .A3(new_n750), .ZN(new_n751));
  NAND2_X1  g565(.A1(new_n751), .A2(new_n261), .ZN(new_n752));
  INV_X1    g566(.A(new_n266), .ZN(new_n753));
  AOI22_X1  g567(.A1(new_n752), .A2(new_n753), .B1(new_n280), .B2(new_n283), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n754), .A2(KEYINPUT45), .ZN(new_n755));
  NAND2_X1  g569(.A1(new_n755), .A2(KEYINPUT104), .ZN(new_n756));
  INV_X1    g570(.A(KEYINPUT104), .ZN(new_n757));
  NAND3_X1  g571(.A1(new_n754), .A2(new_n757), .A3(KEYINPUT45), .ZN(new_n758));
  AND2_X1   g572(.A1(new_n756), .A2(new_n758), .ZN(new_n759));
  OAI21_X1  g573(.A(G469), .B1(new_n754), .B2(KEYINPUT45), .ZN(new_n760));
  OAI211_X1 g574(.A(KEYINPUT46), .B(new_n289), .C1(new_n759), .C2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(KEYINPUT46), .ZN(new_n762));
  AOI21_X1  g576(.A(new_n760), .B1(new_n756), .B2(new_n758), .ZN(new_n763));
  OAI21_X1  g577(.A(new_n762), .B1(new_n763), .B2(new_n288), .ZN(new_n764));
  NAND3_X1  g578(.A1(new_n761), .A2(new_n764), .A3(new_n282), .ZN(new_n765));
  AND2_X1   g579(.A1(new_n765), .A2(new_n679), .ZN(new_n766));
  AOI21_X1  g580(.A(new_n711), .B1(new_n742), .B2(KEYINPUT44), .ZN(new_n767));
  NAND4_X1  g581(.A1(new_n747), .A2(new_n766), .A3(new_n645), .A4(new_n767), .ZN(new_n768));
  XNOR2_X1  g582(.A(new_n768), .B(G137), .ZN(G39));
  NAND2_X1  g583(.A1(new_n765), .A2(new_n679), .ZN(new_n770));
  INV_X1    g584(.A(KEYINPUT109), .ZN(new_n771));
  NOR2_X1   g585(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n772));
  INV_X1    g586(.A(new_n772), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n770), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n771), .A2(KEYINPUT47), .ZN(new_n775));
  OAI211_X1 g589(.A(new_n765), .B(new_n679), .C1(new_n775), .C2(new_n772), .ZN(new_n776));
  NOR4_X1   g590(.A1(new_n554), .A2(new_n587), .A3(new_n711), .A4(new_n664), .ZN(new_n777));
  NAND3_X1  g591(.A1(new_n774), .A2(new_n776), .A3(new_n777), .ZN(new_n778));
  XNOR2_X1  g592(.A(new_n778), .B(G140), .ZN(G42));
  NOR3_X1   g593(.A1(new_n737), .A2(new_n294), .A3(new_n594), .ZN(new_n780));
  NAND4_X1  g594(.A1(new_n587), .A2(new_n733), .A3(new_n734), .A4(new_n780), .ZN(new_n781));
  AOI22_X1  g595(.A1(new_n781), .A2(KEYINPUT110), .B1(new_n671), .B2(KEYINPUT49), .ZN(new_n782));
  OAI21_X1  g596(.A(new_n782), .B1(KEYINPUT110), .B2(new_n781), .ZN(new_n783));
  XNOR2_X1  g597(.A(new_n783), .B(KEYINPUT111), .ZN(new_n784));
  INV_X1    g598(.A(new_n653), .ZN(new_n785));
  OR2_X1    g599(.A1(new_n671), .A2(KEYINPUT49), .ZN(new_n786));
  NAND4_X1  g600(.A1(new_n784), .A2(new_n785), .A3(new_n656), .A4(new_n786), .ZN(new_n787));
  AND4_X1   g601(.A1(new_n282), .A2(new_n712), .A3(new_n376), .A4(new_n670), .ZN(new_n788));
  AND2_X1   g602(.A1(new_n788), .A2(new_n739), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n789), .A2(new_n668), .ZN(new_n790));
  NOR2_X1   g604(.A1(KEYINPUT115), .A2(KEYINPUT48), .ZN(new_n791));
  NAND2_X1  g605(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  XOR2_X1   g606(.A(KEYINPUT115), .B(KEYINPUT48), .Z(new_n793));
  NAND3_X1  g607(.A1(new_n789), .A2(new_n668), .A3(new_n793), .ZN(new_n794));
  AND3_X1   g608(.A1(new_n788), .A2(new_n587), .A3(new_n785), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n795), .A2(new_n663), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n262), .A2(G952), .ZN(new_n797));
  AND3_X1   g611(.A1(new_n697), .A2(new_n376), .A3(new_n739), .ZN(new_n798));
  AOI21_X1  g612(.A(new_n797), .B1(new_n798), .B2(new_n699), .ZN(new_n799));
  NAND4_X1  g613(.A1(new_n792), .A2(new_n794), .A3(new_n796), .A4(new_n799), .ZN(new_n800));
  AND2_X1   g614(.A1(new_n774), .A2(new_n776), .ZN(new_n801));
  NOR2_X1   g615(.A1(new_n671), .A2(new_n295), .ZN(new_n802));
  OAI211_X1 g616(.A(new_n723), .B(new_n798), .C1(new_n801), .C2(new_n802), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n701), .A2(new_n737), .ZN(new_n804));
  INV_X1    g618(.A(new_n804), .ZN(new_n805));
  AND3_X1   g619(.A1(new_n591), .A2(new_n696), .A3(new_n657), .ZN(new_n806));
  AOI22_X1  g620(.A1(new_n795), .A2(new_n805), .B1(new_n789), .B2(new_n806), .ZN(new_n807));
  NOR3_X1   g621(.A1(new_n671), .A2(new_n293), .A3(new_n491), .ZN(new_n808));
  XNOR2_X1  g622(.A(new_n808), .B(KEYINPUT113), .ZN(new_n809));
  NAND3_X1  g623(.A1(new_n809), .A2(new_n656), .A3(new_n798), .ZN(new_n810));
  INV_X1    g624(.A(KEYINPUT50), .ZN(new_n811));
  NAND2_X1  g625(.A1(new_n810), .A2(new_n811), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n809), .A2(KEYINPUT50), .A3(new_n656), .A4(new_n798), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  AND3_X1   g628(.A1(new_n807), .A2(KEYINPUT51), .A3(new_n814), .ZN(new_n815));
  AOI21_X1  g629(.A(new_n800), .B1(new_n803), .B2(new_n815), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n807), .A2(new_n814), .ZN(new_n817));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n817), .A2(new_n818), .ZN(new_n819));
  NAND3_X1  g633(.A1(new_n807), .A2(KEYINPUT114), .A3(new_n814), .ZN(new_n820));
  AND3_X1   g634(.A1(new_n819), .A2(new_n803), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g635(.A(new_n816), .B1(new_n821), .B2(KEYINPUT51), .ZN(new_n822));
  INV_X1    g636(.A(KEYINPUT54), .ZN(new_n823));
  AOI21_X1  g637(.A(new_n636), .B1(new_n610), .B2(KEYINPUT112), .ZN(new_n824));
  OR3_X1    g638(.A1(new_n701), .A2(KEYINPUT112), .A3(new_n737), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n379), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR3_X1   g640(.A1(new_n631), .A2(new_n590), .A3(new_n586), .ZN(new_n827));
  AND3_X1   g641(.A1(new_n374), .A2(new_n491), .A3(new_n493), .ZN(new_n828));
  NAND4_X1  g642(.A1(new_n826), .A2(new_n644), .A3(new_n827), .A4(new_n828), .ZN(new_n829));
  AND4_X1   g643(.A1(new_n588), .A2(new_n633), .A3(new_n705), .A4(new_n829), .ZN(new_n830));
  AND2_X1   g644(.A1(new_n673), .A2(new_n677), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n687), .A2(new_n830), .A3(new_n831), .ZN(new_n832));
  NOR3_X1   g646(.A1(new_n601), .A2(new_n658), .A3(new_n638), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n290), .A2(new_n295), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g648(.A1(new_n684), .A2(new_n834), .A3(new_n630), .ZN(new_n835));
  NAND3_X1  g649(.A1(new_n713), .A2(new_n679), .A3(new_n715), .ZN(new_n836));
  NOR2_X1   g650(.A1(new_n836), .A2(new_n708), .ZN(new_n837));
  OAI21_X1  g651(.A(new_n723), .B1(new_n835), .B2(new_n837), .ZN(new_n838));
  NAND4_X1  g652(.A1(new_n722), .A2(new_n838), .A3(new_n726), .A4(new_n729), .ZN(new_n839));
  NOR2_X1   g653(.A1(new_n832), .A2(new_n839), .ZN(new_n840));
  NAND3_X1  g654(.A1(new_n595), .A2(new_n702), .A3(new_n703), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n626), .A2(new_n679), .A3(new_n639), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n716), .A2(new_n653), .A3(new_n843), .ZN(new_n844));
  INV_X1    g658(.A(new_n709), .ZN(new_n845));
  NAND4_X1  g659(.A1(new_n642), .A2(new_n666), .A3(new_n844), .A4(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n846), .A2(KEYINPUT52), .ZN(new_n847));
  INV_X1    g661(.A(new_n595), .ZN(new_n848));
  NOR3_X1   g662(.A1(new_n684), .A2(new_n848), .A3(new_n630), .ZN(new_n849));
  AOI21_X1  g663(.A(new_n709), .B1(new_n849), .B2(new_n640), .ZN(new_n850));
  INV_X1    g664(.A(KEYINPUT52), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n850), .A2(new_n851), .A3(new_n666), .A4(new_n844), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  AOI21_X1  g667(.A(KEYINPUT53), .B1(new_n840), .B2(new_n853), .ZN(new_n854));
  NAND2_X1  g668(.A1(new_n847), .A2(new_n852), .ZN(new_n855));
  INV_X1    g669(.A(KEYINPUT53), .ZN(new_n856));
  NOR4_X1   g670(.A1(new_n855), .A2(new_n832), .A3(new_n839), .A4(new_n856), .ZN(new_n857));
  OAI21_X1  g671(.A(new_n823), .B1(new_n854), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g672(.A1(new_n722), .A2(new_n726), .A3(new_n729), .ZN(new_n859));
  NAND4_X1  g673(.A1(new_n588), .A2(new_n633), .A3(new_n829), .A4(new_n705), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n673), .A2(new_n677), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n859), .A2(new_n687), .A3(new_n862), .A4(new_n838), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n856), .B1(new_n863), .B2(new_n855), .ZN(new_n864));
  NAND3_X1  g678(.A1(new_n840), .A2(new_n853), .A3(KEYINPUT53), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n864), .A2(KEYINPUT54), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(new_n822), .B1(new_n858), .B2(new_n866), .ZN(new_n867));
  NOR2_X1   g681(.A1(G952), .A2(G953), .ZN(new_n868));
  OAI21_X1  g682(.A(new_n787), .B1(new_n867), .B2(new_n868), .ZN(G75));
  AOI21_X1  g683(.A(new_n188), .B1(new_n864), .B2(new_n865), .ZN(new_n870));
  NAND2_X1  g684(.A1(new_n870), .A2(G210), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n369), .A2(new_n370), .ZN(new_n872));
  XNOR2_X1  g686(.A(new_n872), .B(new_n308), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT55), .ZN(new_n874));
  XOR2_X1   g688(.A(KEYINPUT116), .B(KEYINPUT56), .Z(new_n875));
  AND3_X1   g689(.A1(new_n871), .A2(new_n874), .A3(new_n875), .ZN(new_n876));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n877));
  AOI21_X1  g691(.A(new_n874), .B1(new_n871), .B2(new_n877), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n262), .A2(G952), .ZN(new_n879));
  NOR3_X1   g693(.A1(new_n876), .A2(new_n878), .A3(new_n879), .ZN(G51));
  XNOR2_X1  g694(.A(new_n288), .B(KEYINPUT57), .ZN(new_n881));
  NAND3_X1  g695(.A1(new_n858), .A2(new_n866), .A3(new_n881), .ZN(new_n882));
  INV_X1    g696(.A(KEYINPUT118), .ZN(new_n883));
  XOR2_X1   g697(.A(new_n669), .B(KEYINPUT117), .Z(new_n884));
  NAND3_X1  g698(.A1(new_n882), .A2(new_n883), .A3(new_n884), .ZN(new_n885));
  NAND2_X1  g699(.A1(new_n870), .A2(new_n763), .ZN(new_n886));
  AND2_X1   g700(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  NAND2_X1  g701(.A1(new_n882), .A2(new_n884), .ZN(new_n888));
  NAND2_X1  g702(.A1(new_n888), .A2(KEYINPUT118), .ZN(new_n889));
  AOI21_X1  g703(.A(new_n879), .B1(new_n887), .B2(new_n889), .ZN(G54));
  NAND2_X1  g704(.A1(KEYINPUT58), .A2(G475), .ZN(new_n891));
  XOR2_X1   g705(.A(new_n891), .B(KEYINPUT119), .Z(new_n892));
  AND2_X1   g706(.A1(new_n870), .A2(new_n892), .ZN(new_n893));
  AND2_X1   g707(.A1(new_n893), .A2(new_n598), .ZN(new_n894));
  NOR2_X1   g708(.A1(new_n893), .A2(new_n598), .ZN(new_n895));
  NOR3_X1   g709(.A1(new_n894), .A2(new_n895), .A3(new_n879), .ZN(G60));
  XNOR2_X1  g710(.A(new_n602), .B(KEYINPUT120), .ZN(new_n897));
  XOR2_X1   g711(.A(new_n897), .B(KEYINPUT59), .Z(new_n898));
  NAND3_X1  g712(.A1(new_n858), .A2(new_n866), .A3(new_n898), .ZN(new_n899));
  NAND2_X1  g713(.A1(new_n606), .A2(new_n607), .ZN(new_n900));
  INV_X1    g714(.A(new_n900), .ZN(new_n901));
  AND2_X1   g715(.A1(new_n899), .A2(new_n901), .ZN(new_n902));
  NOR2_X1   g716(.A1(new_n899), .A2(new_n901), .ZN(new_n903));
  NOR3_X1   g717(.A1(new_n902), .A2(new_n903), .A3(new_n879), .ZN(G63));
  NAND2_X1  g718(.A1(G217), .A2(G902), .ZN(new_n905));
  XNOR2_X1  g719(.A(new_n905), .B(KEYINPUT60), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n906), .B1(new_n864), .B2(new_n865), .ZN(new_n907));
  OR2_X1    g721(.A1(new_n907), .A2(new_n577), .ZN(new_n908));
  INV_X1    g722(.A(new_n879), .ZN(new_n909));
  NAND2_X1  g723(.A1(new_n907), .A2(new_n623), .ZN(new_n910));
  NAND3_X1  g724(.A1(new_n908), .A2(new_n909), .A3(new_n910), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT61), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n911), .A2(new_n912), .ZN(new_n913));
  NAND4_X1  g727(.A1(new_n908), .A2(KEYINPUT61), .A3(new_n909), .A4(new_n910), .ZN(new_n914));
  NAND2_X1  g728(.A1(new_n913), .A2(new_n914), .ZN(G66));
  OAI21_X1  g729(.A(G953), .B1(new_n378), .B2(new_n305), .ZN(new_n916));
  INV_X1    g730(.A(new_n832), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n916), .B1(new_n917), .B2(G953), .ZN(new_n918));
  OAI21_X1  g732(.A(new_n872), .B1(G898), .B2(new_n262), .ZN(new_n919));
  XNOR2_X1  g733(.A(new_n918), .B(new_n919), .ZN(G69));
  AOI21_X1  g734(.A(new_n262), .B1(G227), .B2(G900), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n666), .A2(new_n642), .A3(new_n845), .ZN(new_n922));
  XNOR2_X1  g736(.A(new_n922), .B(KEYINPUT122), .ZN(new_n923));
  NAND2_X1  g737(.A1(new_n768), .A2(new_n923), .ZN(new_n924));
  INV_X1    g738(.A(KEYINPUT126), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n924), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n668), .ZN(new_n927));
  NOR2_X1   g741(.A1(new_n927), .A2(new_n841), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n766), .A2(new_n645), .A3(new_n928), .ZN(new_n929));
  AND3_X1   g743(.A1(new_n778), .A2(new_n859), .A3(new_n929), .ZN(new_n930));
  NAND3_X1  g744(.A1(new_n768), .A2(new_n923), .A3(KEYINPUT126), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n926), .A2(new_n930), .A3(new_n262), .A4(new_n931), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n521), .A2(new_n523), .ZN(new_n933));
  XOR2_X1   g747(.A(new_n933), .B(KEYINPUT121), .Z(new_n934));
  XNOR2_X1  g748(.A(new_n934), .B(new_n427), .ZN(new_n935));
  AOI21_X1  g749(.A(new_n935), .B1(G900), .B2(G953), .ZN(new_n936));
  AOI21_X1  g750(.A(KEYINPUT125), .B1(new_n932), .B2(new_n936), .ZN(new_n937));
  INV_X1    g751(.A(new_n935), .ZN(new_n938));
  AND2_X1   g752(.A1(new_n824), .A2(new_n825), .ZN(new_n939));
  NOR4_X1   g753(.A1(new_n927), .A2(new_n646), .A3(new_n939), .A4(new_n711), .ZN(new_n940));
  XNOR2_X1  g754(.A(new_n940), .B(KEYINPUT123), .ZN(new_n941));
  AND3_X1   g755(.A1(new_n768), .A2(new_n778), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g756(.A1(new_n923), .A2(KEYINPUT62), .A3(new_n661), .ZN(new_n943));
  INV_X1    g757(.A(new_n943), .ZN(new_n944));
  AOI21_X1  g758(.A(KEYINPUT62), .B1(new_n923), .B2(new_n661), .ZN(new_n945));
  OAI21_X1  g759(.A(new_n942), .B1(new_n944), .B2(new_n945), .ZN(new_n946));
  AOI21_X1  g760(.A(new_n938), .B1(new_n946), .B2(new_n262), .ZN(new_n947));
  INV_X1    g761(.A(KEYINPUT124), .ZN(new_n948));
  OAI21_X1  g762(.A(new_n937), .B1(new_n947), .B2(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n768), .A2(new_n778), .A3(new_n941), .ZN(new_n950));
  INV_X1    g764(.A(new_n945), .ZN(new_n951));
  AOI21_X1  g765(.A(new_n950), .B1(new_n951), .B2(new_n943), .ZN(new_n952));
  OAI21_X1  g766(.A(new_n935), .B1(new_n952), .B2(G953), .ZN(new_n953));
  NOR2_X1   g767(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n954));
  OAI21_X1  g768(.A(new_n921), .B1(new_n949), .B2(new_n954), .ZN(new_n955));
  NAND2_X1  g769(.A1(new_n953), .A2(KEYINPUT124), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n947), .A2(new_n948), .ZN(new_n957));
  INV_X1    g771(.A(new_n921), .ZN(new_n958));
  NAND4_X1  g772(.A1(new_n956), .A2(new_n957), .A3(new_n958), .A4(new_n937), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n955), .A2(new_n959), .ZN(G72));
  NAND4_X1  g774(.A1(new_n926), .A2(new_n930), .A3(new_n917), .A4(new_n931), .ZN(new_n961));
  NAND2_X1  g775(.A1(G472), .A2(G902), .ZN(new_n962));
  XOR2_X1   g776(.A(new_n962), .B(KEYINPUT63), .Z(new_n963));
  XOR2_X1   g777(.A(new_n963), .B(KEYINPUT127), .Z(new_n964));
  AOI211_X1 g778(.A(new_n500), .B(new_n539), .C1(new_n961), .C2(new_n964), .ZN(new_n965));
  NAND2_X1  g779(.A1(new_n539), .A2(new_n500), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n952), .A2(new_n917), .ZN(new_n967));
  AOI21_X1  g781(.A(new_n966), .B1(new_n967), .B2(new_n964), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n539), .A2(new_n501), .ZN(new_n969));
  NAND2_X1  g783(.A1(new_n648), .A2(new_n969), .ZN(new_n970));
  OAI211_X1 g784(.A(new_n963), .B(new_n970), .C1(new_n854), .C2(new_n857), .ZN(new_n971));
  NAND2_X1  g785(.A1(new_n971), .A2(new_n909), .ZN(new_n972));
  NOR3_X1   g786(.A1(new_n965), .A2(new_n968), .A3(new_n972), .ZN(G57));
endmodule


