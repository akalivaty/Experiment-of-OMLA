//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 1 1 0 1 1 1 0 1 1 1 0 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 1 0 0 1 0 1 0 1 1 0 0 1 1 0 0 0 0 0 1 0 1 1 1 1 1 1 1 1 1 0 0 1 1 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:15 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n436, new_n441, new_n448, new_n452, new_n453, new_n454, new_n455,
    new_n456, new_n459, new_n460, new_n461, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n539, new_n540, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n550,
    new_n552, new_n553, new_n555, new_n556, new_n557, new_n558, new_n559,
    new_n560, new_n561, new_n562, new_n563, new_n567, new_n568, new_n569,
    new_n571, new_n572, new_n573, new_n574, new_n575, new_n576, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n602,
    new_n603, new_n604, new_n605, new_n608, new_n610, new_n611, new_n612,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n641, new_n642, new_n643, new_n644,
    new_n645, new_n646, new_n647, new_n648, new_n649, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n657, new_n658, new_n659,
    new_n660, new_n661, new_n662, new_n663, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n814, new_n815,
    new_n817, new_n818, new_n819, new_n820, new_n821, new_n822, new_n823,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n842, new_n843, new_n844, new_n845,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n911, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n955, new_n956, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1165, new_n1166,
    new_n1167, new_n1168, new_n1169, new_n1170, new_n1171, new_n1172,
    new_n1174, new_n1175, new_n1176;
  BUF_X1    g000(.A(G452), .Z(G350));
  XNOR2_X1  g001(.A(KEYINPUT64), .B(G452), .ZN(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  XOR2_X1   g005(.A(KEYINPUT65), .B(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XOR2_X1   g010(.A(KEYINPUT0), .B(G82), .Z(new_n436));
  INV_X1    g011(.A(new_n436), .ZN(G220));
  INV_X1    g012(.A(G96), .ZN(G221));
  INV_X1    g013(.A(G69), .ZN(G235));
  INV_X1    g014(.A(G120), .ZN(G236));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G57), .ZN(new_n441));
  INV_X1    g016(.A(new_n441), .ZN(G237));
  INV_X1    g017(.A(G108), .ZN(G238));
  NAND4_X1  g018(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g019(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g020(.A(G452), .Z(G391));
  AND2_X1   g021(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g022(.A1(G7), .A2(G661), .ZN(new_n448));
  XOR2_X1   g023(.A(new_n448), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g024(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g025(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NAND4_X1  g026(.A1(new_n436), .A2(G44), .A3(G96), .A4(G132), .ZN(new_n452));
  XNOR2_X1  g027(.A(new_n452), .B(KEYINPUT2), .ZN(new_n453));
  NAND4_X1  g028(.A1(new_n441), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n454));
  XNOR2_X1  g029(.A(KEYINPUT67), .B(KEYINPUT68), .ZN(new_n455));
  XNOR2_X1  g030(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NOR2_X1   g031(.A1(new_n453), .A2(new_n456), .ZN(G325));
  INV_X1    g032(.A(G325), .ZN(G261));
  NAND2_X1  g033(.A1(new_n453), .A2(G2106), .ZN(new_n459));
  NAND2_X1  g034(.A1(new_n456), .A2(G567), .ZN(new_n460));
  NAND2_X1  g035(.A1(new_n459), .A2(new_n460), .ZN(new_n461));
  INV_X1    g036(.A(new_n461), .ZN(G319));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  INV_X1    g038(.A(G2104), .ZN(new_n464));
  NAND2_X1  g039(.A1(new_n464), .A2(KEYINPUT3), .ZN(new_n465));
  INV_X1    g040(.A(KEYINPUT3), .ZN(new_n466));
  NAND2_X1  g041(.A1(new_n466), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n465), .A2(new_n467), .ZN(new_n468));
  INV_X1    g043(.A(G125), .ZN(new_n469));
  OAI21_X1  g044(.A(new_n463), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n470), .A2(G2105), .ZN(new_n471));
  INV_X1    g046(.A(G2105), .ZN(new_n472));
  NAND3_X1  g047(.A1(new_n472), .A2(G101), .A3(G2104), .ZN(new_n473));
  XOR2_X1   g048(.A(new_n473), .B(KEYINPUT69), .Z(new_n474));
  NOR2_X1   g049(.A1(new_n468), .A2(G2105), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n475), .A2(G137), .ZN(new_n476));
  NAND3_X1  g051(.A1(new_n471), .A2(new_n474), .A3(new_n476), .ZN(new_n477));
  INV_X1    g052(.A(new_n477), .ZN(G160));
  NOR2_X1   g053(.A1(new_n468), .A2(new_n472), .ZN(new_n479));
  NAND2_X1  g054(.A1(new_n479), .A2(G124), .ZN(new_n480));
  NAND2_X1  g055(.A1(new_n475), .A2(G136), .ZN(new_n481));
  OR2_X1    g056(.A1(G100), .A2(G2105), .ZN(new_n482));
  OAI211_X1 g057(.A(new_n482), .B(G2104), .C1(G112), .C2(new_n472), .ZN(new_n483));
  NAND3_X1  g058(.A1(new_n480), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  INV_X1    g059(.A(new_n484), .ZN(G162));
  NAND4_X1  g060(.A1(new_n465), .A2(new_n467), .A3(G138), .A4(new_n472), .ZN(new_n486));
  INV_X1    g061(.A(KEYINPUT4), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n486), .A2(new_n487), .ZN(new_n488));
  XNOR2_X1  g063(.A(KEYINPUT3), .B(G2104), .ZN(new_n489));
  NAND4_X1  g064(.A1(new_n489), .A2(KEYINPUT4), .A3(G138), .A4(new_n472), .ZN(new_n490));
  AND2_X1   g065(.A1(new_n488), .A2(new_n490), .ZN(new_n491));
  NAND3_X1  g066(.A1(new_n465), .A2(new_n467), .A3(G126), .ZN(new_n492));
  NAND2_X1  g067(.A1(G114), .A2(G2104), .ZN(new_n493));
  NAND2_X1  g068(.A1(new_n492), .A2(new_n493), .ZN(new_n494));
  NOR2_X1   g069(.A1(new_n464), .A2(G2105), .ZN(new_n495));
  AOI22_X1  g070(.A1(new_n494), .A2(G2105), .B1(G102), .B2(new_n495), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n491), .A2(new_n496), .ZN(new_n497));
  INV_X1    g072(.A(new_n497), .ZN(G164));
  INV_X1    g073(.A(KEYINPUT6), .ZN(new_n499));
  OAI21_X1  g074(.A(KEYINPUT70), .B1(new_n499), .B2(G651), .ZN(new_n500));
  INV_X1    g075(.A(KEYINPUT70), .ZN(new_n501));
  INV_X1    g076(.A(G651), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n501), .A2(new_n502), .A3(KEYINPUT6), .ZN(new_n503));
  AOI22_X1  g078(.A1(new_n500), .A2(new_n503), .B1(new_n499), .B2(G651), .ZN(new_n504));
  AOI22_X1  g079(.A1(new_n504), .A2(G50), .B1(G75), .B2(G651), .ZN(new_n505));
  INV_X1    g080(.A(G543), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n506), .A2(KEYINPUT5), .ZN(new_n508));
  INV_X1    g083(.A(KEYINPUT5), .ZN(new_n509));
  NAND2_X1  g084(.A1(new_n509), .A2(G543), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  XNOR2_X1  g086(.A(KEYINPUT71), .B(G88), .ZN(new_n512));
  NAND2_X1  g087(.A1(new_n504), .A2(new_n512), .ZN(new_n513));
  NAND2_X1  g088(.A1(G62), .A2(G651), .ZN(new_n514));
  AOI21_X1  g089(.A(new_n511), .B1(new_n513), .B2(new_n514), .ZN(new_n515));
  NOR2_X1   g090(.A1(new_n507), .A2(new_n515), .ZN(G166));
  XNOR2_X1  g091(.A(KEYINPUT5), .B(G543), .ZN(new_n517));
  NAND3_X1  g092(.A1(new_n517), .A2(G63), .A3(G651), .ZN(new_n518));
  AND3_X1   g093(.A1(new_n504), .A2(G51), .A3(G543), .ZN(new_n519));
  INV_X1    g094(.A(new_n519), .ZN(new_n520));
  NAND3_X1  g095(.A1(new_n504), .A2(G89), .A3(new_n517), .ZN(new_n521));
  NAND3_X1  g096(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n522));
  XNOR2_X1  g097(.A(new_n522), .B(KEYINPUT7), .ZN(new_n523));
  AND3_X1   g098(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n523), .ZN(new_n524));
  AOI21_X1  g099(.A(KEYINPUT72), .B1(new_n521), .B2(new_n523), .ZN(new_n525));
  OAI211_X1 g100(.A(new_n518), .B(new_n520), .C1(new_n524), .C2(new_n525), .ZN(G286));
  INV_X1    g101(.A(G286), .ZN(G168));
  NAND2_X1  g102(.A1(new_n500), .A2(new_n503), .ZN(new_n528));
  NAND2_X1  g103(.A1(new_n499), .A2(G651), .ZN(new_n529));
  NAND2_X1  g104(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NOR2_X1   g105(.A1(new_n530), .A2(new_n511), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n531), .A2(G90), .ZN(new_n532));
  NOR2_X1   g107(.A1(new_n530), .A2(new_n506), .ZN(new_n533));
  XOR2_X1   g108(.A(KEYINPUT73), .B(G52), .Z(new_n534));
  NAND2_X1  g109(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI22_X1  g110(.A1(new_n517), .A2(G64), .B1(G77), .B2(G543), .ZN(new_n536));
  OR2_X1    g111(.A1(new_n536), .A2(new_n502), .ZN(new_n537));
  AND3_X1   g112(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(G171));
  INV_X1    g113(.A(G56), .ZN(new_n539));
  INV_X1    g114(.A(G68), .ZN(new_n540));
  OAI22_X1  g115(.A1(new_n511), .A2(new_n539), .B1(new_n540), .B2(new_n506), .ZN(new_n541));
  INV_X1    g116(.A(KEYINPUT74), .ZN(new_n542));
  NAND2_X1  g117(.A1(new_n541), .A2(new_n542), .ZN(new_n543));
  OAI221_X1 g118(.A(KEYINPUT74), .B1(new_n540), .B2(new_n506), .C1(new_n511), .C2(new_n539), .ZN(new_n544));
  NAND3_X1  g119(.A1(new_n543), .A2(G651), .A3(new_n544), .ZN(new_n545));
  NAND2_X1  g120(.A1(new_n533), .A2(G43), .ZN(new_n546));
  NAND2_X1  g121(.A1(new_n531), .A2(G81), .ZN(new_n547));
  AND3_X1   g122(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n548));
  NAND2_X1  g123(.A1(new_n548), .A2(G860), .ZN(G153));
  AND3_X1   g124(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n550));
  NAND2_X1  g125(.A1(new_n550), .A2(G36), .ZN(G176));
  NAND2_X1  g126(.A1(G1), .A2(G3), .ZN(new_n552));
  XNOR2_X1  g127(.A(new_n552), .B(KEYINPUT8), .ZN(new_n553));
  NAND2_X1  g128(.A1(new_n550), .A2(new_n553), .ZN(G188));
  AND2_X1   g129(.A1(new_n517), .A2(G65), .ZN(new_n555));
  NAND2_X1  g130(.A1(G78), .A2(G543), .ZN(new_n556));
  XOR2_X1   g131(.A(new_n556), .B(KEYINPUT75), .Z(new_n557));
  OAI21_X1  g132(.A(G651), .B1(new_n555), .B2(new_n557), .ZN(new_n558));
  NAND4_X1  g133(.A1(new_n528), .A2(G53), .A3(G543), .A4(new_n529), .ZN(new_n559));
  INV_X1    g134(.A(KEYINPUT9), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n559), .A2(new_n560), .ZN(new_n561));
  NAND4_X1  g136(.A1(new_n504), .A2(KEYINPUT9), .A3(G53), .A4(G543), .ZN(new_n562));
  NAND3_X1  g137(.A1(new_n504), .A2(G91), .A3(new_n517), .ZN(new_n563));
  NAND4_X1  g138(.A1(new_n558), .A2(new_n561), .A3(new_n562), .A4(new_n563), .ZN(G299));
  NAND3_X1  g139(.A1(new_n532), .A2(new_n535), .A3(new_n537), .ZN(G301));
  OR2_X1    g140(.A1(new_n507), .A2(new_n515), .ZN(G303));
  NAND2_X1  g141(.A1(new_n533), .A2(G49), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n531), .A2(G87), .ZN(new_n568));
  OAI21_X1  g143(.A(G651), .B1(new_n517), .B2(G74), .ZN(new_n569));
  NAND3_X1  g144(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(G288));
  NAND2_X1  g145(.A1(G73), .A2(G543), .ZN(new_n571));
  INV_X1    g146(.A(G61), .ZN(new_n572));
  OAI21_X1  g147(.A(new_n571), .B1(new_n511), .B2(new_n572), .ZN(new_n573));
  NAND2_X1  g148(.A1(new_n573), .A2(G651), .ZN(new_n574));
  NAND3_X1  g149(.A1(new_n504), .A2(G86), .A3(new_n517), .ZN(new_n575));
  NAND3_X1  g150(.A1(new_n504), .A2(G48), .A3(G543), .ZN(new_n576));
  NAND3_X1  g151(.A1(new_n574), .A2(new_n575), .A3(new_n576), .ZN(G305));
  NAND2_X1  g152(.A1(new_n531), .A2(G85), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n533), .A2(G47), .ZN(new_n579));
  AOI22_X1  g154(.A1(new_n517), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n580));
  OR2_X1    g155(.A1(new_n580), .A2(new_n502), .ZN(new_n581));
  NAND3_X1  g156(.A1(new_n578), .A2(new_n579), .A3(new_n581), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n582), .A2(KEYINPUT76), .ZN(new_n583));
  INV_X1    g158(.A(KEYINPUT76), .ZN(new_n584));
  NAND4_X1  g159(.A1(new_n578), .A2(new_n579), .A3(new_n584), .A4(new_n581), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n583), .A2(new_n585), .ZN(G290));
  NAND2_X1  g161(.A1(G301), .A2(G868), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n504), .A2(G92), .A3(new_n517), .ZN(new_n588));
  INV_X1    g163(.A(KEYINPUT10), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NAND4_X1  g165(.A1(new_n504), .A2(KEYINPUT10), .A3(G92), .A4(new_n517), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n590), .A2(new_n591), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n533), .A2(G54), .ZN(new_n593));
  NAND2_X1  g168(.A1(G79), .A2(G543), .ZN(new_n594));
  INV_X1    g169(.A(G66), .ZN(new_n595));
  OAI21_X1  g170(.A(new_n594), .B1(new_n511), .B2(new_n595), .ZN(new_n596));
  NAND2_X1  g171(.A1(new_n596), .A2(G651), .ZN(new_n597));
  NAND3_X1  g172(.A1(new_n592), .A2(new_n593), .A3(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(new_n599));
  OAI21_X1  g174(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G284));
  OAI21_X1  g175(.A(new_n587), .B1(new_n599), .B2(G868), .ZN(G321));
  INV_X1    g176(.A(G868), .ZN(new_n602));
  OR3_X1    g177(.A1(G168), .A2(KEYINPUT77), .A3(new_n602), .ZN(new_n603));
  OAI21_X1  g178(.A(KEYINPUT77), .B1(G168), .B2(new_n602), .ZN(new_n604));
  INV_X1    g179(.A(G299), .ZN(new_n605));
  OAI211_X1 g180(.A(new_n603), .B(new_n604), .C1(G868), .C2(new_n605), .ZN(G297));
  XNOR2_X1  g181(.A(G297), .B(KEYINPUT78), .ZN(G280));
  INV_X1    g182(.A(G559), .ZN(new_n608));
  OAI21_X1  g183(.A(new_n599), .B1(new_n608), .B2(G860), .ZN(G148));
  NAND3_X1  g184(.A1(new_n545), .A2(new_n546), .A3(new_n547), .ZN(new_n610));
  NAND2_X1  g185(.A1(new_n610), .A2(new_n602), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n598), .A2(G559), .ZN(new_n612));
  OAI21_X1  g187(.A(new_n611), .B1(new_n612), .B2(new_n602), .ZN(G323));
  XNOR2_X1  g188(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g189(.A1(new_n479), .A2(G123), .ZN(new_n615));
  XOR2_X1   g190(.A(new_n615), .B(KEYINPUT79), .Z(new_n616));
  OR2_X1    g191(.A1(G99), .A2(G2105), .ZN(new_n617));
  OAI211_X1 g192(.A(new_n617), .B(G2104), .C1(G111), .C2(new_n472), .ZN(new_n618));
  NAND2_X1  g193(.A1(new_n475), .A2(G135), .ZN(new_n619));
  NAND3_X1  g194(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  XOR2_X1   g195(.A(new_n620), .B(G2096), .Z(new_n621));
  NAND2_X1  g196(.A1(new_n489), .A2(new_n495), .ZN(new_n622));
  XNOR2_X1  g197(.A(new_n622), .B(KEYINPUT12), .ZN(new_n623));
  XNOR2_X1  g198(.A(new_n623), .B(KEYINPUT13), .ZN(new_n624));
  XNOR2_X1  g199(.A(new_n624), .B(G2100), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n621), .A2(new_n625), .ZN(G156));
  XNOR2_X1  g201(.A(G2451), .B(G2454), .ZN(new_n627));
  XNOR2_X1  g202(.A(new_n627), .B(KEYINPUT16), .ZN(new_n628));
  XOR2_X1   g203(.A(G2443), .B(G2446), .Z(new_n629));
  XNOR2_X1  g204(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g205(.A(G1341), .B(G1348), .ZN(new_n631));
  XNOR2_X1  g206(.A(new_n630), .B(new_n631), .ZN(new_n632));
  XOR2_X1   g207(.A(KEYINPUT15), .B(G2435), .Z(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(G2438), .ZN(new_n634));
  XOR2_X1   g209(.A(G2427), .B(G2430), .Z(new_n635));
  XNOR2_X1  g210(.A(new_n635), .B(KEYINPUT80), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n634), .B(new_n636), .ZN(new_n637));
  NAND2_X1  g212(.A1(new_n637), .A2(KEYINPUT14), .ZN(new_n638));
  XNOR2_X1  g213(.A(new_n632), .B(new_n638), .ZN(new_n639));
  AND2_X1   g214(.A1(new_n639), .A2(G14), .ZN(G401));
  XOR2_X1   g215(.A(G2084), .B(G2090), .Z(new_n641));
  INV_X1    g216(.A(new_n641), .ZN(new_n642));
  XOR2_X1   g217(.A(G2067), .B(G2678), .Z(new_n643));
  INV_X1    g218(.A(new_n643), .ZN(new_n644));
  XNOR2_X1  g219(.A(G2072), .B(G2078), .ZN(new_n645));
  OR2_X1    g220(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(new_n645), .B(KEYINPUT17), .Z(new_n647));
  OAI211_X1 g222(.A(new_n642), .B(new_n646), .C1(new_n647), .C2(new_n643), .ZN(new_n648));
  XNOR2_X1  g223(.A(new_n648), .B(KEYINPUT81), .ZN(new_n649));
  NAND3_X1  g224(.A1(new_n647), .A2(new_n641), .A3(new_n643), .ZN(new_n650));
  XNOR2_X1  g225(.A(new_n650), .B(KEYINPUT82), .ZN(new_n651));
  NAND3_X1  g226(.A1(new_n644), .A2(new_n641), .A3(new_n645), .ZN(new_n652));
  XOR2_X1   g227(.A(new_n652), .B(KEYINPUT18), .Z(new_n653));
  NAND3_X1  g228(.A1(new_n649), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  XOR2_X1   g229(.A(G2096), .B(G2100), .Z(new_n655));
  XNOR2_X1  g230(.A(new_n654), .B(new_n655), .ZN(G227));
  XNOR2_X1  g231(.A(G1971), .B(G1976), .ZN(new_n657));
  XNOR2_X1  g232(.A(KEYINPUT83), .B(KEYINPUT19), .ZN(new_n658));
  XNOR2_X1  g233(.A(new_n657), .B(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(G1956), .B(G2474), .ZN(new_n660));
  XNOR2_X1  g235(.A(G1961), .B(G1966), .ZN(new_n661));
  NOR3_X1   g236(.A1(new_n659), .A2(new_n660), .A3(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(KEYINPUT20), .ZN(new_n663));
  XNOR2_X1  g238(.A(new_n662), .B(new_n663), .ZN(new_n664));
  AND2_X1   g239(.A1(new_n660), .A2(new_n661), .ZN(new_n665));
  NOR2_X1   g240(.A1(new_n660), .A2(new_n661), .ZN(new_n666));
  AOI21_X1  g241(.A(new_n665), .B1(new_n659), .B2(new_n666), .ZN(new_n667));
  NAND2_X1  g242(.A1(new_n659), .A2(KEYINPUT84), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n667), .B(new_n668), .ZN(new_n669));
  NAND2_X1  g244(.A1(new_n664), .A2(new_n669), .ZN(new_n670));
  XNOR2_X1  g245(.A(new_n670), .B(KEYINPUT21), .ZN(new_n671));
  NAND2_X1  g246(.A1(new_n671), .A2(G1996), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT21), .ZN(new_n673));
  XNOR2_X1  g248(.A(new_n670), .B(new_n673), .ZN(new_n674));
  INV_X1    g249(.A(G1996), .ZN(new_n675));
  NAND2_X1  g250(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(G1981), .B(G1986), .Z(new_n677));
  XNOR2_X1  g252(.A(new_n677), .B(G1991), .ZN(new_n678));
  XNOR2_X1  g253(.A(KEYINPUT85), .B(KEYINPUT86), .ZN(new_n679));
  XNOR2_X1  g254(.A(new_n679), .B(KEYINPUT22), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n678), .B(new_n680), .ZN(new_n681));
  AND3_X1   g256(.A1(new_n672), .A2(new_n676), .A3(new_n681), .ZN(new_n682));
  AOI21_X1  g257(.A(new_n681), .B1(new_n672), .B2(new_n676), .ZN(new_n683));
  NOR2_X1   g258(.A1(new_n682), .A2(new_n683), .ZN(G229));
  NAND2_X1  g259(.A1(G168), .A2(G16), .ZN(new_n685));
  OAI21_X1  g260(.A(new_n685), .B1(G16), .B2(G21), .ZN(new_n686));
  INV_X1    g261(.A(G1966), .ZN(new_n687));
  NAND2_X1  g262(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g263(.A(new_n688), .B(KEYINPUT97), .ZN(new_n689));
  INV_X1    g264(.A(G29), .ZN(new_n690));
  NAND2_X1  g265(.A1(new_n690), .A2(G26), .ZN(new_n691));
  XNOR2_X1  g266(.A(new_n691), .B(KEYINPUT28), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n479), .A2(G128), .ZN(new_n693));
  NAND2_X1  g268(.A1(new_n475), .A2(G140), .ZN(new_n694));
  NOR2_X1   g269(.A1(G104), .A2(G2105), .ZN(new_n695));
  OAI21_X1  g270(.A(G2104), .B1(new_n472), .B2(G116), .ZN(new_n696));
  OAI211_X1 g271(.A(new_n693), .B(new_n694), .C1(new_n695), .C2(new_n696), .ZN(new_n697));
  AND3_X1   g272(.A1(new_n697), .A2(KEYINPUT92), .A3(G29), .ZN(new_n698));
  AOI21_X1  g273(.A(KEYINPUT92), .B1(new_n697), .B2(G29), .ZN(new_n699));
  OAI21_X1  g274(.A(new_n692), .B1(new_n698), .B2(new_n699), .ZN(new_n700));
  XNOR2_X1  g275(.A(new_n700), .B(G2067), .ZN(new_n701));
  NAND2_X1  g276(.A1(new_n479), .A2(G129), .ZN(new_n702));
  NAND2_X1  g277(.A1(new_n475), .A2(G141), .ZN(new_n703));
  NAND2_X1  g278(.A1(new_n495), .A2(G105), .ZN(new_n704));
  NAND3_X1  g279(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n705));
  XOR2_X1   g280(.A(new_n705), .B(KEYINPUT26), .Z(new_n706));
  NAND4_X1  g281(.A1(new_n702), .A2(new_n703), .A3(new_n704), .A4(new_n706), .ZN(new_n707));
  INV_X1    g282(.A(new_n707), .ZN(new_n708));
  NAND2_X1  g283(.A1(new_n708), .A2(G29), .ZN(new_n709));
  OAI21_X1  g284(.A(new_n709), .B1(G29), .B2(G32), .ZN(new_n710));
  XNOR2_X1  g285(.A(KEYINPUT27), .B(G1996), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  INV_X1    g287(.A(G28), .ZN(new_n713));
  OR2_X1    g288(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n714));
  NAND2_X1  g289(.A1(new_n713), .A2(KEYINPUT30), .ZN(new_n715));
  NAND3_X1  g290(.A1(new_n714), .A2(new_n715), .A3(new_n690), .ZN(new_n716));
  OAI211_X1 g291(.A(new_n712), .B(new_n716), .C1(new_n690), .C2(new_n620), .ZN(new_n717));
  XOR2_X1   g292(.A(KEYINPUT31), .B(G11), .Z(new_n718));
  XNOR2_X1  g293(.A(new_n718), .B(KEYINPUT96), .ZN(new_n719));
  OR2_X1    g294(.A1(G29), .A2(G33), .ZN(new_n720));
  NAND2_X1  g295(.A1(new_n495), .A2(G103), .ZN(new_n721));
  XOR2_X1   g296(.A(new_n721), .B(KEYINPUT25), .Z(new_n722));
  NAND2_X1  g297(.A1(new_n475), .A2(G139), .ZN(new_n723));
  AOI22_X1  g298(.A1(new_n489), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n724));
  OAI211_X1 g299(.A(new_n722), .B(new_n723), .C1(new_n472), .C2(new_n724), .ZN(new_n725));
  OAI21_X1  g300(.A(new_n720), .B1(new_n725), .B2(new_n690), .ZN(new_n726));
  INV_X1    g301(.A(G2072), .ZN(new_n727));
  NOR2_X1   g302(.A1(new_n726), .A2(new_n727), .ZN(new_n728));
  OR4_X1    g303(.A1(new_n701), .A2(new_n717), .A3(new_n719), .A4(new_n728), .ZN(new_n729));
  NAND2_X1  g304(.A1(new_n690), .A2(G27), .ZN(new_n730));
  OAI21_X1  g305(.A(new_n730), .B1(G164), .B2(new_n690), .ZN(new_n731));
  XNOR2_X1  g306(.A(new_n731), .B(G2078), .ZN(new_n732));
  INV_X1    g307(.A(G16), .ZN(new_n733));
  NAND2_X1  g308(.A1(new_n733), .A2(G19), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(new_n548), .B2(new_n733), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT91), .B(G1341), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  INV_X1    g312(.A(G1961), .ZN(new_n738));
  NAND2_X1  g313(.A1(G171), .A2(G16), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G5), .B2(G16), .ZN(new_n740));
  INV_X1    g315(.A(G2084), .ZN(new_n741));
  INV_X1    g316(.A(KEYINPUT24), .ZN(new_n742));
  OAI21_X1  g317(.A(new_n690), .B1(new_n742), .B2(G34), .ZN(new_n743));
  INV_X1    g318(.A(KEYINPUT94), .ZN(new_n744));
  OR2_X1    g319(.A1(new_n743), .A2(new_n744), .ZN(new_n745));
  NAND2_X1  g320(.A1(new_n742), .A2(G34), .ZN(new_n746));
  NAND2_X1  g321(.A1(new_n743), .A2(new_n744), .ZN(new_n747));
  NAND3_X1  g322(.A1(new_n745), .A2(new_n746), .A3(new_n747), .ZN(new_n748));
  OAI21_X1  g323(.A(new_n748), .B1(new_n477), .B2(new_n690), .ZN(new_n749));
  XOR2_X1   g324(.A(new_n749), .B(KEYINPUT95), .Z(new_n750));
  OAI221_X1 g325(.A(new_n737), .B1(new_n738), .B2(new_n740), .C1(new_n741), .C2(new_n750), .ZN(new_n751));
  NOR3_X1   g326(.A1(new_n729), .A2(new_n732), .A3(new_n751), .ZN(new_n752));
  NAND2_X1  g327(.A1(new_n750), .A2(new_n741), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n740), .A2(new_n738), .ZN(new_n754));
  OAI211_X1 g329(.A(new_n753), .B(new_n754), .C1(new_n710), .C2(new_n711), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT98), .Z(new_n756));
  NOR2_X1   g331(.A1(G4), .A2(G16), .ZN(new_n757));
  AOI21_X1  g332(.A(new_n757), .B1(new_n599), .B2(G16), .ZN(new_n758));
  XNOR2_X1  g333(.A(KEYINPUT90), .B(G1348), .ZN(new_n759));
  INV_X1    g334(.A(new_n759), .ZN(new_n760));
  XNOR2_X1  g335(.A(new_n758), .B(new_n760), .ZN(new_n761));
  NAND2_X1  g336(.A1(new_n690), .A2(G35), .ZN(new_n762));
  OAI21_X1  g337(.A(new_n762), .B1(G162), .B2(new_n690), .ZN(new_n763));
  XNOR2_X1  g338(.A(new_n763), .B(KEYINPUT29), .ZN(new_n764));
  INV_X1    g339(.A(G2090), .ZN(new_n765));
  XNOR2_X1  g340(.A(new_n764), .B(new_n765), .ZN(new_n766));
  OAI21_X1  g341(.A(new_n766), .B1(new_n687), .B2(new_n686), .ZN(new_n767));
  XNOR2_X1  g342(.A(KEYINPUT99), .B(KEYINPUT23), .ZN(new_n768));
  NAND2_X1  g343(.A1(new_n733), .A2(G20), .ZN(new_n769));
  XNOR2_X1  g344(.A(new_n768), .B(new_n769), .ZN(new_n770));
  AOI21_X1  g345(.A(new_n770), .B1(G299), .B2(G16), .ZN(new_n771));
  XOR2_X1   g346(.A(new_n771), .B(G1956), .Z(new_n772));
  NAND2_X1  g347(.A1(new_n726), .A2(new_n727), .ZN(new_n773));
  XOR2_X1   g348(.A(new_n773), .B(KEYINPUT93), .Z(new_n774));
  NOR3_X1   g349(.A1(new_n767), .A2(new_n772), .A3(new_n774), .ZN(new_n775));
  NAND4_X1  g350(.A1(new_n752), .A2(new_n756), .A3(new_n761), .A4(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n733), .A2(G23), .ZN(new_n777));
  AND3_X1   g352(.A1(new_n567), .A2(new_n568), .A3(new_n569), .ZN(new_n778));
  OAI21_X1  g353(.A(new_n777), .B1(new_n778), .B2(new_n733), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT88), .ZN(new_n780));
  XOR2_X1   g355(.A(KEYINPUT33), .B(G1976), .Z(new_n781));
  XNOR2_X1  g356(.A(new_n780), .B(new_n781), .ZN(new_n782));
  NAND2_X1  g357(.A1(new_n733), .A2(G22), .ZN(new_n783));
  OAI21_X1  g358(.A(new_n783), .B1(G166), .B2(new_n733), .ZN(new_n784));
  MUX2_X1   g359(.A(new_n783), .B(new_n784), .S(KEYINPUT89), .Z(new_n785));
  INV_X1    g360(.A(G1971), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n785), .B(new_n786), .ZN(new_n787));
  NAND2_X1  g362(.A1(new_n733), .A2(G6), .ZN(new_n788));
  INV_X1    g363(.A(G305), .ZN(new_n789));
  OAI21_X1  g364(.A(new_n788), .B1(new_n789), .B2(new_n733), .ZN(new_n790));
  XOR2_X1   g365(.A(KEYINPUT32), .B(G1981), .Z(new_n791));
  XNOR2_X1  g366(.A(new_n790), .B(new_n791), .ZN(new_n792));
  NAND3_X1  g367(.A1(new_n782), .A2(new_n787), .A3(new_n792), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT34), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n690), .A2(G25), .ZN(new_n795));
  NAND2_X1  g370(.A1(new_n479), .A2(G119), .ZN(new_n796));
  NAND2_X1  g371(.A1(new_n475), .A2(G131), .ZN(new_n797));
  OR2_X1    g372(.A1(G95), .A2(G2105), .ZN(new_n798));
  OAI211_X1 g373(.A(new_n798), .B(G2104), .C1(G107), .C2(new_n472), .ZN(new_n799));
  NAND3_X1  g374(.A1(new_n796), .A2(new_n797), .A3(new_n799), .ZN(new_n800));
  INV_X1    g375(.A(new_n800), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n795), .B1(new_n801), .B2(new_n690), .ZN(new_n802));
  XNOR2_X1  g377(.A(KEYINPUT35), .B(G1991), .ZN(new_n803));
  XNOR2_X1  g378(.A(new_n803), .B(KEYINPUT87), .ZN(new_n804));
  XNOR2_X1  g379(.A(new_n802), .B(new_n804), .ZN(new_n805));
  MUX2_X1   g380(.A(G24), .B(G290), .S(G16), .Z(new_n806));
  XNOR2_X1  g381(.A(new_n806), .B(G1986), .ZN(new_n807));
  AOI21_X1  g382(.A(new_n807), .B1(new_n793), .B2(KEYINPUT34), .ZN(new_n808));
  NAND3_X1  g383(.A1(new_n794), .A2(new_n805), .A3(new_n808), .ZN(new_n809));
  NAND2_X1  g384(.A1(new_n809), .A2(KEYINPUT36), .ZN(new_n810));
  INV_X1    g385(.A(KEYINPUT36), .ZN(new_n811));
  NAND4_X1  g386(.A1(new_n794), .A2(new_n808), .A3(new_n811), .A4(new_n805), .ZN(new_n812));
  AOI211_X1 g387(.A(new_n689), .B(new_n776), .C1(new_n810), .C2(new_n812), .ZN(G311));
  AOI21_X1  g388(.A(new_n776), .B1(new_n810), .B2(new_n812), .ZN(new_n814));
  INV_X1    g389(.A(new_n689), .ZN(new_n815));
  NAND2_X1  g390(.A1(new_n814), .A2(new_n815), .ZN(G150));
  NAND3_X1  g391(.A1(new_n508), .A2(new_n510), .A3(G67), .ZN(new_n817));
  NAND2_X1  g392(.A1(G80), .A2(G543), .ZN(new_n818));
  NAND3_X1  g393(.A1(new_n817), .A2(KEYINPUT100), .A3(new_n818), .ZN(new_n819));
  INV_X1    g394(.A(new_n819), .ZN(new_n820));
  AOI21_X1  g395(.A(KEYINPUT100), .B1(new_n817), .B2(new_n818), .ZN(new_n821));
  NOR3_X1   g396(.A1(new_n820), .A2(new_n821), .A3(new_n502), .ZN(new_n822));
  NAND3_X1  g397(.A1(new_n504), .A2(G55), .A3(G543), .ZN(new_n823));
  NAND3_X1  g398(.A1(new_n504), .A2(G93), .A3(new_n517), .ZN(new_n824));
  NAND2_X1  g399(.A1(new_n823), .A2(new_n824), .ZN(new_n825));
  OAI21_X1  g400(.A(G860), .B1(new_n822), .B2(new_n825), .ZN(new_n826));
  XOR2_X1   g401(.A(new_n826), .B(KEYINPUT37), .Z(new_n827));
  NOR2_X1   g402(.A1(new_n598), .A2(new_n608), .ZN(new_n828));
  XNOR2_X1  g403(.A(KEYINPUT38), .B(KEYINPUT39), .ZN(new_n829));
  XNOR2_X1  g404(.A(new_n828), .B(new_n829), .ZN(new_n830));
  NOR2_X1   g405(.A1(new_n822), .A2(new_n825), .ZN(new_n831));
  NAND3_X1  g406(.A1(new_n548), .A2(KEYINPUT101), .A3(new_n831), .ZN(new_n832));
  INV_X1    g407(.A(KEYINPUT101), .ZN(new_n833));
  OAI21_X1  g408(.A(new_n833), .B1(new_n822), .B2(new_n825), .ZN(new_n834));
  INV_X1    g409(.A(new_n821), .ZN(new_n835));
  NAND3_X1  g410(.A1(new_n835), .A2(G651), .A3(new_n819), .ZN(new_n836));
  NAND4_X1  g411(.A1(new_n836), .A2(KEYINPUT101), .A3(new_n823), .A4(new_n824), .ZN(new_n837));
  NAND3_X1  g412(.A1(new_n834), .A2(new_n837), .A3(new_n610), .ZN(new_n838));
  NAND2_X1  g413(.A1(new_n832), .A2(new_n838), .ZN(new_n839));
  XNOR2_X1  g414(.A(new_n830), .B(new_n839), .ZN(new_n840));
  OAI21_X1  g415(.A(new_n827), .B1(new_n840), .B2(G860), .ZN(G145));
  XOR2_X1   g416(.A(new_n725), .B(new_n623), .Z(new_n842));
  XOR2_X1   g417(.A(new_n497), .B(new_n697), .Z(new_n843));
  XOR2_X1   g418(.A(new_n842), .B(new_n843), .Z(new_n844));
  INV_X1    g419(.A(new_n844), .ZN(new_n845));
  NAND2_X1  g420(.A1(new_n479), .A2(G130), .ZN(new_n846));
  INV_X1    g421(.A(KEYINPUT102), .ZN(new_n847));
  XNOR2_X1  g422(.A(new_n846), .B(new_n847), .ZN(new_n848));
  OR2_X1    g423(.A1(G106), .A2(G2105), .ZN(new_n849));
  OAI211_X1 g424(.A(new_n849), .B(G2104), .C1(G118), .C2(new_n472), .ZN(new_n850));
  NAND2_X1  g425(.A1(new_n475), .A2(G142), .ZN(new_n851));
  NAND3_X1  g426(.A1(new_n848), .A2(new_n850), .A3(new_n851), .ZN(new_n852));
  AND2_X1   g427(.A1(new_n852), .A2(new_n708), .ZN(new_n853));
  NOR2_X1   g428(.A1(new_n852), .A2(new_n708), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n477), .B(new_n484), .ZN(new_n855));
  OR3_X1    g430(.A1(new_n853), .A2(new_n854), .A3(new_n855), .ZN(new_n856));
  XNOR2_X1  g431(.A(new_n620), .B(new_n800), .ZN(new_n857));
  OAI21_X1  g432(.A(new_n855), .B1(new_n853), .B2(new_n854), .ZN(new_n858));
  NAND3_X1  g433(.A1(new_n856), .A2(new_n857), .A3(new_n858), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  AOI21_X1  g435(.A(new_n857), .B1(new_n856), .B2(new_n858), .ZN(new_n861));
  OAI21_X1  g436(.A(new_n845), .B1(new_n860), .B2(new_n861), .ZN(new_n862));
  INV_X1    g437(.A(new_n861), .ZN(new_n863));
  NAND3_X1  g438(.A1(new_n863), .A2(new_n844), .A3(new_n859), .ZN(new_n864));
  INV_X1    g439(.A(G37), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n862), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  XNOR2_X1  g441(.A(new_n866), .B(KEYINPUT40), .ZN(G395));
  NAND2_X1  g442(.A1(G166), .A2(G288), .ZN(new_n868));
  INV_X1    g443(.A(new_n868), .ZN(new_n869));
  NOR2_X1   g444(.A1(G166), .A2(G288), .ZN(new_n870));
  NOR3_X1   g445(.A1(new_n869), .A2(new_n870), .A3(new_n789), .ZN(new_n871));
  NAND2_X1  g446(.A1(G303), .A2(new_n778), .ZN(new_n872));
  AOI21_X1  g447(.A(G305), .B1(new_n872), .B2(new_n868), .ZN(new_n873));
  INV_X1    g448(.A(KEYINPUT106), .ZN(new_n874));
  AOI21_X1  g449(.A(new_n874), .B1(new_n583), .B2(new_n585), .ZN(new_n875));
  NAND3_X1  g450(.A1(new_n583), .A2(new_n874), .A3(new_n585), .ZN(new_n876));
  INV_X1    g451(.A(new_n876), .ZN(new_n877));
  OAI22_X1  g452(.A1(new_n871), .A2(new_n873), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n789), .B1(new_n869), .B2(new_n870), .ZN(new_n879));
  INV_X1    g454(.A(new_n875), .ZN(new_n880));
  NAND3_X1  g455(.A1(new_n872), .A2(G305), .A3(new_n868), .ZN(new_n881));
  NAND4_X1  g456(.A1(new_n879), .A2(new_n880), .A3(new_n876), .A4(new_n881), .ZN(new_n882));
  AND2_X1   g457(.A1(new_n878), .A2(new_n882), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(KEYINPUT42), .ZN(new_n884));
  AND2_X1   g459(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n885));
  NOR2_X1   g460(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n886));
  OAI22_X1  g461(.A1(new_n885), .A2(new_n886), .B1(G559), .B2(new_n598), .ZN(new_n887));
  OR2_X1    g462(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n839), .A2(KEYINPUT103), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(new_n612), .A3(new_n889), .ZN(new_n890));
  NAND2_X1  g465(.A1(new_n887), .A2(new_n890), .ZN(new_n891));
  NAND2_X1  g466(.A1(new_n598), .A2(new_n605), .ZN(new_n892));
  NAND4_X1  g467(.A1(G299), .A2(new_n593), .A3(new_n592), .A4(new_n597), .ZN(new_n893));
  NAND3_X1  g468(.A1(new_n892), .A2(KEYINPUT104), .A3(new_n893), .ZN(new_n894));
  INV_X1    g469(.A(KEYINPUT104), .ZN(new_n895));
  NAND3_X1  g470(.A1(new_n599), .A2(new_n895), .A3(G299), .ZN(new_n896));
  NAND3_X1  g471(.A1(new_n894), .A2(KEYINPUT41), .A3(new_n896), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT41), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n892), .A2(new_n898), .A3(new_n893), .ZN(new_n899));
  AND2_X1   g474(.A1(new_n897), .A2(new_n899), .ZN(new_n900));
  NAND2_X1  g475(.A1(new_n891), .A2(new_n900), .ZN(new_n901));
  INV_X1    g476(.A(KEYINPUT105), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n901), .A2(new_n902), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n891), .A2(KEYINPUT105), .A3(new_n900), .ZN(new_n904));
  AND2_X1   g479(.A1(new_n903), .A2(new_n904), .ZN(new_n905));
  NAND2_X1  g480(.A1(new_n894), .A2(new_n896), .ZN(new_n906));
  INV_X1    g481(.A(new_n906), .ZN(new_n907));
  NAND3_X1  g482(.A1(new_n887), .A2(new_n890), .A3(new_n907), .ZN(new_n908));
  AOI21_X1  g483(.A(new_n884), .B1(new_n905), .B2(new_n908), .ZN(new_n909));
  AND4_X1   g484(.A1(new_n908), .A2(new_n884), .A3(new_n903), .A4(new_n904), .ZN(new_n910));
  OAI21_X1  g485(.A(G868), .B1(new_n909), .B2(new_n910), .ZN(new_n911));
  OAI21_X1  g486(.A(new_n911), .B1(G868), .B2(new_n831), .ZN(G295));
  OAI21_X1  g487(.A(new_n911), .B1(G868), .B2(new_n831), .ZN(G331));
  NAND2_X1  g488(.A1(G168), .A2(G301), .ZN(new_n914));
  NAND2_X1  g489(.A1(G286), .A2(G171), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n839), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  NAND2_X1  g491(.A1(new_n521), .A2(new_n523), .ZN(new_n917));
  INV_X1    g492(.A(KEYINPUT72), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n917), .A2(new_n918), .ZN(new_n919));
  NAND3_X1  g494(.A1(new_n521), .A2(KEYINPUT72), .A3(new_n523), .ZN(new_n920));
  AOI21_X1  g495(.A(new_n519), .B1(new_n919), .B2(new_n920), .ZN(new_n921));
  AOI21_X1  g496(.A(G301), .B1(new_n921), .B2(new_n518), .ZN(new_n922));
  NOR2_X1   g497(.A1(G286), .A2(G171), .ZN(new_n923));
  OAI211_X1 g498(.A(new_n832), .B(new_n838), .C1(new_n922), .C2(new_n923), .ZN(new_n924));
  INV_X1    g499(.A(KEYINPUT108), .ZN(new_n925));
  NAND3_X1  g500(.A1(new_n916), .A2(new_n924), .A3(new_n925), .ZN(new_n926));
  INV_X1    g501(.A(new_n839), .ZN(new_n927));
  OAI211_X1 g502(.A(new_n927), .B(KEYINPUT108), .C1(new_n923), .C2(new_n922), .ZN(new_n928));
  NAND3_X1  g503(.A1(new_n900), .A2(new_n926), .A3(new_n928), .ZN(new_n929));
  NAND3_X1  g504(.A1(new_n907), .A2(new_n924), .A3(new_n916), .ZN(new_n930));
  NAND3_X1  g505(.A1(new_n929), .A2(new_n883), .A3(new_n930), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n931), .A2(new_n865), .ZN(new_n932));
  AOI21_X1  g507(.A(new_n883), .B1(new_n929), .B2(new_n930), .ZN(new_n933));
  OAI21_X1  g508(.A(KEYINPUT43), .B1(new_n932), .B2(new_n933), .ZN(new_n934));
  INV_X1    g509(.A(new_n883), .ZN(new_n935));
  NAND2_X1  g510(.A1(new_n916), .A2(new_n924), .ZN(new_n936));
  NAND2_X1  g511(.A1(new_n892), .A2(new_n893), .ZN(new_n937));
  NAND2_X1  g512(.A1(new_n937), .A2(KEYINPUT41), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n906), .A2(new_n898), .ZN(new_n939));
  NAND3_X1  g514(.A1(new_n936), .A2(new_n938), .A3(new_n939), .ZN(new_n940));
  INV_X1    g515(.A(new_n940), .ZN(new_n941));
  AOI21_X1  g516(.A(new_n906), .B1(new_n926), .B2(new_n928), .ZN(new_n942));
  OAI21_X1  g517(.A(new_n935), .B1(new_n941), .B2(new_n942), .ZN(new_n943));
  INV_X1    g518(.A(KEYINPUT43), .ZN(new_n944));
  NAND4_X1  g519(.A1(new_n943), .A2(new_n944), .A3(new_n865), .A4(new_n931), .ZN(new_n945));
  NAND2_X1  g520(.A1(new_n934), .A2(new_n945), .ZN(new_n946));
  XNOR2_X1  g521(.A(KEYINPUT107), .B(KEYINPUT44), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  INV_X1    g523(.A(KEYINPUT44), .ZN(new_n949));
  NAND2_X1  g524(.A1(new_n926), .A2(new_n928), .ZN(new_n950));
  NAND2_X1  g525(.A1(new_n950), .A2(new_n907), .ZN(new_n951));
  AOI21_X1  g526(.A(new_n883), .B1(new_n951), .B2(new_n940), .ZN(new_n952));
  OAI21_X1  g527(.A(KEYINPUT43), .B1(new_n932), .B2(new_n952), .ZN(new_n953));
  AOI21_X1  g528(.A(new_n949), .B1(new_n953), .B2(KEYINPUT109), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n954), .B1(KEYINPUT109), .B2(new_n953), .ZN(new_n955));
  NOR3_X1   g530(.A1(new_n932), .A2(KEYINPUT43), .A3(new_n933), .ZN(new_n956));
  OAI21_X1  g531(.A(new_n948), .B1(new_n955), .B2(new_n956), .ZN(G397));
  INV_X1    g532(.A(G1384), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n495), .A2(G102), .ZN(new_n959));
  INV_X1    g534(.A(new_n493), .ZN(new_n960));
  AOI21_X1  g535(.A(new_n960), .B1(new_n489), .B2(G126), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n959), .B1(new_n961), .B2(new_n472), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n488), .A2(new_n490), .ZN(new_n963));
  OAI21_X1  g538(.A(new_n958), .B1(new_n962), .B2(new_n963), .ZN(new_n964));
  INV_X1    g539(.A(KEYINPUT110), .ZN(new_n965));
  XNOR2_X1  g540(.A(new_n964), .B(new_n965), .ZN(new_n966));
  INV_X1    g541(.A(KEYINPUT45), .ZN(new_n967));
  NAND2_X1  g542(.A1(new_n966), .A2(new_n967), .ZN(new_n968));
  NAND4_X1  g543(.A1(new_n471), .A2(new_n474), .A3(new_n476), .A4(G40), .ZN(new_n969));
  OR3_X1    g544(.A1(new_n968), .A2(KEYINPUT111), .A3(new_n969), .ZN(new_n970));
  OAI21_X1  g545(.A(KEYINPUT111), .B1(new_n968), .B2(new_n969), .ZN(new_n971));
  AND2_X1   g546(.A1(new_n970), .A2(new_n971), .ZN(new_n972));
  XOR2_X1   g547(.A(new_n697), .B(G2067), .Z(new_n973));
  NAND2_X1  g548(.A1(new_n800), .A2(new_n803), .ZN(new_n974));
  XNOR2_X1  g549(.A(new_n707), .B(new_n675), .ZN(new_n975));
  OR2_X1    g550(.A1(new_n800), .A2(new_n803), .ZN(new_n976));
  NAND4_X1  g551(.A1(new_n973), .A2(new_n974), .A3(new_n975), .A4(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(new_n977), .ZN(new_n978));
  NAND2_X1  g553(.A1(G290), .A2(G1986), .ZN(new_n979));
  NOR2_X1   g554(.A1(G290), .A2(G1986), .ZN(new_n980));
  INV_X1    g555(.A(new_n980), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n979), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n972), .A2(new_n982), .ZN(new_n983));
  INV_X1    g558(.A(new_n969), .ZN(new_n984));
  AOI21_X1  g559(.A(G1384), .B1(new_n491), .B2(new_n496), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  NAND2_X1  g561(.A1(new_n986), .A2(G8), .ZN(new_n987));
  OR2_X1    g562(.A1(G305), .A2(KEYINPUT49), .ZN(new_n988));
  NAND2_X1  g563(.A1(G305), .A2(KEYINPUT49), .ZN(new_n989));
  INV_X1    g564(.A(G1981), .ZN(new_n990));
  INV_X1    g565(.A(KEYINPUT115), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n990), .B1(new_n574), .B2(new_n991), .ZN(new_n992));
  AND3_X1   g567(.A1(new_n988), .A2(new_n989), .A3(new_n992), .ZN(new_n993));
  AOI21_X1  g568(.A(new_n992), .B1(new_n988), .B2(new_n989), .ZN(new_n994));
  NOR3_X1   g569(.A1(new_n993), .A2(new_n994), .A3(new_n987), .ZN(new_n995));
  INV_X1    g570(.A(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G1976), .ZN(new_n997));
  NAND3_X1  g572(.A1(new_n996), .A2(new_n997), .A3(new_n778), .ZN(new_n998));
  NAND2_X1  g573(.A1(new_n789), .A2(new_n990), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n987), .B1(new_n998), .B2(new_n999), .ZN(new_n1000));
  OAI211_X1 g575(.A(new_n986), .B(G8), .C1(new_n997), .C2(G288), .ZN(new_n1001));
  INV_X1    g576(.A(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT114), .ZN(new_n1003));
  INV_X1    g578(.A(KEYINPUT52), .ZN(new_n1004));
  NOR2_X1   g579(.A1(new_n778), .A2(G1976), .ZN(new_n1005));
  INV_X1    g580(.A(new_n1005), .ZN(new_n1006));
  NAND4_X1  g581(.A1(new_n1002), .A2(new_n1003), .A3(new_n1004), .A4(new_n1006), .ZN(new_n1007));
  NOR2_X1   g582(.A1(new_n964), .A2(new_n969), .ZN(new_n1008));
  INV_X1    g583(.A(G8), .ZN(new_n1009));
  NOR2_X1   g584(.A1(new_n1008), .A2(new_n1009), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n778), .A2(G1976), .ZN(new_n1011));
  NAND3_X1  g586(.A1(new_n1010), .A2(new_n1004), .A3(new_n1011), .ZN(new_n1012));
  OAI21_X1  g587(.A(KEYINPUT114), .B1(new_n1012), .B2(new_n1005), .ZN(new_n1013));
  NAND2_X1  g588(.A1(new_n1007), .A2(new_n1013), .ZN(new_n1014));
  INV_X1    g589(.A(KEYINPUT113), .ZN(new_n1015));
  AOI21_X1  g590(.A(new_n1004), .B1(new_n1001), .B2(new_n1015), .ZN(new_n1016));
  NAND3_X1  g591(.A1(new_n1010), .A2(KEYINPUT113), .A3(new_n1011), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n1016), .A2(new_n1017), .ZN(new_n1018));
  NAND3_X1  g593(.A1(new_n1014), .A2(new_n1018), .A3(new_n996), .ZN(new_n1019));
  NAND2_X1  g594(.A1(new_n964), .A2(new_n967), .ZN(new_n1020));
  AOI21_X1  g595(.A(new_n969), .B1(new_n1020), .B2(KEYINPUT112), .ZN(new_n1021));
  NAND2_X1  g596(.A1(new_n985), .A2(KEYINPUT45), .ZN(new_n1022));
  AOI21_X1  g597(.A(KEYINPUT45), .B1(new_n497), .B2(new_n958), .ZN(new_n1023));
  INV_X1    g598(.A(KEYINPUT112), .ZN(new_n1024));
  NAND2_X1  g599(.A1(new_n1023), .A2(new_n1024), .ZN(new_n1025));
  NAND3_X1  g600(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .ZN(new_n1026));
  AOI21_X1  g601(.A(new_n969), .B1(new_n964), .B2(KEYINPUT50), .ZN(new_n1027));
  INV_X1    g602(.A(KEYINPUT50), .ZN(new_n1028));
  OAI211_X1 g603(.A(new_n1028), .B(new_n958), .C1(new_n962), .C2(new_n963), .ZN(new_n1029));
  NAND2_X1  g604(.A1(new_n1027), .A2(new_n1029), .ZN(new_n1030));
  INV_X1    g605(.A(new_n1030), .ZN(new_n1031));
  AOI22_X1  g606(.A1(new_n1026), .A2(new_n786), .B1(new_n765), .B2(new_n1031), .ZN(new_n1032));
  INV_X1    g607(.A(new_n1032), .ZN(new_n1033));
  NAND2_X1  g608(.A1(G303), .A2(G8), .ZN(new_n1034));
  XNOR2_X1  g609(.A(new_n1034), .B(KEYINPUT55), .ZN(new_n1035));
  INV_X1    g610(.A(new_n1035), .ZN(new_n1036));
  NAND3_X1  g611(.A1(new_n1033), .A2(G8), .A3(new_n1036), .ZN(new_n1037));
  NOR2_X1   g612(.A1(new_n1019), .A2(new_n1037), .ZN(new_n1038));
  AOI221_X4 g613(.A(new_n995), .B1(new_n1016), .B2(new_n1017), .C1(new_n1007), .C2(new_n1013), .ZN(new_n1039));
  OAI21_X1  g614(.A(KEYINPUT117), .B1(new_n1023), .B2(new_n969), .ZN(new_n1040));
  INV_X1    g615(.A(KEYINPUT117), .ZN(new_n1041));
  NAND3_X1  g616(.A1(new_n1020), .A2(new_n1041), .A3(new_n984), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1040), .A2(new_n1022), .A3(new_n1042), .ZN(new_n1043));
  AOI22_X1  g618(.A1(new_n1043), .A2(new_n687), .B1(new_n741), .B2(new_n1031), .ZN(new_n1044));
  NOR3_X1   g619(.A1(new_n1044), .A2(new_n1009), .A3(G286), .ZN(new_n1045));
  OAI21_X1  g620(.A(new_n1035), .B1(new_n1032), .B2(new_n1009), .ZN(new_n1046));
  NAND4_X1  g621(.A1(new_n1039), .A2(new_n1045), .A3(new_n1037), .A4(new_n1046), .ZN(new_n1047));
  AOI211_X1 g622(.A(new_n1000), .B(new_n1038), .C1(new_n1047), .C2(KEYINPUT63), .ZN(new_n1048));
  XNOR2_X1  g623(.A(KEYINPUT119), .B(KEYINPUT57), .ZN(new_n1049));
  XNOR2_X1  g624(.A(G299), .B(new_n1049), .ZN(new_n1050));
  INV_X1    g625(.A(new_n1050), .ZN(new_n1051));
  INV_X1    g626(.A(KEYINPUT116), .ZN(new_n1052));
  AOI21_X1  g627(.A(new_n1052), .B1(new_n985), .B2(new_n1028), .ZN(new_n1053));
  NOR2_X1   g628(.A1(new_n1029), .A2(KEYINPUT116), .ZN(new_n1054));
  OAI21_X1  g629(.A(new_n1027), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  XNOR2_X1  g630(.A(KEYINPUT118), .B(G1956), .ZN(new_n1056));
  INV_X1    g631(.A(new_n1056), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1055), .A2(new_n1057), .ZN(new_n1058));
  XNOR2_X1  g633(.A(KEYINPUT56), .B(G2072), .ZN(new_n1059));
  NAND4_X1  g634(.A1(new_n1021), .A2(new_n1022), .A3(new_n1025), .A4(new_n1059), .ZN(new_n1060));
  AOI21_X1  g635(.A(new_n1051), .B1(new_n1058), .B2(new_n1060), .ZN(new_n1061));
  NOR3_X1   g636(.A1(new_n964), .A2(new_n969), .A3(G2067), .ZN(new_n1062));
  AOI22_X1  g637(.A1(new_n1030), .A2(new_n760), .B1(KEYINPUT120), .B2(new_n1062), .ZN(new_n1063));
  INV_X1    g638(.A(KEYINPUT120), .ZN(new_n1064));
  OAI21_X1  g639(.A(new_n1064), .B1(new_n986), .B2(G2067), .ZN(new_n1065));
  AOI21_X1  g640(.A(new_n598), .B1(new_n1063), .B2(new_n1065), .ZN(new_n1066));
  OR2_X1    g641(.A1(new_n1061), .A2(new_n1066), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1058), .A2(new_n1051), .A3(new_n1060), .ZN(new_n1068));
  AND2_X1   g643(.A1(new_n1067), .A2(new_n1068), .ZN(new_n1069));
  INV_X1    g644(.A(KEYINPUT61), .ZN(new_n1070));
  NAND2_X1  g645(.A1(new_n1058), .A2(new_n1060), .ZN(new_n1071));
  NAND3_X1  g646(.A1(new_n1071), .A2(KEYINPUT122), .A3(new_n1050), .ZN(new_n1072));
  INV_X1    g647(.A(KEYINPUT122), .ZN(new_n1073));
  NAND2_X1  g648(.A1(new_n1068), .A2(new_n1073), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1070), .B(new_n1072), .C1(new_n1074), .C2(new_n1061), .ZN(new_n1075));
  AND3_X1   g650(.A1(new_n1063), .A2(new_n598), .A3(new_n1065), .ZN(new_n1076));
  OAI21_X1  g651(.A(KEYINPUT60), .B1(new_n1076), .B2(new_n1066), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1030), .A2(new_n760), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT60), .ZN(new_n1079));
  NAND2_X1  g654(.A1(new_n1062), .A2(KEYINPUT120), .ZN(new_n1080));
  NAND4_X1  g655(.A1(new_n1078), .A2(new_n1079), .A3(new_n1065), .A4(new_n1080), .ZN(new_n1081));
  NOR2_X1   g656(.A1(new_n1081), .A2(new_n598), .ZN(new_n1082));
  NAND2_X1  g657(.A1(new_n1068), .A2(KEYINPUT61), .ZN(new_n1083));
  AOI21_X1  g658(.A(new_n1082), .B1(new_n1083), .B2(KEYINPUT123), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT123), .ZN(new_n1085));
  NAND3_X1  g660(.A1(new_n1068), .A2(new_n1085), .A3(KEYINPUT61), .ZN(new_n1086));
  AND4_X1   g661(.A1(new_n1075), .A2(new_n1077), .A3(new_n1084), .A4(new_n1086), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n1025), .A2(new_n1022), .ZN(new_n1088));
  NAND4_X1  g663(.A1(new_n1088), .A2(KEYINPUT121), .A3(new_n675), .A4(new_n1021), .ZN(new_n1089));
  INV_X1    g664(.A(KEYINPUT121), .ZN(new_n1090));
  OAI21_X1  g665(.A(new_n1090), .B1(new_n1026), .B2(G1996), .ZN(new_n1091));
  XNOR2_X1  g666(.A(KEYINPUT58), .B(G1341), .ZN(new_n1092));
  OAI211_X1 g667(.A(new_n1089), .B(new_n1091), .C1(new_n1008), .C2(new_n1092), .ZN(new_n1093));
  AND3_X1   g668(.A1(new_n1093), .A2(KEYINPUT59), .A3(new_n548), .ZN(new_n1094));
  AOI21_X1  g669(.A(KEYINPUT59), .B1(new_n1093), .B2(new_n548), .ZN(new_n1095));
  NOR2_X1   g670(.A1(new_n1094), .A2(new_n1095), .ZN(new_n1096));
  AOI21_X1  g671(.A(new_n1069), .B1(new_n1087), .B2(new_n1096), .ZN(new_n1097));
  NAND2_X1  g672(.A1(new_n1043), .A2(new_n687), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1031), .A2(new_n741), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1098), .A2(G168), .A3(new_n1099), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1100), .A2(G8), .ZN(new_n1101));
  NOR2_X1   g676(.A1(new_n1044), .A2(G168), .ZN(new_n1102));
  OAI21_X1  g677(.A(KEYINPUT51), .B1(new_n1101), .B2(new_n1102), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1009), .B1(new_n1044), .B2(G168), .ZN(new_n1104));
  INV_X1    g679(.A(KEYINPUT51), .ZN(new_n1105));
  NAND2_X1  g680(.A1(new_n1104), .A2(new_n1105), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1103), .A2(new_n1106), .ZN(new_n1107));
  NAND2_X1  g682(.A1(new_n1026), .A2(new_n786), .ZN(new_n1108));
  OAI21_X1  g683(.A(new_n1108), .B1(G2090), .B2(new_n1055), .ZN(new_n1109));
  AOI21_X1  g684(.A(new_n1036), .B1(new_n1109), .B2(G8), .ZN(new_n1110));
  NOR3_X1   g685(.A1(new_n1032), .A2(new_n1009), .A3(new_n1035), .ZN(new_n1111));
  NOR3_X1   g686(.A1(new_n1019), .A2(new_n1110), .A3(new_n1111), .ZN(new_n1112));
  INV_X1    g687(.A(G2078), .ZN(new_n1113));
  NAND4_X1  g688(.A1(new_n1021), .A2(new_n1113), .A3(new_n1025), .A4(new_n1022), .ZN(new_n1114));
  INV_X1    g689(.A(KEYINPUT53), .ZN(new_n1115));
  AOI22_X1  g690(.A1(new_n1114), .A2(new_n1115), .B1(new_n738), .B2(new_n1030), .ZN(new_n1116));
  NOR2_X1   g691(.A1(new_n1115), .A2(G2078), .ZN(new_n1117));
  NAND4_X1  g692(.A1(new_n1040), .A2(new_n1022), .A3(new_n1042), .A4(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1116), .A2(G301), .A3(new_n1118), .ZN(new_n1119));
  NAND4_X1  g694(.A1(new_n968), .A2(new_n984), .A3(new_n1022), .A4(new_n1117), .ZN(new_n1120));
  AND2_X1   g695(.A1(new_n1116), .A2(new_n1120), .ZN(new_n1121));
  OAI211_X1 g696(.A(KEYINPUT54), .B(new_n1119), .C1(new_n1121), .C2(G301), .ZN(new_n1122));
  INV_X1    g697(.A(KEYINPUT54), .ZN(new_n1123));
  AND3_X1   g698(.A1(new_n1116), .A2(G301), .A3(new_n1120), .ZN(new_n1124));
  AOI21_X1  g699(.A(G301), .B1(new_n1116), .B2(new_n1118), .ZN(new_n1125));
  OAI21_X1  g700(.A(new_n1123), .B1(new_n1124), .B2(new_n1125), .ZN(new_n1126));
  NAND4_X1  g701(.A1(new_n1107), .A2(new_n1112), .A3(new_n1122), .A4(new_n1126), .ZN(new_n1127));
  OAI21_X1  g702(.A(new_n1048), .B1(new_n1097), .B2(new_n1127), .ZN(new_n1128));
  INV_X1    g703(.A(new_n1112), .ZN(new_n1129));
  NAND2_X1  g704(.A1(new_n1098), .A2(new_n1099), .ZN(new_n1130));
  NAND2_X1  g705(.A1(new_n1130), .A2(G286), .ZN(new_n1131));
  AOI21_X1  g706(.A(new_n1105), .B1(new_n1104), .B2(new_n1131), .ZN(new_n1132));
  NOR2_X1   g707(.A1(new_n1101), .A2(KEYINPUT51), .ZN(new_n1133));
  OAI21_X1  g708(.A(KEYINPUT62), .B1(new_n1132), .B2(new_n1133), .ZN(new_n1134));
  INV_X1    g709(.A(KEYINPUT62), .ZN(new_n1135));
  NAND3_X1  g710(.A1(new_n1103), .A2(new_n1135), .A3(new_n1106), .ZN(new_n1136));
  NAND3_X1  g711(.A1(new_n1134), .A2(new_n1136), .A3(new_n1125), .ZN(new_n1137));
  INV_X1    g712(.A(KEYINPUT63), .ZN(new_n1138));
  NAND2_X1  g713(.A1(new_n1045), .A2(new_n1138), .ZN(new_n1139));
  AOI21_X1  g714(.A(new_n1129), .B1(new_n1137), .B2(new_n1139), .ZN(new_n1140));
  OAI21_X1  g715(.A(new_n983), .B1(new_n1128), .B2(new_n1140), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT125), .ZN(new_n1142));
  OAI211_X1 g717(.A(new_n972), .B(new_n675), .C1(new_n1142), .C2(KEYINPUT46), .ZN(new_n1143));
  INV_X1    g718(.A(new_n973), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n972), .B1(new_n707), .B2(new_n1144), .ZN(new_n1145));
  XOR2_X1   g720(.A(KEYINPUT125), .B(KEYINPUT46), .Z(new_n1146));
  NAND2_X1  g721(.A1(new_n970), .A2(new_n971), .ZN(new_n1147));
  OAI21_X1  g722(.A(new_n1146), .B1(new_n1147), .B2(G1996), .ZN(new_n1148));
  NAND3_X1  g723(.A1(new_n1143), .A2(new_n1145), .A3(new_n1148), .ZN(new_n1149));
  NAND2_X1  g724(.A1(new_n1149), .A2(KEYINPUT47), .ZN(new_n1150));
  INV_X1    g725(.A(KEYINPUT47), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1143), .A2(new_n1151), .A3(new_n1145), .A4(new_n1148), .ZN(new_n1152));
  NAND2_X1  g727(.A1(new_n972), .A2(new_n980), .ZN(new_n1153));
  XNOR2_X1  g728(.A(new_n1153), .B(KEYINPUT48), .ZN(new_n1154));
  NOR2_X1   g729(.A1(new_n1147), .A2(new_n978), .ZN(new_n1155));
  XNOR2_X1  g730(.A(new_n1155), .B(KEYINPUT126), .ZN(new_n1156));
  AOI22_X1  g731(.A1(new_n1150), .A2(new_n1152), .B1(new_n1154), .B2(new_n1156), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n973), .A2(new_n975), .ZN(new_n1158));
  OAI22_X1  g733(.A1(new_n1158), .A2(new_n976), .B1(G2067), .B2(new_n697), .ZN(new_n1159));
  NAND2_X1  g734(.A1(new_n972), .A2(new_n1159), .ZN(new_n1160));
  XNOR2_X1  g735(.A(new_n1160), .B(KEYINPUT124), .ZN(new_n1161));
  AND2_X1   g736(.A1(new_n1157), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g737(.A1(new_n1141), .A2(new_n1162), .ZN(G329));
  assign    G231 = 1'b0;
  INV_X1    g738(.A(KEYINPUT127), .ZN(new_n1165));
  OAI21_X1  g739(.A(G319), .B1(new_n682), .B2(new_n683), .ZN(new_n1166));
  INV_X1    g740(.A(new_n1166), .ZN(new_n1167));
  NOR2_X1   g741(.A1(G401), .A2(G227), .ZN(new_n1168));
  AND2_X1   g742(.A1(new_n866), .A2(new_n1168), .ZN(new_n1169));
  AND4_X1   g743(.A1(new_n1165), .A2(new_n946), .A3(new_n1167), .A4(new_n1169), .ZN(new_n1170));
  AOI21_X1  g744(.A(new_n1166), .B1(new_n934), .B2(new_n945), .ZN(new_n1171));
  AOI21_X1  g745(.A(new_n1165), .B1(new_n1171), .B2(new_n1169), .ZN(new_n1172));
  NOR2_X1   g746(.A1(new_n1170), .A2(new_n1172), .ZN(G308));
  NAND3_X1  g747(.A1(new_n946), .A2(new_n1167), .A3(new_n1169), .ZN(new_n1174));
  NAND2_X1  g748(.A1(new_n1174), .A2(KEYINPUT127), .ZN(new_n1175));
  NAND3_X1  g749(.A1(new_n1171), .A2(new_n1165), .A3(new_n1169), .ZN(new_n1176));
  NAND2_X1  g750(.A1(new_n1175), .A2(new_n1176), .ZN(G225));
endmodule


