//Secret key is'1 0 0 0 1 0 0 1 0 0 1 1 1 1 0 0 1 1 0 1 0 1 1 0 1 0 0 1 0 0 1 1 0 1 0 1 1 1 0 1 0 1 0 0 0 0 1 1 0 0 1 0 0 0 0 0 1 0 1 1 1 0 0 1 0 1 0 0 1 0 0 0 1 1 0 0 0 0 1 0 0 0 1 1 0 1 0 0 0 1 0 0 1 1 0 0 1 0 1 0 0 1 0 1 0 1 1 0 1 0 0 1 0 0 1 0 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c3540" written by ABC on Sat Dec 16 05:39:03 2023

module locked_locked_c3540 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G13, G20, G33, G41, G45, G50, G58, G68, G77, G87, G97,
    G107, G116, G124, G125, G128, G132, G137, G143, G150, G159, G169, G179,
    G190, G200, G213, G222, G223, G226, G232, G238, G244, G250, G257, G264,
    G270, G274, G283, G294, G303, G311, G317, G322, G326, G329, G330, G343,
    G1698, G2897,
    G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384, G367,
    G387, G393, G390, G378, G375, G381, G407, G409, G405, G402  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G13, G20, G33, G41, G45, G50,
    G58, G68, G77, G87, G97, G107, G116, G124, G125, G128, G132, G137,
    G143, G150, G159, G169, G179, G190, G200, G213, G222, G223, G226, G232,
    G238, G244, G250, G257, G264, G270, G274, G283, G294, G303, G311, G317,
    G322, G326, G329, G330, G343, G1698, G2897;
  output G353, G355, G361, G358, G351, G372, G369, G399, G364, G396, G384,
    G367, G387, G393, G390, G378, G375, G381, G407, G409, G405, G402;
  wire new_n203, new_n204, new_n205, new_n206, new_n207, new_n208, new_n209,
    new_n210, new_n211, new_n212, new_n213, new_n214, new_n215, new_n216,
    new_n217, new_n218, new_n219, new_n220, new_n221, new_n222, new_n223,
    new_n224, new_n225, new_n226, new_n227, new_n228, new_n229, new_n230,
    new_n231, new_n233, new_n234, new_n235, new_n236, new_n237, new_n238,
    new_n239, new_n240, new_n242, new_n243, new_n244, new_n245, new_n246,
    new_n247, new_n249, new_n250, new_n251, new_n252, new_n253, new_n254,
    new_n255, new_n256, new_n257, new_n258, new_n259, new_n260, new_n261,
    new_n262, new_n263, new_n264, new_n265, new_n266, new_n267, new_n268,
    new_n269, new_n270, new_n271, new_n272, new_n273, new_n274, new_n275,
    new_n276, new_n277, new_n278, new_n279, new_n280, new_n281, new_n282,
    new_n283, new_n284, new_n285, new_n286, new_n287, new_n288, new_n289,
    new_n290, new_n291, new_n292, new_n293, new_n294, new_n295, new_n296,
    new_n297, new_n298, new_n299, new_n300, new_n301, new_n302, new_n303,
    new_n304, new_n305, new_n306, new_n307, new_n308, new_n309, new_n310,
    new_n311, new_n312, new_n313, new_n314, new_n315, new_n316, new_n317,
    new_n318, new_n319, new_n320, new_n321, new_n322, new_n323, new_n324,
    new_n325, new_n326, new_n327, new_n328, new_n329, new_n330, new_n331,
    new_n332, new_n333, new_n334, new_n335, new_n336, new_n337, new_n338,
    new_n339, new_n340, new_n341, new_n342, new_n343, new_n344, new_n345,
    new_n346, new_n347, new_n348, new_n349, new_n350, new_n351, new_n352,
    new_n353, new_n354, new_n355, new_n356, new_n357, new_n358, new_n359,
    new_n360, new_n361, new_n362, new_n363, new_n364, new_n365, new_n366,
    new_n367, new_n368, new_n369, new_n370, new_n371, new_n372, new_n373,
    new_n374, new_n375, new_n376, new_n377, new_n378, new_n379, new_n380,
    new_n381, new_n382, new_n383, new_n384, new_n385, new_n386, new_n387,
    new_n388, new_n389, new_n390, new_n391, new_n392, new_n393, new_n394,
    new_n395, new_n396, new_n397, new_n398, new_n399, new_n400, new_n401,
    new_n402, new_n403, new_n404, new_n405, new_n406, new_n407, new_n408,
    new_n409, new_n410, new_n411, new_n412, new_n413, new_n414, new_n415,
    new_n416, new_n417, new_n418, new_n419, new_n420, new_n421, new_n422,
    new_n423, new_n424, new_n425, new_n426, new_n427, new_n428, new_n429,
    new_n430, new_n431, new_n432, new_n433, new_n434, new_n435, new_n436,
    new_n437, new_n438, new_n439, new_n440, new_n441, new_n442, new_n443,
    new_n444, new_n445, new_n446, new_n447, new_n448, new_n449, new_n450,
    new_n451, new_n452, new_n453, new_n454, new_n455, new_n456, new_n457,
    new_n458, new_n459, new_n460, new_n461, new_n462, new_n463, new_n464,
    new_n465, new_n466, new_n467, new_n468, new_n469, new_n470, new_n471,
    new_n472, new_n473, new_n474, new_n475, new_n476, new_n477, new_n478,
    new_n479, new_n480, new_n481, new_n482, new_n483, new_n484, new_n485,
    new_n486, new_n487, new_n488, new_n489, new_n490, new_n491, new_n492,
    new_n493, new_n494, new_n495, new_n496, new_n497, new_n498, new_n499,
    new_n500, new_n501, new_n502, new_n503, new_n504, new_n505, new_n506,
    new_n507, new_n508, new_n509, new_n510, new_n511, new_n512, new_n513,
    new_n514, new_n515, new_n516, new_n517, new_n518, new_n519, new_n520,
    new_n521, new_n522, new_n523, new_n524, new_n525, new_n526, new_n527,
    new_n528, new_n529, new_n530, new_n531, new_n532, new_n533, new_n534,
    new_n535, new_n536, new_n537, new_n538, new_n539, new_n540, new_n541,
    new_n542, new_n543, new_n544, new_n545, new_n546, new_n547, new_n548,
    new_n549, new_n550, new_n551, new_n552, new_n553, new_n554, new_n555,
    new_n556, new_n557, new_n558, new_n559, new_n560, new_n561, new_n562,
    new_n563, new_n564, new_n565, new_n566, new_n567, new_n568, new_n569,
    new_n570, new_n571, new_n572, new_n573, new_n574, new_n575, new_n576,
    new_n577, new_n578, new_n579, new_n580, new_n581, new_n582, new_n583,
    new_n584, new_n585, new_n586, new_n587, new_n588, new_n589, new_n590,
    new_n591, new_n592, new_n593, new_n594, new_n595, new_n596, new_n597,
    new_n598, new_n599, new_n600, new_n601, new_n602, new_n603, new_n604,
    new_n605, new_n606, new_n607, new_n608, new_n609, new_n610, new_n611,
    new_n612, new_n613, new_n614, new_n615, new_n616, new_n617, new_n618,
    new_n619, new_n620, new_n621, new_n622, new_n623, new_n624, new_n625,
    new_n626, new_n627, new_n628, new_n629, new_n630, new_n632, new_n633,
    new_n634, new_n635, new_n636, new_n637, new_n638, new_n639, new_n640,
    new_n641, new_n642, new_n643, new_n644, new_n645, new_n646, new_n647,
    new_n648, new_n649, new_n650, new_n651, new_n652, new_n653, new_n654,
    new_n655, new_n656, new_n657, new_n658, new_n660, new_n661, new_n662,
    new_n663, new_n664, new_n665, new_n666, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n682, new_n683,
    new_n684, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n735, new_n736, new_n737, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n747, new_n748,
    new_n749, new_n750, new_n751, new_n752, new_n753, new_n754, new_n755,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n845, new_n846, new_n847, new_n848,
    new_n849, new_n850, new_n851, new_n852, new_n853, new_n854, new_n855,
    new_n856, new_n857, new_n858, new_n859, new_n860, new_n861, new_n862,
    new_n863, new_n864, new_n865, new_n866, new_n867, new_n868, new_n869,
    new_n870, new_n871, new_n872, new_n873, new_n874, new_n875, new_n876,
    new_n877, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n889, new_n890,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n898, new_n899, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n925, new_n926,
    new_n927, new_n928, new_n929, new_n930, new_n931, new_n932, new_n933,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n940,
    new_n941, new_n942, new_n943, new_n944, new_n945, new_n946, new_n947,
    new_n948, new_n949, new_n950, new_n951, new_n952, new_n953, new_n954,
    new_n955, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n995, new_n996, new_n997,
    new_n998, new_n999, new_n1000, new_n1001, new_n1002, new_n1003,
    new_n1004, new_n1005, new_n1006, new_n1007, new_n1008, new_n1009,
    new_n1010, new_n1011, new_n1012, new_n1013, new_n1014, new_n1015,
    new_n1016, new_n1017, new_n1018, new_n1019, new_n1020, new_n1022,
    new_n1023, new_n1024, new_n1025, new_n1026, new_n1027, new_n1028,
    new_n1029, new_n1030, new_n1031, new_n1032, new_n1033, new_n1034,
    new_n1035, new_n1036, new_n1037, new_n1038, new_n1039, new_n1040,
    new_n1041, new_n1042, new_n1043, new_n1044, new_n1045, new_n1046,
    new_n1047, new_n1048, new_n1049, new_n1051, new_n1052, new_n1053,
    new_n1054, new_n1055, new_n1056, new_n1057, new_n1058, new_n1059,
    new_n1060, new_n1061, new_n1062, new_n1063, new_n1064, new_n1065,
    new_n1066, new_n1067, new_n1068, new_n1069, new_n1070, new_n1071,
    new_n1072, new_n1073, new_n1074, new_n1075, new_n1076, new_n1077,
    new_n1078, new_n1079, new_n1080, new_n1081, new_n1082, new_n1083,
    new_n1084, new_n1085, new_n1086, new_n1087, new_n1088, new_n1089,
    new_n1090, new_n1091, new_n1092, new_n1093, new_n1094, new_n1095,
    new_n1096, new_n1097, new_n1098, new_n1099, new_n1100, new_n1101,
    new_n1102, new_n1103, new_n1104, new_n1105, new_n1106, new_n1107,
    new_n1108, new_n1109, new_n1110, new_n1111, new_n1112, new_n1113,
    new_n1114, new_n1115, new_n1116, new_n1117, new_n1118, new_n1119,
    new_n1120, new_n1121, new_n1122, new_n1123, new_n1124, new_n1125,
    new_n1126, new_n1127, new_n1128, new_n1129, new_n1130, new_n1131,
    new_n1132, new_n1133, new_n1134, new_n1135, new_n1136, new_n1137,
    new_n1138, new_n1139, new_n1140, new_n1141, new_n1142, new_n1143,
    new_n1144, new_n1145, new_n1146, new_n1148, new_n1149, new_n1150,
    new_n1151, new_n1152, new_n1153, new_n1154, new_n1155, new_n1156,
    new_n1157, new_n1158, new_n1159, new_n1160, new_n1161, new_n1162,
    new_n1163, new_n1164, new_n1165, new_n1166, new_n1167, new_n1168,
    new_n1169, new_n1170, new_n1171, new_n1172, new_n1173, new_n1174,
    new_n1175, new_n1176, new_n1177, new_n1178, new_n1179, new_n1180,
    new_n1181, new_n1182, new_n1183, new_n1184, new_n1185, new_n1186,
    new_n1187, new_n1188, new_n1189, new_n1190, new_n1191, new_n1192,
    new_n1193, new_n1194, new_n1195, new_n1196, new_n1197, new_n1198,
    new_n1199, new_n1200, new_n1201, new_n1202, new_n1203, new_n1204,
    new_n1205, new_n1206, new_n1207, new_n1208, new_n1209, new_n1210,
    new_n1211, new_n1212, new_n1213, new_n1214, new_n1215, new_n1216,
    new_n1218, new_n1219, new_n1220, new_n1221, new_n1222, new_n1223,
    new_n1224, new_n1225, new_n1226, new_n1227, new_n1228, new_n1229,
    new_n1230, new_n1231, new_n1232, new_n1233, new_n1234, new_n1235,
    new_n1236, new_n1237, new_n1238, new_n1239, new_n1240, new_n1242,
    new_n1243, new_n1244, new_n1245, new_n1246, new_n1247, new_n1249,
    new_n1250, new_n1251, new_n1253, new_n1254, new_n1255, new_n1256,
    new_n1257, new_n1258, new_n1259, new_n1260, new_n1261, new_n1262,
    new_n1263, new_n1264, new_n1265, new_n1266, new_n1267, new_n1268,
    new_n1269, new_n1270, new_n1271, new_n1272, new_n1273, new_n1274,
    new_n1275, new_n1276, new_n1277, new_n1278, new_n1279, new_n1280,
    new_n1281, new_n1282, new_n1283, new_n1284, new_n1285, new_n1286,
    new_n1287, new_n1288, new_n1289, new_n1290, new_n1291, new_n1292,
    new_n1293, new_n1294, new_n1295, new_n1296, new_n1297, new_n1298,
    new_n1299, new_n1300, new_n1301, new_n1303, new_n1304, new_n1305,
    new_n1306, new_n1307, new_n1308, new_n1309, new_n1310, new_n1311,
    new_n1312, new_n1313, new_n1314, new_n1315;
  NOR4_X1   g0000(.A1(G50), .A2(G58), .A3(G68), .A4(G77), .ZN(G353));
  OAI21_X1  g0001(.A(G87), .B1(G97), .B2(G107), .ZN(G355));
  NAND2_X1  g0002(.A1(G1), .A2(G20), .ZN(new_n203));
  INV_X1    g0003(.A(G87), .ZN(new_n204));
  INV_X1    g0004(.A(G250), .ZN(new_n205));
  INV_X1    g0005(.A(G97), .ZN(new_n206));
  INV_X1    g0006(.A(G257), .ZN(new_n207));
  OAI22_X1  g0007(.A1(new_n204), .A2(new_n205), .B1(new_n206), .B2(new_n207), .ZN(new_n208));
  AOI21_X1  g0008(.A(new_n208), .B1(G68), .B2(G238), .ZN(new_n209));
  INV_X1    g0009(.A(G107), .ZN(new_n210));
  INV_X1    g0010(.A(G264), .ZN(new_n211));
  OAI21_X1  g0011(.A(new_n209), .B1(new_n210), .B2(new_n211), .ZN(new_n212));
  AOI21_X1  g0012(.A(new_n212), .B1(G116), .B2(G270), .ZN(new_n213));
  NAND2_X1  g0013(.A1(G50), .A2(G226), .ZN(new_n214));
  INV_X1    g0014(.A(G77), .ZN(new_n215));
  INV_X1    g0015(.A(G244), .ZN(new_n216));
  OAI211_X1 g0016(.A(new_n213), .B(new_n214), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g0017(.A(G58), .ZN(new_n218));
  INV_X1    g0018(.A(G232), .ZN(new_n219));
  NOR2_X1   g0019(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  OAI21_X1  g0020(.A(new_n203), .B1(new_n217), .B2(new_n220), .ZN(new_n221));
  XNOR2_X1  g0021(.A(new_n221), .B(KEYINPUT1), .ZN(new_n222));
  NOR2_X1   g0022(.A1(new_n203), .A2(G13), .ZN(new_n223));
  OAI211_X1 g0023(.A(new_n223), .B(G250), .C1(G257), .C2(G264), .ZN(new_n224));
  XOR2_X1   g0024(.A(new_n224), .B(KEYINPUT0), .Z(new_n225));
  INV_X1    g0025(.A(G68), .ZN(new_n226));
  NAND2_X1  g0026(.A1(new_n218), .A2(new_n226), .ZN(new_n227));
  NAND2_X1  g0027(.A1(new_n227), .A2(G50), .ZN(new_n228));
  INV_X1    g0028(.A(G20), .ZN(new_n229));
  NAND2_X1  g0029(.A1(G1), .A2(G13), .ZN(new_n230));
  NOR3_X1   g0030(.A1(new_n228), .A2(new_n229), .A3(new_n230), .ZN(new_n231));
  NOR3_X1   g0031(.A1(new_n222), .A2(new_n225), .A3(new_n231), .ZN(G361));
  XNOR2_X1  g0032(.A(G238), .B(G244), .ZN(new_n233));
  XNOR2_X1  g0033(.A(G226), .B(G232), .ZN(new_n234));
  XNOR2_X1  g0034(.A(new_n233), .B(new_n234), .ZN(new_n235));
  XOR2_X1   g0035(.A(KEYINPUT64), .B(KEYINPUT2), .Z(new_n236));
  XNOR2_X1  g0036(.A(new_n235), .B(new_n236), .ZN(new_n237));
  XNOR2_X1  g0037(.A(G250), .B(G257), .ZN(new_n238));
  XNOR2_X1  g0038(.A(new_n238), .B(new_n211), .ZN(new_n239));
  XNOR2_X1  g0039(.A(new_n239), .B(G270), .ZN(new_n240));
  XNOR2_X1  g0040(.A(new_n237), .B(new_n240), .ZN(G358));
  XOR2_X1   g0041(.A(G68), .B(G77), .Z(new_n242));
  XNOR2_X1  g0042(.A(G50), .B(G58), .ZN(new_n243));
  XNOR2_X1  g0043(.A(new_n242), .B(new_n243), .ZN(new_n244));
  XNOR2_X1  g0044(.A(G87), .B(G97), .ZN(new_n245));
  XNOR2_X1  g0045(.A(G107), .B(G116), .ZN(new_n246));
  XNOR2_X1  g0046(.A(new_n245), .B(new_n246), .ZN(new_n247));
  XOR2_X1   g0047(.A(new_n244), .B(new_n247), .Z(G351));
  INV_X1    g0048(.A(KEYINPUT22), .ZN(new_n249));
  NOR3_X1   g0049(.A1(new_n249), .A2(new_n204), .A3(G20), .ZN(new_n250));
  INV_X1    g0050(.A(G33), .ZN(new_n251));
  NAND2_X1  g0051(.A1(new_n251), .A2(KEYINPUT3), .ZN(new_n252));
  INV_X1    g0052(.A(KEYINPUT3), .ZN(new_n253));
  AND3_X1   g0053(.A1(new_n253), .A2(KEYINPUT71), .A3(G33), .ZN(new_n254));
  AOI21_X1  g0054(.A(KEYINPUT71), .B1(new_n253), .B2(G33), .ZN(new_n255));
  OAI211_X1 g0055(.A(new_n250), .B(new_n252), .C1(new_n254), .C2(new_n255), .ZN(new_n256));
  NOR2_X1   g0056(.A1(new_n204), .A2(G20), .ZN(new_n257));
  NAND2_X1  g0057(.A1(new_n253), .A2(G33), .ZN(new_n258));
  NAND3_X1  g0058(.A1(new_n257), .A2(new_n252), .A3(new_n258), .ZN(new_n259));
  NAND2_X1  g0059(.A1(new_n259), .A2(new_n249), .ZN(new_n260));
  INV_X1    g0060(.A(KEYINPUT84), .ZN(new_n261));
  NAND2_X1  g0061(.A1(G33), .A2(G116), .ZN(new_n262));
  OAI21_X1  g0062(.A(new_n261), .B1(new_n262), .B2(G20), .ZN(new_n263));
  NAND4_X1  g0063(.A1(new_n229), .A2(KEYINPUT84), .A3(G33), .A4(G116), .ZN(new_n264));
  NAND2_X1  g0064(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g0065(.A(KEYINPUT23), .ZN(new_n266));
  OAI21_X1  g0066(.A(new_n266), .B1(new_n229), .B2(G107), .ZN(new_n267));
  NAND3_X1  g0067(.A1(new_n210), .A2(KEYINPUT23), .A3(G20), .ZN(new_n268));
  NAND2_X1  g0068(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND4_X1  g0069(.A1(new_n256), .A2(new_n260), .A3(new_n265), .A4(new_n269), .ZN(new_n270));
  NAND2_X1  g0070(.A1(new_n270), .A2(KEYINPUT24), .ZN(new_n271));
  AOI22_X1  g0071(.A1(new_n259), .A2(new_n249), .B1(new_n267), .B2(new_n268), .ZN(new_n272));
  INV_X1    g0072(.A(KEYINPUT24), .ZN(new_n273));
  NAND4_X1  g0073(.A1(new_n272), .A2(new_n273), .A3(new_n256), .A4(new_n265), .ZN(new_n274));
  NAND2_X1  g0074(.A1(new_n271), .A2(new_n274), .ZN(new_n275));
  NAND3_X1  g0075(.A1(G1), .A2(G20), .A3(G33), .ZN(new_n276));
  NAND2_X1  g0076(.A1(new_n276), .A2(new_n230), .ZN(new_n277));
  NAND2_X1  g0077(.A1(new_n275), .A2(new_n277), .ZN(new_n278));
  INV_X1    g0078(.A(KEYINPUT85), .ZN(new_n279));
  NAND2_X1  g0079(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g0080(.A1(new_n275), .A2(KEYINPUT85), .A3(new_n277), .ZN(new_n281));
  INV_X1    g0081(.A(G1), .ZN(new_n282));
  NAND3_X1  g0082(.A1(new_n282), .A2(G13), .A3(G20), .ZN(new_n283));
  INV_X1    g0083(.A(KEYINPUT67), .ZN(new_n284));
  NAND2_X1  g0084(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  NAND4_X1  g0085(.A1(new_n282), .A2(KEYINPUT67), .A3(G13), .A4(G20), .ZN(new_n286));
  AND2_X1   g0086(.A1(new_n285), .A2(new_n286), .ZN(new_n287));
  INV_X1    g0087(.A(KEYINPUT25), .ZN(new_n288));
  OAI211_X1 g0088(.A(new_n287), .B(new_n210), .C1(KEYINPUT86), .C2(new_n288), .ZN(new_n289));
  AOI21_X1  g0089(.A(new_n289), .B1(KEYINPUT86), .B2(new_n288), .ZN(new_n290));
  AOI211_X1 g0090(.A(KEYINPUT86), .B(new_n288), .C1(new_n287), .C2(new_n210), .ZN(new_n291));
  NOR2_X1   g0091(.A1(new_n290), .A2(new_n291), .ZN(new_n292));
  AND3_X1   g0092(.A1(new_n280), .A2(new_n281), .A3(new_n292), .ZN(new_n293));
  INV_X1    g0093(.A(G41), .ZN(new_n294));
  OAI211_X1 g0094(.A(G1), .B(G13), .C1(new_n251), .C2(new_n294), .ZN(new_n295));
  NOR2_X1   g0095(.A1(new_n253), .A2(G33), .ZN(new_n296));
  INV_X1    g0096(.A(KEYINPUT71), .ZN(new_n297));
  OAI21_X1  g0097(.A(new_n297), .B1(new_n251), .B2(KEYINPUT3), .ZN(new_n298));
  NAND3_X1  g0098(.A1(new_n253), .A2(KEYINPUT71), .A3(G33), .ZN(new_n299));
  AOI21_X1  g0099(.A(new_n296), .B1(new_n298), .B2(new_n299), .ZN(new_n300));
  INV_X1    g0100(.A(G1698), .ZN(new_n301));
  NAND2_X1  g0101(.A1(new_n205), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g0102(.A1(new_n207), .A2(G1698), .ZN(new_n303));
  NAND3_X1  g0103(.A1(new_n300), .A2(new_n302), .A3(new_n303), .ZN(new_n304));
  NAND2_X1  g0104(.A1(G33), .A2(G294), .ZN(new_n305));
  AOI21_X1  g0105(.A(new_n295), .B1(new_n304), .B2(new_n305), .ZN(new_n306));
  AND2_X1   g0106(.A1(KEYINPUT5), .A2(G41), .ZN(new_n307));
  NOR2_X1   g0107(.A1(KEYINPUT5), .A2(G41), .ZN(new_n308));
  OAI211_X1 g0108(.A(new_n282), .B(G45), .C1(new_n307), .C2(new_n308), .ZN(new_n309));
  NAND2_X1  g0109(.A1(new_n309), .A2(new_n295), .ZN(new_n310));
  NOR2_X1   g0110(.A1(new_n310), .A2(new_n211), .ZN(new_n311));
  INV_X1    g0111(.A(G274), .ZN(new_n312));
  OR2_X1    g0112(.A1(new_n309), .A2(new_n312), .ZN(new_n313));
  INV_X1    g0113(.A(new_n313), .ZN(new_n314));
  NOR3_X1   g0114(.A1(new_n306), .A2(new_n311), .A3(new_n314), .ZN(new_n315));
  INV_X1    g0115(.A(G200), .ZN(new_n316));
  NOR2_X1   g0116(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g0117(.A(new_n317), .ZN(new_n318));
  INV_X1    g0118(.A(new_n315), .ZN(new_n319));
  INV_X1    g0119(.A(G190), .ZN(new_n320));
  NOR2_X1   g0120(.A1(new_n319), .A2(new_n320), .ZN(new_n321));
  INV_X1    g0121(.A(new_n321), .ZN(new_n322));
  INV_X1    g0122(.A(KEYINPUT66), .ZN(new_n323));
  XNOR2_X1  g0123(.A(new_n277), .B(new_n323), .ZN(new_n324));
  NOR2_X1   g0124(.A1(new_n324), .A2(new_n287), .ZN(new_n325));
  NAND2_X1  g0125(.A1(new_n282), .A2(G33), .ZN(new_n326));
  NAND2_X1  g0126(.A1(new_n325), .A2(new_n326), .ZN(new_n327));
  INV_X1    g0127(.A(new_n327), .ZN(new_n328));
  NAND2_X1  g0128(.A1(new_n328), .A2(G107), .ZN(new_n329));
  NAND4_X1  g0129(.A1(new_n293), .A2(new_n318), .A3(new_n322), .A4(new_n329), .ZN(new_n330));
  INV_X1    g0130(.A(KEYINPUT87), .ZN(new_n331));
  INV_X1    g0131(.A(G169), .ZN(new_n332));
  NOR2_X1   g0132(.A1(new_n315), .A2(new_n332), .ZN(new_n333));
  INV_X1    g0133(.A(G179), .ZN(new_n334));
  NOR4_X1   g0134(.A1(new_n306), .A2(new_n314), .A3(new_n311), .A4(new_n334), .ZN(new_n335));
  OAI21_X1  g0135(.A(new_n331), .B1(new_n333), .B2(new_n335), .ZN(new_n336));
  NAND2_X1  g0136(.A1(new_n315), .A2(G179), .ZN(new_n337));
  OAI211_X1 g0137(.A(new_n337), .B(KEYINPUT87), .C1(new_n315), .C2(new_n332), .ZN(new_n338));
  NAND2_X1  g0138(.A1(new_n336), .A2(new_n338), .ZN(new_n339));
  NAND4_X1  g0139(.A1(new_n280), .A2(new_n329), .A3(new_n281), .A4(new_n292), .ZN(new_n340));
  NAND2_X1  g0140(.A1(new_n339), .A2(new_n340), .ZN(new_n341));
  NAND2_X1  g0141(.A1(new_n298), .A2(new_n299), .ZN(new_n342));
  NAND2_X1  g0142(.A1(new_n207), .A2(new_n301), .ZN(new_n343));
  NAND2_X1  g0143(.A1(new_n211), .A2(G1698), .ZN(new_n344));
  NAND4_X1  g0144(.A1(new_n342), .A2(new_n252), .A3(new_n343), .A4(new_n344), .ZN(new_n345));
  NAND2_X1  g0145(.A1(new_n252), .A2(new_n258), .ZN(new_n346));
  NAND2_X1  g0146(.A1(new_n346), .A2(G303), .ZN(new_n347));
  NAND2_X1  g0147(.A1(new_n345), .A2(new_n347), .ZN(new_n348));
  INV_X1    g0148(.A(new_n295), .ZN(new_n349));
  NAND2_X1  g0149(.A1(new_n348), .A2(new_n349), .ZN(new_n350));
  INV_X1    g0150(.A(new_n310), .ZN(new_n351));
  NAND2_X1  g0151(.A1(new_n351), .A2(G270), .ZN(new_n352));
  NAND2_X1  g0152(.A1(new_n350), .A2(new_n352), .ZN(new_n353));
  INV_X1    g0153(.A(new_n353), .ZN(new_n354));
  NAND2_X1  g0154(.A1(G33), .A2(G283), .ZN(new_n355));
  OAI211_X1 g0155(.A(new_n355), .B(new_n229), .C1(G33), .C2(new_n206), .ZN(new_n356));
  INV_X1    g0156(.A(G116), .ZN(new_n357));
  NAND2_X1  g0157(.A1(new_n357), .A2(G20), .ZN(new_n358));
  NAND3_X1  g0158(.A1(new_n356), .A2(new_n277), .A3(new_n358), .ZN(new_n359));
  INV_X1    g0159(.A(KEYINPUT20), .ZN(new_n360));
  NAND2_X1  g0160(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  NAND4_X1  g0161(.A1(new_n356), .A2(new_n277), .A3(KEYINPUT20), .A4(new_n358), .ZN(new_n362));
  AOI22_X1  g0162(.A1(new_n361), .A2(new_n362), .B1(new_n287), .B2(new_n357), .ZN(new_n363));
  NAND2_X1  g0163(.A1(new_n285), .A2(new_n286), .ZN(new_n364));
  INV_X1    g0164(.A(new_n277), .ZN(new_n365));
  NAND4_X1  g0165(.A1(new_n364), .A2(G116), .A3(new_n365), .A4(new_n326), .ZN(new_n366));
  INV_X1    g0166(.A(KEYINPUT83), .ZN(new_n367));
  NAND2_X1  g0167(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  AOI21_X1  g0168(.A(new_n277), .B1(new_n285), .B2(new_n286), .ZN(new_n369));
  NAND4_X1  g0169(.A1(new_n369), .A2(KEYINPUT83), .A3(G116), .A4(new_n326), .ZN(new_n370));
  NAND3_X1  g0170(.A1(new_n363), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  NAND4_X1  g0171(.A1(new_n354), .A2(G179), .A3(new_n313), .A4(new_n371), .ZN(new_n372));
  NAND3_X1  g0172(.A1(new_n350), .A2(new_n313), .A3(new_n352), .ZN(new_n373));
  NAND2_X1  g0173(.A1(new_n373), .A2(G200), .ZN(new_n374));
  INV_X1    g0174(.A(new_n371), .ZN(new_n375));
  OAI211_X1 g0175(.A(new_n374), .B(new_n375), .C1(new_n320), .C2(new_n373), .ZN(new_n376));
  NAND4_X1  g0176(.A1(new_n373), .A2(new_n371), .A3(KEYINPUT21), .A4(G169), .ZN(new_n377));
  NAND3_X1  g0177(.A1(new_n373), .A2(new_n371), .A3(G169), .ZN(new_n378));
  INV_X1    g0178(.A(KEYINPUT21), .ZN(new_n379));
  NAND2_X1  g0179(.A1(new_n378), .A2(new_n379), .ZN(new_n380));
  AND4_X1   g0180(.A1(new_n372), .A2(new_n376), .A3(new_n377), .A4(new_n380), .ZN(new_n381));
  AND3_X1   g0181(.A1(new_n330), .A2(new_n341), .A3(new_n381), .ZN(new_n382));
  NOR2_X1   g0182(.A1(new_n229), .A2(G1), .ZN(new_n383));
  INV_X1    g0183(.A(new_n383), .ZN(new_n384));
  NAND3_X1  g0184(.A1(new_n325), .A2(G50), .A3(new_n384), .ZN(new_n385));
  INV_X1    g0185(.A(G50), .ZN(new_n386));
  NAND2_X1  g0186(.A1(new_n287), .A2(new_n386), .ZN(new_n387));
  NAND2_X1  g0187(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  INV_X1    g0188(.A(KEYINPUT68), .ZN(new_n389));
  NAND2_X1  g0189(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  NAND3_X1  g0190(.A1(new_n385), .A2(KEYINPUT68), .A3(new_n387), .ZN(new_n391));
  OAI21_X1  g0191(.A(G20), .B1(new_n227), .B2(G50), .ZN(new_n392));
  INV_X1    g0192(.A(G150), .ZN(new_n393));
  NAND2_X1  g0193(.A1(new_n229), .A2(new_n251), .ZN(new_n394));
  NAND2_X1  g0194(.A1(new_n229), .A2(G33), .ZN(new_n395));
  XNOR2_X1  g0195(.A(KEYINPUT8), .B(G58), .ZN(new_n396));
  OAI221_X1 g0196(.A(new_n392), .B1(new_n393), .B2(new_n394), .C1(new_n395), .C2(new_n396), .ZN(new_n397));
  AOI22_X1  g0197(.A1(new_n390), .A2(new_n391), .B1(new_n324), .B2(new_n397), .ZN(new_n398));
  NOR2_X1   g0198(.A1(new_n398), .A2(KEYINPUT9), .ZN(new_n399));
  INV_X1    g0199(.A(new_n399), .ZN(new_n400));
  XNOR2_X1  g0200(.A(KEYINPUT3), .B(G33), .ZN(new_n401));
  NAND3_X1  g0201(.A1(new_n401), .A2(G222), .A3(new_n301), .ZN(new_n402));
  XOR2_X1   g0202(.A(new_n402), .B(KEYINPUT65), .Z(new_n403));
  NAND2_X1  g0203(.A1(new_n401), .A2(G1698), .ZN(new_n404));
  INV_X1    g0204(.A(G223), .ZN(new_n405));
  OAI22_X1  g0205(.A1(new_n404), .A2(new_n405), .B1(new_n215), .B2(new_n401), .ZN(new_n406));
  OAI21_X1  g0206(.A(new_n349), .B1(new_n403), .B2(new_n406), .ZN(new_n407));
  OAI21_X1  g0207(.A(new_n282), .B1(G41), .B2(G45), .ZN(new_n408));
  NAND2_X1  g0208(.A1(new_n295), .A2(new_n408), .ZN(new_n409));
  INV_X1    g0209(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g0210(.A1(new_n410), .A2(G226), .ZN(new_n411));
  NOR2_X1   g0211(.A1(new_n408), .A2(new_n312), .ZN(new_n412));
  INV_X1    g0212(.A(new_n412), .ZN(new_n413));
  NAND3_X1  g0213(.A1(new_n407), .A2(new_n411), .A3(new_n413), .ZN(new_n414));
  NAND2_X1  g0214(.A1(new_n414), .A2(G200), .ZN(new_n415));
  NOR2_X1   g0215(.A1(new_n414), .A2(new_n320), .ZN(new_n416));
  AOI21_X1  g0216(.A(new_n416), .B1(new_n398), .B2(KEYINPUT9), .ZN(new_n417));
  NAND3_X1  g0217(.A1(new_n400), .A2(new_n415), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g0218(.A1(new_n418), .A2(KEYINPUT10), .ZN(new_n419));
  INV_X1    g0219(.A(KEYINPUT10), .ZN(new_n420));
  NAND4_X1  g0220(.A1(new_n400), .A2(new_n417), .A3(new_n420), .A4(new_n415), .ZN(new_n421));
  NAND2_X1  g0221(.A1(new_n419), .A2(new_n421), .ZN(new_n422));
  INV_X1    g0222(.A(new_n398), .ZN(new_n423));
  OR2_X1    g0223(.A1(new_n414), .A2(G179), .ZN(new_n424));
  NAND2_X1  g0224(.A1(new_n414), .A2(new_n332), .ZN(new_n425));
  NAND3_X1  g0225(.A1(new_n423), .A2(new_n424), .A3(new_n425), .ZN(new_n426));
  NAND2_X1  g0226(.A1(new_n422), .A2(new_n426), .ZN(new_n427));
  INV_X1    g0227(.A(G238), .ZN(new_n428));
  NOR2_X1   g0228(.A1(G226), .A2(G1698), .ZN(new_n429));
  AOI21_X1  g0229(.A(new_n429), .B1(new_n219), .B2(G1698), .ZN(new_n430));
  AOI22_X1  g0230(.A1(new_n430), .A2(new_n401), .B1(G33), .B2(G97), .ZN(new_n431));
  OAI221_X1 g0231(.A(new_n413), .B1(new_n428), .B2(new_n409), .C1(new_n431), .C2(new_n295), .ZN(new_n432));
  OR2_X1    g0232(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n433));
  INV_X1    g0233(.A(KEYINPUT70), .ZN(new_n434));
  NAND2_X1  g0234(.A1(new_n432), .A2(KEYINPUT13), .ZN(new_n435));
  NAND3_X1  g0235(.A1(new_n433), .A2(new_n434), .A3(new_n435), .ZN(new_n436));
  NAND3_X1  g0236(.A1(new_n432), .A2(KEYINPUT70), .A3(KEYINPUT13), .ZN(new_n437));
  NAND2_X1  g0237(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  OAI21_X1  g0238(.A(KEYINPUT14), .B1(new_n438), .B2(new_n332), .ZN(new_n439));
  INV_X1    g0239(.A(KEYINPUT14), .ZN(new_n440));
  NAND4_X1  g0240(.A1(new_n436), .A2(new_n440), .A3(G169), .A4(new_n437), .ZN(new_n441));
  NAND3_X1  g0241(.A1(new_n433), .A2(G179), .A3(new_n435), .ZN(new_n442));
  NAND3_X1  g0242(.A1(new_n439), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  NAND2_X1  g0243(.A1(new_n226), .A2(G20), .ZN(new_n444));
  OAI221_X1 g0244(.A(new_n444), .B1(new_n395), .B2(new_n215), .C1(new_n386), .C2(new_n394), .ZN(new_n445));
  AND2_X1   g0245(.A1(new_n324), .A2(new_n445), .ZN(new_n446));
  OR2_X1    g0246(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n447));
  NAND2_X1  g0247(.A1(new_n287), .A2(new_n226), .ZN(new_n448));
  XNOR2_X1  g0248(.A(new_n448), .B(KEYINPUT12), .ZN(new_n449));
  NAND2_X1  g0249(.A1(new_n446), .A2(KEYINPUT11), .ZN(new_n450));
  NAND3_X1  g0250(.A1(new_n369), .A2(G68), .A3(new_n384), .ZN(new_n451));
  NAND4_X1  g0251(.A1(new_n447), .A2(new_n449), .A3(new_n450), .A4(new_n451), .ZN(new_n452));
  NAND2_X1  g0252(.A1(new_n443), .A2(new_n452), .ZN(new_n453));
  INV_X1    g0253(.A(new_n453), .ZN(new_n454));
  NOR2_X1   g0254(.A1(new_n438), .A2(new_n316), .ZN(new_n455));
  AND3_X1   g0255(.A1(new_n433), .A2(G190), .A3(new_n435), .ZN(new_n456));
  NOR3_X1   g0256(.A1(new_n455), .A2(new_n452), .A3(new_n456), .ZN(new_n457));
  NOR3_X1   g0257(.A1(new_n427), .A2(new_n454), .A3(new_n457), .ZN(new_n458));
  XOR2_X1   g0258(.A(KEYINPUT15), .B(G87), .Z(new_n459));
  INV_X1    g0259(.A(new_n459), .ZN(new_n460));
  NOR2_X1   g0260(.A1(new_n460), .A2(new_n395), .ZN(new_n461));
  OAI22_X1  g0261(.A1(new_n396), .A2(new_n394), .B1(new_n229), .B2(new_n215), .ZN(new_n462));
  OAI21_X1  g0262(.A(new_n277), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g0263(.A1(new_n287), .A2(new_n215), .ZN(new_n464));
  NAND3_X1  g0264(.A1(new_n369), .A2(G77), .A3(new_n384), .ZN(new_n465));
  NAND3_X1  g0265(.A1(new_n463), .A2(new_n464), .A3(new_n465), .ZN(new_n466));
  NAND3_X1  g0266(.A1(new_n401), .A2(G232), .A3(new_n301), .ZN(new_n467));
  OAI221_X1 g0267(.A(new_n467), .B1(new_n210), .B2(new_n401), .C1(new_n404), .C2(new_n428), .ZN(new_n468));
  AOI21_X1  g0268(.A(new_n412), .B1(new_n468), .B2(new_n349), .ZN(new_n469));
  INV_X1    g0269(.A(KEYINPUT69), .ZN(new_n470));
  NAND2_X1  g0270(.A1(new_n410), .A2(G244), .ZN(new_n471));
  AND3_X1   g0271(.A1(new_n469), .A2(new_n470), .A3(new_n471), .ZN(new_n472));
  AOI21_X1  g0272(.A(new_n470), .B1(new_n469), .B2(new_n471), .ZN(new_n473));
  NOR2_X1   g0273(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  AOI21_X1  g0274(.A(new_n466), .B1(new_n474), .B2(G200), .ZN(new_n475));
  OAI21_X1  g0275(.A(G190), .B1(new_n472), .B2(new_n473), .ZN(new_n476));
  NAND2_X1  g0276(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  NAND4_X1  g0277(.A1(new_n342), .A2(G223), .A3(new_n301), .A4(new_n252), .ZN(new_n478));
  NAND2_X1  g0278(.A1(new_n478), .A2(KEYINPUT75), .ZN(new_n479));
  OAI21_X1  g0279(.A(new_n301), .B1(new_n405), .B2(KEYINPUT75), .ZN(new_n480));
  OAI211_X1 g0280(.A(new_n300), .B(new_n480), .C1(G226), .C2(new_n301), .ZN(new_n481));
  NOR2_X1   g0281(.A1(new_n251), .A2(new_n204), .ZN(new_n482));
  INV_X1    g0282(.A(new_n482), .ZN(new_n483));
  NAND3_X1  g0283(.A1(new_n479), .A2(new_n481), .A3(new_n483), .ZN(new_n484));
  NAND2_X1  g0284(.A1(new_n484), .A2(new_n349), .ZN(new_n485));
  AOI21_X1  g0285(.A(new_n412), .B1(new_n410), .B2(G232), .ZN(new_n486));
  NAND3_X1  g0286(.A1(new_n485), .A2(G190), .A3(new_n486), .ZN(new_n487));
  AOI21_X1  g0287(.A(new_n482), .B1(new_n478), .B2(KEYINPUT75), .ZN(new_n488));
  AOI21_X1  g0288(.A(new_n295), .B1(new_n488), .B2(new_n481), .ZN(new_n489));
  INV_X1    g0289(.A(new_n486), .ZN(new_n490));
  OAI21_X1  g0290(.A(G200), .B1(new_n489), .B2(new_n490), .ZN(new_n491));
  NOR2_X1   g0291(.A1(new_n396), .A2(new_n383), .ZN(new_n492));
  AOI22_X1  g0292(.A1(new_n325), .A2(new_n492), .B1(new_n287), .B2(new_n396), .ZN(new_n493));
  AND3_X1   g0293(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n494));
  INV_X1    g0294(.A(KEYINPUT17), .ZN(new_n495));
  NOR2_X1   g0295(.A1(new_n495), .A2(KEYINPUT76), .ZN(new_n496));
  NOR2_X1   g0296(.A1(KEYINPUT7), .A2(G20), .ZN(new_n497));
  AOI211_X1 g0297(.A(KEYINPUT72), .B(new_n296), .C1(new_n298), .C2(new_n299), .ZN(new_n498));
  INV_X1    g0298(.A(KEYINPUT72), .ZN(new_n499));
  AOI21_X1  g0299(.A(new_n499), .B1(new_n342), .B2(new_n252), .ZN(new_n500));
  OAI21_X1  g0300(.A(new_n497), .B1(new_n498), .B2(new_n500), .ZN(new_n501));
  OAI21_X1  g0301(.A(KEYINPUT7), .B1(new_n300), .B2(G20), .ZN(new_n502));
  NAND3_X1  g0302(.A1(new_n501), .A2(G68), .A3(new_n502), .ZN(new_n503));
  INV_X1    g0303(.A(G159), .ZN(new_n504));
  NOR2_X1   g0304(.A1(new_n394), .A2(new_n504), .ZN(new_n505));
  NAND2_X1  g0305(.A1(G58), .A2(G68), .ZN(new_n506));
  XNOR2_X1  g0306(.A(new_n506), .B(KEYINPUT73), .ZN(new_n507));
  NAND2_X1  g0307(.A1(new_n507), .A2(new_n227), .ZN(new_n508));
  AOI21_X1  g0308(.A(new_n505), .B1(new_n508), .B2(G20), .ZN(new_n509));
  NAND3_X1  g0309(.A1(new_n503), .A2(KEYINPUT16), .A3(new_n509), .ZN(new_n510));
  AND3_X1   g0310(.A1(new_n346), .A2(KEYINPUT7), .A3(new_n229), .ZN(new_n511));
  AOI21_X1  g0311(.A(KEYINPUT7), .B1(new_n346), .B2(new_n229), .ZN(new_n512));
  OAI21_X1  g0312(.A(G68), .B1(new_n511), .B2(new_n512), .ZN(new_n513));
  NAND2_X1  g0313(.A1(new_n513), .A2(new_n509), .ZN(new_n514));
  INV_X1    g0314(.A(KEYINPUT16), .ZN(new_n515));
  AOI21_X1  g0315(.A(new_n365), .B1(new_n514), .B2(new_n515), .ZN(new_n516));
  NAND3_X1  g0316(.A1(new_n510), .A2(new_n516), .A3(KEYINPUT74), .ZN(new_n517));
  INV_X1    g0317(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g0318(.A(KEYINPUT74), .B1(new_n510), .B2(new_n516), .ZN(new_n519));
  OAI211_X1 g0319(.A(new_n494), .B(new_n496), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  NAND3_X1  g0320(.A1(new_n487), .A2(new_n491), .A3(new_n493), .ZN(new_n521));
  NAND2_X1  g0321(.A1(new_n510), .A2(new_n516), .ZN(new_n522));
  INV_X1    g0322(.A(KEYINPUT74), .ZN(new_n523));
  NAND2_X1  g0323(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  AOI21_X1  g0324(.A(new_n521), .B1(new_n524), .B2(new_n517), .ZN(new_n525));
  XOR2_X1   g0325(.A(KEYINPUT76), .B(KEYINPUT17), .Z(new_n526));
  OAI21_X1  g0326(.A(new_n520), .B1(new_n525), .B2(new_n526), .ZN(new_n527));
  INV_X1    g0327(.A(KEYINPUT77), .ZN(new_n528));
  NAND2_X1  g0328(.A1(new_n527), .A2(new_n528), .ZN(new_n529));
  INV_X1    g0329(.A(KEYINPUT18), .ZN(new_n530));
  INV_X1    g0330(.A(new_n493), .ZN(new_n531));
  AOI21_X1  g0331(.A(new_n531), .B1(new_n524), .B2(new_n517), .ZN(new_n532));
  NAND3_X1  g0332(.A1(new_n485), .A2(G179), .A3(new_n486), .ZN(new_n533));
  OAI21_X1  g0333(.A(G169), .B1(new_n489), .B2(new_n490), .ZN(new_n534));
  NAND2_X1  g0334(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  INV_X1    g0335(.A(new_n535), .ZN(new_n536));
  OAI21_X1  g0336(.A(new_n530), .B1(new_n532), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g0337(.A(new_n493), .B1(new_n518), .B2(new_n519), .ZN(new_n538));
  NAND3_X1  g0338(.A1(new_n538), .A2(KEYINPUT18), .A3(new_n535), .ZN(new_n539));
  NAND2_X1  g0339(.A1(new_n537), .A2(new_n539), .ZN(new_n540));
  OAI211_X1 g0340(.A(new_n520), .B(KEYINPUT77), .C1(new_n525), .C2(new_n526), .ZN(new_n541));
  NAND3_X1  g0341(.A1(new_n529), .A2(new_n540), .A3(new_n541), .ZN(new_n542));
  NAND2_X1  g0342(.A1(new_n474), .A2(new_n332), .ZN(new_n543));
  OAI21_X1  g0343(.A(new_n334), .B1(new_n472), .B2(new_n473), .ZN(new_n544));
  NAND3_X1  g0344(.A1(new_n543), .A2(new_n466), .A3(new_n544), .ZN(new_n545));
  INV_X1    g0345(.A(new_n545), .ZN(new_n546));
  NOR2_X1   g0346(.A1(new_n542), .A2(new_n546), .ZN(new_n547));
  AND3_X1   g0347(.A1(new_n458), .A2(new_n477), .A3(new_n547), .ZN(new_n548));
  NAND3_X1  g0348(.A1(new_n300), .A2(new_n229), .A3(G68), .ZN(new_n549));
  INV_X1    g0349(.A(KEYINPUT19), .ZN(new_n550));
  NAND2_X1  g0350(.A1(G33), .A2(G97), .ZN(new_n551));
  OAI21_X1  g0351(.A(new_n550), .B1(new_n551), .B2(G20), .ZN(new_n552));
  NOR2_X1   g0352(.A1(new_n551), .A2(new_n550), .ZN(new_n553));
  NOR2_X1   g0353(.A1(new_n553), .A2(G20), .ZN(new_n554));
  NOR3_X1   g0354(.A1(G87), .A2(G97), .A3(G107), .ZN(new_n555));
  OAI211_X1 g0355(.A(new_n549), .B(new_n552), .C1(new_n554), .C2(new_n555), .ZN(new_n556));
  NAND2_X1  g0356(.A1(new_n556), .A2(new_n277), .ZN(new_n557));
  NAND2_X1  g0357(.A1(new_n287), .A2(new_n460), .ZN(new_n558));
  NAND2_X1  g0358(.A1(new_n557), .A2(new_n558), .ZN(new_n559));
  INV_X1    g0359(.A(new_n559), .ZN(new_n560));
  NAND2_X1  g0360(.A1(new_n328), .A2(new_n459), .ZN(new_n561));
  NAND2_X1  g0361(.A1(new_n560), .A2(new_n561), .ZN(new_n562));
  INV_X1    g0362(.A(KEYINPUT82), .ZN(new_n563));
  INV_X1    g0363(.A(G45), .ZN(new_n564));
  OAI21_X1  g0364(.A(new_n205), .B1(new_n564), .B2(G1), .ZN(new_n565));
  NAND3_X1  g0365(.A1(new_n282), .A2(new_n312), .A3(G45), .ZN(new_n566));
  NAND3_X1  g0366(.A1(new_n295), .A2(new_n565), .A3(new_n566), .ZN(new_n567));
  INV_X1    g0367(.A(KEYINPUT81), .ZN(new_n568));
  NAND2_X1  g0368(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND4_X1  g0369(.A1(new_n295), .A2(KEYINPUT81), .A3(new_n565), .A4(new_n566), .ZN(new_n570));
  NAND2_X1  g0370(.A1(new_n569), .A2(new_n570), .ZN(new_n571));
  INV_X1    g0371(.A(new_n571), .ZN(new_n572));
  NOR2_X1   g0372(.A1(G238), .A2(G1698), .ZN(new_n573));
  AOI21_X1  g0373(.A(new_n573), .B1(new_n216), .B2(G1698), .ZN(new_n574));
  NAND2_X1  g0374(.A1(new_n300), .A2(new_n574), .ZN(new_n575));
  AOI21_X1  g0375(.A(new_n295), .B1(new_n575), .B2(new_n262), .ZN(new_n576));
  OAI21_X1  g0376(.A(new_n563), .B1(new_n572), .B2(new_n576), .ZN(new_n577));
  AOI22_X1  g0377(.A1(new_n300), .A2(new_n574), .B1(G33), .B2(G116), .ZN(new_n578));
  OAI211_X1 g0378(.A(new_n571), .B(KEYINPUT82), .C1(new_n295), .C2(new_n578), .ZN(new_n579));
  NAND2_X1  g0379(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  NAND2_X1  g0380(.A1(new_n580), .A2(new_n334), .ZN(new_n581));
  NAND3_X1  g0381(.A1(new_n577), .A2(new_n332), .A3(new_n579), .ZN(new_n582));
  NAND3_X1  g0382(.A1(new_n562), .A2(new_n581), .A3(new_n582), .ZN(new_n583));
  NAND2_X1  g0383(.A1(new_n580), .A2(G190), .ZN(new_n584));
  NOR2_X1   g0384(.A1(new_n327), .A2(new_n204), .ZN(new_n585));
  NOR2_X1   g0385(.A1(new_n559), .A2(new_n585), .ZN(new_n586));
  NAND3_X1  g0386(.A1(new_n577), .A2(G200), .A3(new_n579), .ZN(new_n587));
  NAND3_X1  g0387(.A1(new_n584), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  AND2_X1   g0388(.A1(new_n583), .A2(new_n588), .ZN(new_n589));
  NAND4_X1  g0389(.A1(new_n252), .A2(new_n258), .A3(G250), .A4(G1698), .ZN(new_n590));
  NAND2_X1  g0390(.A1(new_n590), .A2(new_n355), .ZN(new_n591));
  AND2_X1   g0391(.A1(KEYINPUT4), .A2(G244), .ZN(new_n592));
  NAND4_X1  g0392(.A1(new_n252), .A2(new_n258), .A3(new_n592), .A4(new_n301), .ZN(new_n593));
  NAND2_X1  g0393(.A1(new_n593), .A2(KEYINPUT78), .ZN(new_n594));
  INV_X1    g0394(.A(KEYINPUT78), .ZN(new_n595));
  NAND4_X1  g0395(.A1(new_n401), .A2(new_n595), .A3(new_n301), .A4(new_n592), .ZN(new_n596));
  AOI21_X1  g0396(.A(new_n591), .B1(new_n594), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g0397(.A1(new_n300), .A2(G244), .A3(new_n301), .ZN(new_n598));
  INV_X1    g0398(.A(KEYINPUT4), .ZN(new_n599));
  NAND2_X1  g0399(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  AND3_X1   g0400(.A1(new_n597), .A2(KEYINPUT79), .A3(new_n600), .ZN(new_n601));
  AOI21_X1  g0401(.A(KEYINPUT79), .B1(new_n597), .B2(new_n600), .ZN(new_n602));
  OAI21_X1  g0402(.A(new_n349), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g0403(.A(new_n314), .B1(new_n351), .B2(G257), .ZN(new_n604));
  NAND2_X1  g0404(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g0405(.A1(new_n605), .A2(new_n320), .ZN(new_n606));
  AND3_X1   g0406(.A1(new_n325), .A2(G97), .A3(new_n326), .ZN(new_n607));
  NOR2_X1   g0407(.A1(new_n394), .A2(new_n215), .ZN(new_n608));
  INV_X1    g0408(.A(new_n608), .ZN(new_n609));
  OAI21_X1  g0409(.A(G107), .B1(new_n511), .B2(new_n512), .ZN(new_n610));
  NOR2_X1   g0410(.A1(new_n206), .A2(new_n210), .ZN(new_n611));
  NOR2_X1   g0411(.A1(G97), .A2(G107), .ZN(new_n612));
  NOR2_X1   g0412(.A1(new_n611), .A2(new_n612), .ZN(new_n613));
  NOR2_X1   g0413(.A1(new_n613), .A2(KEYINPUT6), .ZN(new_n614));
  NOR2_X1   g0414(.A1(new_n206), .A2(G107), .ZN(new_n615));
  AOI21_X1  g0415(.A(new_n614), .B1(KEYINPUT6), .B2(new_n615), .ZN(new_n616));
  OAI211_X1 g0416(.A(new_n609), .B(new_n610), .C1(new_n616), .C2(new_n229), .ZN(new_n617));
  AOI21_X1  g0417(.A(new_n607), .B1(new_n617), .B2(new_n277), .ZN(new_n618));
  NOR2_X1   g0418(.A1(new_n364), .A2(G97), .ZN(new_n619));
  INV_X1    g0419(.A(new_n619), .ZN(new_n620));
  NAND2_X1  g0420(.A1(new_n618), .A2(new_n620), .ZN(new_n621));
  NOR2_X1   g0421(.A1(new_n606), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g0422(.A1(new_n603), .A2(KEYINPUT80), .ZN(new_n623));
  INV_X1    g0423(.A(KEYINPUT80), .ZN(new_n624));
  OAI211_X1 g0424(.A(new_n624), .B(new_n349), .C1(new_n601), .C2(new_n602), .ZN(new_n625));
  NAND3_X1  g0425(.A1(new_n623), .A2(new_n604), .A3(new_n625), .ZN(new_n626));
  NAND2_X1  g0426(.A1(new_n626), .A2(G200), .ZN(new_n627));
  NAND4_X1  g0427(.A1(new_n623), .A2(new_n334), .A3(new_n604), .A4(new_n625), .ZN(new_n628));
  AOI22_X1  g0428(.A1(new_n605), .A2(new_n332), .B1(new_n620), .B2(new_n618), .ZN(new_n629));
  AOI22_X1  g0429(.A1(new_n622), .A2(new_n627), .B1(new_n628), .B2(new_n629), .ZN(new_n630));
  AND4_X1   g0430(.A1(new_n382), .A2(new_n548), .A3(new_n589), .A4(new_n630), .ZN(G372));
  NAND2_X1  g0431(.A1(new_n629), .A2(new_n628), .ZN(new_n632));
  NAND3_X1  g0432(.A1(new_n380), .A2(new_n372), .A3(new_n377), .ZN(new_n633));
  OAI21_X1  g0433(.A(new_n337), .B1(new_n332), .B2(new_n315), .ZN(new_n634));
  AOI21_X1  g0434(.A(new_n633), .B1(new_n340), .B2(new_n634), .ZN(new_n635));
  NOR3_X1   g0435(.A1(new_n340), .A2(new_n317), .A3(new_n321), .ZN(new_n636));
  OAI21_X1  g0436(.A(new_n632), .B1(new_n635), .B2(new_n636), .ZN(new_n637));
  INV_X1    g0437(.A(KEYINPUT26), .ZN(new_n638));
  NAND2_X1  g0438(.A1(new_n622), .A2(new_n627), .ZN(new_n639));
  AOI22_X1  g0439(.A1(new_n560), .A2(new_n561), .B1(new_n580), .B2(new_n334), .ZN(new_n640));
  OAI21_X1  g0440(.A(new_n332), .B1(new_n572), .B2(new_n576), .ZN(new_n641));
  NAND2_X1  g0441(.A1(new_n640), .A2(new_n641), .ZN(new_n642));
  NOR2_X1   g0442(.A1(new_n572), .A2(new_n576), .ZN(new_n643));
  OAI211_X1 g0443(.A(new_n584), .B(new_n586), .C1(new_n316), .C2(new_n643), .ZN(new_n644));
  AND2_X1   g0444(.A1(new_n642), .A2(new_n644), .ZN(new_n645));
  NAND4_X1  g0445(.A1(new_n637), .A2(new_n638), .A3(new_n639), .A4(new_n645), .ZN(new_n646));
  AND3_X1   g0446(.A1(new_n640), .A2(KEYINPUT88), .A3(new_n641), .ZN(new_n647));
  AOI21_X1  g0447(.A(KEYINPUT88), .B1(new_n640), .B2(new_n641), .ZN(new_n648));
  NOR2_X1   g0448(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  NAND4_X1  g0449(.A1(new_n629), .A2(new_n628), .A3(new_n583), .A4(new_n588), .ZN(new_n650));
  AOI21_X1  g0450(.A(new_n649), .B1(KEYINPUT26), .B2(new_n650), .ZN(new_n651));
  NAND2_X1  g0451(.A1(new_n646), .A2(new_n651), .ZN(new_n652));
  NAND2_X1  g0452(.A1(new_n548), .A2(new_n652), .ZN(new_n653));
  INV_X1    g0453(.A(new_n426), .ZN(new_n654));
  OAI21_X1  g0454(.A(new_n453), .B1(new_n545), .B2(new_n457), .ZN(new_n655));
  NAND3_X1  g0455(.A1(new_n655), .A2(new_n541), .A3(new_n529), .ZN(new_n656));
  NAND2_X1  g0456(.A1(new_n656), .A2(new_n540), .ZN(new_n657));
  AOI21_X1  g0457(.A(new_n654), .B1(new_n657), .B2(new_n422), .ZN(new_n658));
  NAND2_X1  g0458(.A1(new_n653), .A2(new_n658), .ZN(G369));
  INV_X1    g0459(.A(new_n381), .ZN(new_n660));
  INV_X1    g0460(.A(G13), .ZN(new_n661));
  NOR2_X1   g0461(.A1(new_n661), .A2(G20), .ZN(new_n662));
  INV_X1    g0462(.A(new_n662), .ZN(new_n663));
  OR3_X1    g0463(.A1(new_n663), .A2(KEYINPUT27), .A3(G1), .ZN(new_n664));
  OAI21_X1  g0464(.A(KEYINPUT27), .B1(new_n663), .B2(G1), .ZN(new_n665));
  NAND3_X1  g0465(.A1(new_n664), .A2(G213), .A3(new_n665), .ZN(new_n666));
  INV_X1    g0466(.A(G343), .ZN(new_n667));
  NOR2_X1   g0467(.A1(new_n666), .A2(new_n667), .ZN(new_n668));
  INV_X1    g0468(.A(new_n668), .ZN(new_n669));
  NOR2_X1   g0469(.A1(new_n375), .A2(new_n669), .ZN(new_n670));
  OAI21_X1  g0470(.A(KEYINPUT89), .B1(new_n660), .B2(new_n670), .ZN(new_n671));
  NAND2_X1  g0471(.A1(new_n633), .A2(new_n670), .ZN(new_n672));
  MUX2_X1   g0472(.A(KEYINPUT89), .B(new_n671), .S(new_n672), .Z(new_n673));
  AND2_X1   g0473(.A1(new_n673), .A2(G330), .ZN(new_n674));
  AND2_X1   g0474(.A1(new_n330), .A2(new_n341), .ZN(new_n675));
  NAND2_X1  g0475(.A1(new_n340), .A2(new_n668), .ZN(new_n676));
  NAND2_X1  g0476(.A1(new_n675), .A2(new_n676), .ZN(new_n677));
  OAI21_X1  g0477(.A(new_n677), .B1(new_n341), .B2(new_n669), .ZN(new_n678));
  NAND2_X1  g0478(.A1(new_n674), .A2(new_n678), .ZN(new_n679));
  INV_X1    g0479(.A(new_n633), .ZN(new_n680));
  NOR2_X1   g0480(.A1(new_n680), .A2(new_n668), .ZN(new_n681));
  AND2_X1   g0481(.A1(new_n675), .A2(new_n681), .ZN(new_n682));
  AND2_X1   g0482(.A1(new_n340), .A2(new_n634), .ZN(new_n683));
  AOI21_X1  g0483(.A(new_n682), .B1(new_n683), .B2(new_n669), .ZN(new_n684));
  NAND2_X1  g0484(.A1(new_n679), .A2(new_n684), .ZN(G399));
  NAND2_X1  g0485(.A1(new_n555), .A2(new_n357), .ZN(new_n686));
  XOR2_X1   g0486(.A(new_n686), .B(KEYINPUT90), .Z(new_n687));
  INV_X1    g0487(.A(new_n223), .ZN(new_n688));
  NOR2_X1   g0488(.A1(new_n688), .A2(G41), .ZN(new_n689));
  OR2_X1    g0489(.A1(new_n687), .A2(new_n689), .ZN(new_n690));
  INV_X1    g0490(.A(new_n689), .ZN(new_n691));
  OAI22_X1  g0491(.A1(new_n690), .A2(new_n282), .B1(new_n228), .B2(new_n691), .ZN(new_n692));
  XNOR2_X1  g0492(.A(new_n692), .B(KEYINPUT28), .ZN(new_n693));
  NAND2_X1  g0493(.A1(new_n652), .A2(new_n669), .ZN(new_n694));
  INV_X1    g0494(.A(KEYINPUT92), .ZN(new_n695));
  NAND2_X1  g0495(.A1(new_n694), .A2(new_n695), .ZN(new_n696));
  INV_X1    g0496(.A(KEYINPUT29), .ZN(new_n697));
  NAND3_X1  g0497(.A1(new_n652), .A2(KEYINPUT92), .A3(new_n669), .ZN(new_n698));
  NAND3_X1  g0498(.A1(new_n696), .A2(new_n697), .A3(new_n698), .ZN(new_n699));
  INV_X1    g0499(.A(KEYINPUT93), .ZN(new_n700));
  NAND2_X1  g0500(.A1(new_n699), .A2(new_n700), .ZN(new_n701));
  INV_X1    g0501(.A(KEYINPUT94), .ZN(new_n702));
  AND3_X1   g0502(.A1(new_n650), .A2(new_n702), .A3(new_n638), .ZN(new_n703));
  AOI21_X1  g0503(.A(new_n702), .B1(new_n650), .B2(new_n638), .ZN(new_n704));
  NAND3_X1  g0504(.A1(new_n642), .A2(KEYINPUT26), .A3(new_n644), .ZN(new_n705));
  NOR2_X1   g0505(.A1(new_n705), .A2(new_n632), .ZN(new_n706));
  NOR3_X1   g0506(.A1(new_n703), .A2(new_n704), .A3(new_n706), .ZN(new_n707));
  INV_X1    g0507(.A(new_n649), .ZN(new_n708));
  NAND2_X1  g0508(.A1(new_n341), .A2(new_n680), .ZN(new_n709));
  NAND3_X1  g0509(.A1(new_n709), .A2(new_n639), .A3(new_n632), .ZN(new_n710));
  NAND2_X1  g0510(.A1(new_n645), .A2(new_n330), .ZN(new_n711));
  OAI21_X1  g0511(.A(new_n708), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  OAI211_X1 g0512(.A(KEYINPUT29), .B(new_n669), .C1(new_n707), .C2(new_n712), .ZN(new_n713));
  NAND4_X1  g0513(.A1(new_n696), .A2(KEYINPUT93), .A3(new_n697), .A4(new_n698), .ZN(new_n714));
  NAND3_X1  g0514(.A1(new_n701), .A2(new_n713), .A3(new_n714), .ZN(new_n715));
  INV_X1    g0515(.A(KEYINPUT91), .ZN(new_n716));
  NAND4_X1  g0516(.A1(new_n603), .A2(new_n580), .A3(new_n335), .A4(new_n604), .ZN(new_n717));
  OAI21_X1  g0517(.A(new_n716), .B1(new_n717), .B2(new_n353), .ZN(new_n718));
  NAND2_X1  g0518(.A1(new_n718), .A2(KEYINPUT30), .ZN(new_n719));
  INV_X1    g0519(.A(KEYINPUT30), .ZN(new_n720));
  OAI211_X1 g0520(.A(new_n716), .B(new_n720), .C1(new_n717), .C2(new_n353), .ZN(new_n721));
  NOR2_X1   g0521(.A1(new_n643), .A2(G179), .ZN(new_n722));
  NAND4_X1  g0522(.A1(new_n626), .A2(new_n319), .A3(new_n373), .A4(new_n722), .ZN(new_n723));
  NAND3_X1  g0523(.A1(new_n719), .A2(new_n721), .A3(new_n723), .ZN(new_n724));
  NAND2_X1  g0524(.A1(new_n724), .A2(new_n668), .ZN(new_n725));
  INV_X1    g0525(.A(KEYINPUT31), .ZN(new_n726));
  NAND2_X1  g0526(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND4_X1  g0527(.A1(new_n382), .A2(new_n589), .A3(new_n630), .A4(new_n669), .ZN(new_n728));
  NAND3_X1  g0528(.A1(new_n724), .A2(KEYINPUT31), .A3(new_n668), .ZN(new_n729));
  NAND3_X1  g0529(.A1(new_n727), .A2(new_n728), .A3(new_n729), .ZN(new_n730));
  AND2_X1   g0530(.A1(new_n730), .A2(G330), .ZN(new_n731));
  INV_X1    g0531(.A(new_n731), .ZN(new_n732));
  AND2_X1   g0532(.A1(new_n715), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g0533(.A(new_n693), .B1(new_n733), .B2(G1), .ZN(G364));
  NOR2_X1   g0534(.A1(new_n673), .A2(G330), .ZN(new_n735));
  INV_X1    g0535(.A(new_n735), .ZN(new_n736));
  AOI21_X1  g0536(.A(new_n674), .B1(new_n736), .B2(KEYINPUT95), .ZN(new_n737));
  AOI21_X1  g0537(.A(new_n282), .B1(new_n662), .B2(G45), .ZN(new_n738));
  INV_X1    g0538(.A(new_n738), .ZN(new_n739));
  NOR2_X1   g0539(.A1(new_n689), .A2(new_n739), .ZN(new_n740));
  INV_X1    g0540(.A(new_n740), .ZN(new_n741));
  OAI211_X1 g0541(.A(new_n737), .B(new_n741), .C1(KEYINPUT95), .C2(new_n736), .ZN(new_n742));
  NOR2_X1   g0542(.A1(new_n229), .A2(new_n334), .ZN(new_n743));
  NAND2_X1  g0543(.A1(new_n743), .A2(G200), .ZN(new_n744));
  NOR2_X1   g0544(.A1(new_n744), .A2(new_n320), .ZN(new_n745));
  INV_X1    g0545(.A(new_n745), .ZN(new_n746));
  NOR3_X1   g0546(.A1(new_n320), .A2(G179), .A3(G200), .ZN(new_n747));
  NOR2_X1   g0547(.A1(new_n747), .A2(new_n229), .ZN(new_n748));
  OAI22_X1  g0548(.A1(new_n746), .A2(new_n386), .B1(new_n206), .B2(new_n748), .ZN(new_n749));
  NAND3_X1  g0549(.A1(new_n743), .A2(G190), .A3(new_n316), .ZN(new_n750));
  OAI21_X1  g0550(.A(new_n401), .B1(new_n750), .B2(new_n218), .ZN(new_n751));
  OR2_X1    g0551(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NOR2_X1   g0552(.A1(new_n316), .A2(G179), .ZN(new_n753));
  XNOR2_X1  g0553(.A(new_n753), .B(KEYINPUT98), .ZN(new_n754));
  NAND2_X1  g0554(.A1(new_n754), .A2(G20), .ZN(new_n755));
  NOR2_X1   g0555(.A1(new_n755), .A2(G190), .ZN(new_n756));
  INV_X1    g0556(.A(new_n756), .ZN(new_n757));
  NOR2_X1   g0557(.A1(new_n757), .A2(new_n210), .ZN(new_n758));
  NOR2_X1   g0558(.A1(new_n755), .A2(new_n320), .ZN(new_n759));
  AOI21_X1  g0559(.A(new_n758), .B1(G87), .B2(new_n759), .ZN(new_n760));
  INV_X1    g0560(.A(KEYINPUT32), .ZN(new_n761));
  NOR2_X1   g0561(.A1(G190), .A2(G200), .ZN(new_n762));
  NAND3_X1  g0562(.A1(new_n762), .A2(G20), .A3(new_n334), .ZN(new_n763));
  NOR2_X1   g0563(.A1(new_n763), .A2(new_n504), .ZN(new_n764));
  OAI21_X1  g0564(.A(new_n760), .B1(new_n761), .B2(new_n764), .ZN(new_n765));
  AOI211_X1 g0565(.A(new_n752), .B(new_n765), .C1(new_n761), .C2(new_n764), .ZN(new_n766));
  NOR2_X1   g0566(.A1(new_n744), .A2(G190), .ZN(new_n767));
  INV_X1    g0567(.A(new_n767), .ZN(new_n768));
  NAND2_X1  g0568(.A1(new_n743), .A2(new_n762), .ZN(new_n769));
  OAI221_X1 g0569(.A(new_n766), .B1(new_n226), .B2(new_n768), .C1(new_n215), .C2(new_n769), .ZN(new_n770));
  INV_X1    g0570(.A(G294), .ZN(new_n771));
  NOR2_X1   g0571(.A1(new_n748), .A2(new_n771), .ZN(new_n772));
  AND2_X1   g0572(.A1(new_n763), .A2(KEYINPUT99), .ZN(new_n773));
  NOR2_X1   g0573(.A1(new_n763), .A2(KEYINPUT99), .ZN(new_n774));
  NOR2_X1   g0574(.A1(new_n773), .A2(new_n774), .ZN(new_n775));
  INV_X1    g0575(.A(new_n775), .ZN(new_n776));
  AOI21_X1  g0576(.A(new_n401), .B1(new_n776), .B2(G329), .ZN(new_n777));
  INV_X1    g0577(.A(G311), .ZN(new_n778));
  OAI21_X1  g0578(.A(new_n777), .B1(new_n778), .B2(new_n769), .ZN(new_n779));
  XNOR2_X1  g0579(.A(KEYINPUT33), .B(G317), .ZN(new_n780));
  AOI21_X1  g0580(.A(new_n779), .B1(new_n767), .B2(new_n780), .ZN(new_n781));
  INV_X1    g0581(.A(new_n750), .ZN(new_n782));
  NAND2_X1  g0582(.A1(new_n782), .A2(G322), .ZN(new_n783));
  AOI22_X1  g0583(.A1(G283), .A2(new_n756), .B1(new_n759), .B2(G303), .ZN(new_n784));
  NAND2_X1  g0584(.A1(new_n745), .A2(G326), .ZN(new_n785));
  NAND4_X1  g0585(.A1(new_n781), .A2(new_n783), .A3(new_n784), .A4(new_n785), .ZN(new_n786));
  OAI21_X1  g0586(.A(new_n770), .B1(new_n772), .B2(new_n786), .ZN(new_n787));
  OAI21_X1  g0587(.A(G20), .B1(KEYINPUT96), .B2(G169), .ZN(new_n788));
  INV_X1    g0588(.A(new_n788), .ZN(new_n789));
  NAND2_X1  g0589(.A1(KEYINPUT96), .A2(G169), .ZN(new_n790));
  AOI21_X1  g0590(.A(new_n230), .B1(new_n789), .B2(new_n790), .ZN(new_n791));
  NAND2_X1  g0591(.A1(new_n787), .A2(new_n791), .ZN(new_n792));
  NOR2_X1   g0592(.A1(new_n688), .A2(new_n346), .ZN(new_n793));
  NAND2_X1  g0593(.A1(new_n793), .A2(G355), .ZN(new_n794));
  OR2_X1    g0594(.A1(new_n498), .A2(new_n500), .ZN(new_n795));
  INV_X1    g0595(.A(new_n795), .ZN(new_n796));
  NOR2_X1   g0596(.A1(new_n796), .A2(new_n688), .ZN(new_n797));
  OAI21_X1  g0597(.A(new_n797), .B1(G45), .B2(new_n228), .ZN(new_n798));
  NOR2_X1   g0598(.A1(new_n244), .A2(new_n564), .ZN(new_n799));
  OAI221_X1 g0599(.A(new_n794), .B1(G116), .B2(new_n223), .C1(new_n798), .C2(new_n799), .ZN(new_n800));
  NOR2_X1   g0600(.A1(G13), .A2(G33), .ZN(new_n801));
  INV_X1    g0601(.A(new_n801), .ZN(new_n802));
  NOR2_X1   g0602(.A1(new_n802), .A2(G20), .ZN(new_n803));
  NOR2_X1   g0603(.A1(new_n791), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g0604(.A(new_n741), .B1(new_n800), .B2(new_n804), .ZN(new_n805));
  XOR2_X1   g0605(.A(new_n805), .B(KEYINPUT97), .Z(new_n806));
  INV_X1    g0606(.A(new_n803), .ZN(new_n807));
  OAI211_X1 g0607(.A(new_n792), .B(new_n806), .C1(new_n673), .C2(new_n807), .ZN(new_n808));
  NAND2_X1  g0608(.A1(new_n742), .A2(new_n808), .ZN(G396));
  NAND4_X1  g0609(.A1(new_n543), .A2(new_n466), .A3(new_n544), .A4(new_n669), .ZN(new_n810));
  AOI22_X1  g0610(.A1(new_n475), .A2(new_n476), .B1(new_n466), .B2(new_n668), .ZN(new_n811));
  OAI21_X1  g0611(.A(new_n810), .B1(new_n811), .B2(new_n546), .ZN(new_n812));
  NAND3_X1  g0612(.A1(new_n696), .A2(new_n698), .A3(new_n812), .ZN(new_n813));
  INV_X1    g0613(.A(new_n812), .ZN(new_n814));
  NAND3_X1  g0614(.A1(new_n652), .A2(new_n814), .A3(new_n669), .ZN(new_n815));
  NAND2_X1  g0615(.A1(new_n813), .A2(new_n815), .ZN(new_n816));
  OAI21_X1  g0616(.A(new_n741), .B1(new_n816), .B2(new_n732), .ZN(new_n817));
  XNOR2_X1  g0617(.A(new_n817), .B(KEYINPUT100), .ZN(new_n818));
  NAND2_X1  g0618(.A1(new_n816), .A2(new_n732), .ZN(new_n819));
  NAND2_X1  g0619(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  AOI22_X1  g0620(.A1(G150), .A2(new_n767), .B1(new_n782), .B2(G143), .ZN(new_n821));
  INV_X1    g0621(.A(G137), .ZN(new_n822));
  OAI221_X1 g0622(.A(new_n821), .B1(new_n822), .B2(new_n746), .C1(new_n504), .C2(new_n769), .ZN(new_n823));
  XNOR2_X1  g0623(.A(new_n823), .B(KEYINPUT34), .ZN(new_n824));
  NAND2_X1  g0624(.A1(new_n776), .A2(G132), .ZN(new_n825));
  INV_X1    g0625(.A(new_n748), .ZN(new_n826));
  AOI22_X1  g0626(.A1(new_n756), .A2(G68), .B1(G58), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g0627(.A1(new_n824), .A2(new_n796), .A3(new_n825), .A4(new_n827), .ZN(new_n828));
  INV_X1    g0628(.A(new_n759), .ZN(new_n829));
  NOR2_X1   g0629(.A1(new_n829), .A2(new_n386), .ZN(new_n830));
  OAI22_X1  g0630(.A1(new_n204), .A2(new_n757), .B1(new_n829), .B2(new_n210), .ZN(new_n831));
  INV_X1    g0631(.A(G303), .ZN(new_n832));
  OAI22_X1  g0632(.A1(new_n746), .A2(new_n832), .B1(new_n206), .B2(new_n748), .ZN(new_n833));
  INV_X1    g0633(.A(G283), .ZN(new_n834));
  OAI221_X1 g0634(.A(new_n346), .B1(new_n768), .B2(new_n834), .C1(new_n775), .C2(new_n778), .ZN(new_n835));
  NOR3_X1   g0635(.A1(new_n831), .A2(new_n833), .A3(new_n835), .ZN(new_n836));
  OAI21_X1  g0636(.A(new_n836), .B1(new_n771), .B2(new_n750), .ZN(new_n837));
  NOR2_X1   g0637(.A1(new_n769), .A2(new_n357), .ZN(new_n838));
  OAI22_X1  g0638(.A1(new_n828), .A2(new_n830), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  AOI21_X1  g0639(.A(new_n741), .B1(new_n839), .B2(new_n791), .ZN(new_n840));
  NOR2_X1   g0640(.A1(new_n791), .A2(new_n801), .ZN(new_n841));
  INV_X1    g0641(.A(new_n841), .ZN(new_n842));
  OAI221_X1 g0642(.A(new_n840), .B1(G77), .B2(new_n842), .C1(new_n814), .C2(new_n802), .ZN(new_n843));
  NAND2_X1  g0643(.A1(new_n820), .A2(new_n843), .ZN(G384));
  INV_X1    g0644(.A(KEYINPUT40), .ZN(new_n845));
  INV_X1    g0645(.A(new_n666), .ZN(new_n846));
  NAND2_X1  g0646(.A1(new_n503), .A2(new_n509), .ZN(new_n847));
  NAND2_X1  g0647(.A1(new_n515), .A2(KEYINPUT103), .ZN(new_n848));
  XNOR2_X1  g0648(.A(new_n847), .B(new_n848), .ZN(new_n849));
  AOI21_X1  g0649(.A(new_n531), .B1(new_n849), .B2(new_n324), .ZN(new_n850));
  INV_X1    g0650(.A(new_n850), .ZN(new_n851));
  NAND3_X1  g0651(.A1(new_n542), .A2(new_n846), .A3(new_n851), .ZN(new_n852));
  OAI21_X1  g0652(.A(new_n494), .B1(new_n518), .B2(new_n519), .ZN(new_n853));
  NOR2_X1   g0653(.A1(new_n535), .A2(new_n846), .ZN(new_n854));
  OAI21_X1  g0654(.A(new_n853), .B1(new_n850), .B2(new_n854), .ZN(new_n855));
  NAND2_X1  g0655(.A1(new_n855), .A2(KEYINPUT37), .ZN(new_n856));
  OAI21_X1  g0656(.A(new_n853), .B1(new_n532), .B2(new_n854), .ZN(new_n857));
  OAI21_X1  g0657(.A(new_n856), .B1(KEYINPUT37), .B2(new_n857), .ZN(new_n858));
  AND3_X1   g0658(.A1(new_n852), .A2(KEYINPUT38), .A3(new_n858), .ZN(new_n859));
  AOI21_X1  g0659(.A(KEYINPUT38), .B1(new_n852), .B2(new_n858), .ZN(new_n860));
  NOR2_X1   g0660(.A1(new_n859), .A2(new_n860), .ZN(new_n861));
  NAND2_X1  g0661(.A1(new_n730), .A2(KEYINPUT104), .ZN(new_n862));
  NAND2_X1  g0662(.A1(new_n454), .A2(new_n668), .ZN(new_n863));
  INV_X1    g0663(.A(new_n457), .ZN(new_n864));
  NAND2_X1  g0664(.A1(new_n452), .A2(new_n668), .ZN(new_n865));
  NAND3_X1  g0665(.A1(new_n453), .A2(new_n864), .A3(new_n865), .ZN(new_n866));
  AOI21_X1  g0666(.A(new_n812), .B1(new_n863), .B2(new_n866), .ZN(new_n867));
  INV_X1    g0667(.A(KEYINPUT104), .ZN(new_n868));
  NAND4_X1  g0668(.A1(new_n727), .A2(new_n728), .A3(new_n868), .A4(new_n729), .ZN(new_n869));
  NAND3_X1  g0669(.A1(new_n862), .A2(new_n867), .A3(new_n869), .ZN(new_n870));
  OAI21_X1  g0670(.A(new_n845), .B1(new_n861), .B2(new_n870), .ZN(new_n871));
  INV_X1    g0671(.A(new_n870), .ZN(new_n872));
  INV_X1    g0672(.A(KEYINPUT38), .ZN(new_n873));
  INV_X1    g0673(.A(new_n527), .ZN(new_n874));
  AOI211_X1 g0674(.A(new_n532), .B(new_n666), .C1(new_n540), .C2(new_n874), .ZN(new_n875));
  XNOR2_X1  g0675(.A(new_n857), .B(KEYINPUT37), .ZN(new_n876));
  INV_X1    g0676(.A(new_n876), .ZN(new_n877));
  OAI21_X1  g0677(.A(new_n873), .B1(new_n875), .B2(new_n877), .ZN(new_n878));
  NAND3_X1  g0678(.A1(new_n852), .A2(new_n858), .A3(KEYINPUT38), .ZN(new_n879));
  AOI21_X1  g0679(.A(new_n845), .B1(new_n878), .B2(new_n879), .ZN(new_n880));
  NAND2_X1  g0680(.A1(new_n872), .A2(new_n880), .ZN(new_n881));
  NAND3_X1  g0681(.A1(new_n871), .A2(new_n881), .A3(G330), .ZN(new_n882));
  AND2_X1   g0682(.A1(new_n862), .A2(new_n869), .ZN(new_n883));
  NAND3_X1  g0683(.A1(new_n548), .A2(G330), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g0684(.A1(new_n882), .A2(new_n884), .ZN(new_n885));
  NAND4_X1  g0685(.A1(new_n871), .A2(new_n548), .A3(new_n883), .A4(new_n881), .ZN(new_n886));
  NAND2_X1  g0686(.A1(new_n885), .A2(new_n886), .ZN(new_n887));
  INV_X1    g0687(.A(KEYINPUT102), .ZN(new_n888));
  AOI211_X1 g0688(.A(new_n668), .B(new_n812), .C1(new_n646), .C2(new_n651), .ZN(new_n889));
  INV_X1    g0689(.A(new_n810), .ZN(new_n890));
  OAI21_X1  g0690(.A(new_n888), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  NAND3_X1  g0691(.A1(new_n815), .A2(KEYINPUT102), .A3(new_n810), .ZN(new_n892));
  NAND2_X1  g0692(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND2_X1  g0693(.A1(new_n852), .A2(new_n858), .ZN(new_n894));
  NAND2_X1  g0694(.A1(new_n894), .A2(new_n873), .ZN(new_n895));
  NAND2_X1  g0695(.A1(new_n895), .A2(new_n879), .ZN(new_n896));
  NAND2_X1  g0696(.A1(new_n863), .A2(new_n866), .ZN(new_n897));
  NAND3_X1  g0697(.A1(new_n893), .A2(new_n896), .A3(new_n897), .ZN(new_n898));
  INV_X1    g0698(.A(KEYINPUT39), .ZN(new_n899));
  INV_X1    g0699(.A(new_n540), .ZN(new_n900));
  OAI211_X1 g0700(.A(new_n538), .B(new_n846), .C1(new_n900), .C2(new_n527), .ZN(new_n901));
  AOI21_X1  g0701(.A(KEYINPUT38), .B1(new_n901), .B2(new_n876), .ZN(new_n902));
  OAI21_X1  g0702(.A(new_n899), .B1(new_n859), .B2(new_n902), .ZN(new_n903));
  NAND3_X1  g0703(.A1(new_n895), .A2(KEYINPUT39), .A3(new_n879), .ZN(new_n904));
  NOR2_X1   g0704(.A1(new_n453), .A2(new_n668), .ZN(new_n905));
  NAND3_X1  g0705(.A1(new_n903), .A2(new_n904), .A3(new_n905), .ZN(new_n906));
  NAND2_X1  g0706(.A1(new_n900), .A2(new_n666), .ZN(new_n907));
  AND3_X1   g0707(.A1(new_n898), .A2(new_n906), .A3(new_n907), .ZN(new_n908));
  NAND4_X1  g0708(.A1(new_n701), .A2(new_n548), .A3(new_n713), .A4(new_n714), .ZN(new_n909));
  NAND2_X1  g0709(.A1(new_n909), .A2(new_n658), .ZN(new_n910));
  XOR2_X1   g0710(.A(new_n908), .B(new_n910), .Z(new_n911));
  OAI21_X1  g0711(.A(new_n887), .B1(new_n911), .B2(KEYINPUT105), .ZN(new_n912));
  NAND2_X1  g0712(.A1(new_n911), .A2(KEYINPUT105), .ZN(new_n913));
  XOR2_X1   g0713(.A(new_n912), .B(new_n913), .Z(new_n914));
  OAI21_X1  g0714(.A(new_n914), .B1(new_n282), .B2(new_n662), .ZN(new_n915));
  INV_X1    g0715(.A(KEYINPUT35), .ZN(new_n916));
  AOI211_X1 g0716(.A(new_n229), .B(new_n230), .C1(new_n616), .C2(new_n916), .ZN(new_n917));
  OAI211_X1 g0717(.A(new_n917), .B(G116), .C1(new_n916), .C2(new_n616), .ZN(new_n918));
  XNOR2_X1  g0718(.A(new_n918), .B(KEYINPUT36), .ZN(new_n919));
  NAND4_X1  g0719(.A1(new_n507), .A2(G50), .A3(G77), .A4(new_n227), .ZN(new_n920));
  XNOR2_X1  g0720(.A(new_n920), .B(KEYINPUT101), .ZN(new_n921));
  OAI21_X1  g0721(.A(new_n921), .B1(G50), .B2(new_n226), .ZN(new_n922));
  NAND3_X1  g0722(.A1(new_n922), .A2(G1), .A3(new_n661), .ZN(new_n923));
  NAND3_X1  g0723(.A1(new_n915), .A2(new_n919), .A3(new_n923), .ZN(G367));
  OAI21_X1  g0724(.A(new_n668), .B1(new_n559), .B2(new_n585), .ZN(new_n925));
  NOR2_X1   g0725(.A1(new_n708), .A2(new_n925), .ZN(new_n926));
  AOI21_X1  g0726(.A(new_n926), .B1(new_n645), .B2(new_n925), .ZN(new_n927));
  NAND2_X1  g0727(.A1(new_n927), .A2(new_n803), .ZN(new_n928));
  INV_X1    g0728(.A(G143), .ZN(new_n929));
  OAI22_X1  g0729(.A1(new_n829), .A2(new_n218), .B1(new_n929), .B2(new_n746), .ZN(new_n930));
  NOR2_X1   g0730(.A1(new_n757), .A2(new_n215), .ZN(new_n931));
  OAI22_X1  g0731(.A1(new_n750), .A2(new_n393), .B1(new_n769), .B2(new_n386), .ZN(new_n932));
  OAI21_X1  g0732(.A(new_n401), .B1(new_n763), .B2(new_n822), .ZN(new_n933));
  NOR4_X1   g0733(.A1(new_n930), .A2(new_n931), .A3(new_n932), .A4(new_n933), .ZN(new_n934));
  OAI221_X1 g0734(.A(new_n934), .B1(new_n226), .B2(new_n748), .C1(new_n504), .C2(new_n768), .ZN(new_n935));
  AOI22_X1  g0735(.A1(G107), .A2(new_n826), .B1(new_n767), .B2(G294), .ZN(new_n936));
  OAI221_X1 g0736(.A(new_n936), .B1(new_n832), .B2(new_n750), .C1(new_n778), .C2(new_n746), .ZN(new_n937));
  AOI21_X1  g0737(.A(new_n937), .B1(G97), .B2(new_n756), .ZN(new_n938));
  INV_X1    g0738(.A(new_n763), .ZN(new_n939));
  AOI21_X1  g0739(.A(new_n796), .B1(G317), .B2(new_n939), .ZN(new_n940));
  OAI211_X1 g0740(.A(new_n938), .B(new_n940), .C1(new_n834), .C2(new_n769), .ZN(new_n941));
  NAND2_X1  g0741(.A1(new_n759), .A2(G116), .ZN(new_n942));
  XOR2_X1   g0742(.A(new_n942), .B(KEYINPUT46), .Z(new_n943));
  OAI21_X1  g0743(.A(new_n935), .B1(new_n941), .B2(new_n943), .ZN(new_n944));
  XNOR2_X1  g0744(.A(new_n944), .B(KEYINPUT47), .ZN(new_n945));
  NAND2_X1  g0745(.A1(new_n945), .A2(new_n791), .ZN(new_n946));
  INV_X1    g0746(.A(new_n797), .ZN(new_n947));
  OAI221_X1 g0747(.A(new_n804), .B1(new_n223), .B2(new_n460), .C1(new_n947), .C2(new_n240), .ZN(new_n948));
  NAND4_X1  g0748(.A1(new_n928), .A2(new_n740), .A3(new_n946), .A4(new_n948), .ZN(new_n949));
  NAND2_X1  g0749(.A1(new_n621), .A2(new_n668), .ZN(new_n950));
  NAND2_X1  g0750(.A1(new_n630), .A2(new_n950), .ZN(new_n951));
  OAI21_X1  g0751(.A(new_n951), .B1(new_n632), .B2(new_n669), .ZN(new_n952));
  NOR2_X1   g0752(.A1(new_n684), .A2(new_n952), .ZN(new_n953));
  XNOR2_X1  g0753(.A(new_n953), .B(KEYINPUT44), .ZN(new_n954));
  NAND2_X1  g0754(.A1(new_n684), .A2(new_n952), .ZN(new_n955));
  INV_X1    g0755(.A(KEYINPUT45), .ZN(new_n956));
  XNOR2_X1  g0756(.A(new_n955), .B(new_n956), .ZN(new_n957));
  NAND2_X1  g0757(.A1(new_n954), .A2(new_n957), .ZN(new_n958));
  INV_X1    g0758(.A(new_n679), .ZN(new_n959));
  NAND2_X1  g0759(.A1(new_n958), .A2(new_n959), .ZN(new_n960));
  NAND3_X1  g0760(.A1(new_n954), .A2(new_n679), .A3(new_n957), .ZN(new_n961));
  NAND2_X1  g0761(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  OR2_X1    g0762(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n963));
  NAND2_X1  g0763(.A1(new_n682), .A2(KEYINPUT106), .ZN(new_n964));
  OAI211_X1 g0764(.A(new_n963), .B(new_n964), .C1(new_n678), .C2(new_n681), .ZN(new_n965));
  XOR2_X1   g0765(.A(new_n965), .B(new_n674), .Z(new_n966));
  OAI21_X1  g0766(.A(new_n733), .B1(new_n962), .B2(new_n966), .ZN(new_n967));
  XNOR2_X1  g0767(.A(new_n689), .B(KEYINPUT41), .ZN(new_n968));
  AOI21_X1  g0768(.A(new_n739), .B1(new_n967), .B2(new_n968), .ZN(new_n969));
  NAND3_X1  g0769(.A1(new_n682), .A2(new_n630), .A3(new_n709), .ZN(new_n970));
  XOR2_X1   g0770(.A(new_n970), .B(KEYINPUT42), .Z(new_n971));
  AOI21_X1  g0771(.A(new_n341), .B1(new_n627), .B2(new_n622), .ZN(new_n972));
  INV_X1    g0772(.A(new_n632), .ZN(new_n973));
  OAI21_X1  g0773(.A(new_n669), .B1(new_n972), .B2(new_n973), .ZN(new_n974));
  NAND2_X1  g0774(.A1(new_n971), .A2(new_n974), .ZN(new_n975));
  INV_X1    g0775(.A(new_n927), .ZN(new_n976));
  NOR3_X1   g0776(.A1(new_n975), .A2(KEYINPUT43), .A3(new_n976), .ZN(new_n977));
  NOR2_X1   g0777(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n978));
  AND2_X1   g0778(.A1(new_n976), .A2(KEYINPUT43), .ZN(new_n979));
  AOI211_X1 g0779(.A(new_n978), .B(new_n979), .C1(new_n971), .C2(new_n974), .ZN(new_n980));
  NAND2_X1  g0780(.A1(new_n959), .A2(new_n952), .ZN(new_n981));
  OR3_X1    g0781(.A1(new_n977), .A2(new_n980), .A3(new_n981), .ZN(new_n982));
  OAI21_X1  g0782(.A(new_n981), .B1(new_n977), .B2(new_n980), .ZN(new_n983));
  NAND2_X1  g0783(.A1(new_n982), .A2(new_n983), .ZN(new_n984));
  OAI21_X1  g0784(.A(new_n949), .B1(new_n969), .B2(new_n984), .ZN(G387));
  INV_X1    g0785(.A(new_n966), .ZN(new_n986));
  NOR2_X1   g0786(.A1(new_n733), .A2(new_n986), .ZN(new_n987));
  NAND2_X1  g0787(.A1(new_n733), .A2(new_n986), .ZN(new_n988));
  NAND2_X1  g0788(.A1(new_n988), .A2(new_n689), .ZN(new_n989));
  AOI21_X1  g0789(.A(new_n987), .B1(new_n989), .B2(KEYINPUT108), .ZN(new_n990));
  OAI21_X1  g0790(.A(new_n990), .B1(KEYINPUT108), .B2(new_n989), .ZN(new_n991));
  NAND2_X1  g0791(.A1(new_n986), .A2(new_n739), .ZN(new_n992));
  OAI22_X1  g0792(.A1(new_n829), .A2(new_n215), .B1(new_n504), .B2(new_n746), .ZN(new_n993));
  OAI22_X1  g0793(.A1(new_n757), .A2(new_n206), .B1(new_n396), .B2(new_n768), .ZN(new_n994));
  NAND2_X1  g0794(.A1(new_n826), .A2(new_n459), .ZN(new_n995));
  OAI21_X1  g0795(.A(new_n995), .B1(new_n226), .B2(new_n769), .ZN(new_n996));
  NOR4_X1   g0796(.A1(new_n993), .A2(new_n994), .A3(new_n795), .A4(new_n996), .ZN(new_n997));
  OAI221_X1 g0797(.A(new_n997), .B1(new_n386), .B2(new_n750), .C1(new_n393), .C2(new_n763), .ZN(new_n998));
  AOI22_X1  g0798(.A1(G311), .A2(new_n767), .B1(new_n782), .B2(G317), .ZN(new_n999));
  NAND2_X1  g0799(.A1(new_n745), .A2(G322), .ZN(new_n1000));
  OAI211_X1 g0800(.A(new_n999), .B(new_n1000), .C1(new_n832), .C2(new_n769), .ZN(new_n1001));
  XNOR2_X1  g0801(.A(new_n1001), .B(KEYINPUT48), .ZN(new_n1002));
  OAI221_X1 g0802(.A(new_n1002), .B1(new_n834), .B2(new_n748), .C1(new_n771), .C2(new_n829), .ZN(new_n1003));
  XNOR2_X1  g0803(.A(new_n1003), .B(KEYINPUT49), .ZN(new_n1004));
  NAND2_X1  g0804(.A1(new_n939), .A2(G326), .ZN(new_n1005));
  NAND3_X1  g0805(.A1(new_n1004), .A2(new_n795), .A3(new_n1005), .ZN(new_n1006));
  NOR2_X1   g0806(.A1(new_n757), .A2(new_n357), .ZN(new_n1007));
  OAI21_X1  g0807(.A(new_n998), .B1(new_n1006), .B2(new_n1007), .ZN(new_n1008));
  NAND2_X1  g0808(.A1(new_n1008), .A2(new_n791), .ZN(new_n1009));
  OR2_X1    g0809(.A1(new_n237), .A2(new_n564), .ZN(new_n1010));
  AOI22_X1  g0810(.A1(new_n1010), .A2(new_n797), .B1(new_n687), .B2(new_n793), .ZN(new_n1011));
  INV_X1    g0811(.A(new_n396), .ZN(new_n1012));
  NAND2_X1  g0812(.A1(new_n1012), .A2(new_n386), .ZN(new_n1013));
  XNOR2_X1  g0813(.A(new_n1013), .B(KEYINPUT50), .ZN(new_n1014));
  NOR2_X1   g0814(.A1(new_n226), .A2(new_n215), .ZN(new_n1015));
  NOR4_X1   g0815(.A1(new_n1014), .A2(new_n687), .A3(G45), .A4(new_n1015), .ZN(new_n1016));
  OAI22_X1  g0816(.A1(new_n1011), .A2(new_n1016), .B1(G107), .B2(new_n223), .ZN(new_n1017));
  AOI21_X1  g0817(.A(new_n741), .B1(new_n1017), .B2(new_n804), .ZN(new_n1018));
  XOR2_X1   g0818(.A(new_n1018), .B(KEYINPUT107), .Z(new_n1019));
  OAI211_X1 g0819(.A(new_n1009), .B(new_n1019), .C1(new_n678), .C2(new_n807), .ZN(new_n1020));
  NAND3_X1  g0820(.A1(new_n991), .A2(new_n992), .A3(new_n1020), .ZN(G393));
  NAND3_X1  g0821(.A1(new_n960), .A2(new_n739), .A3(new_n961), .ZN(new_n1022));
  INV_X1    g0822(.A(new_n791), .ZN(new_n1023));
  INV_X1    g0823(.A(new_n769), .ZN(new_n1024));
  AOI22_X1  g0824(.A1(new_n767), .A2(G50), .B1(new_n1024), .B2(new_n1012), .ZN(new_n1025));
  AOI22_X1  g0825(.A1(G150), .A2(new_n745), .B1(new_n782), .B2(G159), .ZN(new_n1026));
  OAI221_X1 g0826(.A(new_n1025), .B1(new_n215), .B2(new_n748), .C1(new_n1026), .C2(KEYINPUT51), .ZN(new_n1027));
  OAI21_X1  g0827(.A(new_n796), .B1(new_n829), .B2(new_n226), .ZN(new_n1028));
  AOI211_X1 g0828(.A(new_n1027), .B(new_n1028), .C1(G87), .C2(new_n756), .ZN(new_n1029));
  OAI21_X1  g0829(.A(new_n1029), .B1(new_n929), .B2(new_n763), .ZN(new_n1030));
  AOI21_X1  g0830(.A(new_n1030), .B1(KEYINPUT51), .B2(new_n1026), .ZN(new_n1031));
  XNOR2_X1  g0831(.A(new_n1031), .B(KEYINPUT109), .ZN(new_n1032));
  AOI22_X1  g0832(.A1(G317), .A2(new_n745), .B1(new_n782), .B2(G311), .ZN(new_n1033));
  AOI21_X1  g0833(.A(new_n758), .B1(KEYINPUT52), .B2(new_n1033), .ZN(new_n1034));
  NAND2_X1  g0834(.A1(new_n1034), .A2(new_n346), .ZN(new_n1035));
  AOI22_X1  g0835(.A1(G116), .A2(new_n826), .B1(new_n767), .B2(G303), .ZN(new_n1036));
  XNOR2_X1  g0836(.A(new_n1036), .B(KEYINPUT110), .ZN(new_n1037));
  OAI22_X1  g0837(.A1(new_n829), .A2(new_n834), .B1(new_n1033), .B2(KEYINPUT52), .ZN(new_n1038));
  NOR3_X1   g0838(.A1(new_n1035), .A2(new_n1037), .A3(new_n1038), .ZN(new_n1039));
  NAND2_X1  g0839(.A1(new_n939), .A2(G322), .ZN(new_n1040));
  OAI211_X1 g0840(.A(new_n1039), .B(new_n1040), .C1(new_n771), .C2(new_n769), .ZN(new_n1041));
  AOI21_X1  g0841(.A(new_n1023), .B1(new_n1032), .B2(new_n1041), .ZN(new_n1042));
  OAI21_X1  g0842(.A(new_n804), .B1(new_n206), .B2(new_n223), .ZN(new_n1043));
  AOI21_X1  g0843(.A(new_n1043), .B1(new_n797), .B2(new_n247), .ZN(new_n1044));
  NOR3_X1   g0844(.A1(new_n1042), .A2(new_n741), .A3(new_n1044), .ZN(new_n1045));
  OAI21_X1  g0845(.A(new_n1045), .B1(new_n807), .B2(new_n952), .ZN(new_n1046));
  NAND2_X1  g0846(.A1(new_n988), .A2(new_n962), .ZN(new_n1047));
  NAND2_X1  g0847(.A1(new_n1047), .A2(new_n689), .ZN(new_n1048));
  NOR2_X1   g0848(.A1(new_n988), .A2(new_n962), .ZN(new_n1049));
  OAI211_X1 g0849(.A(new_n1022), .B(new_n1046), .C1(new_n1048), .C2(new_n1049), .ZN(G390));
  INV_X1    g0850(.A(new_n905), .ZN(new_n1051));
  OAI21_X1  g0851(.A(new_n1051), .B1(new_n859), .B2(new_n902), .ZN(new_n1052));
  INV_X1    g0852(.A(new_n897), .ZN(new_n1053));
  INV_X1    g0853(.A(new_n811), .ZN(new_n1054));
  NAND2_X1  g0854(.A1(new_n1054), .A2(new_n545), .ZN(new_n1055));
  OAI211_X1 g0855(.A(new_n669), .B(new_n1055), .C1(new_n707), .C2(new_n712), .ZN(new_n1056));
  AOI21_X1  g0856(.A(new_n1053), .B1(new_n1056), .B2(new_n810), .ZN(new_n1057));
  OAI21_X1  g0857(.A(KEYINPUT111), .B1(new_n1052), .B2(new_n1057), .ZN(new_n1058));
  NAND2_X1  g0858(.A1(new_n1056), .A2(new_n810), .ZN(new_n1059));
  NAND2_X1  g0859(.A1(new_n1059), .A2(new_n897), .ZN(new_n1060));
  INV_X1    g0860(.A(KEYINPUT111), .ZN(new_n1061));
  AOI21_X1  g0861(.A(new_n905), .B1(new_n878), .B2(new_n879), .ZN(new_n1062));
  NAND3_X1  g0862(.A1(new_n1060), .A2(new_n1061), .A3(new_n1062), .ZN(new_n1063));
  NAND2_X1  g0863(.A1(new_n1058), .A2(new_n1063), .ZN(new_n1064));
  AOI21_X1  g0864(.A(new_n1053), .B1(new_n891), .B2(new_n892), .ZN(new_n1065));
  NOR3_X1   g0865(.A1(new_n859), .A2(new_n860), .A3(new_n899), .ZN(new_n1066));
  AOI21_X1  g0866(.A(KEYINPUT39), .B1(new_n878), .B2(new_n879), .ZN(new_n1067));
  OAI22_X1  g0867(.A1(new_n1065), .A2(new_n905), .B1(new_n1066), .B2(new_n1067), .ZN(new_n1068));
  AND4_X1   g0868(.A1(G330), .A2(new_n730), .A3(new_n897), .A4(new_n814), .ZN(new_n1069));
  NAND4_X1  g0869(.A1(new_n862), .A2(G330), .A3(new_n867), .A4(new_n869), .ZN(new_n1070));
  INV_X1    g0870(.A(KEYINPUT112), .ZN(new_n1071));
  OAI21_X1  g0871(.A(new_n1069), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND3_X1  g0872(.A1(new_n1064), .A2(new_n1068), .A3(new_n1072), .ZN(new_n1073));
  NOR3_X1   g0873(.A1(new_n889), .A2(new_n888), .A3(new_n890), .ZN(new_n1074));
  AOI21_X1  g0874(.A(KEYINPUT102), .B1(new_n815), .B2(new_n810), .ZN(new_n1075));
  OAI21_X1  g0875(.A(new_n897), .B1(new_n1074), .B2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g0876(.A1(new_n1076), .A2(new_n1051), .ZN(new_n1077));
  NAND2_X1  g0877(.A1(new_n903), .A2(new_n904), .ZN(new_n1078));
  AOI22_X1  g0878(.A1(new_n1077), .A2(new_n1078), .B1(new_n1058), .B2(new_n1063), .ZN(new_n1079));
  NOR2_X1   g0879(.A1(new_n1070), .A2(KEYINPUT112), .ZN(new_n1080));
  INV_X1    g0880(.A(new_n1080), .ZN(new_n1081));
  OAI211_X1 g0881(.A(new_n1073), .B(new_n739), .C1(new_n1079), .C2(new_n1081), .ZN(new_n1082));
  AOI21_X1  g0882(.A(new_n802), .B1(new_n903), .B2(new_n904), .ZN(new_n1083));
  INV_X1    g0883(.A(KEYINPUT115), .ZN(new_n1084));
  INV_X1    g0884(.A(G128), .ZN(new_n1085));
  NOR2_X1   g0885(.A1(new_n746), .A2(new_n1085), .ZN(new_n1086));
  AOI211_X1 g0886(.A(new_n346), .B(new_n1086), .C1(new_n776), .C2(G125), .ZN(new_n1087));
  INV_X1    g0887(.A(G132), .ZN(new_n1088));
  OAI221_X1 g0888(.A(new_n1087), .B1(new_n386), .B2(new_n757), .C1(new_n1088), .C2(new_n750), .ZN(new_n1089));
  NOR2_X1   g0889(.A1(new_n748), .A2(new_n504), .ZN(new_n1090));
  XOR2_X1   g0890(.A(KEYINPUT114), .B(KEYINPUT53), .Z(new_n1091));
  INV_X1    g0891(.A(new_n1091), .ZN(new_n1092));
  OAI21_X1  g0892(.A(new_n1092), .B1(new_n829), .B2(new_n393), .ZN(new_n1093));
  NAND3_X1  g0893(.A1(new_n759), .A2(G150), .A3(new_n1091), .ZN(new_n1094));
  XOR2_X1   g0894(.A(KEYINPUT54), .B(G143), .Z(new_n1095));
  INV_X1    g0895(.A(new_n1095), .ZN(new_n1096));
  OAI211_X1 g0896(.A(new_n1093), .B(new_n1094), .C1(new_n769), .C2(new_n1096), .ZN(new_n1097));
  NOR2_X1   g0897(.A1(new_n768), .A2(new_n822), .ZN(new_n1098));
  NOR4_X1   g0898(.A1(new_n1089), .A2(new_n1090), .A3(new_n1097), .A4(new_n1098), .ZN(new_n1099));
  OAI22_X1  g0899(.A1(new_n226), .A2(new_n757), .B1(new_n829), .B2(new_n204), .ZN(new_n1100));
  AOI21_X1  g0900(.A(new_n401), .B1(new_n776), .B2(G294), .ZN(new_n1101));
  AOI22_X1  g0901(.A1(new_n826), .A2(G77), .B1(new_n782), .B2(G116), .ZN(new_n1102));
  OAI211_X1 g0902(.A(new_n1101), .B(new_n1102), .C1(new_n210), .C2(new_n768), .ZN(new_n1103));
  NOR2_X1   g0903(.A1(new_n769), .A2(new_n206), .ZN(new_n1104));
  NOR2_X1   g0904(.A1(new_n746), .A2(new_n834), .ZN(new_n1105));
  NOR4_X1   g0905(.A1(new_n1100), .A2(new_n1103), .A3(new_n1104), .A4(new_n1105), .ZN(new_n1106));
  OAI21_X1  g0906(.A(new_n791), .B1(new_n1099), .B2(new_n1106), .ZN(new_n1107));
  OAI211_X1 g0907(.A(new_n1107), .B(new_n740), .C1(new_n1012), .C2(new_n842), .ZN(new_n1108));
  OR3_X1    g0908(.A1(new_n1083), .A2(new_n1084), .A3(new_n1108), .ZN(new_n1109));
  OAI21_X1  g0909(.A(new_n1084), .B1(new_n1083), .B2(new_n1108), .ZN(new_n1110));
  NAND2_X1  g0910(.A1(new_n1109), .A2(new_n1110), .ZN(new_n1111));
  NAND2_X1  g0911(.A1(new_n1082), .A2(new_n1111), .ZN(new_n1112));
  NAND2_X1  g0912(.A1(new_n1112), .A2(KEYINPUT116), .ZN(new_n1113));
  AND3_X1   g0913(.A1(new_n1064), .A2(new_n1072), .A3(new_n1068), .ZN(new_n1114));
  AOI21_X1  g0914(.A(new_n1081), .B1(new_n1064), .B2(new_n1068), .ZN(new_n1115));
  NAND4_X1  g0915(.A1(new_n862), .A2(G330), .A3(new_n814), .A4(new_n869), .ZN(new_n1116));
  AOI211_X1 g0916(.A(new_n1059), .B(new_n1069), .C1(new_n1053), .C2(new_n1116), .ZN(new_n1117));
  NAND3_X1  g0917(.A1(new_n730), .A2(G330), .A3(new_n814), .ZN(new_n1118));
  NAND2_X1  g0918(.A1(new_n1118), .A2(new_n1053), .ZN(new_n1119));
  NAND2_X1  g0919(.A1(new_n1070), .A2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g0920(.A1(new_n1120), .A2(new_n893), .ZN(new_n1121));
  INV_X1    g0921(.A(KEYINPUT113), .ZN(new_n1122));
  NAND2_X1  g0922(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g0923(.A1(new_n1120), .A2(KEYINPUT113), .A3(new_n893), .ZN(new_n1124));
  AOI21_X1  g0924(.A(new_n1117), .B1(new_n1123), .B2(new_n1124), .ZN(new_n1125));
  NAND3_X1  g0925(.A1(new_n909), .A2(new_n658), .A3(new_n884), .ZN(new_n1126));
  OAI22_X1  g0926(.A1(new_n1114), .A2(new_n1115), .B1(new_n1125), .B2(new_n1126), .ZN(new_n1127));
  NOR3_X1   g0927(.A1(new_n1052), .A2(KEYINPUT111), .A3(new_n1057), .ZN(new_n1128));
  AOI21_X1  g0928(.A(new_n1061), .B1(new_n1060), .B2(new_n1062), .ZN(new_n1129));
  NOR2_X1   g0929(.A1(new_n1128), .A2(new_n1129), .ZN(new_n1130));
  AOI22_X1  g0930(.A1(new_n1076), .A2(new_n1051), .B1(new_n903), .B2(new_n904), .ZN(new_n1131));
  OAI21_X1  g0931(.A(new_n1080), .B1(new_n1130), .B2(new_n1131), .ZN(new_n1132));
  INV_X1    g0932(.A(new_n1126), .ZN(new_n1133));
  AOI21_X1  g0933(.A(new_n1069), .B1(new_n1116), .B2(new_n1053), .ZN(new_n1134));
  NAND3_X1  g0934(.A1(new_n1134), .A2(new_n810), .A3(new_n1056), .ZN(new_n1135));
  INV_X1    g0935(.A(new_n1124), .ZN(new_n1136));
  AOI21_X1  g0936(.A(KEYINPUT113), .B1(new_n1120), .B2(new_n893), .ZN(new_n1137));
  OAI21_X1  g0937(.A(new_n1135), .B1(new_n1136), .B2(new_n1137), .ZN(new_n1138));
  NAND4_X1  g0938(.A1(new_n1132), .A2(new_n1073), .A3(new_n1133), .A4(new_n1138), .ZN(new_n1139));
  NAND3_X1  g0939(.A1(new_n1127), .A2(new_n1139), .A3(new_n689), .ZN(new_n1140));
  INV_X1    g0940(.A(KEYINPUT116), .ZN(new_n1141));
  NAND3_X1  g0941(.A1(new_n1082), .A2(new_n1141), .A3(new_n1111), .ZN(new_n1142));
  NAND3_X1  g0942(.A1(new_n1113), .A2(new_n1140), .A3(new_n1142), .ZN(new_n1143));
  NAND2_X1  g0943(.A1(new_n1143), .A2(KEYINPUT117), .ZN(new_n1144));
  INV_X1    g0944(.A(KEYINPUT117), .ZN(new_n1145));
  NAND4_X1  g0945(.A1(new_n1113), .A2(new_n1140), .A3(new_n1145), .A4(new_n1142), .ZN(new_n1146));
  NAND2_X1  g0946(.A1(new_n1144), .A2(new_n1146), .ZN(G378));
  NAND2_X1  g0947(.A1(new_n427), .A2(KEYINPUT55), .ZN(new_n1148));
  INV_X1    g0948(.A(KEYINPUT55), .ZN(new_n1149));
  NAND3_X1  g0949(.A1(new_n422), .A2(new_n1149), .A3(new_n426), .ZN(new_n1150));
  NOR2_X1   g0950(.A1(new_n398), .A2(new_n666), .ZN(new_n1151));
  INV_X1    g0951(.A(new_n1151), .ZN(new_n1152));
  NAND3_X1  g0952(.A1(new_n1148), .A2(new_n1150), .A3(new_n1152), .ZN(new_n1153));
  AOI21_X1  g0953(.A(new_n1149), .B1(new_n422), .B2(new_n426), .ZN(new_n1154));
  AOI211_X1 g0954(.A(KEYINPUT55), .B(new_n654), .C1(new_n419), .C2(new_n421), .ZN(new_n1155));
  OAI21_X1  g0955(.A(new_n1151), .B1(new_n1154), .B2(new_n1155), .ZN(new_n1156));
  NAND2_X1  g0956(.A1(new_n1153), .A2(new_n1156), .ZN(new_n1157));
  XNOR2_X1  g0957(.A(KEYINPUT120), .B(KEYINPUT56), .ZN(new_n1158));
  INV_X1    g0958(.A(new_n1158), .ZN(new_n1159));
  NAND2_X1  g0959(.A1(new_n1157), .A2(new_n1159), .ZN(new_n1160));
  NAND3_X1  g0960(.A1(new_n1153), .A2(new_n1156), .A3(new_n1158), .ZN(new_n1161));
  AND2_X1   g0961(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1162));
  NAND2_X1  g0962(.A1(new_n882), .A2(new_n1162), .ZN(new_n1163));
  NAND2_X1  g0963(.A1(new_n1160), .A2(new_n1161), .ZN(new_n1164));
  NAND4_X1  g0964(.A1(new_n1164), .A2(new_n871), .A3(new_n881), .A4(G330), .ZN(new_n1165));
  NAND2_X1  g0965(.A1(new_n1163), .A2(new_n1165), .ZN(new_n1166));
  INV_X1    g0966(.A(new_n908), .ZN(new_n1167));
  NAND2_X1  g0967(.A1(new_n1166), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g0968(.A1(new_n1168), .A2(KEYINPUT121), .ZN(new_n1169));
  NAND3_X1  g0969(.A1(new_n1163), .A2(new_n908), .A3(new_n1165), .ZN(new_n1170));
  NAND2_X1  g0970(.A1(new_n1170), .A2(KEYINPUT122), .ZN(new_n1171));
  INV_X1    g0971(.A(KEYINPUT122), .ZN(new_n1172));
  NAND4_X1  g0972(.A1(new_n1163), .A2(new_n908), .A3(new_n1165), .A4(new_n1172), .ZN(new_n1173));
  AOI21_X1  g0973(.A(new_n908), .B1(new_n1163), .B2(new_n1165), .ZN(new_n1174));
  INV_X1    g0974(.A(KEYINPUT121), .ZN(new_n1175));
  NAND2_X1  g0975(.A1(new_n1174), .A2(new_n1175), .ZN(new_n1176));
  NAND4_X1  g0976(.A1(new_n1169), .A2(new_n1171), .A3(new_n1173), .A4(new_n1176), .ZN(new_n1177));
  NAND2_X1  g0977(.A1(new_n1177), .A2(new_n739), .ZN(new_n1178));
  NOR2_X1   g0978(.A1(new_n750), .A2(new_n1085), .ZN(new_n1179));
  OAI22_X1  g0979(.A1(new_n829), .A2(new_n1096), .B1(new_n822), .B2(new_n769), .ZN(new_n1180));
  AOI211_X1 g0980(.A(new_n1179), .B(new_n1180), .C1(G125), .C2(new_n745), .ZN(new_n1181));
  OAI221_X1 g0981(.A(new_n1181), .B1(new_n1088), .B2(new_n768), .C1(new_n393), .C2(new_n748), .ZN(new_n1182));
  XOR2_X1   g0982(.A(KEYINPUT119), .B(KEYINPUT59), .Z(new_n1183));
  XNOR2_X1  g0983(.A(new_n1182), .B(new_n1183), .ZN(new_n1184));
  OAI211_X1 g0984(.A(new_n251), .B(new_n294), .C1(new_n757), .C2(new_n504), .ZN(new_n1185));
  AOI21_X1  g0985(.A(new_n1185), .B1(G124), .B2(new_n939), .ZN(new_n1186));
  NAND2_X1  g0986(.A1(new_n1184), .A2(new_n1186), .ZN(new_n1187));
  OAI221_X1 g0987(.A(new_n294), .B1(new_n210), .B2(new_n750), .C1(new_n829), .C2(new_n215), .ZN(new_n1188));
  AOI22_X1  g0988(.A1(new_n776), .A2(G283), .B1(G68), .B2(new_n826), .ZN(new_n1189));
  NAND2_X1  g0989(.A1(new_n756), .A2(G58), .ZN(new_n1190));
  NAND2_X1  g0990(.A1(new_n745), .A2(G116), .ZN(new_n1191));
  NAND4_X1  g0991(.A1(new_n1189), .A2(new_n1190), .A3(new_n795), .A4(new_n1191), .ZN(new_n1192));
  AOI22_X1  g0992(.A1(new_n767), .A2(G97), .B1(new_n1024), .B2(new_n459), .ZN(new_n1193));
  XOR2_X1   g0993(.A(new_n1193), .B(KEYINPUT118), .Z(new_n1194));
  NOR3_X1   g0994(.A1(new_n1188), .A2(new_n1192), .A3(new_n1194), .ZN(new_n1195));
  XOR2_X1   g0995(.A(new_n1195), .B(KEYINPUT58), .Z(new_n1196));
  AOI21_X1  g0996(.A(G41), .B1(new_n796), .B2(G33), .ZN(new_n1197));
  OAI211_X1 g0997(.A(new_n1187), .B(new_n1196), .C1(G50), .C2(new_n1197), .ZN(new_n1198));
  AOI21_X1  g0998(.A(new_n741), .B1(new_n1198), .B2(new_n791), .ZN(new_n1199));
  OAI221_X1 g0999(.A(new_n1199), .B1(G50), .B2(new_n842), .C1(new_n1164), .C2(new_n802), .ZN(new_n1200));
  NAND2_X1  g1000(.A1(new_n1178), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g1001(.A1(new_n1139), .A2(new_n1133), .ZN(new_n1202));
  NAND2_X1  g1002(.A1(new_n1177), .A2(new_n1202), .ZN(new_n1203));
  INV_X1    g1003(.A(KEYINPUT57), .ZN(new_n1204));
  AOI21_X1  g1004(.A(new_n691), .B1(new_n1203), .B2(new_n1204), .ZN(new_n1205));
  AOI21_X1  g1005(.A(new_n1204), .B1(new_n1168), .B2(new_n1170), .ZN(new_n1206));
  AND3_X1   g1006(.A1(new_n1206), .A2(new_n1202), .A3(KEYINPUT123), .ZN(new_n1207));
  AOI21_X1  g1007(.A(KEYINPUT123), .B1(new_n1206), .B2(new_n1202), .ZN(new_n1208));
  NOR2_X1   g1008(.A1(new_n1207), .A2(new_n1208), .ZN(new_n1209));
  AOI211_X1 g1009(.A(KEYINPUT124), .B(new_n1201), .C1(new_n1205), .C2(new_n1209), .ZN(new_n1210));
  INV_X1    g1010(.A(KEYINPUT124), .ZN(new_n1211));
  NAND2_X1  g1011(.A1(new_n1203), .A2(new_n1204), .ZN(new_n1212));
  NAND3_X1  g1012(.A1(new_n1209), .A2(new_n1212), .A3(new_n689), .ZN(new_n1213));
  AND2_X1   g1013(.A1(new_n1178), .A2(new_n1200), .ZN(new_n1214));
  AOI21_X1  g1014(.A(new_n1211), .B1(new_n1213), .B2(new_n1214), .ZN(new_n1215));
  NOR2_X1   g1015(.A1(new_n1210), .A2(new_n1215), .ZN(new_n1216));
  INV_X1    g1016(.A(new_n1216), .ZN(G375));
  NOR2_X1   g1017(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1218));
  INV_X1    g1018(.A(new_n1218), .ZN(new_n1219));
  NAND2_X1  g1019(.A1(new_n1125), .A2(new_n1126), .ZN(new_n1220));
  NAND3_X1  g1020(.A1(new_n1219), .A2(new_n968), .A3(new_n1220), .ZN(new_n1221));
  NAND2_X1  g1021(.A1(new_n1053), .A2(new_n801), .ZN(new_n1222));
  OAI21_X1  g1022(.A(new_n1190), .B1(new_n1085), .B2(new_n775), .ZN(new_n1223));
  AOI211_X1 g1023(.A(new_n795), .B(new_n1223), .C1(G159), .C2(new_n759), .ZN(new_n1224));
  OAI221_X1 g1024(.A(new_n1224), .B1(new_n386), .B2(new_n748), .C1(new_n393), .C2(new_n769), .ZN(new_n1225));
  XOR2_X1   g1025(.A(new_n1225), .B(KEYINPUT127), .Z(new_n1226));
  AOI22_X1  g1026(.A1(new_n767), .A2(new_n1095), .B1(new_n782), .B2(G137), .ZN(new_n1227));
  OAI21_X1  g1027(.A(new_n1227), .B1(new_n1088), .B2(new_n746), .ZN(new_n1228));
  XNOR2_X1  g1028(.A(new_n1228), .B(KEYINPUT126), .ZN(new_n1229));
  NAND2_X1  g1029(.A1(new_n1226), .A2(new_n1229), .ZN(new_n1230));
  OAI221_X1 g1030(.A(new_n995), .B1(new_n746), .B2(new_n771), .C1(new_n357), .C2(new_n768), .ZN(new_n1231));
  AOI22_X1  g1031(.A1(new_n759), .A2(G97), .B1(new_n776), .B2(G303), .ZN(new_n1232));
  XNOR2_X1  g1032(.A(new_n1232), .B(KEYINPUT125), .ZN(new_n1233));
  AOI211_X1 g1033(.A(new_n1231), .B(new_n1233), .C1(G107), .C2(new_n1024), .ZN(new_n1234));
  INV_X1    g1034(.A(new_n931), .ZN(new_n1235));
  NAND2_X1  g1035(.A1(new_n782), .A2(G283), .ZN(new_n1236));
  NAND4_X1  g1036(.A1(new_n1234), .A2(new_n346), .A3(new_n1235), .A4(new_n1236), .ZN(new_n1237));
  AOI21_X1  g1037(.A(new_n1023), .B1(new_n1230), .B2(new_n1237), .ZN(new_n1238));
  AOI211_X1 g1038(.A(new_n741), .B(new_n1238), .C1(new_n226), .C2(new_n841), .ZN(new_n1239));
  AOI22_X1  g1039(.A1(new_n1138), .A2(new_n739), .B1(new_n1222), .B2(new_n1239), .ZN(new_n1240));
  NAND2_X1  g1040(.A1(new_n1221), .A2(new_n1240), .ZN(G381));
  NOR2_X1   g1041(.A1(G375), .A2(new_n1143), .ZN(new_n1242));
  INV_X1    g1042(.A(G384), .ZN(new_n1243));
  INV_X1    g1043(.A(G381), .ZN(new_n1244));
  INV_X1    g1044(.A(G396), .ZN(new_n1245));
  NAND4_X1  g1045(.A1(new_n991), .A2(new_n1245), .A3(new_n992), .A4(new_n1020), .ZN(new_n1246));
  NOR3_X1   g1046(.A1(new_n1246), .A2(G387), .A3(G390), .ZN(new_n1247));
  NAND4_X1  g1047(.A1(new_n1242), .A2(new_n1243), .A3(new_n1244), .A4(new_n1247), .ZN(G407));
  INV_X1    g1048(.A(new_n1143), .ZN(new_n1249));
  NAND3_X1  g1049(.A1(new_n1216), .A2(new_n667), .A3(new_n1249), .ZN(new_n1250));
  AND2_X1   g1050(.A1(new_n1250), .A2(G213), .ZN(new_n1251));
  NAND2_X1  g1051(.A1(G407), .A2(new_n1251), .ZN(G409));
  XNOR2_X1  g1052(.A(G387), .B(G390), .ZN(new_n1253));
  INV_X1    g1053(.A(new_n1253), .ZN(new_n1254));
  NAND2_X1  g1054(.A1(G393), .A2(G396), .ZN(new_n1255));
  NAND2_X1  g1055(.A1(new_n1255), .A2(new_n1246), .ZN(new_n1256));
  XNOR2_X1  g1056(.A(new_n1254), .B(new_n1256), .ZN(new_n1257));
  INV_X1    g1057(.A(G213), .ZN(new_n1258));
  NOR2_X1   g1058(.A1(new_n1258), .A2(G343), .ZN(new_n1259));
  INV_X1    g1059(.A(KEYINPUT60), .ZN(new_n1260));
  AOI21_X1  g1060(.A(new_n691), .B1(new_n1220), .B2(new_n1260), .ZN(new_n1261));
  OAI211_X1 g1061(.A(new_n1261), .B(new_n1219), .C1(new_n1260), .C2(new_n1220), .ZN(new_n1262));
  AOI21_X1  g1062(.A(G384), .B1(new_n1262), .B2(new_n1240), .ZN(new_n1263));
  INV_X1    g1063(.A(new_n1263), .ZN(new_n1264));
  NAND3_X1  g1064(.A1(new_n1262), .A2(G384), .A3(new_n1240), .ZN(new_n1265));
  NAND2_X1  g1065(.A1(new_n1264), .A2(new_n1265), .ZN(new_n1266));
  NOR2_X1   g1066(.A1(new_n1114), .A2(new_n1115), .ZN(new_n1267));
  AOI21_X1  g1067(.A(new_n1126), .B1(new_n1267), .B2(new_n1218), .ZN(new_n1268));
  XNOR2_X1  g1068(.A(new_n1174), .B(KEYINPUT121), .ZN(new_n1269));
  AND2_X1   g1069(.A1(new_n1171), .A2(new_n1173), .ZN(new_n1270));
  AOI21_X1  g1070(.A(new_n1268), .B1(new_n1269), .B2(new_n1270), .ZN(new_n1271));
  OAI21_X1  g1071(.A(new_n689), .B1(new_n1271), .B2(KEYINPUT57), .ZN(new_n1272));
  INV_X1    g1072(.A(new_n1208), .ZN(new_n1273));
  NAND3_X1  g1073(.A1(new_n1206), .A2(new_n1202), .A3(KEYINPUT123), .ZN(new_n1274));
  NAND2_X1  g1074(.A1(new_n1273), .A2(new_n1274), .ZN(new_n1275));
  OAI211_X1 g1075(.A(G378), .B(new_n1214), .C1(new_n1272), .C2(new_n1275), .ZN(new_n1276));
  NAND2_X1  g1076(.A1(new_n1168), .A2(new_n1170), .ZN(new_n1277));
  NAND2_X1  g1077(.A1(new_n1277), .A2(new_n739), .ZN(new_n1278));
  INV_X1    g1078(.A(new_n968), .ZN(new_n1279));
  OAI211_X1 g1079(.A(new_n1200), .B(new_n1278), .C1(new_n1203), .C2(new_n1279), .ZN(new_n1280));
  NAND2_X1  g1080(.A1(new_n1280), .A2(new_n1249), .ZN(new_n1281));
  AOI211_X1 g1081(.A(new_n1259), .B(new_n1266), .C1(new_n1276), .C2(new_n1281), .ZN(new_n1282));
  INV_X1    g1082(.A(KEYINPUT62), .ZN(new_n1283));
  AOI21_X1  g1083(.A(new_n1259), .B1(new_n1276), .B2(new_n1281), .ZN(new_n1284));
  NAND3_X1  g1084(.A1(new_n1266), .A2(G2897), .A3(new_n1259), .ZN(new_n1285));
  NAND2_X1  g1085(.A1(new_n1259), .A2(G2897), .ZN(new_n1286));
  NAND3_X1  g1086(.A1(new_n1264), .A2(new_n1265), .A3(new_n1286), .ZN(new_n1287));
  NAND2_X1  g1087(.A1(new_n1285), .A2(new_n1287), .ZN(new_n1288));
  OAI22_X1  g1088(.A1(new_n1282), .A2(new_n1283), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1289));
  NAND2_X1  g1089(.A1(new_n1276), .A2(new_n1281), .ZN(new_n1290));
  INV_X1    g1090(.A(new_n1259), .ZN(new_n1291));
  INV_X1    g1091(.A(new_n1266), .ZN(new_n1292));
  NAND4_X1  g1092(.A1(new_n1290), .A2(new_n1283), .A3(new_n1291), .A4(new_n1292), .ZN(new_n1293));
  INV_X1    g1093(.A(KEYINPUT61), .ZN(new_n1294));
  NAND2_X1  g1094(.A1(new_n1293), .A2(new_n1294), .ZN(new_n1295));
  OAI21_X1  g1095(.A(new_n1257), .B1(new_n1289), .B2(new_n1295), .ZN(new_n1296));
  OAI21_X1  g1096(.A(KEYINPUT63), .B1(new_n1284), .B2(new_n1288), .ZN(new_n1297));
  NAND2_X1  g1097(.A1(new_n1284), .A2(new_n1292), .ZN(new_n1298));
  NAND2_X1  g1098(.A1(new_n1297), .A2(new_n1298), .ZN(new_n1299));
  AOI21_X1  g1099(.A(new_n1257), .B1(new_n1282), .B2(KEYINPUT63), .ZN(new_n1300));
  NAND3_X1  g1100(.A1(new_n1299), .A2(new_n1300), .A3(new_n1294), .ZN(new_n1301));
  NAND2_X1  g1101(.A1(new_n1296), .A2(new_n1301), .ZN(G405));
  OAI21_X1  g1102(.A(new_n1214), .B1(new_n1272), .B2(new_n1275), .ZN(new_n1303));
  NAND2_X1  g1103(.A1(new_n1303), .A2(KEYINPUT124), .ZN(new_n1304));
  NAND3_X1  g1104(.A1(new_n1213), .A2(new_n1211), .A3(new_n1214), .ZN(new_n1305));
  AOI21_X1  g1105(.A(new_n1143), .B1(new_n1304), .B2(new_n1305), .ZN(new_n1306));
  XNOR2_X1  g1106(.A(new_n1256), .B(new_n1253), .ZN(new_n1307));
  INV_X1    g1107(.A(new_n1276), .ZN(new_n1308));
  NOR3_X1   g1108(.A1(new_n1306), .A2(new_n1307), .A3(new_n1308), .ZN(new_n1309));
  OAI21_X1  g1109(.A(new_n1249), .B1(new_n1210), .B2(new_n1215), .ZN(new_n1310));
  AOI21_X1  g1110(.A(new_n1257), .B1(new_n1310), .B2(new_n1276), .ZN(new_n1311));
  OAI21_X1  g1111(.A(new_n1266), .B1(new_n1309), .B2(new_n1311), .ZN(new_n1312));
  OAI21_X1  g1112(.A(new_n1307), .B1(new_n1306), .B2(new_n1308), .ZN(new_n1313));
  NAND3_X1  g1113(.A1(new_n1310), .A2(new_n1257), .A3(new_n1276), .ZN(new_n1314));
  NAND3_X1  g1114(.A1(new_n1313), .A2(new_n1292), .A3(new_n1314), .ZN(new_n1315));
  NAND2_X1  g1115(.A1(new_n1312), .A2(new_n1315), .ZN(G402));
endmodule


