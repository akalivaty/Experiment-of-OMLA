//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 1 0 1 1 0 0 1 1 1 1 1 0 1 1 0 0 1 0 1 0 1 0 0 1 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 1 1 0 1 0 1 0 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:26 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n664,
    new_n665, new_n666, new_n667, new_n669, new_n670, new_n671, new_n672,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n729, new_n730, new_n731, new_n732, new_n734, new_n735,
    new_n736, new_n737, new_n739, new_n740, new_n741, new_n742, new_n743,
    new_n745, new_n747, new_n748, new_n749, new_n750, new_n751, new_n752,
    new_n753, new_n754, new_n755, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n828, new_n829, new_n831, new_n832, new_n833, new_n835, new_n836,
    new_n837, new_n838, new_n839, new_n840, new_n841, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n897, new_n898, new_n900, new_n901, new_n903, new_n904,
    new_n905, new_n906, new_n907, new_n908, new_n909, new_n910, new_n912,
    new_n913, new_n914, new_n916, new_n917, new_n918, new_n919, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n934, new_n935, new_n936, new_n938,
    new_n939, new_n940, new_n941, new_n942, new_n944, new_n945, new_n946,
    new_n947;
  XNOR2_X1  g000(.A(G57gat), .B(G64gat), .ZN(new_n202));
  AOI21_X1  g001(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n203));
  NOR2_X1   g002(.A1(new_n202), .A2(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(G71gat), .ZN(new_n205));
  INV_X1    g004(.A(G78gat), .ZN(new_n206));
  NAND3_X1  g005(.A1(new_n205), .A2(new_n206), .A3(KEYINPUT91), .ZN(new_n207));
  NAND2_X1  g006(.A1(G71gat), .A2(G78gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n208), .A2(KEYINPUT90), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT91), .ZN(new_n210));
  OAI21_X1  g009(.A(new_n210), .B1(G71gat), .B2(G78gat), .ZN(new_n211));
  INV_X1    g010(.A(KEYINPUT90), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n212), .A2(G71gat), .A3(G78gat), .ZN(new_n213));
  NAND4_X1  g012(.A1(new_n207), .A2(new_n209), .A3(new_n211), .A4(new_n213), .ZN(new_n214));
  NOR2_X1   g013(.A1(new_n204), .A2(new_n214), .ZN(new_n215));
  INV_X1    g014(.A(KEYINPUT92), .ZN(new_n216));
  OAI211_X1 g015(.A(new_n205), .B(new_n206), .C1(new_n216), .C2(KEYINPUT9), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n217), .A2(new_n208), .ZN(new_n218));
  XOR2_X1   g017(.A(G57gat), .B(G64gat), .Z(new_n219));
  INV_X1    g018(.A(KEYINPUT9), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n208), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(new_n216), .ZN(new_n222));
  NAND3_X1  g021(.A1(new_n218), .A2(new_n219), .A3(new_n222), .ZN(new_n223));
  INV_X1    g022(.A(KEYINPUT93), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n223), .A2(new_n224), .ZN(new_n225));
  NAND4_X1  g024(.A1(new_n218), .A2(new_n219), .A3(KEYINPUT93), .A4(new_n222), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n215), .B1(new_n225), .B2(new_n226), .ZN(new_n227));
  XOR2_X1   g026(.A(KEYINPUT94), .B(KEYINPUT21), .Z(new_n228));
  NOR2_X1   g027(.A1(new_n227), .A2(new_n228), .ZN(new_n229));
  NAND2_X1  g028(.A1(G231gat), .A2(G233gat), .ZN(new_n230));
  XOR2_X1   g029(.A(new_n229), .B(new_n230), .Z(new_n231));
  INV_X1    g030(.A(G127gat), .ZN(new_n232));
  XNOR2_X1  g031(.A(new_n231), .B(new_n232), .ZN(new_n233));
  OR2_X1    g032(.A1(new_n227), .A2(KEYINPUT96), .ZN(new_n234));
  NAND2_X1  g033(.A1(new_n227), .A2(KEYINPUT96), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n234), .A2(KEYINPUT21), .A3(new_n235), .ZN(new_n236));
  XNOR2_X1  g035(.A(G15gat), .B(G22gat), .ZN(new_n237));
  NAND2_X1  g036(.A1(new_n237), .A2(KEYINPUT87), .ZN(new_n238));
  INV_X1    g037(.A(G1gat), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n238), .A2(new_n239), .ZN(new_n240));
  NAND3_X1  g039(.A1(new_n237), .A2(KEYINPUT87), .A3(G1gat), .ZN(new_n241));
  INV_X1    g040(.A(KEYINPUT16), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n237), .A2(new_n242), .ZN(new_n243));
  NAND3_X1  g042(.A1(new_n240), .A2(new_n241), .A3(new_n243), .ZN(new_n244));
  INV_X1    g043(.A(G8gat), .ZN(new_n245));
  XNOR2_X1  g044(.A(new_n244), .B(new_n245), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n236), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(new_n233), .B(new_n247), .ZN(new_n248));
  XNOR2_X1  g047(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(KEYINPUT95), .ZN(new_n250));
  XNOR2_X1  g049(.A(new_n250), .B(G155gat), .ZN(new_n251));
  XOR2_X1   g050(.A(G183gat), .B(G211gat), .Z(new_n252));
  XNOR2_X1  g051(.A(new_n251), .B(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(new_n248), .B(new_n253), .ZN(new_n254));
  AND2_X1   g053(.A1(G232gat), .A2(G233gat), .ZN(new_n255));
  NOR2_X1   g054(.A1(new_n255), .A2(KEYINPUT41), .ZN(new_n256));
  XNOR2_X1  g055(.A(new_n256), .B(G134gat), .ZN(new_n257));
  INV_X1    g056(.A(G162gat), .ZN(new_n258));
  XNOR2_X1  g057(.A(new_n257), .B(new_n258), .ZN(new_n259));
  AND2_X1   g058(.A1(G99gat), .A2(G106gat), .ZN(new_n260));
  NOR2_X1   g059(.A1(G99gat), .A2(G106gat), .ZN(new_n261));
  OAI21_X1  g060(.A(KEYINPUT97), .B1(new_n260), .B2(new_n261), .ZN(new_n262));
  INV_X1    g061(.A(G99gat), .ZN(new_n263));
  INV_X1    g062(.A(G106gat), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n263), .A2(new_n264), .ZN(new_n265));
  INV_X1    g064(.A(KEYINPUT97), .ZN(new_n266));
  NAND2_X1  g065(.A1(G99gat), .A2(G106gat), .ZN(new_n267));
  NAND3_X1  g066(.A1(new_n265), .A2(new_n266), .A3(new_n267), .ZN(new_n268));
  AND2_X1   g067(.A1(new_n262), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n267), .A2(KEYINPUT8), .ZN(new_n270));
  NAND2_X1  g069(.A1(G85gat), .A2(G92gat), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT7), .ZN(new_n272));
  NAND2_X1  g071(.A1(new_n271), .A2(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(G85gat), .ZN(new_n274));
  INV_X1    g073(.A(G92gat), .ZN(new_n275));
  NAND2_X1  g074(.A1(new_n274), .A2(new_n275), .ZN(new_n276));
  NAND3_X1  g075(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n277));
  NAND4_X1  g076(.A1(new_n270), .A2(new_n273), .A3(new_n276), .A4(new_n277), .ZN(new_n278));
  NAND2_X1  g077(.A1(new_n269), .A2(new_n278), .ZN(new_n279));
  AND4_X1   g078(.A1(new_n270), .A2(new_n273), .A3(new_n276), .A4(new_n277), .ZN(new_n280));
  NAND2_X1  g079(.A1(new_n262), .A2(new_n268), .ZN(new_n281));
  AND3_X1   g080(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT98), .ZN(new_n282));
  AOI21_X1  g081(.A(KEYINPUT98), .B1(new_n280), .B2(new_n281), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n279), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  INV_X1    g083(.A(G50gat), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(G43gat), .ZN(new_n286));
  INV_X1    g085(.A(G43gat), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n287), .A2(G50gat), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n286), .A2(new_n288), .A3(KEYINPUT15), .ZN(new_n289));
  INV_X1    g088(.A(G29gat), .ZN(new_n290));
  INV_X1    g089(.A(G36gat), .ZN(new_n291));
  NAND3_X1  g090(.A1(new_n290), .A2(new_n291), .A3(KEYINPUT14), .ZN(new_n292));
  INV_X1    g091(.A(KEYINPUT14), .ZN(new_n293));
  OAI21_X1  g092(.A(new_n293), .B1(G29gat), .B2(G36gat), .ZN(new_n294));
  AND2_X1   g093(.A1(new_n292), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G29gat), .A2(G36gat), .ZN(new_n296));
  AOI21_X1  g095(.A(new_n289), .B1(new_n295), .B2(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(KEYINPUT85), .ZN(new_n299));
  INV_X1    g098(.A(new_n289), .ZN(new_n300));
  AOI21_X1  g099(.A(KEYINPUT15), .B1(new_n286), .B2(new_n288), .ZN(new_n301));
  NOR2_X1   g100(.A1(new_n300), .A2(new_n301), .ZN(new_n302));
  NAND2_X1  g101(.A1(new_n296), .A2(KEYINPUT84), .ZN(new_n303));
  INV_X1    g102(.A(KEYINPUT84), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n304), .A2(G29gat), .A3(G36gat), .ZN(new_n305));
  NAND4_X1  g104(.A1(new_n292), .A2(new_n303), .A3(new_n294), .A4(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(new_n306), .ZN(new_n307));
  AOI21_X1  g106(.A(new_n299), .B1(new_n302), .B2(new_n307), .ZN(new_n308));
  INV_X1    g107(.A(KEYINPUT15), .ZN(new_n309));
  NOR2_X1   g108(.A1(new_n287), .A2(G50gat), .ZN(new_n310));
  NOR2_X1   g109(.A1(new_n285), .A2(G43gat), .ZN(new_n311));
  OAI21_X1  g110(.A(new_n309), .B1(new_n310), .B2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n312), .A2(new_n289), .ZN(new_n313));
  NOR3_X1   g112(.A1(new_n313), .A2(KEYINPUT85), .A3(new_n306), .ZN(new_n314));
  OAI21_X1  g113(.A(new_n298), .B1(new_n308), .B2(new_n314), .ZN(new_n315));
  AOI21_X1  g114(.A(KEYINPUT17), .B1(new_n315), .B2(KEYINPUT86), .ZN(new_n316));
  OAI21_X1  g115(.A(KEYINPUT85), .B1(new_n313), .B2(new_n306), .ZN(new_n317));
  NAND4_X1  g116(.A1(new_n307), .A2(new_n299), .A3(new_n289), .A4(new_n312), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n297), .B1(new_n317), .B2(new_n318), .ZN(new_n319));
  INV_X1    g118(.A(KEYINPUT86), .ZN(new_n320));
  INV_X1    g119(.A(KEYINPUT17), .ZN(new_n321));
  NOR3_X1   g120(.A1(new_n319), .A2(new_n320), .A3(new_n321), .ZN(new_n322));
  OAI21_X1  g121(.A(new_n284), .B1(new_n316), .B2(new_n322), .ZN(new_n323));
  NOR2_X1   g122(.A1(new_n280), .A2(new_n281), .ZN(new_n324));
  INV_X1    g123(.A(KEYINPUT98), .ZN(new_n325));
  OAI21_X1  g124(.A(new_n325), .B1(new_n269), .B2(new_n278), .ZN(new_n326));
  NAND3_X1  g125(.A1(new_n280), .A2(new_n281), .A3(KEYINPUT98), .ZN(new_n327));
  AOI21_X1  g126(.A(new_n324), .B1(new_n326), .B2(new_n327), .ZN(new_n328));
  AOI22_X1  g127(.A1(new_n315), .A2(new_n328), .B1(KEYINPUT41), .B2(new_n255), .ZN(new_n329));
  AND2_X1   g128(.A1(new_n323), .A2(new_n329), .ZN(new_n330));
  XNOR2_X1  g129(.A(G190gat), .B(G218gat), .ZN(new_n331));
  INV_X1    g130(.A(new_n331), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n330), .A2(new_n332), .ZN(new_n333));
  OAI21_X1  g132(.A(new_n259), .B1(new_n333), .B2(KEYINPUT99), .ZN(new_n334));
  XNOR2_X1  g133(.A(new_n330), .B(new_n332), .ZN(new_n335));
  AND2_X1   g134(.A1(new_n334), .A2(new_n335), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n334), .A2(new_n335), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  NOR2_X1   g137(.A1(new_n254), .A2(new_n338), .ZN(new_n339));
  XNOR2_X1  g138(.A(G120gat), .B(G148gat), .ZN(new_n340));
  XNOR2_X1  g139(.A(G176gat), .B(G204gat), .ZN(new_n341));
  XOR2_X1   g140(.A(new_n340), .B(new_n341), .Z(new_n342));
  INV_X1    g141(.A(new_n342), .ZN(new_n343));
  OR2_X1    g142(.A1(new_n269), .A2(KEYINPUT101), .ZN(new_n344));
  NAND2_X1  g143(.A1(new_n269), .A2(KEYINPUT101), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n344), .A2(new_n278), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g145(.A1(new_n326), .A2(new_n327), .ZN(new_n347));
  NAND3_X1  g146(.A1(new_n346), .A2(new_n347), .A3(new_n227), .ZN(new_n348));
  INV_X1    g147(.A(new_n348), .ZN(new_n349));
  INV_X1    g148(.A(new_n215), .ZN(new_n350));
  AOI21_X1  g149(.A(new_n202), .B1(new_n208), .B2(new_n217), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT93), .B1(new_n351), .B2(new_n222), .ZN(new_n352));
  INV_X1    g151(.A(new_n226), .ZN(new_n353));
  OAI21_X1  g152(.A(new_n350), .B1(new_n352), .B2(new_n353), .ZN(new_n354));
  AOI21_X1  g153(.A(KEYINPUT100), .B1(new_n284), .B2(new_n354), .ZN(new_n355));
  INV_X1    g154(.A(new_n355), .ZN(new_n356));
  NAND3_X1  g155(.A1(new_n284), .A2(new_n354), .A3(KEYINPUT100), .ZN(new_n357));
  AOI21_X1  g156(.A(new_n349), .B1(new_n356), .B2(new_n357), .ZN(new_n358));
  NAND2_X1  g157(.A1(G230gat), .A2(G233gat), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n358), .A2(new_n359), .ZN(new_n360));
  AOI21_X1  g159(.A(new_n343), .B1(new_n360), .B2(KEYINPUT102), .ZN(new_n361));
  INV_X1    g160(.A(KEYINPUT10), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT100), .ZN(new_n363));
  NOR3_X1   g162(.A1(new_n328), .A2(new_n363), .A3(new_n227), .ZN(new_n364));
  OAI211_X1 g163(.A(new_n362), .B(new_n348), .C1(new_n364), .C2(new_n355), .ZN(new_n365));
  NAND4_X1  g164(.A1(new_n234), .A2(KEYINPUT10), .A3(new_n235), .A4(new_n328), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n365), .A2(new_n366), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n367), .A2(new_n359), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT102), .ZN(new_n369));
  OAI21_X1  g168(.A(new_n369), .B1(new_n358), .B2(new_n359), .ZN(new_n370));
  NAND3_X1  g169(.A1(new_n361), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  INV_X1    g170(.A(new_n359), .ZN(new_n372));
  AOI21_X1  g171(.A(new_n372), .B1(new_n365), .B2(new_n366), .ZN(new_n373));
  OAI21_X1  g172(.A(new_n343), .B1(new_n360), .B2(new_n373), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n371), .A2(new_n374), .ZN(new_n375));
  INV_X1    g174(.A(new_n375), .ZN(new_n376));
  NAND2_X1  g175(.A1(new_n339), .A2(new_n376), .ZN(new_n377));
  OAI21_X1  g176(.A(new_n246), .B1(new_n316), .B2(new_n322), .ZN(new_n378));
  NAND2_X1  g177(.A1(G229gat), .A2(G233gat), .ZN(new_n379));
  OR2_X1    g178(.A1(new_n246), .A2(new_n319), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n378), .A2(new_n379), .A3(new_n380), .ZN(new_n381));
  INV_X1    g180(.A(KEYINPUT18), .ZN(new_n382));
  XNOR2_X1  g181(.A(new_n246), .B(new_n319), .ZN(new_n383));
  XOR2_X1   g182(.A(new_n379), .B(KEYINPUT13), .Z(new_n384));
  AOI22_X1  g183(.A1(new_n381), .A2(new_n382), .B1(new_n383), .B2(new_n384), .ZN(new_n385));
  NAND4_X1  g184(.A1(new_n378), .A2(KEYINPUT18), .A3(new_n379), .A4(new_n380), .ZN(new_n386));
  AND2_X1   g185(.A1(new_n386), .A2(KEYINPUT88), .ZN(new_n387));
  NOR2_X1   g186(.A1(new_n386), .A2(KEYINPUT88), .ZN(new_n388));
  OAI21_X1  g187(.A(new_n385), .B1(new_n387), .B2(new_n388), .ZN(new_n389));
  XNOR2_X1  g188(.A(G113gat), .B(G141gat), .ZN(new_n390));
  XNOR2_X1  g189(.A(new_n390), .B(G197gat), .ZN(new_n391));
  XOR2_X1   g190(.A(KEYINPUT11), .B(G169gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  XOR2_X1   g192(.A(new_n393), .B(KEYINPUT12), .Z(new_n394));
  NAND2_X1  g193(.A1(new_n389), .A2(new_n394), .ZN(new_n395));
  INV_X1    g194(.A(new_n394), .ZN(new_n396));
  OAI211_X1 g195(.A(new_n396), .B(new_n385), .C1(new_n387), .C2(new_n388), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n395), .A2(new_n397), .ZN(new_n398));
  XNOR2_X1  g197(.A(G8gat), .B(G36gat), .ZN(new_n399));
  XNOR2_X1  g198(.A(G64gat), .B(G92gat), .ZN(new_n400));
  XOR2_X1   g199(.A(new_n399), .B(new_n400), .Z(new_n401));
  INV_X1    g200(.A(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT74), .ZN(new_n403));
  XNOR2_X1  g202(.A(G197gat), .B(G204gat), .ZN(new_n404));
  NAND2_X1  g203(.A1(G211gat), .A2(G218gat), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT22), .ZN(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NAND2_X1  g206(.A1(new_n404), .A2(new_n407), .ZN(new_n408));
  INV_X1    g207(.A(KEYINPUT73), .ZN(new_n409));
  OAI21_X1  g208(.A(new_n403), .B1(new_n408), .B2(new_n409), .ZN(new_n410));
  XOR2_X1   g209(.A(G211gat), .B(G218gat), .Z(new_n411));
  OAI21_X1  g210(.A(KEYINPUT73), .B1(new_n411), .B2(KEYINPUT74), .ZN(new_n412));
  AOI22_X1  g211(.A1(new_n410), .A2(new_n411), .B1(new_n412), .B2(new_n408), .ZN(new_n413));
  INV_X1    g212(.A(G226gat), .ZN(new_n414));
  INV_X1    g213(.A(G233gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  INV_X1    g215(.A(G183gat), .ZN(new_n417));
  INV_X1    g216(.A(G190gat), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n417), .A2(new_n418), .ZN(new_n419));
  NAND2_X1  g218(.A1(G183gat), .A2(G190gat), .ZN(new_n420));
  INV_X1    g219(.A(KEYINPUT66), .ZN(new_n421));
  OAI211_X1 g220(.A(new_n419), .B(new_n420), .C1(new_n421), .C2(KEYINPUT24), .ZN(new_n422));
  OR2_X1    g221(.A1(new_n421), .A2(KEYINPUT24), .ZN(new_n423));
  OAI211_X1 g222(.A(new_n422), .B(KEYINPUT25), .C1(new_n420), .C2(new_n423), .ZN(new_n424));
  NOR2_X1   g223(.A1(G169gat), .A2(G176gat), .ZN(new_n425));
  OR3_X1    g224(.A1(new_n425), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n426));
  OAI21_X1  g225(.A(KEYINPUT65), .B1(new_n425), .B2(KEYINPUT23), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n425), .A2(KEYINPUT23), .ZN(new_n428));
  INV_X1    g227(.A(G169gat), .ZN(new_n429));
  INV_X1    g228(.A(G176gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(new_n431), .ZN(new_n432));
  NAND4_X1  g231(.A1(new_n426), .A2(new_n427), .A3(new_n428), .A4(new_n432), .ZN(new_n433));
  OR2_X1    g232(.A1(new_n424), .A2(new_n433), .ZN(new_n434));
  INV_X1    g233(.A(KEYINPUT25), .ZN(new_n435));
  OAI211_X1 g234(.A(KEYINPUT64), .B(KEYINPUT24), .C1(G183gat), .C2(G190gat), .ZN(new_n436));
  INV_X1    g235(.A(new_n420), .ZN(new_n437));
  OAI211_X1 g236(.A(new_n436), .B(new_n437), .C1(KEYINPUT64), .C2(KEYINPUT24), .ZN(new_n438));
  OAI21_X1  g237(.A(new_n438), .B1(new_n436), .B2(new_n437), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n435), .B1(new_n433), .B2(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n434), .A2(new_n440), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT67), .ZN(new_n442));
  XNOR2_X1  g241(.A(KEYINPUT27), .B(G183gat), .ZN(new_n443));
  AOI21_X1  g242(.A(new_n442), .B1(new_n443), .B2(new_n418), .ZN(new_n444));
  OR2_X1    g243(.A1(new_n444), .A2(KEYINPUT28), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n425), .A2(KEYINPUT26), .ZN(new_n446));
  INV_X1    g245(.A(KEYINPUT26), .ZN(new_n447));
  OAI21_X1  g246(.A(new_n447), .B1(G169gat), .B2(G176gat), .ZN(new_n448));
  OAI211_X1 g247(.A(new_n446), .B(new_n420), .C1(new_n431), .C2(new_n448), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n449), .B1(new_n444), .B2(KEYINPUT28), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n445), .A2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n441), .A2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT29), .ZN(new_n453));
  AOI21_X1  g252(.A(new_n416), .B1(new_n452), .B2(new_n453), .ZN(new_n454));
  AOI22_X1  g253(.A1(new_n434), .A2(new_n440), .B1(new_n450), .B2(new_n445), .ZN(new_n455));
  NOR3_X1   g254(.A1(new_n455), .A2(new_n414), .A3(new_n415), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n413), .B1(new_n454), .B2(new_n456), .ZN(new_n457));
  OAI22_X1  g256(.A1(new_n455), .A2(KEYINPUT29), .B1(new_n414), .B2(new_n415), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n412), .A2(new_n408), .ZN(new_n459));
  XNOR2_X1  g258(.A(G211gat), .B(G218gat), .ZN(new_n460));
  INV_X1    g259(.A(G197gat), .ZN(new_n461));
  INV_X1    g260(.A(G204gat), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n461), .A2(new_n462), .ZN(new_n463));
  NAND2_X1  g262(.A1(G197gat), .A2(G204gat), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n463), .A2(new_n464), .B1(new_n406), .B2(new_n405), .ZN(new_n465));
  AOI21_X1  g264(.A(KEYINPUT74), .B1(new_n465), .B2(KEYINPUT73), .ZN(new_n466));
  OAI21_X1  g265(.A(new_n459), .B1(new_n460), .B2(new_n466), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n452), .A2(new_n416), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n458), .A2(new_n467), .A3(new_n468), .ZN(new_n469));
  AOI21_X1  g268(.A(new_n402), .B1(new_n457), .B2(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT75), .ZN(new_n471));
  OAI21_X1  g270(.A(KEYINPUT30), .B1(new_n470), .B2(new_n471), .ZN(new_n472));
  AND3_X1   g271(.A1(new_n458), .A2(new_n467), .A3(new_n468), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n467), .B1(new_n458), .B2(new_n468), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n401), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT30), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT75), .A3(new_n476), .ZN(new_n477));
  NAND3_X1  g276(.A1(new_n457), .A2(new_n402), .A3(new_n469), .ZN(new_n478));
  AND3_X1   g277(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n479));
  XNOR2_X1  g278(.A(G1gat), .B(G29gat), .ZN(new_n480));
  XNOR2_X1  g279(.A(new_n480), .B(KEYINPUT0), .ZN(new_n481));
  XNOR2_X1  g280(.A(G57gat), .B(G85gat), .ZN(new_n482));
  XOR2_X1   g281(.A(new_n481), .B(new_n482), .Z(new_n483));
  NAND2_X1  g282(.A1(G225gat), .A2(G233gat), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  INV_X1    g284(.A(G120gat), .ZN(new_n486));
  NAND2_X1  g285(.A1(new_n486), .A2(G113gat), .ZN(new_n487));
  INV_X1    g286(.A(G113gat), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G120gat), .ZN(new_n489));
  AOI21_X1  g288(.A(KEYINPUT1), .B1(new_n487), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(G134gat), .ZN(new_n491));
  OR2_X1    g290(.A1(new_n491), .A2(KEYINPUT68), .ZN(new_n492));
  NOR2_X1   g291(.A1(new_n490), .A2(new_n492), .ZN(new_n493));
  AOI211_X1 g292(.A(KEYINPUT1), .B(G134gat), .C1(new_n487), .C2(new_n489), .ZN(new_n494));
  OAI21_X1  g293(.A(G127gat), .B1(new_n493), .B2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n490), .A2(new_n491), .ZN(new_n496));
  OAI211_X1 g295(.A(new_n496), .B(new_n232), .C1(new_n490), .C2(new_n492), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n495), .A2(new_n497), .ZN(new_n498));
  XOR2_X1   g297(.A(G141gat), .B(G148gat), .Z(new_n499));
  INV_X1    g298(.A(G155gat), .ZN(new_n500));
  OAI21_X1  g299(.A(KEYINPUT2), .B1(new_n500), .B2(new_n258), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n499), .A2(new_n501), .ZN(new_n502));
  XNOR2_X1  g301(.A(G155gat), .B(G162gat), .ZN(new_n503));
  INV_X1    g302(.A(new_n503), .ZN(new_n504));
  NAND2_X1  g303(.A1(new_n502), .A2(new_n504), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n499), .A2(new_n503), .A3(new_n501), .ZN(new_n506));
  AND2_X1   g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NOR2_X1   g306(.A1(new_n498), .A2(new_n507), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n505), .A2(new_n506), .ZN(new_n509));
  AOI21_X1  g308(.A(new_n509), .B1(new_n495), .B2(new_n497), .ZN(new_n510));
  OAI21_X1  g309(.A(new_n485), .B1(new_n508), .B2(new_n510), .ZN(new_n511));
  NAND2_X1  g310(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  AND2_X1   g311(.A1(new_n495), .A2(new_n497), .ZN(new_n513));
  NAND2_X1  g312(.A1(new_n509), .A2(KEYINPUT3), .ZN(new_n514));
  INV_X1    g313(.A(KEYINPUT3), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n505), .A2(new_n515), .A3(new_n506), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n513), .A2(new_n514), .A3(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT4), .ZN(new_n518));
  AND3_X1   g317(.A1(new_n498), .A2(new_n518), .A3(new_n507), .ZN(new_n519));
  AOI21_X1  g318(.A(new_n518), .B1(new_n498), .B2(new_n507), .ZN(new_n520));
  OAI211_X1 g319(.A(new_n517), .B(new_n484), .C1(new_n519), .C2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n512), .A2(new_n521), .A3(KEYINPUT76), .ZN(new_n522));
  INV_X1    g321(.A(new_n522), .ZN(new_n523));
  AOI21_X1  g322(.A(new_n512), .B1(new_n521), .B2(KEYINPUT76), .ZN(new_n524));
  OAI21_X1  g323(.A(new_n483), .B1(new_n523), .B2(new_n524), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n521), .A2(KEYINPUT76), .ZN(new_n526));
  NAND3_X1  g325(.A1(new_n526), .A2(KEYINPUT5), .A3(new_n511), .ZN(new_n527));
  INV_X1    g326(.A(new_n483), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n527), .A2(new_n522), .A3(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(KEYINPUT6), .ZN(new_n530));
  NAND3_X1  g329(.A1(new_n525), .A2(new_n529), .A3(new_n530), .ZN(new_n531));
  NOR2_X1   g330(.A1(new_n523), .A2(new_n524), .ZN(new_n532));
  NAND3_X1  g331(.A1(new_n532), .A2(KEYINPUT6), .A3(new_n528), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n531), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n479), .A2(new_n534), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT82), .ZN(new_n536));
  XNOR2_X1  g335(.A(G78gat), .B(G106gat), .ZN(new_n537));
  XNOR2_X1  g336(.A(KEYINPUT31), .B(G50gat), .ZN(new_n538));
  XNOR2_X1  g337(.A(new_n537), .B(new_n538), .ZN(new_n539));
  INV_X1    g338(.A(KEYINPUT79), .ZN(new_n540));
  INV_X1    g339(.A(G22gat), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g341(.A1(G228gat), .A2(G233gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n516), .A2(new_n453), .ZN(new_n544));
  AOI21_X1  g343(.A(new_n543), .B1(new_n544), .B2(new_n467), .ZN(new_n545));
  OAI211_X1 g344(.A(new_n459), .B(new_n453), .C1(new_n460), .C2(new_n466), .ZN(new_n546));
  AOI21_X1  g345(.A(new_n507), .B1(new_n546), .B2(new_n515), .ZN(new_n547));
  OAI21_X1  g346(.A(new_n545), .B1(new_n547), .B2(KEYINPUT78), .ZN(new_n548));
  AOI21_X1  g347(.A(KEYINPUT3), .B1(new_n413), .B2(new_n453), .ZN(new_n549));
  INV_X1    g348(.A(KEYINPUT78), .ZN(new_n550));
  NOR3_X1   g349(.A1(new_n549), .A2(new_n550), .A3(new_n507), .ZN(new_n551));
  NOR2_X1   g350(.A1(new_n548), .A2(new_n551), .ZN(new_n552));
  OAI21_X1  g351(.A(new_n453), .B1(new_n465), .B2(new_n411), .ZN(new_n553));
  NOR2_X1   g352(.A1(new_n408), .A2(new_n460), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n515), .B1(new_n553), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n555), .A2(new_n509), .ZN(new_n556));
  AOI22_X1  g355(.A1(KEYINPUT77), .A2(new_n556), .B1(new_n544), .B2(new_n467), .ZN(new_n557));
  INV_X1    g356(.A(KEYINPUT77), .ZN(new_n558));
  NAND3_X1  g357(.A1(new_n555), .A2(new_n558), .A3(new_n509), .ZN(new_n559));
  AOI22_X1  g358(.A1(new_n557), .A2(new_n559), .B1(G228gat), .B2(G233gat), .ZN(new_n560));
  OAI21_X1  g359(.A(new_n542), .B1(new_n552), .B2(new_n560), .ZN(new_n561));
  NOR2_X1   g360(.A1(new_n540), .A2(new_n541), .ZN(new_n562));
  INV_X1    g361(.A(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n561), .A2(new_n563), .ZN(new_n564));
  NAND2_X1  g363(.A1(new_n547), .A2(KEYINPUT78), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n550), .B1(new_n549), .B2(new_n507), .ZN(new_n566));
  NAND3_X1  g365(.A1(new_n565), .A2(new_n566), .A3(new_n545), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n556), .A2(KEYINPUT77), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n544), .A2(new_n467), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n568), .A2(new_n569), .A3(new_n559), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n570), .A2(new_n543), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  NAND3_X1  g371(.A1(new_n572), .A2(KEYINPUT79), .A3(G22gat), .ZN(new_n573));
  AOI21_X1  g372(.A(new_n539), .B1(new_n564), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n539), .ZN(new_n575));
  NOR2_X1   g374(.A1(new_n541), .A2(KEYINPUT80), .ZN(new_n576));
  AOI21_X1  g375(.A(new_n576), .B1(new_n567), .B2(new_n571), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n567), .A2(new_n571), .A3(new_n576), .ZN(new_n579));
  AOI21_X1  g378(.A(new_n575), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  OAI21_X1  g379(.A(KEYINPUT81), .B1(new_n574), .B2(new_n580), .ZN(new_n581));
  AOI21_X1  g380(.A(new_n562), .B1(new_n572), .B2(new_n542), .ZN(new_n582));
  AOI211_X1 g381(.A(new_n540), .B(new_n541), .C1(new_n567), .C2(new_n571), .ZN(new_n583));
  OAI21_X1  g382(.A(new_n575), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT81), .ZN(new_n585));
  INV_X1    g384(.A(new_n579), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n539), .B1(new_n586), .B2(new_n577), .ZN(new_n587));
  NAND3_X1  g386(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n588));
  AOI21_X1  g387(.A(KEYINPUT35), .B1(new_n581), .B2(new_n588), .ZN(new_n589));
  INV_X1    g388(.A(KEYINPUT82), .ZN(new_n590));
  NAND3_X1  g389(.A1(new_n479), .A2(new_n534), .A3(new_n590), .ZN(new_n591));
  XNOR2_X1  g390(.A(G15gat), .B(G43gat), .ZN(new_n592));
  XNOR2_X1  g391(.A(new_n592), .B(KEYINPUT70), .ZN(new_n593));
  XNOR2_X1  g392(.A(G71gat), .B(G99gat), .ZN(new_n594));
  XNOR2_X1  g393(.A(new_n593), .B(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n595), .A2(KEYINPUT33), .ZN(new_n596));
  NOR2_X1   g395(.A1(new_n596), .A2(KEYINPUT69), .ZN(new_n597));
  NAND2_X1  g396(.A1(new_n452), .A2(new_n498), .ZN(new_n598));
  NAND2_X1  g397(.A1(new_n455), .A2(new_n513), .ZN(new_n599));
  NAND2_X1  g398(.A1(new_n598), .A2(new_n599), .ZN(new_n600));
  INV_X1    g399(.A(G227gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(new_n415), .ZN(new_n602));
  INV_X1    g401(.A(new_n602), .ZN(new_n603));
  OAI211_X1 g402(.A(KEYINPUT32), .B(new_n597), .C1(new_n600), .C2(new_n603), .ZN(new_n604));
  INV_X1    g403(.A(KEYINPUT32), .ZN(new_n605));
  AND2_X1   g404(.A1(new_n598), .A2(new_n599), .ZN(new_n606));
  AOI21_X1  g405(.A(new_n605), .B1(new_n606), .B2(new_n602), .ZN(new_n607));
  NAND4_X1  g406(.A1(new_n598), .A2(new_n602), .A3(new_n599), .A4(new_n595), .ZN(new_n608));
  AOI21_X1  g407(.A(KEYINPUT69), .B1(new_n608), .B2(new_n596), .ZN(new_n609));
  OAI21_X1  g408(.A(new_n604), .B1(new_n607), .B2(new_n609), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n600), .A2(new_n603), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT34), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT34), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n600), .A2(new_n613), .A3(new_n603), .ZN(new_n614));
  AND2_X1   g413(.A1(new_n612), .A2(new_n614), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n610), .A2(new_n615), .ZN(new_n616));
  NAND2_X1  g415(.A1(new_n612), .A2(new_n614), .ZN(new_n617));
  OAI211_X1 g416(.A(new_n617), .B(new_n604), .C1(new_n607), .C2(new_n609), .ZN(new_n618));
  INV_X1    g417(.A(KEYINPUT72), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n616), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  NAND3_X1  g419(.A1(new_n610), .A2(new_n615), .A3(KEYINPUT72), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n620), .A2(new_n621), .ZN(new_n622));
  NAND4_X1  g421(.A1(new_n536), .A2(new_n589), .A3(new_n591), .A4(new_n622), .ZN(new_n623));
  AND2_X1   g422(.A1(new_n616), .A2(new_n618), .ZN(new_n624));
  AND3_X1   g423(.A1(new_n584), .A2(new_n585), .A3(new_n587), .ZN(new_n625));
  AOI21_X1  g424(.A(new_n585), .B1(new_n584), .B2(new_n587), .ZN(new_n626));
  OAI21_X1  g425(.A(new_n624), .B1(new_n625), .B2(new_n626), .ZN(new_n627));
  OAI21_X1  g426(.A(KEYINPUT35), .B1(new_n627), .B2(new_n535), .ZN(new_n628));
  NAND2_X1  g427(.A1(new_n623), .A2(new_n628), .ZN(new_n629));
  NAND2_X1  g428(.A1(new_n581), .A2(new_n588), .ZN(new_n630));
  OAI21_X1  g429(.A(new_n517), .B1(new_n519), .B2(new_n520), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n631), .A2(new_n485), .ZN(new_n632));
  OR2_X1    g431(.A1(new_n508), .A2(new_n510), .ZN(new_n633));
  OAI211_X1 g432(.A(new_n632), .B(KEYINPUT39), .C1(new_n485), .C2(new_n633), .ZN(new_n634));
  OAI211_X1 g433(.A(new_n634), .B(new_n483), .C1(KEYINPUT39), .C2(new_n632), .ZN(new_n635));
  INV_X1    g434(.A(KEYINPUT40), .ZN(new_n636));
  AOI22_X1  g435(.A1(new_n635), .A2(new_n636), .B1(new_n532), .B2(new_n528), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n472), .A2(new_n477), .A3(new_n478), .ZN(new_n638));
  OAI211_X1 g437(.A(new_n637), .B(new_n638), .C1(new_n636), .C2(new_n635), .ZN(new_n639));
  OAI21_X1  g438(.A(KEYINPUT37), .B1(new_n473), .B2(new_n474), .ZN(new_n640));
  INV_X1    g439(.A(KEYINPUT37), .ZN(new_n641));
  NAND3_X1  g440(.A1(new_n457), .A2(new_n641), .A3(new_n469), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n401), .B1(new_n640), .B2(new_n642), .ZN(new_n643));
  INV_X1    g442(.A(KEYINPUT38), .ZN(new_n644));
  AOI21_X1  g443(.A(new_n470), .B1(new_n643), .B2(new_n644), .ZN(new_n645));
  OAI21_X1  g444(.A(new_n645), .B1(new_n644), .B2(new_n643), .ZN(new_n646));
  OAI211_X1 g445(.A(new_n630), .B(new_n639), .C1(new_n646), .C2(new_n534), .ZN(new_n647));
  NAND2_X1  g446(.A1(new_n624), .A2(KEYINPUT36), .ZN(new_n648));
  XNOR2_X1  g447(.A(KEYINPUT71), .B(KEYINPUT36), .ZN(new_n649));
  INV_X1    g448(.A(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n648), .B1(new_n622), .B2(new_n650), .ZN(new_n651));
  NAND3_X1  g450(.A1(new_n535), .A2(new_n581), .A3(new_n588), .ZN(new_n652));
  NAND3_X1  g451(.A1(new_n647), .A2(new_n651), .A3(new_n652), .ZN(new_n653));
  AND3_X1   g452(.A1(new_n629), .A2(KEYINPUT83), .A3(new_n653), .ZN(new_n654));
  AOI21_X1  g453(.A(KEYINPUT83), .B1(new_n629), .B2(new_n653), .ZN(new_n655));
  OAI21_X1  g454(.A(new_n398), .B1(new_n654), .B2(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT89), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n656), .A2(new_n657), .ZN(new_n658));
  OAI211_X1 g457(.A(KEYINPUT89), .B(new_n398), .C1(new_n654), .C2(new_n655), .ZN(new_n659));
  AOI21_X1  g458(.A(new_n377), .B1(new_n658), .B2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n534), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  XNOR2_X1  g461(.A(new_n662), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g462(.A(KEYINPUT16), .B(G8gat), .Z(new_n664));
  AND3_X1   g463(.A1(new_n660), .A2(new_n638), .A3(new_n664), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n245), .B1(new_n660), .B2(new_n638), .ZN(new_n666));
  OAI21_X1  g465(.A(KEYINPUT42), .B1(new_n665), .B2(new_n666), .ZN(new_n667));
  OAI21_X1  g466(.A(new_n667), .B1(KEYINPUT42), .B2(new_n665), .ZN(G1325gat));
  INV_X1    g467(.A(G15gat), .ZN(new_n669));
  NAND3_X1  g468(.A1(new_n660), .A2(new_n669), .A3(new_n622), .ZN(new_n670));
  INV_X1    g469(.A(new_n651), .ZN(new_n671));
  AND2_X1   g470(.A1(new_n660), .A2(new_n671), .ZN(new_n672));
  OAI21_X1  g471(.A(new_n670), .B1(new_n672), .B2(new_n669), .ZN(G1326gat));
  INV_X1    g472(.A(new_n630), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n660), .A2(new_n674), .ZN(new_n675));
  XNOR2_X1  g474(.A(KEYINPUT43), .B(G22gat), .ZN(new_n676));
  XNOR2_X1  g475(.A(new_n675), .B(new_n676), .ZN(G1327gat));
  NAND3_X1  g476(.A1(new_n254), .A2(new_n376), .A3(new_n338), .ZN(new_n678));
  AOI21_X1  g477(.A(new_n678), .B1(new_n658), .B2(new_n659), .ZN(new_n679));
  NAND3_X1  g478(.A1(new_n679), .A2(new_n290), .A3(new_n661), .ZN(new_n680));
  XNOR2_X1  g479(.A(new_n680), .B(KEYINPUT45), .ZN(new_n681));
  INV_X1    g480(.A(KEYINPUT105), .ZN(new_n682));
  INV_X1    g481(.A(new_n338), .ZN(new_n683));
  AOI21_X1  g482(.A(new_n683), .B1(new_n629), .B2(new_n653), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT44), .ZN(new_n685));
  AOI21_X1  g484(.A(new_n682), .B1(new_n684), .B2(new_n685), .ZN(new_n686));
  NAND2_X1  g485(.A1(new_n629), .A2(new_n653), .ZN(new_n687));
  INV_X1    g486(.A(KEYINPUT83), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n687), .A2(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n629), .A2(KEYINPUT83), .A3(new_n653), .ZN(new_n690));
  AOI21_X1  g489(.A(new_n683), .B1(new_n689), .B2(new_n690), .ZN(new_n691));
  OAI21_X1  g490(.A(new_n686), .B1(new_n691), .B2(new_n685), .ZN(new_n692));
  OAI21_X1  g491(.A(new_n338), .B1(new_n654), .B2(new_n655), .ZN(new_n693));
  NAND3_X1  g492(.A1(new_n693), .A2(new_n682), .A3(KEYINPUT44), .ZN(new_n694));
  XNOR2_X1  g493(.A(new_n375), .B(KEYINPUT103), .ZN(new_n695));
  NAND3_X1  g494(.A1(new_n254), .A2(new_n398), .A3(new_n695), .ZN(new_n696));
  XNOR2_X1  g495(.A(new_n696), .B(KEYINPUT104), .ZN(new_n697));
  NAND4_X1  g496(.A1(new_n692), .A2(new_n661), .A3(new_n694), .A4(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n290), .B1(new_n698), .B2(KEYINPUT106), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n699), .B1(KEYINPUT106), .B2(new_n698), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n681), .A2(new_n700), .ZN(G1328gat));
  NAND3_X1  g500(.A1(new_n679), .A2(new_n291), .A3(new_n638), .ZN(new_n702));
  OR2_X1    g501(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n703));
  NAND3_X1  g502(.A1(new_n692), .A2(new_n694), .A3(new_n697), .ZN(new_n704));
  OAI21_X1  g503(.A(G36gat), .B1(new_n704), .B2(new_n479), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(KEYINPUT46), .ZN(new_n706));
  NAND3_X1  g505(.A1(new_n703), .A2(new_n705), .A3(new_n706), .ZN(G1329gat));
  NAND4_X1  g506(.A1(new_n692), .A2(new_n671), .A3(new_n694), .A4(new_n697), .ZN(new_n708));
  NAND2_X1  g507(.A1(new_n708), .A2(G43gat), .ZN(new_n709));
  NAND3_X1  g508(.A1(new_n679), .A2(new_n287), .A3(new_n622), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(new_n710), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT47), .B1(new_n711), .B2(KEYINPUT107), .ZN(new_n712));
  INV_X1    g511(.A(KEYINPUT107), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT47), .ZN(new_n714));
  AOI211_X1 g513(.A(new_n713), .B(new_n714), .C1(new_n709), .C2(new_n710), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n712), .A2(new_n715), .ZN(G1330gat));
  NAND3_X1  g515(.A1(new_n679), .A2(new_n285), .A3(new_n674), .ZN(new_n717));
  NAND4_X1  g516(.A1(new_n692), .A2(new_n674), .A3(new_n694), .A4(new_n697), .ZN(new_n718));
  INV_X1    g517(.A(KEYINPUT108), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g519(.A1(new_n720), .A2(G50gat), .ZN(new_n721));
  NOR2_X1   g520(.A1(new_n718), .A2(new_n719), .ZN(new_n722));
  OAI211_X1 g521(.A(KEYINPUT48), .B(new_n717), .C1(new_n721), .C2(new_n722), .ZN(new_n723));
  NAND2_X1  g522(.A1(new_n718), .A2(G50gat), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n724), .A2(new_n717), .ZN(new_n725));
  INV_X1    g524(.A(KEYINPUT48), .ZN(new_n726));
  NAND2_X1  g525(.A1(new_n725), .A2(new_n726), .ZN(new_n727));
  NAND2_X1  g526(.A1(new_n723), .A2(new_n727), .ZN(G1331gat));
  NOR4_X1   g527(.A1(new_n254), .A2(new_n695), .A3(new_n398), .A4(new_n338), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n687), .A2(new_n729), .ZN(new_n730));
  INV_X1    g529(.A(new_n730), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n731), .A2(new_n661), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n732), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g532(.A1(new_n730), .A2(new_n479), .ZN(new_n734));
  NOR2_X1   g533(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n735));
  AND2_X1   g534(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(new_n737));
  OAI21_X1  g536(.A(new_n737), .B1(new_n734), .B2(new_n735), .ZN(G1333gat));
  OAI21_X1  g537(.A(G71gat), .B1(new_n730), .B2(new_n651), .ZN(new_n739));
  NAND2_X1  g538(.A1(new_n622), .A2(new_n205), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n739), .B1(new_n730), .B2(new_n740), .ZN(new_n741));
  XNOR2_X1  g540(.A(new_n741), .B(KEYINPUT110), .ZN(new_n742));
  XOR2_X1   g541(.A(KEYINPUT109), .B(KEYINPUT50), .Z(new_n743));
  XNOR2_X1  g542(.A(new_n742), .B(new_n743), .ZN(G1334gat));
  NOR2_X1   g543(.A1(new_n730), .A2(new_n630), .ZN(new_n745));
  XNOR2_X1  g544(.A(new_n745), .B(new_n206), .ZN(G1335gat));
  AND2_X1   g545(.A1(new_n395), .A2(new_n397), .ZN(new_n747));
  NAND3_X1  g546(.A1(new_n684), .A2(new_n747), .A3(new_n254), .ZN(new_n748));
  XNOR2_X1  g547(.A(new_n748), .B(KEYINPUT51), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n749), .A2(new_n376), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n750), .A2(new_n274), .A3(new_n661), .ZN(new_n751));
  INV_X1    g550(.A(new_n254), .ZN(new_n752));
  NOR3_X1   g551(.A1(new_n752), .A2(new_n398), .A3(new_n376), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n692), .A2(new_n694), .A3(new_n753), .ZN(new_n754));
  OAI21_X1  g553(.A(G85gat), .B1(new_n754), .B2(new_n534), .ZN(new_n755));
  NAND2_X1  g554(.A1(new_n751), .A2(new_n755), .ZN(G1336gat));
  NOR2_X1   g555(.A1(new_n749), .A2(new_n695), .ZN(new_n757));
  NAND3_X1  g556(.A1(new_n757), .A2(new_n275), .A3(new_n638), .ZN(new_n758));
  OAI21_X1  g557(.A(G92gat), .B1(new_n754), .B2(new_n479), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n758), .A2(new_n759), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(KEYINPUT52), .ZN(new_n761));
  INV_X1    g560(.A(KEYINPUT52), .ZN(new_n762));
  NAND3_X1  g561(.A1(new_n758), .A2(new_n759), .A3(new_n762), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n761), .A2(new_n763), .ZN(G1337gat));
  NAND3_X1  g563(.A1(new_n750), .A2(new_n263), .A3(new_n622), .ZN(new_n765));
  OAI21_X1  g564(.A(G99gat), .B1(new_n754), .B2(new_n651), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n765), .A2(new_n766), .ZN(new_n767));
  INV_X1    g566(.A(KEYINPUT111), .ZN(new_n768));
  NAND2_X1  g567(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n765), .A2(new_n766), .A3(KEYINPUT111), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(G1338gat));
  NAND3_X1  g570(.A1(new_n757), .A2(new_n264), .A3(new_n674), .ZN(new_n772));
  XOR2_X1   g571(.A(KEYINPUT112), .B(G106gat), .Z(new_n773));
  OAI21_X1  g572(.A(new_n773), .B1(new_n754), .B2(new_n630), .ZN(new_n774));
  NAND2_X1  g573(.A1(new_n772), .A2(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n775), .A2(KEYINPUT53), .ZN(new_n776));
  INV_X1    g575(.A(KEYINPUT53), .ZN(new_n777));
  NAND3_X1  g576(.A1(new_n772), .A2(new_n774), .A3(new_n777), .ZN(new_n778));
  NAND2_X1  g577(.A1(new_n776), .A2(new_n778), .ZN(G1339gat));
  NOR4_X1   g578(.A1(new_n254), .A2(new_n338), .A3(new_n398), .A4(new_n375), .ZN(new_n780));
  AOI21_X1  g579(.A(new_n379), .B1(new_n378), .B2(new_n380), .ZN(new_n781));
  NOR2_X1   g580(.A1(new_n383), .A2(new_n384), .ZN(new_n782));
  OAI21_X1  g581(.A(new_n393), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n397), .A2(new_n783), .ZN(new_n784));
  INV_X1    g583(.A(new_n784), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n785), .A2(new_n375), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n365), .A2(new_n372), .A3(new_n366), .ZN(new_n787));
  NAND3_X1  g586(.A1(new_n368), .A2(KEYINPUT54), .A3(new_n787), .ZN(new_n788));
  INV_X1    g587(.A(KEYINPUT54), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n342), .B1(new_n373), .B2(new_n789), .ZN(new_n790));
  NAND3_X1  g589(.A1(new_n788), .A2(KEYINPUT55), .A3(new_n790), .ZN(new_n791));
  NAND2_X1  g590(.A1(new_n791), .A2(new_n371), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  INV_X1    g592(.A(KEYINPUT55), .ZN(new_n794));
  AND3_X1   g593(.A1(new_n365), .A2(new_n372), .A3(new_n366), .ZN(new_n795));
  NOR3_X1   g594(.A1(new_n795), .A2(new_n373), .A3(new_n789), .ZN(new_n796));
  NAND3_X1  g595(.A1(new_n367), .A2(new_n789), .A3(new_n359), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n797), .A2(new_n343), .ZN(new_n798));
  OAI21_X1  g597(.A(new_n794), .B1(new_n796), .B2(new_n798), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n793), .A2(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(new_n786), .B1(new_n800), .B2(new_n747), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n801), .A2(new_n683), .ZN(new_n802));
  NAND4_X1  g601(.A1(new_n338), .A2(new_n785), .A3(new_n793), .A4(new_n799), .ZN(new_n803));
  NAND2_X1  g602(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n780), .B1(new_n804), .B2(new_n254), .ZN(new_n805));
  NOR3_X1   g604(.A1(new_n805), .A2(new_n534), .A3(new_n627), .ZN(new_n806));
  AND2_X1   g605(.A1(new_n806), .A2(new_n479), .ZN(new_n807));
  AOI21_X1  g606(.A(G113gat), .B1(new_n807), .B2(new_n398), .ZN(new_n808));
  NOR2_X1   g607(.A1(new_n534), .A2(new_n638), .ZN(new_n809));
  AND2_X1   g608(.A1(new_n622), .A2(new_n809), .ZN(new_n810));
  INV_X1    g609(.A(new_n780), .ZN(new_n811));
  INV_X1    g610(.A(new_n803), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n683), .B2(new_n801), .ZN(new_n813));
  OAI21_X1  g612(.A(new_n811), .B1(new_n813), .B2(new_n752), .ZN(new_n814));
  AOI21_X1  g613(.A(KEYINPUT113), .B1(new_n814), .B2(new_n630), .ZN(new_n815));
  INV_X1    g614(.A(KEYINPUT113), .ZN(new_n816));
  NOR3_X1   g615(.A1(new_n805), .A2(new_n816), .A3(new_n674), .ZN(new_n817));
  OAI21_X1  g616(.A(new_n810), .B1(new_n815), .B2(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n818), .A2(KEYINPUT114), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n816), .B1(new_n805), .B2(new_n674), .ZN(new_n820));
  NAND3_X1  g619(.A1(new_n814), .A2(KEYINPUT113), .A3(new_n630), .ZN(new_n821));
  NAND2_X1  g620(.A1(new_n820), .A2(new_n821), .ZN(new_n822));
  INV_X1    g621(.A(KEYINPUT114), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n822), .A2(new_n823), .A3(new_n810), .ZN(new_n824));
  AND2_X1   g623(.A1(new_n819), .A2(new_n824), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n747), .A2(new_n488), .ZN(new_n826));
  AOI21_X1  g625(.A(new_n808), .B1(new_n825), .B2(new_n826), .ZN(G1340gat));
  AOI21_X1  g626(.A(G120gat), .B1(new_n807), .B2(new_n375), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n695), .A2(new_n486), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n828), .B1(new_n825), .B2(new_n829), .ZN(G1341gat));
  XNOR2_X1  g629(.A(KEYINPUT68), .B(G127gat), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n254), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n807), .A2(new_n752), .ZN(new_n833));
  AOI22_X1  g632(.A1(new_n825), .A2(new_n832), .B1(new_n833), .B2(new_n831), .ZN(G1342gat));
  NAND2_X1  g633(.A1(new_n338), .A2(new_n479), .ZN(new_n835));
  XNOR2_X1  g634(.A(new_n835), .B(KEYINPUT115), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n806), .A2(new_n491), .A3(new_n836), .ZN(new_n837));
  XOR2_X1   g636(.A(new_n837), .B(KEYINPUT56), .Z(new_n838));
  NAND3_X1  g637(.A1(new_n819), .A2(new_n338), .A3(new_n824), .ZN(new_n839));
  AND3_X1   g638(.A1(new_n839), .A2(KEYINPUT116), .A3(G134gat), .ZN(new_n840));
  AOI21_X1  g639(.A(KEYINPUT116), .B1(new_n839), .B2(G134gat), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n838), .B1(new_n840), .B2(new_n841), .ZN(G1343gat));
  INV_X1    g641(.A(KEYINPUT119), .ZN(new_n843));
  INV_X1    g642(.A(KEYINPUT57), .ZN(new_n844));
  NAND3_X1  g643(.A1(new_n814), .A2(new_n844), .A3(new_n674), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n651), .A2(new_n809), .ZN(new_n846));
  INV_X1    g645(.A(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n845), .A2(new_n847), .ZN(new_n848));
  XOR2_X1   g647(.A(KEYINPUT117), .B(KEYINPUT55), .Z(new_n849));
  INV_X1    g648(.A(new_n849), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n850), .B1(new_n788), .B2(new_n790), .ZN(new_n851));
  OAI21_X1  g650(.A(KEYINPUT118), .B1(new_n792), .B2(new_n851), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n849), .B1(new_n796), .B2(new_n798), .ZN(new_n853));
  INV_X1    g652(.A(KEYINPUT118), .ZN(new_n854));
  NAND4_X1  g653(.A1(new_n853), .A2(new_n854), .A3(new_n371), .A4(new_n791), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n852), .A2(new_n398), .A3(new_n855), .ZN(new_n856));
  AOI21_X1  g655(.A(new_n338), .B1(new_n856), .B2(new_n786), .ZN(new_n857));
  OAI21_X1  g656(.A(new_n254), .B1(new_n857), .B2(new_n812), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n630), .B1(new_n858), .B2(new_n811), .ZN(new_n859));
  NOR2_X1   g658(.A1(new_n859), .A2(new_n844), .ZN(new_n860));
  NOR3_X1   g659(.A1(new_n848), .A2(new_n747), .A3(new_n860), .ZN(new_n861));
  INV_X1    g660(.A(G141gat), .ZN(new_n862));
  OAI21_X1  g661(.A(new_n843), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n671), .A2(new_n630), .ZN(new_n864));
  AND3_X1   g663(.A1(new_n814), .A2(new_n661), .A3(new_n864), .ZN(new_n865));
  NAND4_X1  g664(.A1(new_n865), .A2(new_n862), .A3(new_n398), .A4(new_n479), .ZN(new_n866));
  OAI21_X1  g665(.A(new_n866), .B1(new_n861), .B2(new_n862), .ZN(new_n867));
  INV_X1    g666(.A(KEYINPUT58), .ZN(new_n868));
  AND3_X1   g667(.A1(new_n863), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n867), .B1(new_n868), .B2(new_n863), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n869), .A2(new_n870), .ZN(G1344gat));
  INV_X1    g670(.A(KEYINPUT122), .ZN(new_n872));
  NOR2_X1   g671(.A1(new_n376), .A2(new_n784), .ZN(new_n873));
  AND2_X1   g672(.A1(new_n398), .A2(new_n855), .ZN(new_n874));
  AOI21_X1  g673(.A(new_n873), .B1(new_n874), .B2(new_n852), .ZN(new_n875));
  OAI21_X1  g674(.A(new_n803), .B1(new_n875), .B2(new_n338), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n780), .B1(new_n876), .B2(new_n254), .ZN(new_n877));
  OAI211_X1 g676(.A(new_n872), .B(new_n844), .C1(new_n877), .C2(new_n630), .ZN(new_n878));
  OAI21_X1  g677(.A(KEYINPUT122), .B1(new_n859), .B2(KEYINPUT57), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n814), .A2(KEYINPUT57), .A3(new_n674), .ZN(new_n880));
  NAND3_X1  g679(.A1(new_n878), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  OAI21_X1  g680(.A(new_n375), .B1(new_n846), .B2(KEYINPUT121), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n882), .B1(KEYINPUT121), .B2(new_n846), .ZN(new_n883));
  NAND3_X1  g682(.A1(new_n881), .A2(KEYINPUT123), .A3(new_n883), .ZN(new_n884));
  NAND2_X1  g683(.A1(new_n884), .A2(G148gat), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT123), .B1(new_n881), .B2(new_n883), .ZN(new_n886));
  OAI21_X1  g685(.A(KEYINPUT59), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  INV_X1    g686(.A(G148gat), .ZN(new_n888));
  NOR2_X1   g687(.A1(new_n888), .A2(KEYINPUT59), .ZN(new_n889));
  OR2_X1    g688(.A1(new_n848), .A2(new_n860), .ZN(new_n890));
  OAI21_X1  g689(.A(new_n889), .B1(new_n890), .B2(new_n376), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n887), .A2(new_n891), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n865), .A2(new_n479), .ZN(new_n893));
  NOR3_X1   g692(.A1(new_n893), .A2(G148gat), .A3(new_n376), .ZN(new_n894));
  XNOR2_X1  g693(.A(new_n894), .B(KEYINPUT120), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n892), .A2(new_n895), .ZN(G1345gat));
  OAI21_X1  g695(.A(G155gat), .B1(new_n890), .B2(new_n254), .ZN(new_n897));
  NAND2_X1  g696(.A1(new_n752), .A2(new_n500), .ZN(new_n898));
  OAI21_X1  g697(.A(new_n897), .B1(new_n893), .B2(new_n898), .ZN(G1346gat));
  OAI21_X1  g698(.A(G162gat), .B1(new_n890), .B2(new_n683), .ZN(new_n900));
  NAND3_X1  g699(.A1(new_n865), .A2(new_n258), .A3(new_n836), .ZN(new_n901));
  NAND2_X1  g700(.A1(new_n900), .A2(new_n901), .ZN(G1347gat));
  NOR4_X1   g701(.A1(new_n805), .A2(new_n661), .A3(new_n479), .A4(new_n627), .ZN(new_n903));
  NAND3_X1  g702(.A1(new_n903), .A2(new_n429), .A3(new_n398), .ZN(new_n904));
  NOR2_X1   g703(.A1(new_n661), .A2(new_n479), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n905), .A2(new_n622), .ZN(new_n906));
  AOI21_X1  g705(.A(new_n906), .B1(new_n820), .B2(new_n821), .ZN(new_n907));
  NAND2_X1  g706(.A1(new_n907), .A2(new_n398), .ZN(new_n908));
  AND3_X1   g707(.A1(new_n908), .A2(KEYINPUT124), .A3(G169gat), .ZN(new_n909));
  AOI21_X1  g708(.A(KEYINPUT124), .B1(new_n908), .B2(G169gat), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n904), .B1(new_n909), .B2(new_n910), .ZN(G1348gat));
  INV_X1    g710(.A(new_n907), .ZN(new_n912));
  OAI21_X1  g711(.A(G176gat), .B1(new_n912), .B2(new_n695), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n903), .A2(new_n430), .A3(new_n375), .ZN(new_n914));
  NAND2_X1  g713(.A1(new_n913), .A2(new_n914), .ZN(G1349gat));
  AOI21_X1  g714(.A(new_n417), .B1(new_n907), .B2(new_n752), .ZN(new_n916));
  AND3_X1   g715(.A1(new_n903), .A2(new_n443), .A3(new_n752), .ZN(new_n917));
  NOR3_X1   g716(.A1(new_n916), .A2(KEYINPUT125), .A3(new_n917), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT60), .ZN(new_n919));
  XNOR2_X1  g718(.A(new_n918), .B(new_n919), .ZN(G1350gat));
  NAND3_X1  g719(.A1(new_n903), .A2(new_n418), .A3(new_n338), .ZN(new_n921));
  INV_X1    g720(.A(KEYINPUT61), .ZN(new_n922));
  NAND2_X1  g721(.A1(new_n907), .A2(new_n338), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n922), .B1(new_n923), .B2(G190gat), .ZN(new_n924));
  AOI211_X1 g723(.A(KEYINPUT61), .B(new_n418), .C1(new_n907), .C2(new_n338), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n921), .B1(new_n924), .B2(new_n925), .ZN(G1351gat));
  AND4_X1   g725(.A1(new_n534), .A2(new_n814), .A3(new_n638), .A4(new_n864), .ZN(new_n927));
  NAND3_X1  g726(.A1(new_n927), .A2(new_n461), .A3(new_n398), .ZN(new_n928));
  XOR2_X1   g727(.A(new_n928), .B(KEYINPUT126), .Z(new_n929));
  AND2_X1   g728(.A1(new_n651), .A2(new_n905), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n881), .A2(new_n930), .ZN(new_n931));
  OAI21_X1  g730(.A(G197gat), .B1(new_n931), .B2(new_n747), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n929), .A2(new_n932), .ZN(G1352gat));
  NAND3_X1  g732(.A1(new_n927), .A2(new_n462), .A3(new_n375), .ZN(new_n934));
  XOR2_X1   g733(.A(new_n934), .B(KEYINPUT62), .Z(new_n935));
  OAI21_X1  g734(.A(G204gat), .B1(new_n931), .B2(new_n695), .ZN(new_n936));
  NAND2_X1  g735(.A1(new_n935), .A2(new_n936), .ZN(G1353gat));
  INV_X1    g736(.A(G211gat), .ZN(new_n938));
  NAND3_X1  g737(.A1(new_n927), .A2(new_n938), .A3(new_n752), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n881), .A2(new_n752), .A3(new_n930), .ZN(new_n940));
  AND3_X1   g739(.A1(new_n940), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n941));
  AOI21_X1  g740(.A(KEYINPUT63), .B1(new_n940), .B2(G211gat), .ZN(new_n942));
  OAI21_X1  g741(.A(new_n939), .B1(new_n941), .B2(new_n942), .ZN(G1354gat));
  AOI21_X1  g742(.A(G218gat), .B1(new_n927), .B2(new_n338), .ZN(new_n944));
  XNOR2_X1  g743(.A(new_n944), .B(KEYINPUT127), .ZN(new_n945));
  INV_X1    g744(.A(G218gat), .ZN(new_n946));
  NOR3_X1   g745(.A1(new_n931), .A2(new_n946), .A3(new_n683), .ZN(new_n947));
  NOR2_X1   g746(.A1(new_n945), .A2(new_n947), .ZN(G1355gat));
endmodule


