

module locked_locked_c1355 ( G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, 
        G43GAT, G50GAT, G57GAT, G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, 
        G106GAT, G113GAT, G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, 
        G162GAT, G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT, 
        G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT, G231GAT, 
        G232GAT, G233GAT, G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, 
        G1329GAT, G1330GAT, G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, 
        G1336GAT, G1337GAT, G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, 
        G1343GAT, G1344GAT, G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, 
        G1350GAT, G1351GAT, G1352GAT, G1353GAT, G1354GAT, G1355GAT, KEYINPUT63, 
        KEYINPUT62, KEYINPUT61, KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, 
        KEYINPUT56, KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51, 
        KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46, KEYINPUT45, 
        KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41, KEYINPUT40, KEYINPUT39, 
        KEYINPUT38, KEYINPUT37, KEYINPUT36, KEYINPUT35, KEYINPUT34, KEYINPUT33, 
        KEYINPUT32, KEYINPUT31, KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, 
        KEYINPUT26, KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21, 
        KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16, KEYINPUT15, 
        KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11, KEYINPUT10, KEYINPUT9, 
        KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5, KEYINPUT4, KEYINPUT3, 
        KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127, KEYINPUT126, KEYINPUT125, 
        KEYINPUT124, KEYINPUT123, KEYINPUT122, KEYINPUT121, KEYINPUT120, 
        KEYINPUT119, KEYINPUT118, KEYINPUT117, KEYINPUT116, KEYINPUT115, 
        KEYINPUT114, KEYINPUT113, KEYINPUT112, KEYINPUT111, KEYINPUT110, 
        KEYINPUT109, KEYINPUT108, KEYINPUT107, KEYINPUT106, KEYINPUT105, 
        KEYINPUT104, KEYINPUT103, KEYINPUT102, KEYINPUT101, KEYINPUT100, 
        KEYINPUT99, KEYINPUT98, KEYINPUT97, KEYINPUT96, KEYINPUT95, KEYINPUT94, 
        KEYINPUT93, KEYINPUT92, KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, 
        KEYINPUT87, KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82, 
        KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77, KEYINPUT76, 
        KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72, KEYINPUT71, KEYINPUT70, 
        KEYINPUT69, KEYINPUT68, KEYINPUT67, KEYINPUT66, KEYINPUT65, KEYINPUT64
 );
  input G1GAT, G8GAT, G15GAT, G22GAT, G29GAT, G36GAT, G43GAT, G50GAT, G57GAT,
         G64GAT, G71GAT, G78GAT, G85GAT, G92GAT, G99GAT, G106GAT, G113GAT,
         G120GAT, G127GAT, G134GAT, G141GAT, G148GAT, G155GAT, G162GAT,
         G169GAT, G176GAT, G183GAT, G190GAT, G197GAT, G204GAT, G211GAT,
         G218GAT, G225GAT, G226GAT, G227GAT, G228GAT, G229GAT, G230GAT,
         G231GAT, G232GAT, G233GAT, KEYINPUT63, KEYINPUT62, KEYINPUT61,
         KEYINPUT60, KEYINPUT59, KEYINPUT58, KEYINPUT57, KEYINPUT56,
         KEYINPUT55, KEYINPUT54, KEYINPUT53, KEYINPUT52, KEYINPUT51,
         KEYINPUT50, KEYINPUT49, KEYINPUT48, KEYINPUT47, KEYINPUT46,
         KEYINPUT45, KEYINPUT44, KEYINPUT43, KEYINPUT42, KEYINPUT41,
         KEYINPUT40, KEYINPUT39, KEYINPUT38, KEYINPUT37, KEYINPUT36,
         KEYINPUT35, KEYINPUT34, KEYINPUT33, KEYINPUT32, KEYINPUT31,
         KEYINPUT30, KEYINPUT29, KEYINPUT28, KEYINPUT27, KEYINPUT26,
         KEYINPUT25, KEYINPUT24, KEYINPUT23, KEYINPUT22, KEYINPUT21,
         KEYINPUT20, KEYINPUT19, KEYINPUT18, KEYINPUT17, KEYINPUT16,
         KEYINPUT15, KEYINPUT14, KEYINPUT13, KEYINPUT12, KEYINPUT11,
         KEYINPUT10, KEYINPUT9, KEYINPUT8, KEYINPUT7, KEYINPUT6, KEYINPUT5,
         KEYINPUT4, KEYINPUT3, KEYINPUT2, KEYINPUT1, KEYINPUT0, KEYINPUT127,
         KEYINPUT126, KEYINPUT125, KEYINPUT124, KEYINPUT123, KEYINPUT122,
         KEYINPUT121, KEYINPUT120, KEYINPUT119, KEYINPUT118, KEYINPUT117,
         KEYINPUT116, KEYINPUT115, KEYINPUT114, KEYINPUT113, KEYINPUT112,
         KEYINPUT111, KEYINPUT110, KEYINPUT109, KEYINPUT108, KEYINPUT107,
         KEYINPUT106, KEYINPUT105, KEYINPUT104, KEYINPUT103, KEYINPUT102,
         KEYINPUT101, KEYINPUT100, KEYINPUT99, KEYINPUT98, KEYINPUT97,
         KEYINPUT96, KEYINPUT95, KEYINPUT94, KEYINPUT93, KEYINPUT92,
         KEYINPUT91, KEYINPUT90, KEYINPUT89, KEYINPUT88, KEYINPUT87,
         KEYINPUT86, KEYINPUT85, KEYINPUT84, KEYINPUT83, KEYINPUT82,
         KEYINPUT81, KEYINPUT80, KEYINPUT79, KEYINPUT78, KEYINPUT77,
         KEYINPUT76, KEYINPUT75, KEYINPUT74, KEYINPUT73, KEYINPUT72,
         KEYINPUT71, KEYINPUT70, KEYINPUT69, KEYINPUT68, KEYINPUT67,
         KEYINPUT66, KEYINPUT65, KEYINPUT64;
  output G1324GAT, G1325GAT, G1326GAT, G1327GAT, G1328GAT, G1329GAT, G1330GAT,
         G1331GAT, G1332GAT, G1333GAT, G1334GAT, G1335GAT, G1336GAT, G1337GAT,
         G1338GAT, G1339GAT, G1340GAT, G1341GAT, G1342GAT, G1343GAT, G1344GAT,
         G1345GAT, G1346GAT, G1347GAT, G1348GAT, G1349GAT, G1350GAT, G1351GAT,
         G1352GAT, G1353GAT, G1354GAT, G1355GAT;
  wire   n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578;

  XNOR2_X1 U321 ( .A(n376), .B(KEYINPUT46), .ZN(n377) );
  INV_X1 U322 ( .A(KEYINPUT54), .ZN(n403) );
  XNOR2_X1 U323 ( .A(n373), .B(n372), .ZN(n374) );
  XNOR2_X1 U324 ( .A(n419), .B(KEYINPUT55), .ZN(n439) );
  XNOR2_X1 U325 ( .A(n375), .B(n374), .ZN(n444) );
  INV_X1 U326 ( .A(G190GAT), .ZN(n440) );
  XNOR2_X1 U327 ( .A(n441), .B(n440), .ZN(n442) );
  XNOR2_X1 U328 ( .A(n443), .B(n442), .ZN(G1351GAT) );
  XOR2_X1 U329 ( .A(KEYINPUT9), .B(G218GAT), .Z(n290) );
  XNOR2_X1 U330 ( .A(G162GAT), .B(G106GAT), .ZN(n289) );
  XNOR2_X1 U331 ( .A(n290), .B(n289), .ZN(n293) );
  XOR2_X1 U332 ( .A(KEYINPUT72), .B(G92GAT), .Z(n292) );
  XNOR2_X1 U333 ( .A(G99GAT), .B(G85GAT), .ZN(n291) );
  XNOR2_X1 U334 ( .A(n292), .B(n291), .ZN(n364) );
  XOR2_X1 U335 ( .A(n293), .B(n364), .Z(n295) );
  XOR2_X1 U336 ( .A(G29GAT), .B(G134GAT), .Z(n308) );
  XOR2_X1 U337 ( .A(G36GAT), .B(G190GAT), .Z(n400) );
  XNOR2_X1 U338 ( .A(n308), .B(n400), .ZN(n294) );
  XNOR2_X1 U339 ( .A(n295), .B(n294), .ZN(n299) );
  XOR2_X1 U340 ( .A(KEYINPUT11), .B(KEYINPUT10), .Z(n297) );
  NAND2_X1 U341 ( .A1(G232GAT), .A2(G233GAT), .ZN(n296) );
  XNOR2_X1 U342 ( .A(n297), .B(n296), .ZN(n298) );
  XOR2_X1 U343 ( .A(n299), .B(n298), .Z(n304) );
  XOR2_X1 U344 ( .A(KEYINPUT7), .B(KEYINPUT68), .Z(n301) );
  XNOR2_X1 U345 ( .A(G50GAT), .B(G43GAT), .ZN(n300) );
  XNOR2_X1 U346 ( .A(n301), .B(n300), .ZN(n302) );
  XOR2_X1 U347 ( .A(KEYINPUT8), .B(n302), .Z(n357) );
  XNOR2_X1 U348 ( .A(n357), .B(KEYINPUT74), .ZN(n303) );
  XOR2_X1 U349 ( .A(n304), .B(n303), .Z(n533) );
  INV_X1 U350 ( .A(n533), .ZN(n549) );
  XOR2_X1 U351 ( .A(KEYINPUT88), .B(KEYINPUT89), .Z(n306) );
  XNOR2_X1 U352 ( .A(G85GAT), .B(KEYINPUT5), .ZN(n305) );
  XNOR2_X1 U353 ( .A(n306), .B(n305), .ZN(n307) );
  XOR2_X1 U354 ( .A(n307), .B(KEYINPUT90), .Z(n310) );
  XNOR2_X1 U355 ( .A(G1GAT), .B(n308), .ZN(n309) );
  XNOR2_X1 U356 ( .A(n310), .B(n309), .ZN(n320) );
  XOR2_X1 U357 ( .A(KEYINPUT1), .B(KEYINPUT6), .Z(n312) );
  NAND2_X1 U358 ( .A1(G225GAT), .A2(G233GAT), .ZN(n311) );
  XNOR2_X1 U359 ( .A(n312), .B(n311), .ZN(n313) );
  XOR2_X1 U360 ( .A(n313), .B(KEYINPUT4), .Z(n318) );
  XOR2_X1 U361 ( .A(G127GAT), .B(KEYINPUT80), .Z(n315) );
  XNOR2_X1 U362 ( .A(G113GAT), .B(KEYINPUT0), .ZN(n314) );
  XNOR2_X1 U363 ( .A(n315), .B(n314), .ZN(n436) );
  XNOR2_X1 U364 ( .A(G120GAT), .B(G148GAT), .ZN(n316) );
  XNOR2_X1 U365 ( .A(n316), .B(G57GAT), .ZN(n369) );
  XNOR2_X1 U366 ( .A(n436), .B(n369), .ZN(n317) );
  XNOR2_X1 U367 ( .A(n318), .B(n317), .ZN(n319) );
  XNOR2_X1 U368 ( .A(n320), .B(n319), .ZN(n325) );
  XOR2_X1 U369 ( .A(KEYINPUT3), .B(KEYINPUT86), .Z(n322) );
  XNOR2_X1 U370 ( .A(G141GAT), .B(G155GAT), .ZN(n321) );
  XNOR2_X1 U371 ( .A(n322), .B(n321), .ZN(n324) );
  XOR2_X1 U372 ( .A(G162GAT), .B(KEYINPUT2), .Z(n323) );
  XNOR2_X1 U373 ( .A(n324), .B(n323), .ZN(n417) );
  XNOR2_X1 U374 ( .A(n325), .B(n417), .ZN(n456) );
  XNOR2_X1 U375 ( .A(KEYINPUT91), .B(n456), .ZN(n505) );
  XOR2_X1 U376 ( .A(G57GAT), .B(G211GAT), .Z(n327) );
  XNOR2_X1 U377 ( .A(G155GAT), .B(G78GAT), .ZN(n326) );
  XNOR2_X1 U378 ( .A(n327), .B(n326), .ZN(n328) );
  XOR2_X1 U379 ( .A(G71GAT), .B(KEYINPUT13), .Z(n367) );
  XOR2_X1 U380 ( .A(n328), .B(n367), .Z(n330) );
  XNOR2_X1 U381 ( .A(G127GAT), .B(G183GAT), .ZN(n329) );
  XNOR2_X1 U382 ( .A(n330), .B(n329), .ZN(n335) );
  XNOR2_X1 U383 ( .A(G15GAT), .B(G22GAT), .ZN(n331) );
  XNOR2_X1 U384 ( .A(n331), .B(G1GAT), .ZN(n349) );
  XOR2_X1 U385 ( .A(n349), .B(KEYINPUT12), .Z(n333) );
  NAND2_X1 U386 ( .A1(G231GAT), .A2(G233GAT), .ZN(n332) );
  XNOR2_X1 U387 ( .A(n333), .B(n332), .ZN(n334) );
  XOR2_X1 U388 ( .A(n335), .B(n334), .Z(n343) );
  XOR2_X1 U389 ( .A(KEYINPUT78), .B(KEYINPUT75), .Z(n337) );
  XNOR2_X1 U390 ( .A(G8GAT), .B(G64GAT), .ZN(n336) );
  XNOR2_X1 U391 ( .A(n337), .B(n336), .ZN(n341) );
  XOR2_X1 U392 ( .A(KEYINPUT77), .B(KEYINPUT76), .Z(n339) );
  XNOR2_X1 U393 ( .A(KEYINPUT15), .B(KEYINPUT14), .ZN(n338) );
  XNOR2_X1 U394 ( .A(n339), .B(n338), .ZN(n340) );
  XNOR2_X1 U395 ( .A(n341), .B(n340), .ZN(n342) );
  XOR2_X1 U396 ( .A(n343), .B(n342), .Z(n572) );
  INV_X1 U397 ( .A(n572), .ZN(n526) );
  XOR2_X1 U398 ( .A(KEYINPUT66), .B(G197GAT), .Z(n345) );
  XNOR2_X1 U399 ( .A(G113GAT), .B(G141GAT), .ZN(n344) );
  XNOR2_X1 U400 ( .A(n345), .B(n344), .ZN(n346) );
  XOR2_X1 U401 ( .A(n346), .B(G36GAT), .Z(n348) );
  XOR2_X1 U402 ( .A(G169GAT), .B(G8GAT), .Z(n396) );
  XNOR2_X1 U403 ( .A(n396), .B(G29GAT), .ZN(n347) );
  XNOR2_X1 U404 ( .A(n348), .B(n347), .ZN(n353) );
  XOR2_X1 U405 ( .A(n349), .B(KEYINPUT64), .Z(n351) );
  NAND2_X1 U406 ( .A1(G229GAT), .A2(G233GAT), .ZN(n350) );
  XNOR2_X1 U407 ( .A(n351), .B(n350), .ZN(n352) );
  XOR2_X1 U408 ( .A(n353), .B(n352), .Z(n359) );
  XOR2_X1 U409 ( .A(KEYINPUT30), .B(KEYINPUT67), .Z(n355) );
  XNOR2_X1 U410 ( .A(KEYINPUT29), .B(KEYINPUT65), .ZN(n354) );
  XNOR2_X1 U411 ( .A(n355), .B(n354), .ZN(n356) );
  XNOR2_X1 U412 ( .A(n357), .B(n356), .ZN(n358) );
  XOR2_X1 U413 ( .A(n359), .B(n358), .Z(n522) );
  XOR2_X1 U414 ( .A(KEYINPUT32), .B(KEYINPUT69), .Z(n361) );
  NAND2_X1 U415 ( .A1(G230GAT), .A2(G233GAT), .ZN(n360) );
  XNOR2_X1 U416 ( .A(n361), .B(n360), .ZN(n362) );
  XOR2_X1 U417 ( .A(n362), .B(KEYINPUT73), .Z(n366) );
  XNOR2_X1 U418 ( .A(G106GAT), .B(G78GAT), .ZN(n363) );
  XNOR2_X1 U419 ( .A(n363), .B(G204GAT), .ZN(n412) );
  XNOR2_X1 U420 ( .A(n364), .B(n412), .ZN(n365) );
  XNOR2_X1 U421 ( .A(n366), .B(n365), .ZN(n368) );
  XOR2_X1 U422 ( .A(n368), .B(n367), .Z(n375) );
  XOR2_X1 U423 ( .A(G176GAT), .B(G64GAT), .Z(n401) );
  XNOR2_X1 U424 ( .A(n369), .B(n401), .ZN(n373) );
  XOR2_X1 U425 ( .A(KEYINPUT31), .B(KEYINPUT71), .Z(n371) );
  XNOR2_X1 U426 ( .A(KEYINPUT33), .B(KEYINPUT70), .ZN(n370) );
  XNOR2_X1 U427 ( .A(n371), .B(n370), .ZN(n372) );
  XOR2_X1 U428 ( .A(n444), .B(KEYINPUT41), .Z(n543) );
  NAND2_X1 U429 ( .A1(n522), .A2(n543), .ZN(n376) );
  NAND2_X1 U430 ( .A1(n377), .A2(n549), .ZN(n378) );
  NOR2_X1 U431 ( .A1(n526), .A2(n378), .ZN(n379) );
  XNOR2_X1 U432 ( .A(n379), .B(KEYINPUT47), .ZN(n384) );
  XOR2_X1 U433 ( .A(KEYINPUT36), .B(n533), .Z(n575) );
  NOR2_X1 U434 ( .A1(n575), .A2(n572), .ZN(n380) );
  XOR2_X1 U435 ( .A(KEYINPUT45), .B(n380), .Z(n381) );
  NOR2_X1 U436 ( .A1(n444), .A2(n381), .ZN(n382) );
  INV_X1 U437 ( .A(n522), .ZN(n565) );
  NAND2_X1 U438 ( .A1(n382), .A2(n565), .ZN(n383) );
  NAND2_X1 U439 ( .A1(n384), .A2(n383), .ZN(n385) );
  XOR2_X1 U440 ( .A(KEYINPUT48), .B(n385), .Z(n537) );
  XOR2_X1 U441 ( .A(KEYINPUT75), .B(KEYINPUT92), .Z(n387) );
  NAND2_X1 U442 ( .A1(G226GAT), .A2(G233GAT), .ZN(n386) );
  XNOR2_X1 U443 ( .A(n387), .B(n386), .ZN(n388) );
  XOR2_X1 U444 ( .A(n388), .B(KEYINPUT93), .Z(n394) );
  XOR2_X1 U445 ( .A(G183GAT), .B(KEYINPUT18), .Z(n390) );
  XNOR2_X1 U446 ( .A(KEYINPUT19), .B(KEYINPUT17), .ZN(n389) );
  XNOR2_X1 U447 ( .A(n390), .B(n389), .ZN(n435) );
  XOR2_X1 U448 ( .A(G211GAT), .B(KEYINPUT21), .Z(n392) );
  XNOR2_X1 U449 ( .A(G197GAT), .B(G218GAT), .ZN(n391) );
  XNOR2_X1 U450 ( .A(n392), .B(n391), .ZN(n410) );
  XNOR2_X1 U451 ( .A(n435), .B(n410), .ZN(n393) );
  XNOR2_X1 U452 ( .A(n394), .B(n393), .ZN(n395) );
  XOR2_X1 U453 ( .A(n395), .B(G92GAT), .Z(n398) );
  XNOR2_X1 U454 ( .A(n396), .B(G204GAT), .ZN(n397) );
  XNOR2_X1 U455 ( .A(n398), .B(n397), .ZN(n399) );
  XNOR2_X1 U456 ( .A(n400), .B(n399), .ZN(n402) );
  XOR2_X1 U457 ( .A(n402), .B(n401), .Z(n447) );
  NOR2_X1 U458 ( .A1(n537), .A2(n447), .ZN(n404) );
  XNOR2_X1 U459 ( .A(n404), .B(n403), .ZN(n405) );
  NOR2_X1 U460 ( .A1(n505), .A2(n405), .ZN(n563) );
  XOR2_X1 U461 ( .A(KEYINPUT22), .B(KEYINPUT23), .Z(n407) );
  XNOR2_X1 U462 ( .A(G50GAT), .B(KEYINPUT24), .ZN(n406) );
  XNOR2_X1 U463 ( .A(n407), .B(n406), .ZN(n416) );
  XOR2_X1 U464 ( .A(KEYINPUT87), .B(G148GAT), .Z(n409) );
  NAND2_X1 U465 ( .A1(G228GAT), .A2(G233GAT), .ZN(n408) );
  XNOR2_X1 U466 ( .A(n409), .B(n408), .ZN(n411) );
  XOR2_X1 U467 ( .A(n411), .B(n410), .Z(n414) );
  XNOR2_X1 U468 ( .A(G22GAT), .B(n412), .ZN(n413) );
  XNOR2_X1 U469 ( .A(n414), .B(n413), .ZN(n415) );
  XNOR2_X1 U470 ( .A(n416), .B(n415), .ZN(n418) );
  XNOR2_X1 U471 ( .A(n418), .B(n417), .ZN(n459) );
  NAND2_X1 U472 ( .A1(n563), .A2(n459), .ZN(n419) );
  XOR2_X1 U473 ( .A(G99GAT), .B(G190GAT), .Z(n421) );
  XNOR2_X1 U474 ( .A(G43GAT), .B(G134GAT), .ZN(n420) );
  XNOR2_X1 U475 ( .A(n421), .B(n420), .ZN(n425) );
  XOR2_X1 U476 ( .A(KEYINPUT84), .B(G120GAT), .Z(n423) );
  XNOR2_X1 U477 ( .A(G169GAT), .B(G15GAT), .ZN(n422) );
  XNOR2_X1 U478 ( .A(n423), .B(n422), .ZN(n424) );
  XOR2_X1 U479 ( .A(n425), .B(n424), .Z(n430) );
  XOR2_X1 U480 ( .A(KEYINPUT20), .B(G176GAT), .Z(n427) );
  NAND2_X1 U481 ( .A1(G227GAT), .A2(G233GAT), .ZN(n426) );
  XNOR2_X1 U482 ( .A(n427), .B(n426), .ZN(n428) );
  XNOR2_X1 U483 ( .A(KEYINPUT82), .B(n428), .ZN(n429) );
  XNOR2_X1 U484 ( .A(n430), .B(n429), .ZN(n434) );
  XOR2_X1 U485 ( .A(KEYINPUT81), .B(G71GAT), .Z(n432) );
  XNOR2_X1 U486 ( .A(KEYINPUT83), .B(KEYINPUT85), .ZN(n431) );
  XNOR2_X1 U487 ( .A(n432), .B(n431), .ZN(n433) );
  XOR2_X1 U488 ( .A(n434), .B(n433), .Z(n438) );
  XNOR2_X1 U489 ( .A(n436), .B(n435), .ZN(n437) );
  XOR2_X1 U490 ( .A(n438), .B(n437), .Z(n460) );
  INV_X1 U491 ( .A(n460), .ZN(n520) );
  NAND2_X1 U492 ( .A1(n439), .A2(n520), .ZN(n558) );
  NOR2_X1 U493 ( .A1(n549), .A2(n558), .ZN(n443) );
  XNOR2_X1 U494 ( .A(KEYINPUT124), .B(KEYINPUT58), .ZN(n441) );
  INV_X1 U495 ( .A(n444), .ZN(n569) );
  NAND2_X1 U496 ( .A1(n569), .A2(n522), .ZN(n480) );
  NAND2_X1 U497 ( .A1(n526), .A2(n549), .ZN(n445) );
  XNOR2_X1 U498 ( .A(n445), .B(KEYINPUT79), .ZN(n446) );
  XNOR2_X1 U499 ( .A(n446), .B(KEYINPUT16), .ZN(n463) );
  INV_X1 U500 ( .A(n447), .ZN(n509) );
  NAND2_X1 U501 ( .A1(n509), .A2(n520), .ZN(n448) );
  NAND2_X1 U502 ( .A1(n448), .A2(n459), .ZN(n449) );
  XNOR2_X1 U503 ( .A(n449), .B(KEYINPUT96), .ZN(n450) );
  XNOR2_X1 U504 ( .A(KEYINPUT25), .B(n450), .ZN(n451) );
  XNOR2_X1 U505 ( .A(n451), .B(KEYINPUT95), .ZN(n455) );
  NOR2_X1 U506 ( .A1(n520), .A2(n459), .ZN(n453) );
  XNOR2_X1 U507 ( .A(KEYINPUT26), .B(KEYINPUT94), .ZN(n452) );
  XNOR2_X1 U508 ( .A(n453), .B(n452), .ZN(n562) );
  XNOR2_X1 U509 ( .A(KEYINPUT27), .B(n509), .ZN(n458) );
  NAND2_X1 U510 ( .A1(n562), .A2(n458), .ZN(n454) );
  NAND2_X1 U511 ( .A1(n455), .A2(n454), .ZN(n457) );
  NAND2_X1 U512 ( .A1(n457), .A2(n456), .ZN(n462) );
  NAND2_X1 U513 ( .A1(n505), .A2(n458), .ZN(n536) );
  XOR2_X1 U514 ( .A(KEYINPUT28), .B(n459), .Z(n514) );
  NOR2_X1 U515 ( .A1(n536), .A2(n514), .ZN(n519) );
  NAND2_X1 U516 ( .A1(n519), .A2(n460), .ZN(n461) );
  NAND2_X1 U517 ( .A1(n462), .A2(n461), .ZN(n477) );
  NAND2_X1 U518 ( .A1(n463), .A2(n477), .ZN(n492) );
  NOR2_X1 U519 ( .A1(n480), .A2(n492), .ZN(n464) );
  XOR2_X1 U520 ( .A(KEYINPUT97), .B(n464), .Z(n474) );
  NAND2_X1 U521 ( .A1(n474), .A2(n505), .ZN(n468) );
  XOR2_X1 U522 ( .A(KEYINPUT99), .B(KEYINPUT34), .Z(n466) );
  XNOR2_X1 U523 ( .A(G1GAT), .B(KEYINPUT98), .ZN(n465) );
  XNOR2_X1 U524 ( .A(n466), .B(n465), .ZN(n467) );
  XNOR2_X1 U525 ( .A(n468), .B(n467), .ZN(G1324GAT) );
  XOR2_X1 U526 ( .A(KEYINPUT100), .B(KEYINPUT101), .Z(n470) );
  NAND2_X1 U527 ( .A1(n474), .A2(n509), .ZN(n469) );
  XNOR2_X1 U528 ( .A(n470), .B(n469), .ZN(n471) );
  XNOR2_X1 U529 ( .A(G8GAT), .B(n471), .ZN(G1325GAT) );
  XOR2_X1 U530 ( .A(G15GAT), .B(KEYINPUT35), .Z(n473) );
  NAND2_X1 U531 ( .A1(n474), .A2(n520), .ZN(n472) );
  XNOR2_X1 U532 ( .A(n473), .B(n472), .ZN(G1326GAT) );
  NAND2_X1 U533 ( .A1(n514), .A2(n474), .ZN(n475) );
  XNOR2_X1 U534 ( .A(n475), .B(KEYINPUT102), .ZN(n476) );
  XNOR2_X1 U535 ( .A(G22GAT), .B(n476), .ZN(G1327GAT) );
  XOR2_X1 U536 ( .A(KEYINPUT39), .B(KEYINPUT103), .Z(n483) );
  NAND2_X1 U537 ( .A1(n572), .A2(n477), .ZN(n478) );
  NOR2_X1 U538 ( .A1(n575), .A2(n478), .ZN(n479) );
  XNOR2_X1 U539 ( .A(KEYINPUT37), .B(n479), .ZN(n504) );
  NOR2_X1 U540 ( .A1(n504), .A2(n480), .ZN(n481) );
  XNOR2_X1 U541 ( .A(KEYINPUT38), .B(n481), .ZN(n490) );
  NAND2_X1 U542 ( .A1(n505), .A2(n490), .ZN(n482) );
  XNOR2_X1 U543 ( .A(n483), .B(n482), .ZN(n484) );
  XOR2_X1 U544 ( .A(G29GAT), .B(n484), .Z(G1328GAT) );
  NAND2_X1 U545 ( .A1(n490), .A2(n509), .ZN(n485) );
  XNOR2_X1 U546 ( .A(n485), .B(KEYINPUT104), .ZN(n486) );
  XNOR2_X1 U547 ( .A(G36GAT), .B(n486), .ZN(G1329GAT) );
  XOR2_X1 U548 ( .A(KEYINPUT105), .B(KEYINPUT40), .Z(n488) );
  NAND2_X1 U549 ( .A1(n520), .A2(n490), .ZN(n487) );
  XNOR2_X1 U550 ( .A(n488), .B(n487), .ZN(n489) );
  XNOR2_X1 U551 ( .A(G43GAT), .B(n489), .ZN(G1330GAT) );
  NAND2_X1 U552 ( .A1(n490), .A2(n514), .ZN(n491) );
  XNOR2_X1 U553 ( .A(n491), .B(G50GAT), .ZN(G1331GAT) );
  XNOR2_X1 U554 ( .A(G57GAT), .B(KEYINPUT42), .ZN(n495) );
  NAND2_X1 U555 ( .A1(n565), .A2(n543), .ZN(n503) );
  NOR2_X1 U556 ( .A1(n503), .A2(n492), .ZN(n493) );
  XNOR2_X1 U557 ( .A(n493), .B(KEYINPUT106), .ZN(n499) );
  NAND2_X1 U558 ( .A1(n505), .A2(n499), .ZN(n494) );
  XNOR2_X1 U559 ( .A(n495), .B(n494), .ZN(G1332GAT) );
  XOR2_X1 U560 ( .A(G64GAT), .B(KEYINPUT107), .Z(n497) );
  NAND2_X1 U561 ( .A1(n509), .A2(n499), .ZN(n496) );
  XNOR2_X1 U562 ( .A(n497), .B(n496), .ZN(G1333GAT) );
  NAND2_X1 U563 ( .A1(n499), .A2(n520), .ZN(n498) );
  XNOR2_X1 U564 ( .A(n498), .B(G71GAT), .ZN(G1334GAT) );
  XOR2_X1 U565 ( .A(KEYINPUT43), .B(KEYINPUT108), .Z(n501) );
  NAND2_X1 U566 ( .A1(n499), .A2(n514), .ZN(n500) );
  XNOR2_X1 U567 ( .A(n501), .B(n500), .ZN(n502) );
  XNOR2_X1 U568 ( .A(G78GAT), .B(n502), .ZN(G1335GAT) );
  XOR2_X1 U569 ( .A(KEYINPUT109), .B(KEYINPUT110), .Z(n507) );
  NOR2_X1 U570 ( .A1(n504), .A2(n503), .ZN(n515) );
  NAND2_X1 U571 ( .A1(n515), .A2(n505), .ZN(n506) );
  XNOR2_X1 U572 ( .A(n507), .B(n506), .ZN(n508) );
  XNOR2_X1 U573 ( .A(G85GAT), .B(n508), .ZN(G1336GAT) );
  XOR2_X1 U574 ( .A(G92GAT), .B(KEYINPUT111), .Z(n511) );
  NAND2_X1 U575 ( .A1(n515), .A2(n509), .ZN(n510) );
  XNOR2_X1 U576 ( .A(n511), .B(n510), .ZN(G1337GAT) );
  NAND2_X1 U577 ( .A1(n515), .A2(n520), .ZN(n512) );
  XNOR2_X1 U578 ( .A(n512), .B(KEYINPUT112), .ZN(n513) );
  XNOR2_X1 U579 ( .A(G99GAT), .B(n513), .ZN(G1338GAT) );
  XOR2_X1 U580 ( .A(KEYINPUT113), .B(KEYINPUT44), .Z(n517) );
  NAND2_X1 U581 ( .A1(n515), .A2(n514), .ZN(n516) );
  XNOR2_X1 U582 ( .A(n517), .B(n516), .ZN(n518) );
  XNOR2_X1 U583 ( .A(G106GAT), .B(n518), .ZN(G1339GAT) );
  NAND2_X1 U584 ( .A1(n520), .A2(n519), .ZN(n521) );
  NOR2_X1 U585 ( .A1(n537), .A2(n521), .ZN(n532) );
  NAND2_X1 U586 ( .A1(n522), .A2(n532), .ZN(n523) );
  XNOR2_X1 U587 ( .A(n523), .B(G113GAT), .ZN(G1340GAT) );
  XOR2_X1 U588 ( .A(G120GAT), .B(KEYINPUT49), .Z(n525) );
  NAND2_X1 U589 ( .A1(n532), .A2(n543), .ZN(n524) );
  XNOR2_X1 U590 ( .A(n525), .B(n524), .ZN(G1341GAT) );
  XOR2_X1 U591 ( .A(KEYINPUT50), .B(KEYINPUT114), .Z(n528) );
  NAND2_X1 U592 ( .A1(n532), .A2(n526), .ZN(n527) );
  XNOR2_X1 U593 ( .A(n528), .B(n527), .ZN(n529) );
  XOR2_X1 U594 ( .A(G127GAT), .B(n529), .Z(G1342GAT) );
  XOR2_X1 U595 ( .A(KEYINPUT115), .B(KEYINPUT51), .Z(n531) );
  XNOR2_X1 U596 ( .A(G134GAT), .B(KEYINPUT116), .ZN(n530) );
  XNOR2_X1 U597 ( .A(n531), .B(n530), .ZN(n535) );
  NAND2_X1 U598 ( .A1(n533), .A2(n532), .ZN(n534) );
  XOR2_X1 U599 ( .A(n535), .B(n534), .Z(G1343GAT) );
  NOR2_X1 U600 ( .A1(n537), .A2(n536), .ZN(n538) );
  NAND2_X1 U601 ( .A1(n562), .A2(n538), .ZN(n548) );
  NOR2_X1 U602 ( .A1(n565), .A2(n548), .ZN(n540) );
  XNOR2_X1 U603 ( .A(G141GAT), .B(KEYINPUT117), .ZN(n539) );
  XNOR2_X1 U604 ( .A(n540), .B(n539), .ZN(G1344GAT) );
  XOR2_X1 U605 ( .A(KEYINPUT53), .B(KEYINPUT52), .Z(n542) );
  XNOR2_X1 U606 ( .A(G148GAT), .B(KEYINPUT118), .ZN(n541) );
  XNOR2_X1 U607 ( .A(n542), .B(n541), .ZN(n545) );
  INV_X1 U608 ( .A(n543), .ZN(n553) );
  NOR2_X1 U609 ( .A1(n553), .A2(n548), .ZN(n544) );
  XOR2_X1 U610 ( .A(n545), .B(n544), .Z(G1345GAT) );
  NOR2_X1 U611 ( .A1(n572), .A2(n548), .ZN(n547) );
  XNOR2_X1 U612 ( .A(G155GAT), .B(KEYINPUT119), .ZN(n546) );
  XNOR2_X1 U613 ( .A(n547), .B(n546), .ZN(G1346GAT) );
  NOR2_X1 U614 ( .A1(n549), .A2(n548), .ZN(n550) );
  XOR2_X1 U615 ( .A(KEYINPUT120), .B(n550), .Z(n551) );
  XNOR2_X1 U616 ( .A(G162GAT), .B(n551), .ZN(G1347GAT) );
  NOR2_X1 U617 ( .A1(n565), .A2(n558), .ZN(n552) );
  XOR2_X1 U618 ( .A(G169GAT), .B(n552), .Z(G1348GAT) );
  NOR2_X1 U619 ( .A1(n558), .A2(n553), .ZN(n557) );
  XOR2_X1 U620 ( .A(KEYINPUT56), .B(KEYINPUT121), .Z(n555) );
  XNOR2_X1 U621 ( .A(G176GAT), .B(KEYINPUT57), .ZN(n554) );
  XNOR2_X1 U622 ( .A(n555), .B(n554), .ZN(n556) );
  XNOR2_X1 U623 ( .A(n557), .B(n556), .ZN(G1349GAT) );
  NOR2_X1 U624 ( .A1(n572), .A2(n558), .ZN(n560) );
  XNOR2_X1 U625 ( .A(KEYINPUT122), .B(KEYINPUT123), .ZN(n559) );
  XNOR2_X1 U626 ( .A(n560), .B(n559), .ZN(n561) );
  XNOR2_X1 U627 ( .A(G183GAT), .B(n561), .ZN(G1350GAT) );
  NAND2_X1 U628 ( .A1(n563), .A2(n562), .ZN(n564) );
  XOR2_X1 U629 ( .A(KEYINPUT125), .B(n564), .Z(n574) );
  NOR2_X1 U630 ( .A1(n565), .A2(n574), .ZN(n567) );
  XNOR2_X1 U631 ( .A(KEYINPUT60), .B(KEYINPUT59), .ZN(n566) );
  XNOR2_X1 U632 ( .A(n567), .B(n566), .ZN(n568) );
  XNOR2_X1 U633 ( .A(G197GAT), .B(n568), .ZN(G1352GAT) );
  NOR2_X1 U634 ( .A1(n569), .A2(n574), .ZN(n571) );
  XNOR2_X1 U635 ( .A(G204GAT), .B(KEYINPUT61), .ZN(n570) );
  XNOR2_X1 U636 ( .A(n571), .B(n570), .ZN(G1353GAT) );
  NOR2_X1 U637 ( .A1(n572), .A2(n574), .ZN(n573) );
  XOR2_X1 U638 ( .A(G211GAT), .B(n573), .Z(G1354GAT) );
  NOR2_X1 U639 ( .A1(n575), .A2(n574), .ZN(n577) );
  XNOR2_X1 U640 ( .A(KEYINPUT62), .B(KEYINPUT126), .ZN(n576) );
  XNOR2_X1 U641 ( .A(n577), .B(n576), .ZN(n578) );
  XOR2_X1 U642 ( .A(G218GAT), .B(n578), .Z(G1355GAT) );
endmodule

