//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 0 1 1 0 1 0 1 1 0 0 1 1 0 0 0 1 1 0 1 1 1 0 1 1 1 0 1 0 1 1 0 1 1 1 0 0 1 1 1 0 1 1 1 1 1 0 0 1 1 0 0 0 0 0 1 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:25:36 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n599,
    new_n600, new_n601, new_n602, new_n603, new_n604, new_n605, new_n606,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n633, new_n634, new_n635, new_n636,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n650, new_n651,
    new_n652, new_n653, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n664, new_n665, new_n666,
    new_n667, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n700, new_n701, new_n702, new_n703,
    new_n704, new_n705, new_n706, new_n707, new_n708, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n725, new_n726, new_n727,
    new_n728, new_n729, new_n731, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n742,
    new_n743, new_n745, new_n746, new_n747, new_n748, new_n749, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n759,
    new_n760, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n778, new_n779, new_n780, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n790, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n914, new_n915, new_n916, new_n917,
    new_n918, new_n919, new_n920, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n934, new_n935, new_n936, new_n937, new_n938, new_n939, new_n941,
    new_n942, new_n943, new_n944, new_n945, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n954, new_n955, new_n956,
    new_n957, new_n958, new_n959, new_n960, new_n961, new_n962, new_n963,
    new_n964, new_n966, new_n967, new_n968, new_n969, new_n970, new_n971,
    new_n972, new_n973, new_n975, new_n976, new_n977, new_n978, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n986,
    new_n987, new_n988, new_n989, new_n990, new_n991, new_n992, new_n993,
    new_n994, new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006;
  INV_X1    g000(.A(G128), .ZN(new_n187));
  INV_X1    g001(.A(G146), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G143), .ZN(new_n189));
  AOI21_X1  g003(.A(new_n187), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n190));
  XNOR2_X1  g004(.A(G143), .B(G146), .ZN(new_n191));
  XNOR2_X1  g005(.A(new_n190), .B(new_n191), .ZN(new_n192));
  XNOR2_X1  g006(.A(KEYINPUT70), .B(G125), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G143), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n195), .A2(G146), .ZN(new_n196));
  NAND4_X1  g010(.A1(new_n189), .A2(new_n196), .A3(KEYINPUT0), .A4(G128), .ZN(new_n197));
  XNOR2_X1  g011(.A(KEYINPUT0), .B(G128), .ZN(new_n198));
  OAI21_X1  g012(.A(new_n197), .B1(new_n191), .B2(new_n198), .ZN(new_n199));
  INV_X1    g013(.A(new_n199), .ZN(new_n200));
  INV_X1    g014(.A(G125), .ZN(new_n201));
  NAND2_X1  g015(.A1(new_n201), .A2(KEYINPUT70), .ZN(new_n202));
  INV_X1    g016(.A(KEYINPUT70), .ZN(new_n203));
  NAND2_X1  g017(.A1(new_n203), .A2(G125), .ZN(new_n204));
  NAND2_X1  g018(.A1(new_n202), .A2(new_n204), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n200), .A2(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n194), .A2(new_n206), .ZN(new_n207));
  INV_X1    g021(.A(G953), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n208), .A2(G224), .ZN(new_n209));
  XNOR2_X1  g023(.A(new_n209), .B(KEYINPUT82), .ZN(new_n210));
  XNOR2_X1  g024(.A(new_n207), .B(new_n210), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT73), .ZN(new_n212));
  INV_X1    g026(.A(G104), .ZN(new_n213));
  OAI21_X1  g027(.A(KEYINPUT3), .B1(new_n213), .B2(G107), .ZN(new_n214));
  INV_X1    g028(.A(KEYINPUT3), .ZN(new_n215));
  INV_X1    g029(.A(G107), .ZN(new_n216));
  NAND3_X1  g030(.A1(new_n215), .A2(new_n216), .A3(G104), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n213), .A2(G107), .ZN(new_n218));
  NAND3_X1  g032(.A1(new_n214), .A2(new_n217), .A3(new_n218), .ZN(new_n219));
  AND2_X1   g033(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n220));
  INV_X1    g034(.A(KEYINPUT72), .ZN(new_n221));
  NAND4_X1  g035(.A1(new_n214), .A2(new_n217), .A3(new_n221), .A4(new_n218), .ZN(new_n222));
  NAND2_X1  g036(.A1(new_n222), .A2(G101), .ZN(new_n223));
  OAI21_X1  g037(.A(new_n212), .B1(new_n220), .B2(new_n223), .ZN(new_n224));
  NAND2_X1  g038(.A1(new_n219), .A2(KEYINPUT72), .ZN(new_n225));
  NAND4_X1  g039(.A1(new_n225), .A2(KEYINPUT73), .A3(G101), .A4(new_n222), .ZN(new_n226));
  INV_X1    g040(.A(KEYINPUT4), .ZN(new_n227));
  AOI21_X1  g041(.A(G101), .B1(new_n213), .B2(G107), .ZN(new_n228));
  NAND3_X1  g042(.A1(new_n214), .A2(new_n228), .A3(new_n217), .ZN(new_n229));
  NAND2_X1  g043(.A1(new_n229), .A2(KEYINPUT74), .ZN(new_n230));
  INV_X1    g044(.A(KEYINPUT74), .ZN(new_n231));
  NAND4_X1  g045(.A1(new_n214), .A2(new_n228), .A3(new_n217), .A4(new_n231), .ZN(new_n232));
  AOI21_X1  g046(.A(new_n227), .B1(new_n230), .B2(new_n232), .ZN(new_n233));
  NAND3_X1  g047(.A1(new_n224), .A2(new_n226), .A3(new_n233), .ZN(new_n234));
  INV_X1    g048(.A(G116), .ZN(new_n235));
  OAI21_X1  g049(.A(KEYINPUT65), .B1(new_n235), .B2(G119), .ZN(new_n236));
  INV_X1    g050(.A(KEYINPUT65), .ZN(new_n237));
  INV_X1    g051(.A(G119), .ZN(new_n238));
  NAND3_X1  g052(.A1(new_n237), .A2(new_n238), .A3(G116), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n235), .A2(G119), .ZN(new_n240));
  AND3_X1   g054(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT2), .B(G113), .ZN(new_n242));
  INV_X1    g056(.A(new_n242), .ZN(new_n243));
  NAND2_X1  g057(.A1(new_n241), .A2(new_n243), .ZN(new_n244));
  NAND3_X1  g058(.A1(new_n236), .A2(new_n239), .A3(new_n240), .ZN(new_n245));
  NAND2_X1  g059(.A1(new_n245), .A2(new_n242), .ZN(new_n246));
  NAND2_X1  g060(.A1(new_n244), .A2(new_n246), .ZN(new_n247));
  NAND4_X1  g061(.A1(new_n225), .A2(new_n227), .A3(G101), .A4(new_n222), .ZN(new_n248));
  AND2_X1   g062(.A1(new_n247), .A2(new_n248), .ZN(new_n249));
  NAND2_X1  g063(.A1(new_n234), .A2(new_n249), .ZN(new_n250));
  NAND2_X1  g064(.A1(new_n241), .A2(KEYINPUT5), .ZN(new_n251));
  NOR3_X1   g065(.A1(new_n235), .A2(KEYINPUT5), .A3(G119), .ZN(new_n252));
  INV_X1    g066(.A(G113), .ZN(new_n253));
  NOR2_X1   g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  AOI22_X1  g068(.A1(new_n251), .A2(new_n254), .B1(new_n243), .B2(new_n241), .ZN(new_n255));
  INV_X1    g069(.A(KEYINPUT75), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n230), .A2(new_n232), .ZN(new_n257));
  INV_X1    g071(.A(G101), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n216), .A2(G104), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n258), .B1(new_n218), .B2(new_n259), .ZN(new_n260));
  INV_X1    g074(.A(new_n260), .ZN(new_n261));
  AOI21_X1  g075(.A(new_n256), .B1(new_n257), .B2(new_n261), .ZN(new_n262));
  AOI211_X1 g076(.A(KEYINPUT75), .B(new_n260), .C1(new_n230), .C2(new_n232), .ZN(new_n263));
  OAI21_X1  g077(.A(new_n255), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  NAND2_X1  g078(.A1(new_n250), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n265), .A2(KEYINPUT80), .ZN(new_n266));
  INV_X1    g080(.A(KEYINPUT80), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n250), .A2(new_n264), .A3(new_n267), .ZN(new_n268));
  XNOR2_X1  g082(.A(G110), .B(G122), .ZN(new_n269));
  INV_X1    g083(.A(new_n269), .ZN(new_n270));
  XNOR2_X1  g084(.A(KEYINPUT81), .B(KEYINPUT6), .ZN(new_n271));
  NAND4_X1  g085(.A1(new_n266), .A2(new_n268), .A3(new_n270), .A4(new_n271), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n250), .A2(new_n264), .A3(new_n267), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n267), .B1(new_n250), .B2(new_n264), .ZN(new_n274));
  NOR3_X1   g088(.A1(new_n273), .A2(new_n274), .A3(new_n269), .ZN(new_n275));
  NAND3_X1  g089(.A1(new_n250), .A2(new_n264), .A3(new_n269), .ZN(new_n276));
  NAND2_X1  g090(.A1(new_n276), .A2(KEYINPUT6), .ZN(new_n277));
  OAI211_X1 g091(.A(new_n211), .B(new_n272), .C1(new_n275), .C2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT85), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n210), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n194), .A2(new_n206), .A3(new_n280), .ZN(new_n281));
  AND2_X1   g095(.A1(new_n210), .A2(KEYINPUT7), .ZN(new_n282));
  XNOR2_X1  g096(.A(new_n281), .B(new_n282), .ZN(new_n283));
  XOR2_X1   g097(.A(new_n254), .B(KEYINPUT84), .Z(new_n284));
  INV_X1    g098(.A(KEYINPUT83), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n251), .A2(new_n285), .ZN(new_n286));
  NAND2_X1  g100(.A1(new_n284), .A2(new_n286), .ZN(new_n287));
  NOR2_X1   g101(.A1(new_n251), .A2(new_n285), .ZN(new_n288));
  OAI21_X1  g102(.A(new_n244), .B1(new_n287), .B2(new_n288), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n262), .A2(new_n263), .ZN(new_n290));
  AOI21_X1  g104(.A(new_n260), .B1(new_n230), .B2(new_n232), .ZN(new_n291));
  OAI22_X1  g105(.A1(new_n289), .A2(new_n290), .B1(new_n291), .B2(new_n255), .ZN(new_n292));
  XNOR2_X1  g106(.A(new_n269), .B(KEYINPUT8), .ZN(new_n293));
  AOI21_X1  g107(.A(new_n283), .B1(new_n292), .B2(new_n293), .ZN(new_n294));
  AOI21_X1  g108(.A(G902), .B1(new_n294), .B2(new_n276), .ZN(new_n295));
  OAI21_X1  g109(.A(G210), .B1(G237), .B2(G902), .ZN(new_n296));
  AND3_X1   g110(.A1(new_n278), .A2(new_n295), .A3(new_n296), .ZN(new_n297));
  AOI21_X1  g111(.A(new_n296), .B1(new_n278), .B2(new_n295), .ZN(new_n298));
  NOR2_X1   g112(.A1(new_n297), .A2(new_n298), .ZN(new_n299));
  INV_X1    g113(.A(new_n299), .ZN(new_n300));
  OAI21_X1  g114(.A(G214), .B1(G237), .B2(G902), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n301), .B(KEYINPUT79), .ZN(new_n302));
  INV_X1    g116(.A(new_n302), .ZN(new_n303));
  XOR2_X1   g117(.A(KEYINPUT86), .B(KEYINPUT20), .Z(new_n304));
  INV_X1    g118(.A(new_n304), .ZN(new_n305));
  XNOR2_X1  g119(.A(G125), .B(G140), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n306), .A2(new_n188), .ZN(new_n307));
  NOR2_X1   g121(.A1(new_n201), .A2(G140), .ZN(new_n308));
  AOI21_X1  g122(.A(new_n308), .B1(new_n193), .B2(G140), .ZN(new_n309));
  OAI211_X1 g123(.A(KEYINPUT87), .B(new_n307), .C1(new_n309), .C2(new_n188), .ZN(new_n310));
  NAND2_X1  g124(.A1(KEYINPUT18), .A2(G131), .ZN(new_n311));
  INV_X1    g125(.A(G237), .ZN(new_n312));
  NAND3_X1  g126(.A1(new_n312), .A2(new_n208), .A3(G214), .ZN(new_n313));
  NOR2_X1   g127(.A1(new_n313), .A2(new_n195), .ZN(new_n314));
  NOR2_X1   g128(.A1(G237), .A2(G953), .ZN(new_n315));
  AOI21_X1  g129(.A(G143), .B1(new_n315), .B2(G214), .ZN(new_n316));
  OAI21_X1  g130(.A(new_n311), .B1(new_n314), .B2(new_n316), .ZN(new_n317));
  NAND2_X1  g131(.A1(new_n313), .A2(new_n195), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(G143), .A3(G214), .ZN(new_n319));
  NAND4_X1  g133(.A1(new_n318), .A2(KEYINPUT18), .A3(G131), .A4(new_n319), .ZN(new_n320));
  NAND2_X1  g134(.A1(new_n317), .A2(new_n320), .ZN(new_n321));
  NAND3_X1  g135(.A1(new_n202), .A2(new_n204), .A3(G140), .ZN(new_n322));
  INV_X1    g136(.A(new_n308), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT87), .ZN(new_n325));
  NAND3_X1  g139(.A1(new_n324), .A2(new_n325), .A3(G146), .ZN(new_n326));
  NAND3_X1  g140(.A1(new_n310), .A2(new_n321), .A3(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(new_n327), .ZN(new_n328));
  OAI21_X1  g142(.A(G131), .B1(new_n314), .B2(new_n316), .ZN(new_n329));
  INV_X1    g143(.A(G131), .ZN(new_n330));
  NAND3_X1  g144(.A1(new_n318), .A2(new_n330), .A3(new_n319), .ZN(new_n331));
  NAND2_X1  g145(.A1(new_n329), .A2(new_n331), .ZN(new_n332));
  NOR2_X1   g146(.A1(new_n332), .A2(KEYINPUT17), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n322), .A2(KEYINPUT16), .A3(new_n323), .ZN(new_n334));
  NOR2_X1   g148(.A1(KEYINPUT16), .A2(G140), .ZN(new_n335));
  NAND2_X1  g149(.A1(new_n205), .A2(new_n335), .ZN(new_n336));
  NAND3_X1  g150(.A1(new_n334), .A2(new_n336), .A3(G146), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n334), .A2(new_n336), .ZN(new_n338));
  NAND2_X1  g152(.A1(new_n338), .A2(new_n188), .ZN(new_n339));
  OAI211_X1 g153(.A(KEYINPUT17), .B(G131), .C1(new_n314), .C2(new_n316), .ZN(new_n340));
  NOR2_X1   g154(.A1(new_n340), .A2(KEYINPUT90), .ZN(new_n341));
  INV_X1    g155(.A(KEYINPUT90), .ZN(new_n342));
  AOI21_X1  g156(.A(new_n330), .B1(new_n318), .B2(new_n319), .ZN(new_n343));
  AOI21_X1  g157(.A(new_n342), .B1(new_n343), .B2(KEYINPUT17), .ZN(new_n344));
  OAI211_X1 g158(.A(new_n337), .B(new_n339), .C1(new_n341), .C2(new_n344), .ZN(new_n345));
  AOI21_X1  g159(.A(new_n333), .B1(new_n345), .B2(KEYINPUT91), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n340), .A2(KEYINPUT90), .ZN(new_n347));
  NAND3_X1  g161(.A1(new_n343), .A2(new_n342), .A3(KEYINPUT17), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  INV_X1    g163(.A(KEYINPUT91), .ZN(new_n350));
  NAND4_X1  g164(.A1(new_n349), .A2(new_n350), .A3(new_n337), .A4(new_n339), .ZN(new_n351));
  AOI21_X1  g165(.A(new_n328), .B1(new_n346), .B2(new_n351), .ZN(new_n352));
  XOR2_X1   g166(.A(G113), .B(G122), .Z(new_n353));
  XOR2_X1   g167(.A(KEYINPUT88), .B(G104), .Z(new_n354));
  XOR2_X1   g168(.A(new_n353), .B(new_n354), .Z(new_n355));
  INV_X1    g169(.A(new_n355), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n306), .A2(KEYINPUT19), .ZN(new_n357));
  AOI21_X1  g171(.A(new_n357), .B1(new_n309), .B2(KEYINPUT19), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n332), .B(new_n337), .C1(new_n358), .C2(G146), .ZN(new_n359));
  NAND2_X1  g173(.A1(new_n359), .A2(new_n327), .ZN(new_n360));
  NAND2_X1  g174(.A1(new_n360), .A2(new_n355), .ZN(new_n361));
  NAND2_X1  g175(.A1(new_n361), .A2(KEYINPUT89), .ZN(new_n362));
  INV_X1    g176(.A(KEYINPUT89), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n360), .A2(new_n363), .A3(new_n355), .ZN(new_n364));
  AOI22_X1  g178(.A1(new_n352), .A2(new_n356), .B1(new_n362), .B2(new_n364), .ZN(new_n365));
  NOR2_X1   g179(.A1(G475), .A2(G902), .ZN(new_n366));
  INV_X1    g180(.A(new_n366), .ZN(new_n367));
  OAI21_X1  g181(.A(new_n305), .B1(new_n365), .B2(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n345), .A2(KEYINPUT91), .ZN(new_n369));
  INV_X1    g183(.A(new_n333), .ZN(new_n370));
  NAND3_X1  g184(.A1(new_n369), .A2(new_n351), .A3(new_n370), .ZN(new_n371));
  NAND3_X1  g185(.A1(new_n371), .A2(new_n327), .A3(new_n356), .ZN(new_n372));
  NAND2_X1  g186(.A1(new_n362), .A2(new_n364), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  INV_X1    g188(.A(KEYINPUT20), .ZN(new_n375));
  NAND3_X1  g189(.A1(new_n374), .A2(new_n375), .A3(new_n366), .ZN(new_n376));
  INV_X1    g190(.A(G902), .ZN(new_n377));
  AOI211_X1 g191(.A(new_n328), .B(new_n355), .C1(new_n346), .C2(new_n351), .ZN(new_n378));
  AOI21_X1  g192(.A(new_n356), .B1(new_n371), .B2(new_n327), .ZN(new_n379));
  OAI21_X1  g193(.A(new_n377), .B1(new_n378), .B2(new_n379), .ZN(new_n380));
  AOI22_X1  g194(.A1(new_n368), .A2(new_n376), .B1(G475), .B2(new_n380), .ZN(new_n381));
  NAND2_X1  g195(.A1(new_n195), .A2(G128), .ZN(new_n382));
  INV_X1    g196(.A(KEYINPUT13), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n382), .A2(new_n383), .ZN(new_n384));
  NAND3_X1  g198(.A1(new_n195), .A2(KEYINPUT13), .A3(G128), .ZN(new_n385));
  NAND2_X1  g199(.A1(new_n187), .A2(G143), .ZN(new_n386));
  NAND3_X1  g200(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n387), .A2(G134), .ZN(new_n388));
  INV_X1    g202(.A(G122), .ZN(new_n389));
  NAND2_X1  g203(.A1(new_n389), .A2(G116), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n235), .A2(G122), .ZN(new_n391));
  NAND2_X1  g205(.A1(new_n390), .A2(new_n391), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n392), .A2(G107), .ZN(new_n393));
  NAND3_X1  g207(.A1(new_n390), .A2(new_n391), .A3(new_n216), .ZN(new_n394));
  NAND2_X1  g208(.A1(new_n393), .A2(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(G134), .ZN(new_n396));
  NAND3_X1  g210(.A1(new_n382), .A2(new_n386), .A3(new_n396), .ZN(new_n397));
  NAND3_X1  g211(.A1(new_n388), .A2(new_n395), .A3(new_n397), .ZN(new_n398));
  NAND2_X1  g212(.A1(new_n398), .A2(KEYINPUT92), .ZN(new_n399));
  INV_X1    g213(.A(KEYINPUT92), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n388), .A2(new_n395), .A3(new_n400), .A4(new_n397), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n382), .A2(new_n386), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n402), .A2(G134), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n403), .A2(new_n397), .ZN(new_n404));
  NAND3_X1  g218(.A1(new_n235), .A2(KEYINPUT14), .A3(G122), .ZN(new_n405));
  OAI211_X1 g219(.A(G107), .B(new_n405), .C1(new_n392), .C2(KEYINPUT14), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(new_n394), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n399), .A2(new_n401), .A3(new_n407), .ZN(new_n408));
  XNOR2_X1  g222(.A(KEYINPUT9), .B(G234), .ZN(new_n409));
  INV_X1    g223(.A(G217), .ZN(new_n410));
  NOR3_X1   g224(.A1(new_n409), .A2(new_n410), .A3(G953), .ZN(new_n411));
  XNOR2_X1  g225(.A(new_n411), .B(KEYINPUT93), .ZN(new_n412));
  INV_X1    g226(.A(new_n412), .ZN(new_n413));
  NAND2_X1  g227(.A1(new_n408), .A2(new_n413), .ZN(new_n414));
  NAND4_X1  g228(.A1(new_n399), .A2(new_n412), .A3(new_n401), .A4(new_n407), .ZN(new_n415));
  AOI21_X1  g229(.A(G902), .B1(new_n414), .B2(new_n415), .ZN(new_n416));
  INV_X1    g230(.A(new_n416), .ZN(new_n417));
  INV_X1    g231(.A(G478), .ZN(new_n418));
  NOR2_X1   g232(.A1(new_n418), .A2(KEYINPUT15), .ZN(new_n419));
  NAND2_X1  g233(.A1(new_n417), .A2(new_n419), .ZN(new_n420));
  AOI211_X1 g234(.A(G902), .B(new_n419), .C1(new_n414), .C2(new_n415), .ZN(new_n421));
  INV_X1    g235(.A(new_n421), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n420), .A2(new_n422), .A3(KEYINPUT94), .ZN(new_n423));
  INV_X1    g237(.A(KEYINPUT94), .ZN(new_n424));
  INV_X1    g238(.A(new_n419), .ZN(new_n425));
  NOR2_X1   g239(.A1(new_n416), .A2(new_n425), .ZN(new_n426));
  OAI21_X1  g240(.A(new_n424), .B1(new_n426), .B2(new_n421), .ZN(new_n427));
  INV_X1    g241(.A(G952), .ZN(new_n428));
  AOI211_X1 g242(.A(G953), .B(new_n428), .C1(G234), .C2(G237), .ZN(new_n429));
  AOI211_X1 g243(.A(new_n377), .B(new_n208), .C1(G234), .C2(G237), .ZN(new_n430));
  XNOR2_X1  g244(.A(KEYINPUT21), .B(G898), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n429), .B1(new_n430), .B2(new_n431), .ZN(new_n432));
  INV_X1    g246(.A(new_n432), .ZN(new_n433));
  AND3_X1   g247(.A1(new_n423), .A2(new_n427), .A3(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n381), .A2(new_n434), .A3(KEYINPUT95), .ZN(new_n435));
  AOI21_X1  g249(.A(KEYINPUT95), .B1(new_n381), .B2(new_n434), .ZN(new_n436));
  OAI211_X1 g250(.A(new_n300), .B(new_n303), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g251(.A(G221), .B1(new_n409), .B2(G902), .ZN(new_n438));
  INV_X1    g252(.A(new_n438), .ZN(new_n439));
  AND2_X1   g253(.A1(new_n248), .A2(new_n200), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n234), .A2(new_n440), .ZN(new_n441));
  NAND2_X1  g255(.A1(new_n189), .A2(new_n196), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n190), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n190), .A2(new_n442), .ZN(new_n444));
  NAND2_X1  g258(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT10), .ZN(new_n446));
  NOR2_X1   g260(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n447), .B1(new_n262), .B2(new_n263), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n291), .A2(new_n192), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n449), .A2(new_n446), .ZN(new_n450));
  NAND3_X1  g264(.A1(new_n441), .A2(new_n448), .A3(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(KEYINPUT11), .ZN(new_n452));
  OAI21_X1  g266(.A(new_n452), .B1(new_n396), .B2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT11), .A3(G134), .ZN(new_n455));
  NAND2_X1  g269(.A1(new_n396), .A2(G137), .ZN(new_n456));
  NAND3_X1  g270(.A1(new_n453), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g271(.A1(new_n457), .A2(G131), .ZN(new_n458));
  NAND4_X1  g272(.A1(new_n453), .A2(new_n455), .A3(new_n330), .A4(new_n456), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n458), .A2(KEYINPUT64), .A3(new_n459), .ZN(new_n460));
  INV_X1    g274(.A(KEYINPUT64), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n457), .A2(new_n461), .A3(G131), .ZN(new_n462));
  NAND2_X1  g276(.A1(new_n460), .A2(new_n462), .ZN(new_n463));
  INV_X1    g277(.A(new_n463), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n451), .A2(new_n464), .ZN(new_n465));
  NAND4_X1  g279(.A1(new_n441), .A2(new_n448), .A3(new_n463), .A4(new_n450), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XNOR2_X1  g281(.A(G110), .B(G140), .ZN(new_n468));
  INV_X1    g282(.A(G227), .ZN(new_n469));
  NOR2_X1   g283(.A1(new_n469), .A2(G953), .ZN(new_n470));
  XNOR2_X1  g284(.A(new_n468), .B(new_n470), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n467), .A2(new_n471), .ZN(new_n472));
  INV_X1    g286(.A(KEYINPUT78), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(KEYINPUT12), .ZN(new_n475));
  INV_X1    g289(.A(new_n449), .ZN(new_n476));
  AOI21_X1  g290(.A(new_n476), .B1(new_n290), .B2(new_n445), .ZN(new_n477));
  OAI21_X1  g291(.A(new_n475), .B1(new_n477), .B2(new_n463), .ZN(new_n478));
  NAND2_X1  g292(.A1(new_n257), .A2(new_n261), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n479), .A2(KEYINPUT75), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n291), .A2(new_n256), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n480), .A2(new_n481), .A3(new_n445), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n482), .A2(new_n449), .ZN(new_n483));
  NAND3_X1  g297(.A1(new_n483), .A2(KEYINPUT12), .A3(new_n464), .ZN(new_n484));
  NAND2_X1  g298(.A1(new_n478), .A2(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n471), .ZN(new_n486));
  NAND2_X1  g300(.A1(new_n466), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g301(.A1(new_n487), .A2(KEYINPUT77), .ZN(new_n488));
  INV_X1    g302(.A(KEYINPUT77), .ZN(new_n489));
  NAND3_X1  g303(.A1(new_n466), .A2(new_n489), .A3(new_n486), .ZN(new_n490));
  NAND3_X1  g304(.A1(new_n485), .A2(new_n488), .A3(new_n490), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n467), .A2(KEYINPUT78), .A3(new_n471), .ZN(new_n492));
  NAND3_X1  g306(.A1(new_n474), .A2(new_n491), .A3(new_n492), .ZN(new_n493));
  INV_X1    g307(.A(G469), .ZN(new_n494));
  NAND3_X1  g308(.A1(new_n493), .A2(new_n494), .A3(new_n377), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n494), .A2(new_n377), .ZN(new_n496));
  NAND3_X1  g310(.A1(new_n466), .A2(KEYINPUT76), .A3(new_n486), .ZN(new_n497));
  NAND2_X1  g311(.A1(new_n497), .A2(new_n465), .ZN(new_n498));
  INV_X1    g312(.A(new_n498), .ZN(new_n499));
  AOI21_X1  g313(.A(KEYINPUT76), .B1(new_n466), .B2(new_n486), .ZN(new_n500));
  INV_X1    g314(.A(new_n500), .ZN(new_n501));
  AOI21_X1  g315(.A(KEYINPUT12), .B1(new_n483), .B2(new_n464), .ZN(new_n502));
  AOI211_X1 g316(.A(new_n475), .B(new_n463), .C1(new_n482), .C2(new_n449), .ZN(new_n503));
  OAI21_X1  g317(.A(new_n466), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  AOI22_X1  g318(.A1(new_n499), .A2(new_n501), .B1(new_n504), .B2(new_n471), .ZN(new_n505));
  AOI21_X1  g319(.A(new_n496), .B1(new_n505), .B2(G469), .ZN(new_n506));
  AOI21_X1  g320(.A(new_n439), .B1(new_n495), .B2(new_n506), .ZN(new_n507));
  INV_X1    g321(.A(new_n507), .ZN(new_n508));
  OAI21_X1  g322(.A(KEYINPUT96), .B1(new_n437), .B2(new_n508), .ZN(new_n509));
  INV_X1    g323(.A(new_n436), .ZN(new_n510));
  NAND3_X1  g324(.A1(new_n381), .A2(new_n434), .A3(KEYINPUT95), .ZN(new_n511));
  NAND2_X1  g325(.A1(new_n510), .A2(new_n511), .ZN(new_n512));
  INV_X1    g326(.A(KEYINPUT96), .ZN(new_n513));
  NOR2_X1   g327(.A1(new_n299), .A2(new_n302), .ZN(new_n514));
  NAND4_X1  g328(.A1(new_n512), .A2(new_n513), .A3(new_n507), .A4(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT69), .ZN(new_n516));
  INV_X1    g330(.A(KEYINPUT23), .ZN(new_n517));
  NOR2_X1   g331(.A1(new_n516), .A2(new_n517), .ZN(new_n518));
  NOR2_X1   g332(.A1(KEYINPUT69), .A2(KEYINPUT23), .ZN(new_n519));
  OAI211_X1 g333(.A(G119), .B(new_n187), .C1(new_n518), .C2(new_n519), .ZN(new_n520));
  OAI22_X1  g334(.A1(new_n516), .A2(new_n517), .B1(new_n238), .B2(G128), .ZN(new_n521));
  OAI211_X1 g335(.A(new_n520), .B(new_n521), .C1(G119), .C2(new_n187), .ZN(new_n522));
  XNOR2_X1  g336(.A(KEYINPUT71), .B(G110), .ZN(new_n523));
  XNOR2_X1  g337(.A(G119), .B(G128), .ZN(new_n524));
  XOR2_X1   g338(.A(KEYINPUT24), .B(G110), .Z(new_n525));
  OAI22_X1  g339(.A1(new_n522), .A2(new_n523), .B1(new_n524), .B2(new_n525), .ZN(new_n526));
  NAND3_X1  g340(.A1(new_n526), .A2(new_n307), .A3(new_n337), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n339), .A2(new_n337), .ZN(new_n528));
  AOI22_X1  g342(.A1(new_n522), .A2(G110), .B1(new_n524), .B2(new_n525), .ZN(new_n529));
  NAND2_X1  g343(.A1(new_n528), .A2(new_n529), .ZN(new_n530));
  NAND2_X1  g344(.A1(new_n527), .A2(new_n530), .ZN(new_n531));
  XNOR2_X1  g345(.A(KEYINPUT22), .B(G137), .ZN(new_n532));
  NAND3_X1  g346(.A1(new_n208), .A2(G221), .A3(G234), .ZN(new_n533));
  XNOR2_X1  g347(.A(new_n532), .B(new_n533), .ZN(new_n534));
  INV_X1    g348(.A(new_n534), .ZN(new_n535));
  NAND2_X1  g349(.A1(new_n531), .A2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n527), .A2(new_n530), .A3(new_n534), .ZN(new_n537));
  AND2_X1   g351(.A1(new_n536), .A2(new_n537), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n538), .A2(KEYINPUT25), .A3(new_n377), .ZN(new_n539));
  NAND3_X1  g353(.A1(new_n536), .A2(new_n377), .A3(new_n537), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT25), .ZN(new_n541));
  NAND2_X1  g355(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  NAND2_X1  g356(.A1(new_n539), .A2(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n410), .B1(G234), .B2(new_n377), .ZN(new_n544));
  NAND2_X1  g358(.A1(new_n543), .A2(new_n544), .ZN(new_n545));
  NOR2_X1   g359(.A1(new_n544), .A2(G902), .ZN(new_n546));
  NAND2_X1  g360(.A1(new_n538), .A2(new_n546), .ZN(new_n547));
  NAND2_X1  g361(.A1(new_n545), .A2(new_n547), .ZN(new_n548));
  NAND3_X1  g362(.A1(new_n460), .A2(new_n462), .A3(new_n200), .ZN(new_n549));
  INV_X1    g363(.A(KEYINPUT30), .ZN(new_n550));
  INV_X1    g364(.A(new_n456), .ZN(new_n551));
  NOR2_X1   g365(.A1(new_n396), .A2(G137), .ZN(new_n552));
  OAI21_X1  g366(.A(G131), .B1(new_n551), .B2(new_n552), .ZN(new_n553));
  NAND4_X1  g367(.A1(new_n443), .A2(new_n444), .A3(new_n459), .A4(new_n553), .ZN(new_n554));
  AND3_X1   g368(.A1(new_n549), .A2(new_n550), .A3(new_n554), .ZN(new_n555));
  AOI21_X1  g369(.A(new_n550), .B1(new_n549), .B2(new_n554), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n247), .B1(new_n555), .B2(new_n556), .ZN(new_n557));
  NAND2_X1  g371(.A1(new_n315), .A2(G210), .ZN(new_n558));
  XNOR2_X1  g372(.A(new_n558), .B(KEYINPUT27), .ZN(new_n559));
  XNOR2_X1  g373(.A(KEYINPUT26), .B(G101), .ZN(new_n560));
  XNOR2_X1  g374(.A(new_n559), .B(new_n560), .ZN(new_n561));
  INV_X1    g375(.A(new_n247), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n549), .A2(new_n562), .A3(new_n554), .ZN(new_n563));
  NAND3_X1  g377(.A1(new_n557), .A2(new_n561), .A3(new_n563), .ZN(new_n564));
  NAND2_X1  g378(.A1(new_n564), .A2(KEYINPUT31), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n565), .A2(KEYINPUT66), .ZN(new_n566));
  INV_X1    g380(.A(new_n561), .ZN(new_n567));
  INV_X1    g381(.A(KEYINPUT67), .ZN(new_n568));
  AND3_X1   g382(.A1(new_n549), .A2(new_n562), .A3(new_n554), .ZN(new_n569));
  AOI21_X1  g383(.A(new_n562), .B1(new_n549), .B2(new_n554), .ZN(new_n570));
  OAI211_X1 g384(.A(new_n568), .B(KEYINPUT28), .C1(new_n569), .C2(new_n570), .ZN(new_n571));
  INV_X1    g385(.A(KEYINPUT28), .ZN(new_n572));
  NAND2_X1  g386(.A1(new_n563), .A2(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g388(.A1(new_n549), .A2(new_n554), .ZN(new_n575));
  NAND2_X1  g389(.A1(new_n575), .A2(new_n247), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n576), .A2(new_n563), .ZN(new_n577));
  AOI21_X1  g391(.A(new_n568), .B1(new_n577), .B2(KEYINPUT28), .ZN(new_n578));
  OAI21_X1  g392(.A(new_n567), .B1(new_n574), .B2(new_n578), .ZN(new_n579));
  INV_X1    g393(.A(KEYINPUT31), .ZN(new_n580));
  NAND4_X1  g394(.A1(new_n557), .A2(new_n580), .A3(new_n561), .A4(new_n563), .ZN(new_n581));
  INV_X1    g395(.A(KEYINPUT66), .ZN(new_n582));
  NAND3_X1  g396(.A1(new_n564), .A2(new_n582), .A3(KEYINPUT31), .ZN(new_n583));
  NAND4_X1  g397(.A1(new_n566), .A2(new_n579), .A3(new_n581), .A4(new_n583), .ZN(new_n584));
  NOR2_X1   g398(.A1(G472), .A2(G902), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n584), .A2(new_n585), .ZN(new_n586));
  NAND2_X1  g400(.A1(new_n586), .A2(KEYINPUT32), .ZN(new_n587));
  INV_X1    g401(.A(KEYINPUT32), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n589));
  NAND2_X1  g403(.A1(new_n587), .A2(new_n589), .ZN(new_n590));
  NOR3_X1   g404(.A1(new_n574), .A2(new_n578), .A3(new_n567), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n557), .A2(new_n563), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(new_n567), .ZN(new_n593));
  INV_X1    g407(.A(new_n593), .ZN(new_n594));
  NOR3_X1   g408(.A1(new_n591), .A2(new_n594), .A3(KEYINPUT29), .ZN(new_n595));
  INV_X1    g409(.A(KEYINPUT68), .ZN(new_n596));
  NAND2_X1  g410(.A1(new_n563), .A2(new_n596), .ZN(new_n597));
  INV_X1    g411(.A(new_n597), .ZN(new_n598));
  AOI21_X1  g412(.A(new_n598), .B1(new_n577), .B2(KEYINPUT68), .ZN(new_n599));
  OAI21_X1  g413(.A(new_n573), .B1(new_n599), .B2(new_n572), .ZN(new_n600));
  NAND2_X1  g414(.A1(new_n561), .A2(KEYINPUT29), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n377), .B1(new_n600), .B2(new_n601), .ZN(new_n602));
  OAI21_X1  g416(.A(G472), .B1(new_n595), .B2(new_n602), .ZN(new_n603));
  AOI21_X1  g417(.A(new_n548), .B1(new_n590), .B2(new_n603), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n509), .A2(new_n515), .A3(new_n604), .ZN(new_n605));
  XOR2_X1   g419(.A(KEYINPUT97), .B(G101), .Z(new_n606));
  XNOR2_X1  g420(.A(new_n605), .B(new_n606), .ZN(G3));
  NOR2_X1   g421(.A1(new_n508), .A2(new_n548), .ZN(new_n608));
  OAI21_X1  g422(.A(new_n301), .B1(new_n297), .B2(new_n298), .ZN(new_n609));
  NAND2_X1  g423(.A1(new_n380), .A2(G475), .ZN(new_n610));
  AOI21_X1  g424(.A(new_n304), .B1(new_n374), .B2(new_n366), .ZN(new_n611));
  AOI211_X1 g425(.A(KEYINPUT20), .B(new_n367), .C1(new_n372), .C2(new_n373), .ZN(new_n612));
  OAI21_X1  g426(.A(new_n610), .B1(new_n611), .B2(new_n612), .ZN(new_n613));
  NOR2_X1   g427(.A1(new_n418), .A2(new_n377), .ZN(new_n614));
  INV_X1    g428(.A(new_n614), .ZN(new_n615));
  OAI21_X1  g429(.A(new_n615), .B1(new_n417), .B2(G478), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n414), .A2(new_n415), .ZN(new_n617));
  INV_X1    g431(.A(KEYINPUT33), .ZN(new_n618));
  NAND2_X1  g432(.A1(new_n617), .A2(new_n618), .ZN(new_n619));
  NAND3_X1  g433(.A1(new_n414), .A2(KEYINPUT33), .A3(new_n415), .ZN(new_n620));
  AOI21_X1  g434(.A(new_n418), .B1(new_n619), .B2(new_n620), .ZN(new_n621));
  NOR2_X1   g435(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g436(.A1(new_n613), .A2(new_n622), .ZN(new_n623));
  NOR3_X1   g437(.A1(new_n609), .A2(new_n623), .A3(new_n432), .ZN(new_n624));
  INV_X1    g438(.A(G472), .ZN(new_n625));
  AOI21_X1  g439(.A(new_n625), .B1(new_n584), .B2(new_n377), .ZN(new_n626));
  AOI21_X1  g440(.A(new_n626), .B1(new_n585), .B2(new_n584), .ZN(new_n627));
  NAND3_X1  g441(.A1(new_n608), .A2(new_n624), .A3(new_n627), .ZN(new_n628));
  XOR2_X1   g442(.A(KEYINPUT34), .B(G104), .Z(new_n629));
  XNOR2_X1  g443(.A(new_n628), .B(new_n629), .ZN(new_n630));
  XNOR2_X1  g444(.A(KEYINPUT98), .B(KEYINPUT99), .ZN(new_n631));
  XNOR2_X1  g445(.A(new_n630), .B(new_n631), .ZN(G6));
  INV_X1    g446(.A(new_n301), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n278), .A2(new_n295), .ZN(new_n634));
  INV_X1    g448(.A(new_n296), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  NAND3_X1  g450(.A1(new_n278), .A2(new_n295), .A3(new_n296), .ZN(new_n637));
  AOI21_X1  g451(.A(new_n633), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND2_X1  g452(.A1(new_n423), .A2(new_n427), .ZN(new_n639));
  NAND3_X1  g453(.A1(new_n374), .A2(new_n366), .A3(new_n304), .ZN(new_n640));
  NAND2_X1  g454(.A1(new_n368), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g455(.A1(new_n641), .A2(new_n610), .ZN(new_n642));
  INV_X1    g456(.A(new_n642), .ZN(new_n643));
  NAND4_X1  g457(.A1(new_n638), .A2(new_n433), .A3(new_n639), .A4(new_n643), .ZN(new_n644));
  INV_X1    g458(.A(new_n644), .ZN(new_n645));
  NAND3_X1  g459(.A1(new_n608), .A2(new_n627), .A3(new_n645), .ZN(new_n646));
  XOR2_X1   g460(.A(new_n646), .B(KEYINPUT100), .Z(new_n647));
  XNOR2_X1  g461(.A(KEYINPUT35), .B(G107), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n647), .B(new_n648), .ZN(G9));
  INV_X1    g463(.A(KEYINPUT101), .ZN(new_n650));
  NOR2_X1   g464(.A1(new_n535), .A2(KEYINPUT36), .ZN(new_n651));
  XNOR2_X1  g465(.A(new_n531), .B(new_n651), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n652), .A2(new_n546), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n545), .A2(new_n650), .A3(new_n653), .ZN(new_n654));
  INV_X1    g468(.A(new_n544), .ZN(new_n655));
  AOI21_X1  g469(.A(new_n655), .B1(new_n539), .B2(new_n542), .ZN(new_n656));
  INV_X1    g470(.A(new_n653), .ZN(new_n657));
  OAI21_X1  g471(.A(KEYINPUT101), .B1(new_n656), .B2(new_n657), .ZN(new_n658));
  AND2_X1   g472(.A1(new_n654), .A2(new_n658), .ZN(new_n659));
  AND2_X1   g473(.A1(new_n627), .A2(new_n659), .ZN(new_n660));
  NAND3_X1  g474(.A1(new_n509), .A2(new_n515), .A3(new_n660), .ZN(new_n661));
  XOR2_X1   g475(.A(KEYINPUT37), .B(G110), .Z(new_n662));
  XNOR2_X1  g476(.A(new_n661), .B(new_n662), .ZN(G12));
  AND3_X1   g477(.A1(new_n584), .A2(new_n588), .A3(new_n585), .ZN(new_n664));
  AOI21_X1  g478(.A(new_n588), .B1(new_n584), .B2(new_n585), .ZN(new_n665));
  OAI21_X1  g479(.A(new_n603), .B1(new_n664), .B2(new_n665), .ZN(new_n666));
  NAND3_X1  g480(.A1(new_n666), .A2(new_n507), .A3(new_n659), .ZN(new_n667));
  INV_X1    g481(.A(new_n639), .ZN(new_n668));
  INV_X1    g482(.A(G900), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n430), .A2(new_n669), .ZN(new_n670));
  INV_X1    g484(.A(new_n429), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  INV_X1    g486(.A(new_n672), .ZN(new_n673));
  NOR3_X1   g487(.A1(new_n642), .A2(new_n668), .A3(new_n673), .ZN(new_n674));
  NAND2_X1  g488(.A1(new_n674), .A2(new_n638), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n667), .A2(new_n675), .ZN(new_n676));
  XNOR2_X1  g490(.A(new_n676), .B(new_n187), .ZN(G30));
  NAND2_X1  g491(.A1(new_n599), .A2(new_n567), .ZN(new_n678));
  NAND2_X1  g492(.A1(new_n678), .A2(new_n377), .ZN(new_n679));
  AOI21_X1  g493(.A(new_n567), .B1(new_n557), .B2(new_n563), .ZN(new_n680));
  OAI21_X1  g494(.A(G472), .B1(new_n679), .B2(new_n680), .ZN(new_n681));
  AOI21_X1  g495(.A(KEYINPUT102), .B1(new_n590), .B2(new_n681), .ZN(new_n682));
  OAI211_X1 g496(.A(KEYINPUT102), .B(new_n681), .C1(new_n664), .C2(new_n665), .ZN(new_n683));
  INV_X1    g497(.A(new_n683), .ZN(new_n684));
  OR2_X1    g498(.A1(new_n682), .A2(new_n684), .ZN(new_n685));
  XNOR2_X1  g499(.A(new_n672), .B(KEYINPUT39), .ZN(new_n686));
  NAND2_X1  g500(.A1(new_n507), .A2(new_n686), .ZN(new_n687));
  NAND2_X1  g501(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n688));
  OR2_X1    g502(.A1(new_n687), .A2(KEYINPUT40), .ZN(new_n689));
  INV_X1    g503(.A(KEYINPUT38), .ZN(new_n690));
  OAI21_X1  g504(.A(new_n690), .B1(new_n297), .B2(new_n298), .ZN(new_n691));
  NAND3_X1  g505(.A1(new_n636), .A2(KEYINPUT38), .A3(new_n637), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n691), .A2(new_n692), .ZN(new_n693));
  NOR2_X1   g507(.A1(new_n656), .A2(new_n657), .ZN(new_n694));
  INV_X1    g508(.A(new_n694), .ZN(new_n695));
  NAND3_X1  g509(.A1(new_n613), .A2(new_n639), .A3(new_n301), .ZN(new_n696));
  NOR3_X1   g510(.A1(new_n693), .A2(new_n695), .A3(new_n696), .ZN(new_n697));
  NAND4_X1  g511(.A1(new_n685), .A2(new_n688), .A3(new_n689), .A4(new_n697), .ZN(new_n698));
  XNOR2_X1  g512(.A(new_n698), .B(G143), .ZN(G45));
  NAND3_X1  g513(.A1(new_n613), .A2(new_n622), .A3(new_n672), .ZN(new_n700));
  NOR2_X1   g514(.A1(new_n609), .A2(new_n700), .ZN(new_n701));
  INV_X1    g515(.A(new_n701), .ZN(new_n702));
  OAI21_X1  g516(.A(KEYINPUT103), .B1(new_n667), .B2(new_n702), .ZN(new_n703));
  NAND2_X1  g517(.A1(new_n654), .A2(new_n658), .ZN(new_n704));
  AOI21_X1  g518(.A(new_n704), .B1(new_n590), .B2(new_n603), .ZN(new_n705));
  INV_X1    g519(.A(KEYINPUT103), .ZN(new_n706));
  NAND4_X1  g520(.A1(new_n705), .A2(new_n706), .A3(new_n507), .A4(new_n701), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G146), .ZN(G48));
  AND3_X1   g523(.A1(new_n493), .A2(new_n494), .A3(new_n377), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n494), .B1(new_n493), .B2(new_n377), .ZN(new_n711));
  NOR3_X1   g525(.A1(new_n710), .A2(new_n711), .A3(new_n439), .ZN(new_n712));
  NAND3_X1  g526(.A1(new_n604), .A2(new_n624), .A3(new_n712), .ZN(new_n713));
  XNOR2_X1  g527(.A(KEYINPUT41), .B(G113), .ZN(new_n714));
  XNOR2_X1  g528(.A(new_n714), .B(KEYINPUT104), .ZN(new_n715));
  XNOR2_X1  g529(.A(new_n713), .B(new_n715), .ZN(G15));
  NOR2_X1   g530(.A1(new_n710), .A2(new_n711), .ZN(new_n717));
  INV_X1    g531(.A(new_n548), .ZN(new_n718));
  NAND4_X1  g532(.A1(new_n717), .A2(new_n666), .A3(new_n438), .A4(new_n718), .ZN(new_n719));
  OAI21_X1  g533(.A(KEYINPUT105), .B1(new_n719), .B2(new_n644), .ZN(new_n720));
  INV_X1    g534(.A(KEYINPUT105), .ZN(new_n721));
  NAND4_X1  g535(.A1(new_n645), .A2(new_n604), .A3(new_n721), .A4(new_n712), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  XNOR2_X1  g537(.A(new_n723), .B(G116), .ZN(G18));
  NAND2_X1  g538(.A1(new_n493), .A2(new_n377), .ZN(new_n725));
  NAND2_X1  g539(.A1(new_n725), .A2(G469), .ZN(new_n726));
  NAND4_X1  g540(.A1(new_n638), .A2(new_n726), .A3(new_n438), .A4(new_n495), .ZN(new_n727));
  INV_X1    g541(.A(new_n727), .ZN(new_n728));
  NAND3_X1  g542(.A1(new_n728), .A2(new_n512), .A3(new_n705), .ZN(new_n729));
  XNOR2_X1  g543(.A(new_n729), .B(G119), .ZN(G21));
  NOR2_X1   g544(.A1(new_n696), .A2(new_n299), .ZN(new_n731));
  INV_X1    g545(.A(new_n585), .ZN(new_n732));
  INV_X1    g546(.A(KEYINPUT106), .ZN(new_n733));
  OAI211_X1 g547(.A(new_n733), .B(new_n573), .C1(new_n599), .C2(new_n572), .ZN(new_n734));
  OAI21_X1  g548(.A(KEYINPUT68), .B1(new_n569), .B2(new_n570), .ZN(new_n735));
  AOI21_X1  g549(.A(new_n572), .B1(new_n735), .B2(new_n597), .ZN(new_n736));
  INV_X1    g550(.A(new_n573), .ZN(new_n737));
  OAI21_X1  g551(.A(KEYINPUT106), .B1(new_n736), .B2(new_n737), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n734), .A2(new_n738), .A3(new_n567), .ZN(new_n739));
  AND2_X1   g553(.A1(new_n565), .A2(new_n581), .ZN(new_n740));
  AOI21_X1  g554(.A(new_n732), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NOR3_X1   g555(.A1(new_n626), .A2(new_n548), .A3(new_n741), .ZN(new_n742));
  NAND4_X1  g556(.A1(new_n712), .A2(new_n731), .A3(new_n433), .A4(new_n742), .ZN(new_n743));
  XNOR2_X1  g557(.A(new_n743), .B(G122), .ZN(G24));
  NOR2_X1   g558(.A1(new_n626), .A2(new_n741), .ZN(new_n745));
  INV_X1    g559(.A(new_n622), .ZN(new_n746));
  NOR3_X1   g560(.A1(new_n381), .A2(new_n746), .A3(new_n673), .ZN(new_n747));
  NAND3_X1  g561(.A1(new_n745), .A2(new_n695), .A3(new_n747), .ZN(new_n748));
  NOR2_X1   g562(.A1(new_n727), .A2(new_n748), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n749), .B(new_n201), .ZN(G27));
  INV_X1    g564(.A(KEYINPUT42), .ZN(new_n751));
  NOR3_X1   g565(.A1(new_n297), .A2(new_n298), .A3(new_n633), .ZN(new_n752));
  NAND4_X1  g566(.A1(new_n666), .A2(new_n507), .A3(new_n718), .A4(new_n752), .ZN(new_n753));
  OAI21_X1  g567(.A(new_n751), .B1(new_n753), .B2(new_n700), .ZN(new_n754));
  AND2_X1   g568(.A1(new_n507), .A2(new_n752), .ZN(new_n755));
  NAND4_X1  g569(.A1(new_n755), .A2(new_n604), .A3(KEYINPUT42), .A4(new_n747), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n754), .A2(new_n756), .ZN(new_n757));
  XNOR2_X1  g571(.A(new_n757), .B(G131), .ZN(G33));
  XNOR2_X1  g572(.A(new_n674), .B(KEYINPUT107), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n759), .A2(new_n604), .A3(new_n755), .ZN(new_n760));
  XNOR2_X1  g574(.A(new_n760), .B(G134), .ZN(G36));
  NOR2_X1   g575(.A1(new_n627), .A2(new_n694), .ZN(new_n762));
  INV_X1    g576(.A(KEYINPUT108), .ZN(new_n763));
  OAI211_X1 g577(.A(new_n610), .B(new_n763), .C1(new_n611), .C2(new_n612), .ZN(new_n764));
  OAI211_X1 g578(.A(new_n610), .B(new_n622), .C1(new_n611), .C2(new_n612), .ZN(new_n765));
  INV_X1    g579(.A(KEYINPUT43), .ZN(new_n766));
  NAND3_X1  g580(.A1(new_n764), .A2(new_n765), .A3(new_n766), .ZN(new_n767));
  OAI211_X1 g581(.A(new_n381), .B(new_n622), .C1(new_n763), .C2(KEYINPUT43), .ZN(new_n768));
  NAND2_X1  g582(.A1(new_n767), .A2(new_n768), .ZN(new_n769));
  AND2_X1   g583(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n770));
  NOR2_X1   g584(.A1(new_n769), .A2(KEYINPUT109), .ZN(new_n771));
  OAI21_X1  g585(.A(new_n762), .B1(new_n770), .B2(new_n771), .ZN(new_n772));
  INV_X1    g586(.A(KEYINPUT44), .ZN(new_n773));
  OR2_X1    g587(.A1(new_n772), .A2(new_n773), .ZN(new_n774));
  AND2_X1   g588(.A1(new_n774), .A2(new_n752), .ZN(new_n775));
  INV_X1    g589(.A(new_n686), .ZN(new_n776));
  INV_X1    g590(.A(new_n466), .ZN(new_n777));
  AOI21_X1  g591(.A(new_n777), .B1(new_n478), .B2(new_n484), .ZN(new_n778));
  OAI22_X1  g592(.A1(new_n778), .A2(new_n486), .B1(new_n498), .B2(new_n500), .ZN(new_n779));
  INV_X1    g593(.A(KEYINPUT45), .ZN(new_n780));
  AOI21_X1  g594(.A(new_n494), .B1(new_n779), .B2(new_n780), .ZN(new_n781));
  NAND2_X1  g595(.A1(new_n505), .A2(KEYINPUT45), .ZN(new_n782));
  AOI21_X1  g596(.A(new_n496), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g597(.A1(new_n783), .A2(KEYINPUT46), .ZN(new_n784));
  OAI21_X1  g598(.A(new_n495), .B1(new_n783), .B2(KEYINPUT46), .ZN(new_n785));
  OAI21_X1  g599(.A(new_n438), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  AOI211_X1 g600(.A(new_n776), .B(new_n786), .C1(new_n772), .C2(new_n773), .ZN(new_n787));
  NAND2_X1  g601(.A1(new_n775), .A2(new_n787), .ZN(new_n788));
  XNOR2_X1  g602(.A(new_n788), .B(G137), .ZN(G39));
  INV_X1    g603(.A(KEYINPUT47), .ZN(new_n790));
  NAND2_X1  g604(.A1(new_n786), .A2(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(KEYINPUT47), .B(new_n438), .C1(new_n784), .C2(new_n785), .ZN(new_n792));
  NAND2_X1  g606(.A1(new_n791), .A2(new_n792), .ZN(new_n793));
  NAND3_X1  g607(.A1(new_n636), .A2(new_n637), .A3(new_n301), .ZN(new_n794));
  NOR4_X1   g608(.A1(new_n666), .A2(new_n700), .A3(new_n794), .A4(new_n718), .ZN(new_n795));
  NAND2_X1  g609(.A1(new_n793), .A2(new_n795), .ZN(new_n796));
  XNOR2_X1  g610(.A(new_n796), .B(G140), .ZN(G42));
  INV_X1    g611(.A(KEYINPUT118), .ZN(new_n798));
  NAND2_X1  g612(.A1(new_n717), .A2(new_n439), .ZN(new_n799));
  NAND3_X1  g613(.A1(new_n791), .A2(new_n792), .A3(new_n799), .ZN(new_n800));
  AND3_X1   g614(.A1(new_n769), .A2(new_n429), .A3(new_n742), .ZN(new_n801));
  AND2_X1   g615(.A1(new_n801), .A2(new_n752), .ZN(new_n802));
  NAND2_X1  g616(.A1(new_n800), .A2(new_n802), .ZN(new_n803));
  INV_X1    g617(.A(new_n803), .ZN(new_n804));
  INV_X1    g618(.A(KEYINPUT113), .ZN(new_n805));
  AND2_X1   g619(.A1(new_n691), .A2(new_n692), .ZN(new_n806));
  NAND4_X1  g620(.A1(new_n726), .A2(new_n438), .A3(new_n495), .A4(new_n633), .ZN(new_n807));
  OAI21_X1  g621(.A(new_n805), .B1(new_n806), .B2(new_n807), .ZN(new_n808));
  NAND4_X1  g622(.A1(new_n712), .A2(KEYINPUT113), .A3(new_n633), .A4(new_n693), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n808), .A2(new_n801), .A3(new_n809), .A4(KEYINPUT114), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n810), .A2(KEYINPUT115), .ZN(new_n811));
  INV_X1    g625(.A(KEYINPUT50), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n811), .A2(new_n812), .ZN(new_n813));
  NAND3_X1  g627(.A1(new_n808), .A2(new_n801), .A3(new_n809), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT115), .ZN(new_n815));
  OAI21_X1  g629(.A(KEYINPUT114), .B1(new_n815), .B2(new_n812), .ZN(new_n816));
  NAND2_X1  g630(.A1(new_n814), .A2(new_n816), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n712), .A2(new_n752), .ZN(new_n818));
  NAND2_X1  g632(.A1(new_n769), .A2(new_n429), .ZN(new_n819));
  NAND2_X1  g633(.A1(new_n745), .A2(new_n695), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n818), .A2(new_n819), .A3(new_n820), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n548), .A2(new_n671), .ZN(new_n822));
  NAND3_X1  g636(.A1(new_n712), .A2(new_n752), .A3(new_n822), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n823), .A2(new_n682), .A3(new_n684), .ZN(new_n824));
  NOR2_X1   g638(.A1(new_n613), .A2(new_n622), .ZN(new_n825));
  AOI21_X1  g639(.A(new_n821), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NAND3_X1  g640(.A1(new_n813), .A2(new_n817), .A3(new_n826), .ZN(new_n827));
  INV_X1    g641(.A(KEYINPUT116), .ZN(new_n828));
  AOI21_X1  g642(.A(new_n804), .B1(new_n827), .B2(new_n828), .ZN(new_n829));
  NAND4_X1  g643(.A1(new_n813), .A2(KEYINPUT116), .A3(new_n817), .A4(new_n826), .ZN(new_n830));
  AOI21_X1  g644(.A(KEYINPUT51), .B1(new_n829), .B2(new_n830), .ZN(new_n831));
  NAND3_X1  g645(.A1(new_n824), .A2(new_n613), .A3(new_n622), .ZN(new_n832));
  NAND2_X1  g646(.A1(new_n666), .A2(new_n718), .ZN(new_n833));
  OR2_X1    g647(.A1(new_n818), .A2(new_n819), .ZN(new_n834));
  NOR2_X1   g648(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n835));
  AND2_X1   g649(.A1(KEYINPUT117), .A2(KEYINPUT48), .ZN(new_n836));
  OR4_X1    g650(.A1(new_n833), .A2(new_n834), .A3(new_n835), .A4(new_n836), .ZN(new_n837));
  AOI211_X1 g651(.A(new_n428), .B(G953), .C1(new_n801), .C2(new_n728), .ZN(new_n838));
  OAI21_X1  g652(.A(new_n835), .B1(new_n834), .B2(new_n833), .ZN(new_n839));
  AND4_X1   g653(.A1(new_n832), .A2(new_n837), .A3(new_n838), .A4(new_n839), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n826), .A2(new_n817), .ZN(new_n841));
  AOI21_X1  g655(.A(KEYINPUT50), .B1(new_n810), .B2(KEYINPUT115), .ZN(new_n842));
  NOR2_X1   g656(.A1(new_n841), .A2(new_n842), .ZN(new_n843));
  NAND3_X1  g657(.A1(new_n843), .A2(KEYINPUT51), .A3(new_n803), .ZN(new_n844));
  NAND2_X1  g658(.A1(new_n840), .A2(new_n844), .ZN(new_n845));
  OAI21_X1  g659(.A(new_n798), .B1(new_n831), .B2(new_n845), .ZN(new_n846));
  OAI21_X1  g660(.A(new_n828), .B1(new_n841), .B2(new_n842), .ZN(new_n847));
  NAND3_X1  g661(.A1(new_n847), .A2(new_n830), .A3(new_n803), .ZN(new_n848));
  INV_X1    g662(.A(KEYINPUT51), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n848), .A2(new_n849), .ZN(new_n850));
  NAND4_X1  g664(.A1(new_n850), .A2(KEYINPUT118), .A3(new_n844), .A4(new_n840), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT53), .ZN(new_n852));
  AND2_X1   g666(.A1(new_n720), .A2(new_n722), .ZN(new_n853));
  NAND3_X1  g667(.A1(new_n729), .A2(new_n713), .A3(new_n743), .ZN(new_n854));
  OAI21_X1  g668(.A(KEYINPUT111), .B1(new_n853), .B2(new_n854), .ZN(new_n855));
  AND3_X1   g669(.A1(new_n729), .A2(new_n713), .A3(new_n743), .ZN(new_n856));
  INV_X1    g670(.A(KEYINPUT111), .ZN(new_n857));
  NAND3_X1  g671(.A1(new_n856), .A2(new_n857), .A3(new_n723), .ZN(new_n858));
  NOR2_X1   g672(.A1(new_n426), .A2(new_n421), .ZN(new_n859));
  NOR2_X1   g673(.A1(new_n613), .A2(new_n859), .ZN(new_n860));
  AOI21_X1  g674(.A(new_n860), .B1(new_n613), .B2(new_n622), .ZN(new_n861));
  NOR2_X1   g675(.A1(new_n861), .A2(new_n432), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n608), .A3(new_n514), .A4(new_n627), .ZN(new_n863));
  AND3_X1   g677(.A1(new_n605), .A2(new_n661), .A3(new_n863), .ZN(new_n864));
  NAND4_X1  g678(.A1(new_n641), .A2(new_n610), .A3(new_n859), .A4(new_n672), .ZN(new_n865));
  INV_X1    g679(.A(new_n865), .ZN(new_n866));
  AOI21_X1  g680(.A(KEYINPUT112), .B1(new_n752), .B2(new_n866), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT112), .ZN(new_n868));
  NOR3_X1   g682(.A1(new_n794), .A2(new_n868), .A3(new_n865), .ZN(new_n869));
  NOR2_X1   g683(.A1(new_n867), .A2(new_n869), .ZN(new_n870));
  INV_X1    g684(.A(new_n667), .ZN(new_n871));
  NOR2_X1   g685(.A1(new_n820), .A2(new_n700), .ZN(new_n872));
  AOI22_X1  g686(.A1(new_n870), .A2(new_n871), .B1(new_n872), .B2(new_n755), .ZN(new_n873));
  AND3_X1   g687(.A1(new_n757), .A2(new_n873), .A3(new_n760), .ZN(new_n874));
  NAND4_X1  g688(.A1(new_n855), .A2(new_n858), .A3(new_n864), .A4(new_n874), .ZN(new_n875));
  OAI22_X1  g689(.A1(new_n667), .A2(new_n675), .B1(new_n727), .B2(new_n748), .ZN(new_n876));
  AOI21_X1  g690(.A(new_n876), .B1(new_n707), .B2(new_n703), .ZN(new_n877));
  NAND2_X1  g691(.A1(new_n590), .A2(new_n681), .ZN(new_n878));
  NOR2_X1   g692(.A1(new_n695), .A2(new_n673), .ZN(new_n879));
  NAND4_X1  g693(.A1(new_n878), .A2(new_n731), .A3(new_n507), .A4(new_n879), .ZN(new_n880));
  AOI21_X1  g694(.A(KEYINPUT52), .B1(new_n877), .B2(new_n880), .ZN(new_n881));
  INV_X1    g695(.A(new_n876), .ZN(new_n882));
  AND4_X1   g696(.A1(KEYINPUT52), .A2(new_n708), .A3(new_n882), .A4(new_n880), .ZN(new_n883));
  NOR2_X1   g697(.A1(new_n881), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g698(.A(new_n852), .B1(new_n875), .B2(new_n884), .ZN(new_n885));
  AND3_X1   g699(.A1(new_n856), .A2(new_n857), .A3(new_n723), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n857), .B1(new_n856), .B2(new_n723), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n886), .A2(new_n887), .ZN(new_n888));
  NAND3_X1  g702(.A1(new_n708), .A2(new_n882), .A3(new_n880), .ZN(new_n889));
  INV_X1    g703(.A(KEYINPUT52), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g705(.A1(new_n877), .A2(KEYINPUT52), .A3(new_n880), .ZN(new_n892));
  NAND2_X1  g706(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NAND3_X1  g707(.A1(new_n605), .A2(new_n661), .A3(new_n863), .ZN(new_n894));
  NAND3_X1  g708(.A1(new_n757), .A2(new_n873), .A3(new_n760), .ZN(new_n895));
  NOR2_X1   g709(.A1(new_n894), .A2(new_n895), .ZN(new_n896));
  NAND4_X1  g710(.A1(new_n888), .A2(KEYINPUT53), .A3(new_n893), .A4(new_n896), .ZN(new_n897));
  NAND2_X1  g711(.A1(new_n885), .A2(new_n897), .ZN(new_n898));
  NAND2_X1  g712(.A1(new_n898), .A2(KEYINPUT54), .ZN(new_n899));
  INV_X1    g713(.A(KEYINPUT54), .ZN(new_n900));
  NOR3_X1   g714(.A1(new_n853), .A2(new_n852), .A3(new_n854), .ZN(new_n901));
  NAND3_X1  g715(.A1(new_n893), .A2(new_n896), .A3(new_n901), .ZN(new_n902));
  NAND3_X1  g716(.A1(new_n885), .A2(new_n900), .A3(new_n902), .ZN(new_n903));
  NAND4_X1  g717(.A1(new_n846), .A2(new_n851), .A3(new_n899), .A4(new_n903), .ZN(new_n904));
  NAND2_X1  g718(.A1(new_n428), .A2(new_n208), .ZN(new_n905));
  NAND2_X1  g719(.A1(new_n904), .A2(new_n905), .ZN(new_n906));
  NOR4_X1   g720(.A1(new_n548), .A2(new_n765), .A3(new_n439), .A4(new_n302), .ZN(new_n907));
  XOR2_X1   g721(.A(new_n907), .B(KEYINPUT110), .Z(new_n908));
  XOR2_X1   g722(.A(new_n717), .B(KEYINPUT49), .Z(new_n909));
  OR4_X1    g723(.A1(new_n685), .A2(new_n908), .A3(new_n806), .A4(new_n909), .ZN(new_n910));
  NAND2_X1  g724(.A1(new_n906), .A2(new_n910), .ZN(G75));
  NOR2_X1   g725(.A1(new_n275), .A2(new_n277), .ZN(new_n912));
  AOI21_X1  g726(.A(new_n912), .B1(new_n275), .B2(new_n271), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(new_n211), .ZN(new_n914));
  XNOR2_X1  g728(.A(new_n914), .B(KEYINPUT55), .ZN(new_n915));
  INV_X1    g729(.A(G210), .ZN(new_n916));
  AOI211_X1 g730(.A(new_n916), .B(new_n377), .C1(new_n885), .C2(new_n902), .ZN(new_n917));
  OAI21_X1  g731(.A(new_n915), .B1(new_n917), .B2(KEYINPUT56), .ZN(new_n918));
  INV_X1    g732(.A(KEYINPUT56), .ZN(new_n919));
  INV_X1    g733(.A(new_n915), .ZN(new_n920));
  NAND2_X1  g734(.A1(new_n885), .A2(new_n902), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n921), .A2(G902), .ZN(new_n922));
  OAI211_X1 g736(.A(new_n919), .B(new_n920), .C1(new_n922), .C2(new_n916), .ZN(new_n923));
  NOR2_X1   g737(.A1(new_n208), .A2(G952), .ZN(new_n924));
  INV_X1    g738(.A(new_n924), .ZN(new_n925));
  AND3_X1   g739(.A1(new_n918), .A2(new_n923), .A3(new_n925), .ZN(G51));
  XNOR2_X1  g740(.A(new_n496), .B(KEYINPUT57), .ZN(new_n927));
  AND3_X1   g741(.A1(new_n885), .A2(new_n900), .A3(new_n902), .ZN(new_n928));
  AOI21_X1  g742(.A(new_n900), .B1(new_n885), .B2(new_n902), .ZN(new_n929));
  OAI21_X1  g743(.A(new_n927), .B1(new_n928), .B2(new_n929), .ZN(new_n930));
  NAND2_X1  g744(.A1(new_n930), .A2(new_n493), .ZN(new_n931));
  NAND4_X1  g745(.A1(new_n921), .A2(G902), .A3(new_n782), .A4(new_n781), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n924), .B1(new_n931), .B2(new_n932), .ZN(G54));
  NAND2_X1  g747(.A1(KEYINPUT58), .A2(G475), .ZN(new_n934));
  AOI211_X1 g748(.A(new_n377), .B(new_n934), .C1(new_n885), .C2(new_n902), .ZN(new_n935));
  OAI21_X1  g749(.A(KEYINPUT119), .B1(new_n935), .B2(new_n374), .ZN(new_n936));
  AOI21_X1  g750(.A(new_n924), .B1(new_n935), .B2(new_n374), .ZN(new_n937));
  INV_X1    g751(.A(KEYINPUT119), .ZN(new_n938));
  OAI211_X1 g752(.A(new_n938), .B(new_n365), .C1(new_n922), .C2(new_n934), .ZN(new_n939));
  AND3_X1   g753(.A1(new_n936), .A2(new_n937), .A3(new_n939), .ZN(G60));
  AND2_X1   g754(.A1(new_n619), .A2(new_n620), .ZN(new_n941));
  NAND2_X1  g755(.A1(new_n899), .A2(new_n903), .ZN(new_n942));
  XNOR2_X1  g756(.A(KEYINPUT120), .B(KEYINPUT59), .ZN(new_n943));
  XNOR2_X1  g757(.A(new_n943), .B(new_n614), .ZN(new_n944));
  AOI21_X1  g758(.A(new_n941), .B1(new_n942), .B2(new_n944), .ZN(new_n945));
  AND2_X1   g759(.A1(new_n941), .A2(new_n944), .ZN(new_n946));
  OAI21_X1  g760(.A(new_n946), .B1(new_n928), .B2(new_n929), .ZN(new_n947));
  NAND2_X1  g761(.A1(new_n947), .A2(new_n925), .ZN(new_n948));
  NOR2_X1   g762(.A1(new_n945), .A2(new_n948), .ZN(G63));
  XOR2_X1   g763(.A(KEYINPUT121), .B(KEYINPUT61), .Z(new_n950));
  NAND2_X1  g764(.A1(G217), .A2(G902), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n951), .B(KEYINPUT123), .ZN(new_n952));
  XNOR2_X1  g766(.A(KEYINPUT122), .B(KEYINPUT60), .ZN(new_n953));
  XOR2_X1   g767(.A(new_n952), .B(new_n953), .Z(new_n954));
  INV_X1    g768(.A(new_n954), .ZN(new_n955));
  AOI21_X1  g769(.A(new_n955), .B1(new_n885), .B2(new_n902), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n956), .A2(new_n652), .ZN(new_n957));
  INV_X1    g771(.A(new_n957), .ZN(new_n958));
  OAI21_X1  g772(.A(new_n925), .B1(new_n956), .B2(new_n538), .ZN(new_n959));
  OAI21_X1  g773(.A(new_n950), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND2_X1  g774(.A1(new_n921), .A2(new_n954), .ZN(new_n961));
  INV_X1    g775(.A(new_n538), .ZN(new_n962));
  NAND2_X1  g776(.A1(new_n961), .A2(new_n962), .ZN(new_n963));
  NAND4_X1  g777(.A1(new_n963), .A2(KEYINPUT61), .A3(new_n925), .A4(new_n957), .ZN(new_n964));
  NAND2_X1  g778(.A1(new_n960), .A2(new_n964), .ZN(G66));
  NAND2_X1  g779(.A1(new_n888), .A2(new_n864), .ZN(new_n966));
  NAND2_X1  g780(.A1(new_n966), .A2(new_n208), .ZN(new_n967));
  INV_X1    g781(.A(G224), .ZN(new_n968));
  OAI21_X1  g782(.A(G953), .B1(new_n431), .B2(new_n968), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n969), .B(KEYINPUT124), .Z(new_n970));
  NAND2_X1  g784(.A1(new_n967), .A2(new_n970), .ZN(new_n971));
  INV_X1    g785(.A(G898), .ZN(new_n972));
  AOI21_X1  g786(.A(new_n913), .B1(new_n972), .B2(G953), .ZN(new_n973));
  XOR2_X1   g787(.A(new_n971), .B(new_n973), .Z(G69));
  NOR2_X1   g788(.A1(new_n555), .A2(new_n556), .ZN(new_n975));
  XOR2_X1   g789(.A(new_n975), .B(KEYINPUT125), .Z(new_n976));
  XNOR2_X1  g790(.A(new_n976), .B(new_n358), .ZN(new_n977));
  AOI22_X1  g791(.A1(new_n775), .A2(new_n787), .B1(new_n793), .B2(new_n795), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n877), .A2(new_n698), .ZN(new_n979));
  NAND2_X1  g793(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n980));
  OR2_X1    g794(.A1(new_n979), .A2(KEYINPUT62), .ZN(new_n981));
  OR4_X1    g795(.A1(new_n833), .A2(new_n687), .A3(new_n861), .A4(new_n794), .ZN(new_n982));
  NAND4_X1  g796(.A1(new_n978), .A2(new_n980), .A3(new_n981), .A4(new_n982), .ZN(new_n983));
  AOI21_X1  g797(.A(new_n977), .B1(new_n983), .B2(new_n208), .ZN(new_n984));
  OAI21_X1  g798(.A(new_n977), .B1(new_n669), .B2(new_n208), .ZN(new_n985));
  AND2_X1   g799(.A1(new_n757), .A2(new_n760), .ZN(new_n986));
  NAND2_X1  g800(.A1(new_n604), .A2(new_n731), .ZN(new_n987));
  OR3_X1    g801(.A1(new_n786), .A2(new_n987), .A3(new_n776), .ZN(new_n988));
  AND2_X1   g802(.A1(new_n988), .A2(new_n877), .ZN(new_n989));
  AND4_X1   g803(.A1(new_n788), .A2(new_n796), .A3(new_n986), .A4(new_n989), .ZN(new_n990));
  AOI21_X1  g804(.A(new_n985), .B1(new_n990), .B2(new_n208), .ZN(new_n991));
  AOI21_X1  g805(.A(new_n208), .B1(G227), .B2(G900), .ZN(new_n992));
  OR3_X1    g806(.A1(new_n984), .A2(new_n991), .A3(new_n992), .ZN(new_n993));
  OAI21_X1  g807(.A(new_n992), .B1(new_n984), .B2(new_n991), .ZN(new_n994));
  NAND2_X1  g808(.A1(new_n993), .A2(new_n994), .ZN(G72));
  XNOR2_X1  g809(.A(KEYINPUT126), .B(KEYINPUT63), .ZN(new_n996));
  NOR2_X1   g810(.A1(new_n625), .A2(new_n377), .ZN(new_n997));
  XNOR2_X1  g811(.A(new_n996), .B(new_n997), .ZN(new_n998));
  OAI21_X1  g812(.A(new_n998), .B1(new_n983), .B2(new_n966), .ZN(new_n999));
  NAND2_X1  g813(.A1(new_n999), .A2(new_n680), .ZN(new_n1000));
  NAND2_X1  g814(.A1(new_n593), .A2(new_n564), .ZN(new_n1001));
  NAND3_X1  g815(.A1(new_n898), .A2(new_n998), .A3(new_n1001), .ZN(new_n1002));
  NAND4_X1  g816(.A1(new_n788), .A2(new_n796), .A3(new_n986), .A4(new_n989), .ZN(new_n1003));
  OAI21_X1  g817(.A(new_n998), .B1(new_n1003), .B2(new_n966), .ZN(new_n1004));
  NOR2_X1   g818(.A1(new_n592), .A2(new_n561), .ZN(new_n1005));
  NAND2_X1  g819(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1006));
  AND4_X1   g820(.A1(new_n925), .A2(new_n1000), .A3(new_n1002), .A4(new_n1006), .ZN(G57));
endmodule


