//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 1 1 0 1 0 0 1 1 1 0 0 0 1 1 0 1 1 0 0 0 0 0 0 0 0 1 1 0 1 1 0 1 1 0 0 0 0 1 0 1 1 0 1 1 0 0 0 0 0 1 0 1 0 0 1 1 0 0 0 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:51 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n693, new_n694, new_n695, new_n696, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n748, new_n749, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n760, new_n761,
    new_n762, new_n763, new_n764, new_n765, new_n766, new_n767, new_n768,
    new_n769, new_n770, new_n771, new_n772, new_n773, new_n774, new_n775,
    new_n776, new_n777, new_n778, new_n779, new_n781, new_n782, new_n783,
    new_n784, new_n786, new_n787, new_n788, new_n789, new_n790, new_n792,
    new_n793, new_n794, new_n795, new_n796, new_n797, new_n798, new_n799,
    new_n801, new_n803, new_n804, new_n805, new_n806, new_n807, new_n808,
    new_n809, new_n810, new_n811, new_n812, new_n813, new_n814, new_n815,
    new_n816, new_n818, new_n819, new_n820, new_n821, new_n822, new_n824,
    new_n825, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n857, new_n858, new_n859, new_n860, new_n861,
    new_n862, new_n863, new_n864, new_n865, new_n866, new_n867, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n884, new_n885, new_n887, new_n888, new_n890, new_n891, new_n892,
    new_n893, new_n894, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n913, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n930,
    new_n931, new_n932, new_n933, new_n935, new_n936, new_n937, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n960, new_n961, new_n962,
    new_n963, new_n964, new_n965, new_n967, new_n968, new_n969, new_n970,
    new_n972, new_n973, new_n974, new_n975, new_n976, new_n977, new_n979,
    new_n980, new_n981, new_n982, new_n983, new_n984, new_n985, new_n987,
    new_n988, new_n989, new_n990, new_n991, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999;
  XNOR2_X1  g000(.A(G113gat), .B(G141gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(G197gat), .ZN(new_n203));
  XOR2_X1   g002(.A(KEYINPUT11), .B(G169gat), .Z(new_n204));
  XNOR2_X1  g003(.A(new_n203), .B(new_n204), .ZN(new_n205));
  XOR2_X1   g004(.A(new_n205), .B(KEYINPUT12), .Z(new_n206));
  INV_X1    g005(.A(KEYINPUT94), .ZN(new_n207));
  OR2_X1    g006(.A1(G43gat), .A2(G50gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G43gat), .A2(G50gat), .ZN(new_n209));
  NAND2_X1  g008(.A1(new_n208), .A2(new_n209), .ZN(new_n210));
  NAND2_X1  g009(.A1(new_n210), .A2(KEYINPUT15), .ZN(new_n211));
  NAND2_X1  g010(.A1(G29gat), .A2(G36gat), .ZN(new_n212));
  INV_X1    g011(.A(KEYINPUT14), .ZN(new_n213));
  INV_X1    g012(.A(G29gat), .ZN(new_n214));
  INV_X1    g013(.A(G36gat), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n213), .A2(new_n214), .A3(new_n215), .ZN(new_n216));
  OAI21_X1  g015(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n217));
  NAND2_X1  g016(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND3_X1  g017(.A1(new_n211), .A2(new_n212), .A3(new_n218), .ZN(new_n219));
  AOI21_X1  g018(.A(KEYINPUT15), .B1(G43gat), .B2(G50gat), .ZN(new_n220));
  INV_X1    g019(.A(new_n220), .ZN(new_n221));
  XNOR2_X1  g020(.A(KEYINPUT93), .B(G50gat), .ZN(new_n222));
  INV_X1    g021(.A(G43gat), .ZN(new_n223));
  AOI21_X1  g022(.A(new_n221), .B1(new_n222), .B2(new_n223), .ZN(new_n224));
  NOR2_X1   g023(.A1(new_n219), .A2(new_n224), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT92), .ZN(new_n226));
  NAND2_X1  g025(.A1(new_n216), .A2(new_n226), .ZN(new_n227));
  NAND4_X1  g026(.A1(new_n213), .A2(new_n214), .A3(new_n215), .A4(KEYINPUT92), .ZN(new_n228));
  NAND3_X1  g027(.A1(new_n227), .A2(new_n228), .A3(new_n217), .ZN(new_n229));
  AOI21_X1  g028(.A(new_n211), .B1(new_n229), .B2(new_n212), .ZN(new_n230));
  OAI21_X1  g029(.A(new_n207), .B1(new_n225), .B2(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n229), .A2(new_n212), .ZN(new_n232));
  INV_X1    g031(.A(new_n211), .ZN(new_n233));
  NAND2_X1  g032(.A1(new_n232), .A2(new_n233), .ZN(new_n234));
  XOR2_X1   g033(.A(KEYINPUT93), .B(G50gat), .Z(new_n235));
  OAI21_X1  g034(.A(new_n220), .B1(new_n235), .B2(G43gat), .ZN(new_n236));
  NAND4_X1  g035(.A1(new_n236), .A2(new_n211), .A3(new_n212), .A4(new_n218), .ZN(new_n237));
  NAND3_X1  g036(.A1(new_n234), .A2(new_n237), .A3(KEYINPUT94), .ZN(new_n238));
  INV_X1    g037(.A(G8gat), .ZN(new_n239));
  XNOR2_X1  g038(.A(G15gat), .B(G22gat), .ZN(new_n240));
  INV_X1    g039(.A(KEYINPUT16), .ZN(new_n241));
  OAI21_X1  g040(.A(new_n240), .B1(new_n241), .B2(G1gat), .ZN(new_n242));
  AOI21_X1  g041(.A(new_n239), .B1(new_n242), .B2(KEYINPUT96), .ZN(new_n243));
  OAI21_X1  g042(.A(new_n242), .B1(G1gat), .B2(new_n240), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n243), .A2(new_n244), .ZN(new_n245));
  OAI221_X1 g044(.A(new_n242), .B1(KEYINPUT96), .B2(new_n239), .C1(G1gat), .C2(new_n240), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n231), .A2(new_n238), .A3(new_n247), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n248), .A2(KEYINPUT97), .ZN(new_n249));
  INV_X1    g048(.A(KEYINPUT97), .ZN(new_n250));
  NAND4_X1  g049(.A1(new_n231), .A2(new_n238), .A3(new_n247), .A4(new_n250), .ZN(new_n251));
  NAND2_X1  g050(.A1(new_n249), .A2(new_n251), .ZN(new_n252));
  NOR2_X1   g051(.A1(new_n225), .A2(new_n230), .ZN(new_n253));
  AOI21_X1  g052(.A(new_n247), .B1(new_n253), .B2(KEYINPUT17), .ZN(new_n254));
  XNOR2_X1  g053(.A(KEYINPUT95), .B(KEYINPUT17), .ZN(new_n255));
  INV_X1    g054(.A(new_n255), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n231), .A2(new_n238), .A3(new_n256), .ZN(new_n257));
  AOI22_X1  g056(.A1(new_n254), .A2(new_n257), .B1(G229gat), .B2(G233gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n252), .A2(new_n258), .A3(KEYINPUT18), .ZN(new_n259));
  NAND2_X1  g058(.A1(new_n231), .A2(new_n238), .ZN(new_n260));
  INV_X1    g059(.A(new_n247), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n260), .A2(new_n261), .ZN(new_n262));
  AND2_X1   g061(.A1(new_n252), .A2(new_n262), .ZN(new_n263));
  NAND2_X1  g062(.A1(G229gat), .A2(G233gat), .ZN(new_n264));
  XNOR2_X1  g063(.A(new_n264), .B(KEYINPUT13), .ZN(new_n265));
  OAI21_X1  g064(.A(new_n259), .B1(new_n263), .B2(new_n265), .ZN(new_n266));
  AOI21_X1  g065(.A(KEYINPUT18), .B1(new_n252), .B2(new_n258), .ZN(new_n267));
  OAI21_X1  g066(.A(new_n206), .B1(new_n266), .B2(new_n267), .ZN(new_n268));
  XNOR2_X1  g067(.A(new_n267), .B(KEYINPUT98), .ZN(new_n269));
  INV_X1    g068(.A(new_n206), .ZN(new_n270));
  OAI211_X1 g069(.A(new_n259), .B(new_n270), .C1(new_n263), .C2(new_n265), .ZN(new_n271));
  INV_X1    g070(.A(KEYINPUT99), .ZN(new_n272));
  NOR3_X1   g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  INV_X1    g072(.A(KEYINPUT98), .ZN(new_n274));
  XNOR2_X1  g073(.A(new_n267), .B(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(new_n259), .ZN(new_n276));
  AOI21_X1  g075(.A(new_n265), .B1(new_n252), .B2(new_n262), .ZN(new_n277));
  NOR3_X1   g076(.A1(new_n276), .A2(new_n277), .A3(new_n206), .ZN(new_n278));
  AOI21_X1  g077(.A(KEYINPUT99), .B1(new_n275), .B2(new_n278), .ZN(new_n279));
  OAI21_X1  g078(.A(new_n268), .B1(new_n273), .B2(new_n279), .ZN(new_n280));
  INV_X1    g079(.A(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(KEYINPUT40), .ZN(new_n282));
  XNOR2_X1  g081(.A(G127gat), .B(G134gat), .ZN(new_n283));
  INV_X1    g082(.A(KEYINPUT71), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n283), .A2(new_n284), .ZN(new_n285));
  INV_X1    g084(.A(KEYINPUT1), .ZN(new_n286));
  INV_X1    g085(.A(G113gat), .ZN(new_n287));
  NOR2_X1   g086(.A1(new_n287), .A2(G120gat), .ZN(new_n288));
  INV_X1    g087(.A(G120gat), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n289), .A2(G113gat), .ZN(new_n290));
  OAI21_X1  g089(.A(new_n286), .B1(new_n288), .B2(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(G127gat), .ZN(new_n292));
  NOR2_X1   g091(.A1(new_n292), .A2(G134gat), .ZN(new_n293));
  INV_X1    g092(.A(G134gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n294), .A2(G127gat), .ZN(new_n295));
  OAI21_X1  g094(.A(KEYINPUT71), .B1(new_n293), .B2(new_n295), .ZN(new_n296));
  NAND3_X1  g095(.A1(new_n285), .A2(new_n291), .A3(new_n296), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT72), .ZN(new_n298));
  OAI21_X1  g097(.A(new_n298), .B1(new_n287), .B2(G120gat), .ZN(new_n299));
  NAND3_X1  g098(.A1(new_n289), .A2(KEYINPUT72), .A3(G113gat), .ZN(new_n300));
  OAI211_X1 g099(.A(new_n299), .B(new_n300), .C1(G113gat), .C2(new_n289), .ZN(new_n301));
  XOR2_X1   g100(.A(KEYINPUT73), .B(KEYINPUT1), .Z(new_n302));
  NAND3_X1  g101(.A1(new_n301), .A2(new_n283), .A3(new_n302), .ZN(new_n303));
  AND2_X1   g102(.A1(new_n297), .A2(new_n303), .ZN(new_n304));
  AND2_X1   g103(.A1(G155gat), .A2(G162gat), .ZN(new_n305));
  NOR2_X1   g104(.A1(G155gat), .A2(G162gat), .ZN(new_n306));
  NOR2_X1   g105(.A1(new_n305), .A2(new_n306), .ZN(new_n307));
  INV_X1    g106(.A(new_n307), .ZN(new_n308));
  NAND2_X1  g107(.A1(G155gat), .A2(G162gat), .ZN(new_n309));
  NAND2_X1  g108(.A1(new_n309), .A2(KEYINPUT2), .ZN(new_n310));
  OR2_X1    g109(.A1(G141gat), .A2(G148gat), .ZN(new_n311));
  NAND2_X1  g110(.A1(G141gat), .A2(G148gat), .ZN(new_n312));
  NAND3_X1  g111(.A1(new_n310), .A2(new_n311), .A3(new_n312), .ZN(new_n313));
  NAND3_X1  g112(.A1(new_n311), .A2(KEYINPUT77), .A3(new_n312), .ZN(new_n314));
  NAND3_X1  g113(.A1(new_n308), .A2(new_n313), .A3(new_n314), .ZN(new_n315));
  AND2_X1   g114(.A1(G141gat), .A2(G148gat), .ZN(new_n316));
  NOR2_X1   g115(.A1(G141gat), .A2(G148gat), .ZN(new_n317));
  NOR2_X1   g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  OAI211_X1 g117(.A(new_n310), .B(new_n318), .C1(new_n307), .C2(KEYINPUT77), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(new_n304), .A2(new_n320), .ZN(new_n321));
  NAND2_X1  g120(.A1(G225gat), .A2(G233gat), .ZN(new_n322));
  AND2_X1   g121(.A1(new_n315), .A2(new_n319), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n297), .A2(new_n303), .ZN(new_n324));
  NAND2_X1  g123(.A1(new_n323), .A2(new_n324), .ZN(new_n325));
  NAND3_X1  g124(.A1(new_n321), .A2(new_n322), .A3(new_n325), .ZN(new_n326));
  OR2_X1    g125(.A1(new_n326), .A2(KEYINPUT84), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(KEYINPUT84), .ZN(new_n328));
  NAND3_X1  g127(.A1(new_n327), .A2(KEYINPUT39), .A3(new_n328), .ZN(new_n329));
  INV_X1    g128(.A(KEYINPUT85), .ZN(new_n330));
  OR2_X1    g129(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  INV_X1    g130(.A(KEYINPUT4), .ZN(new_n332));
  NAND3_X1  g131(.A1(new_n304), .A2(new_n332), .A3(new_n320), .ZN(new_n333));
  NAND2_X1  g132(.A1(new_n333), .A2(KEYINPUT82), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n321), .A2(KEYINPUT4), .ZN(new_n335));
  XNOR2_X1  g134(.A(new_n334), .B(new_n335), .ZN(new_n336));
  OAI21_X1  g135(.A(KEYINPUT78), .B1(new_n323), .B2(KEYINPUT3), .ZN(new_n337));
  INV_X1    g136(.A(KEYINPUT78), .ZN(new_n338));
  INV_X1    g137(.A(KEYINPUT3), .ZN(new_n339));
  NAND3_X1  g138(.A1(new_n320), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n337), .A2(new_n340), .ZN(new_n341));
  INV_X1    g140(.A(KEYINPUT79), .ZN(new_n342));
  NAND3_X1  g141(.A1(new_n315), .A2(new_n319), .A3(KEYINPUT3), .ZN(new_n343));
  NAND2_X1  g142(.A1(new_n324), .A2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n344), .ZN(new_n345));
  NAND3_X1  g144(.A1(new_n341), .A2(new_n342), .A3(new_n345), .ZN(new_n346));
  AOI21_X1  g145(.A(new_n338), .B1(new_n320), .B2(new_n339), .ZN(new_n347));
  AOI211_X1 g146(.A(KEYINPUT78), .B(KEYINPUT3), .C1(new_n315), .C2(new_n319), .ZN(new_n348));
  NOR2_X1   g147(.A1(new_n347), .A2(new_n348), .ZN(new_n349));
  OAI21_X1  g148(.A(KEYINPUT79), .B1(new_n349), .B2(new_n344), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n346), .A2(new_n350), .ZN(new_n351));
  NAND2_X1  g150(.A1(new_n336), .A2(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n322), .ZN(new_n353));
  NAND2_X1  g152(.A1(new_n352), .A2(new_n353), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n329), .A2(new_n330), .ZN(new_n355));
  NAND3_X1  g154(.A1(new_n331), .A2(new_n354), .A3(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357));
  XNOR2_X1  g156(.A(G57gat), .B(G85gat), .ZN(new_n358));
  XNOR2_X1  g157(.A(new_n357), .B(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(KEYINPUT81), .B(KEYINPUT0), .ZN(new_n360));
  XNOR2_X1  g159(.A(new_n359), .B(new_n360), .ZN(new_n361));
  OAI211_X1 g160(.A(new_n356), .B(new_n361), .C1(KEYINPUT39), .C2(new_n354), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT86), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n282), .B1(new_n362), .B2(new_n363), .ZN(new_n364));
  INV_X1    g163(.A(new_n361), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT5), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n321), .A2(new_n325), .ZN(new_n367));
  AOI21_X1  g166(.A(new_n366), .B1(new_n367), .B2(new_n353), .ZN(new_n368));
  INV_X1    g167(.A(new_n368), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n353), .B1(new_n335), .B2(new_n333), .ZN(new_n370));
  AOI21_X1  g169(.A(new_n342), .B1(new_n341), .B2(new_n345), .ZN(new_n371));
  NOR3_X1   g170(.A1(new_n349), .A2(KEYINPUT79), .A3(new_n344), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n370), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(KEYINPUT80), .ZN(new_n374));
  NAND2_X1  g173(.A1(new_n373), .A2(new_n374), .ZN(new_n375));
  NAND3_X1  g174(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n370), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n369), .B1(new_n375), .B2(new_n376), .ZN(new_n377));
  NAND2_X1  g176(.A1(new_n322), .A2(new_n366), .ZN(new_n378));
  NOR2_X1   g177(.A1(new_n352), .A2(new_n378), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n365), .B1(new_n377), .B2(new_n379), .ZN(new_n380));
  INV_X1    g179(.A(new_n380), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n364), .A2(new_n381), .ZN(new_n382));
  XNOR2_X1  g181(.A(G8gat), .B(G36gat), .ZN(new_n383));
  XNOR2_X1  g182(.A(G64gat), .B(G92gat), .ZN(new_n384));
  XOR2_X1   g183(.A(new_n383), .B(new_n384), .Z(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  XNOR2_X1  g185(.A(G197gat), .B(G204gat), .ZN(new_n387));
  INV_X1    g186(.A(G211gat), .ZN(new_n388));
  INV_X1    g187(.A(G218gat), .ZN(new_n389));
  NOR2_X1   g188(.A1(new_n388), .A2(new_n389), .ZN(new_n390));
  OAI21_X1  g189(.A(new_n387), .B1(KEYINPUT22), .B2(new_n390), .ZN(new_n391));
  XOR2_X1   g190(.A(G211gat), .B(G218gat), .Z(new_n392));
  XNOR2_X1  g191(.A(new_n391), .B(new_n392), .ZN(new_n393));
  NAND2_X1  g192(.A1(G183gat), .A2(G190gat), .ZN(new_n394));
  INV_X1    g193(.A(KEYINPUT24), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n394), .A2(new_n395), .ZN(new_n396));
  NAND3_X1  g195(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n396), .B(new_n397), .C1(G183gat), .C2(G190gat), .ZN(new_n398));
  INV_X1    g197(.A(G169gat), .ZN(new_n399));
  INV_X1    g198(.A(G176gat), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n399), .A2(new_n400), .A3(KEYINPUT23), .ZN(new_n401));
  NAND2_X1  g200(.A1(G169gat), .A2(G176gat), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT23), .ZN(new_n403));
  OAI21_X1  g202(.A(new_n403), .B1(G169gat), .B2(G176gat), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n398), .A2(new_n401), .A3(new_n402), .A4(new_n404), .ZN(new_n405));
  XOR2_X1   g204(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n406));
  NAND2_X1  g205(.A1(new_n405), .A2(new_n406), .ZN(new_n407));
  NOR2_X1   g206(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n408));
  INV_X1    g207(.A(new_n408), .ZN(new_n409));
  INV_X1    g208(.A(G183gat), .ZN(new_n410));
  NAND2_X1  g209(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n409), .A2(new_n410), .A3(new_n411), .ZN(new_n412));
  INV_X1    g211(.A(KEYINPUT65), .ZN(new_n413));
  OR2_X1    g212(.A1(new_n397), .A2(new_n413), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n397), .A2(new_n413), .ZN(new_n415));
  NAND4_X1  g214(.A1(new_n412), .A2(new_n414), .A3(new_n396), .A4(new_n415), .ZN(new_n416));
  AND4_X1   g215(.A1(KEYINPUT25), .A2(new_n401), .A3(new_n404), .A4(new_n402), .ZN(new_n417));
  NAND2_X1  g216(.A1(new_n416), .A2(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n407), .A2(new_n418), .ZN(new_n419));
  INV_X1    g218(.A(KEYINPUT28), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n410), .A2(KEYINPUT27), .ZN(new_n421));
  INV_X1    g220(.A(KEYINPUT27), .ZN(new_n422));
  NOR2_X1   g221(.A1(new_n422), .A2(G183gat), .ZN(new_n423));
  OAI21_X1  g222(.A(KEYINPUT68), .B1(new_n421), .B2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n422), .A2(G183gat), .ZN(new_n425));
  NAND2_X1  g224(.A1(new_n410), .A2(KEYINPUT27), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT68), .ZN(new_n427));
  NAND3_X1  g226(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  AND2_X1   g228(.A1(KEYINPUT66), .A2(G190gat), .ZN(new_n430));
  NOR2_X1   g229(.A1(new_n430), .A2(new_n408), .ZN(new_n431));
  AOI21_X1  g230(.A(new_n420), .B1(new_n429), .B2(new_n431), .ZN(new_n432));
  AOI21_X1  g231(.A(KEYINPUT28), .B1(new_n422), .B2(G183gat), .ZN(new_n433));
  INV_X1    g232(.A(KEYINPUT67), .ZN(new_n434));
  AOI21_X1  g233(.A(new_n434), .B1(KEYINPUT27), .B2(new_n410), .ZN(new_n435));
  NOR3_X1   g234(.A1(new_n422), .A2(KEYINPUT67), .A3(G183gat), .ZN(new_n436));
  OAI211_X1 g235(.A(new_n431), .B(new_n433), .C1(new_n435), .C2(new_n436), .ZN(new_n437));
  OAI21_X1  g236(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n438));
  INV_X1    g237(.A(KEYINPUT69), .ZN(new_n439));
  NAND2_X1  g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  OAI211_X1 g239(.A(KEYINPUT69), .B(KEYINPUT26), .C1(G169gat), .C2(G176gat), .ZN(new_n441));
  INV_X1    g240(.A(KEYINPUT26), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n442), .A2(new_n399), .A3(new_n400), .ZN(new_n443));
  NAND4_X1  g242(.A1(new_n440), .A2(new_n402), .A3(new_n441), .A4(new_n443), .ZN(new_n444));
  NAND3_X1  g243(.A1(new_n437), .A2(new_n394), .A3(new_n444), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT70), .ZN(new_n446));
  NOR3_X1   g245(.A1(new_n432), .A2(new_n445), .A3(new_n446), .ZN(new_n447));
  AND3_X1   g246(.A1(new_n437), .A2(new_n394), .A3(new_n444), .ZN(new_n448));
  AND3_X1   g247(.A1(new_n425), .A2(new_n426), .A3(new_n427), .ZN(new_n449));
  AOI21_X1  g248(.A(new_n427), .B1(new_n425), .B2(new_n426), .ZN(new_n450));
  OAI21_X1  g249(.A(new_n431), .B1(new_n449), .B2(new_n450), .ZN(new_n451));
  NAND2_X1  g250(.A1(new_n451), .A2(KEYINPUT28), .ZN(new_n452));
  AOI21_X1  g251(.A(KEYINPUT70), .B1(new_n448), .B2(new_n452), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n419), .B1(new_n447), .B2(new_n453), .ZN(new_n454));
  NAND2_X1  g253(.A1(new_n454), .A2(KEYINPUT75), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT29), .ZN(new_n456));
  OAI21_X1  g255(.A(new_n446), .B1(new_n432), .B2(new_n445), .ZN(new_n457));
  NAND3_X1  g256(.A1(new_n448), .A2(new_n452), .A3(KEYINPUT70), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(KEYINPUT75), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n459), .A2(new_n460), .A3(new_n419), .ZN(new_n461));
  NAND3_X1  g260(.A1(new_n455), .A2(new_n456), .A3(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(G226gat), .A2(G233gat), .ZN(new_n463));
  NAND2_X1  g262(.A1(new_n462), .A2(new_n463), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n419), .B1(new_n432), .B2(new_n445), .ZN(new_n465));
  INV_X1    g264(.A(new_n463), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  XOR2_X1   g266(.A(new_n467), .B(KEYINPUT76), .Z(new_n468));
  AOI21_X1  g267(.A(new_n393), .B1(new_n464), .B2(new_n468), .ZN(new_n469));
  INV_X1    g268(.A(new_n393), .ZN(new_n470));
  NAND2_X1  g269(.A1(new_n455), .A2(new_n461), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n471), .A2(new_n466), .ZN(new_n472));
  NAND3_X1  g271(.A1(new_n465), .A2(new_n456), .A3(new_n463), .ZN(new_n473));
  AOI21_X1  g272(.A(new_n470), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  OAI21_X1  g273(.A(new_n386), .B1(new_n469), .B2(new_n474), .ZN(new_n475));
  AOI21_X1  g274(.A(new_n463), .B1(new_n455), .B2(new_n461), .ZN(new_n476));
  INV_X1    g275(.A(new_n473), .ZN(new_n477));
  OAI21_X1  g276(.A(new_n393), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  XNOR2_X1  g277(.A(new_n467), .B(KEYINPUT76), .ZN(new_n479));
  AOI21_X1  g278(.A(new_n479), .B1(new_n463), .B2(new_n462), .ZN(new_n480));
  OAI211_X1 g279(.A(new_n385), .B(new_n478), .C1(new_n480), .C2(new_n393), .ZN(new_n481));
  NAND3_X1  g280(.A1(new_n475), .A2(KEYINPUT30), .A3(new_n481), .ZN(new_n482));
  NOR2_X1   g281(.A1(new_n469), .A2(new_n474), .ZN(new_n483));
  INV_X1    g282(.A(KEYINPUT30), .ZN(new_n484));
  NAND3_X1  g283(.A1(new_n483), .A2(new_n484), .A3(new_n385), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n482), .A2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n362), .A2(new_n363), .ZN(new_n488));
  OAI211_X1 g287(.A(new_n382), .B(new_n487), .C1(KEYINPUT40), .C2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT37), .ZN(new_n490));
  AOI21_X1  g289(.A(new_n385), .B1(new_n483), .B2(new_n490), .ZN(new_n491));
  INV_X1    g290(.A(new_n491), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n472), .A2(new_n473), .ZN(new_n493));
  AOI21_X1  g292(.A(new_n490), .B1(new_n493), .B2(new_n470), .ZN(new_n494));
  OAI21_X1  g293(.A(new_n494), .B1(new_n470), .B2(new_n480), .ZN(new_n495));
  XNOR2_X1  g294(.A(KEYINPUT87), .B(KEYINPUT38), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n495), .A2(new_n496), .ZN(new_n497));
  OAI21_X1  g296(.A(KEYINPUT88), .B1(new_n492), .B2(new_n497), .ZN(new_n498));
  INV_X1    g297(.A(new_n496), .ZN(new_n499));
  NOR2_X1   g298(.A1(new_n483), .A2(new_n490), .ZN(new_n500));
  OAI21_X1  g299(.A(new_n499), .B1(new_n492), .B2(new_n500), .ZN(new_n501));
  AND3_X1   g300(.A1(new_n351), .A2(KEYINPUT80), .A3(new_n370), .ZN(new_n502));
  AOI21_X1  g301(.A(KEYINPUT80), .B1(new_n351), .B2(new_n370), .ZN(new_n503));
  OAI21_X1  g302(.A(new_n368), .B1(new_n502), .B2(new_n503), .ZN(new_n504));
  OR2_X1    g303(.A1(new_n352), .A2(new_n378), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n504), .A2(new_n505), .A3(new_n361), .ZN(new_n506));
  INV_X1    g305(.A(KEYINPUT6), .ZN(new_n507));
  NAND3_X1  g306(.A1(new_n380), .A2(new_n506), .A3(new_n507), .ZN(new_n508));
  OAI211_X1 g307(.A(KEYINPUT6), .B(new_n365), .C1(new_n377), .C2(new_n379), .ZN(new_n509));
  AND3_X1   g308(.A1(new_n508), .A2(new_n509), .A3(new_n481), .ZN(new_n510));
  INV_X1    g309(.A(KEYINPUT88), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n491), .A2(new_n511), .A3(new_n496), .A4(new_n495), .ZN(new_n512));
  NAND4_X1  g311(.A1(new_n498), .A2(new_n501), .A3(new_n510), .A4(new_n512), .ZN(new_n513));
  NAND2_X1  g312(.A1(G228gat), .A2(G233gat), .ZN(new_n514));
  OAI21_X1  g313(.A(new_n470), .B1(new_n349), .B2(KEYINPUT29), .ZN(new_n515));
  AOI21_X1  g314(.A(new_n514), .B1(new_n515), .B2(KEYINPUT83), .ZN(new_n516));
  INV_X1    g315(.A(new_n516), .ZN(new_n517));
  OAI21_X1  g316(.A(new_n339), .B1(new_n470), .B2(KEYINPUT29), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n518), .A2(new_n323), .ZN(new_n519));
  NAND2_X1  g318(.A1(new_n515), .A2(new_n519), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n520), .A2(G22gat), .ZN(new_n521));
  INV_X1    g320(.A(G22gat), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n515), .A2(new_n519), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n517), .A2(new_n521), .A3(new_n523), .ZN(new_n524));
  XNOR2_X1  g323(.A(G78gat), .B(G106gat), .ZN(new_n525));
  XNOR2_X1  g324(.A(KEYINPUT31), .B(G50gat), .ZN(new_n526));
  XNOR2_X1  g325(.A(new_n525), .B(new_n526), .ZN(new_n527));
  AND3_X1   g326(.A1(new_n515), .A2(new_n522), .A3(new_n519), .ZN(new_n528));
  AOI21_X1  g327(.A(new_n522), .B1(new_n515), .B2(new_n519), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n516), .B1(new_n528), .B2(new_n529), .ZN(new_n530));
  AND3_X1   g329(.A1(new_n524), .A2(new_n527), .A3(new_n530), .ZN(new_n531));
  AOI21_X1  g330(.A(new_n527), .B1(new_n524), .B2(new_n530), .ZN(new_n532));
  NOR2_X1   g331(.A1(new_n531), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n489), .A2(new_n513), .A3(new_n533), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT36), .ZN(new_n535));
  NAND2_X1  g334(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n536));
  OR2_X1    g335(.A1(new_n535), .A2(KEYINPUT74), .ZN(new_n537));
  AOI21_X1  g336(.A(new_n324), .B1(new_n459), .B2(new_n419), .ZN(new_n538));
  AOI22_X1  g337(.A1(new_n405), .A2(new_n406), .B1(new_n416), .B2(new_n417), .ZN(new_n539));
  AOI211_X1 g338(.A(new_n304), .B(new_n539), .C1(new_n457), .C2(new_n458), .ZN(new_n540));
  NOR2_X1   g339(.A1(new_n538), .A2(new_n540), .ZN(new_n541));
  INV_X1    g340(.A(G227gat), .ZN(new_n542));
  INV_X1    g341(.A(G233gat), .ZN(new_n543));
  NOR2_X1   g342(.A1(new_n542), .A2(new_n543), .ZN(new_n544));
  OAI21_X1  g343(.A(KEYINPUT34), .B1(new_n541), .B2(new_n544), .ZN(new_n545));
  NAND2_X1  g344(.A1(new_n454), .A2(new_n304), .ZN(new_n546));
  NAND3_X1  g345(.A1(new_n459), .A2(new_n324), .A3(new_n419), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(KEYINPUT34), .ZN(new_n549));
  INV_X1    g348(.A(new_n544), .ZN(new_n550));
  NAND3_X1  g349(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  AOI21_X1  g350(.A(KEYINPUT33), .B1(new_n541), .B2(new_n544), .ZN(new_n552));
  XNOR2_X1  g351(.A(G15gat), .B(G43gat), .ZN(new_n553));
  XNOR2_X1  g352(.A(G71gat), .B(G99gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n553), .B(new_n554), .ZN(new_n555));
  OAI211_X1 g354(.A(new_n545), .B(new_n551), .C1(new_n552), .C2(new_n555), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n546), .A2(new_n544), .A3(new_n547), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n557), .A2(KEYINPUT32), .ZN(new_n558));
  INV_X1    g357(.A(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT33), .ZN(new_n560));
  AOI21_X1  g359(.A(new_n555), .B1(new_n557), .B2(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n562));
  AOI211_X1 g361(.A(KEYINPUT34), .B(new_n544), .C1(new_n546), .C2(new_n547), .ZN(new_n563));
  OAI21_X1  g362(.A(new_n561), .B1(new_n562), .B2(new_n563), .ZN(new_n564));
  AND3_X1   g363(.A1(new_n556), .A2(new_n559), .A3(new_n564), .ZN(new_n565));
  AOI21_X1  g364(.A(new_n559), .B1(new_n556), .B2(new_n564), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n536), .B(new_n537), .C1(new_n565), .C2(new_n566), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n556), .A2(new_n564), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n568), .A2(new_n558), .ZN(new_n569));
  NAND3_X1  g368(.A1(new_n556), .A2(new_n564), .A3(new_n559), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(KEYINPUT74), .A3(new_n535), .A4(new_n570), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n567), .A2(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n533), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n508), .A2(new_n509), .ZN(new_n574));
  NAND2_X1  g373(.A1(new_n574), .A2(new_n486), .ZN(new_n575));
  AOI21_X1  g374(.A(new_n572), .B1(new_n573), .B2(new_n575), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n534), .A2(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(KEYINPUT89), .ZN(new_n578));
  OAI21_X1  g377(.A(new_n578), .B1(new_n565), .B2(new_n566), .ZN(new_n579));
  NAND3_X1  g378(.A1(new_n569), .A2(KEYINPUT89), .A3(new_n570), .ZN(new_n580));
  AND2_X1   g379(.A1(new_n579), .A2(new_n580), .ZN(new_n581));
  AOI22_X1  g380(.A1(new_n509), .A2(new_n508), .B1(new_n482), .B2(new_n485), .ZN(new_n582));
  NOR3_X1   g381(.A1(new_n531), .A2(new_n532), .A3(KEYINPUT35), .ZN(new_n583));
  NAND4_X1  g382(.A1(new_n581), .A2(KEYINPUT90), .A3(new_n582), .A4(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(KEYINPUT90), .ZN(new_n585));
  NAND3_X1  g384(.A1(new_n579), .A2(new_n580), .A3(new_n583), .ZN(new_n586));
  OAI21_X1  g385(.A(new_n585), .B1(new_n586), .B2(new_n575), .ZN(new_n587));
  NAND2_X1  g386(.A1(new_n584), .A2(new_n587), .ZN(new_n588));
  NAND3_X1  g387(.A1(new_n569), .A2(new_n533), .A3(new_n570), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n589), .A2(KEYINPUT91), .ZN(new_n590));
  INV_X1    g389(.A(KEYINPUT91), .ZN(new_n591));
  NAND4_X1  g390(.A1(new_n569), .A2(new_n533), .A3(new_n591), .A4(new_n570), .ZN(new_n592));
  NAND3_X1  g391(.A1(new_n582), .A2(new_n590), .A3(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n593), .A2(KEYINPUT35), .ZN(new_n594));
  NAND2_X1  g393(.A1(new_n588), .A2(new_n594), .ZN(new_n595));
  AOI21_X1  g394(.A(new_n281), .B1(new_n577), .B2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(G57gat), .ZN(new_n597));
  NOR2_X1   g396(.A1(new_n597), .A2(KEYINPUT100), .ZN(new_n598));
  INV_X1    g397(.A(G64gat), .ZN(new_n599));
  XNOR2_X1  g398(.A(new_n598), .B(new_n599), .ZN(new_n600));
  NAND2_X1  g399(.A1(G71gat), .A2(G78gat), .ZN(new_n601));
  OR2_X1    g400(.A1(G71gat), .A2(G78gat), .ZN(new_n602));
  INV_X1    g401(.A(KEYINPUT9), .ZN(new_n603));
  OAI21_X1  g402(.A(new_n601), .B1(new_n602), .B2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n600), .A2(new_n604), .ZN(new_n605));
  NOR2_X1   g404(.A1(new_n597), .A2(new_n599), .ZN(new_n606));
  OAI21_X1  g405(.A(KEYINPUT9), .B1(G57gat), .B2(G64gat), .ZN(new_n607));
  OAI211_X1 g406(.A(new_n601), .B(new_n602), .C1(new_n606), .C2(new_n607), .ZN(new_n608));
  NAND2_X1  g407(.A1(new_n605), .A2(new_n608), .ZN(new_n609));
  INV_X1    g408(.A(KEYINPUT21), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n609), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(G231gat), .A2(G233gat), .ZN(new_n612));
  XNOR2_X1  g411(.A(new_n611), .B(new_n612), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(G127gat), .ZN(new_n614));
  XNOR2_X1  g413(.A(G183gat), .B(G211gat), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n614), .B(new_n615), .ZN(new_n616));
  OAI21_X1  g415(.A(new_n261), .B1(new_n610), .B2(new_n609), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT101), .ZN(new_n618));
  XNOR2_X1  g417(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n619), .B(G155gat), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n618), .B(new_n620), .ZN(new_n621));
  OR2_X1    g420(.A1(new_n616), .A2(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n616), .A2(new_n621), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  XOR2_X1   g423(.A(G190gat), .B(G218gat), .Z(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(KEYINPUT104), .ZN(new_n626));
  AOI21_X1  g425(.A(KEYINPUT41), .B1(G232gat), .B2(G233gat), .ZN(new_n627));
  XNOR2_X1  g426(.A(new_n626), .B(new_n627), .ZN(new_n628));
  INV_X1    g427(.A(new_n628), .ZN(new_n629));
  NAND3_X1  g428(.A1(KEYINPUT41), .A2(G232gat), .A3(G233gat), .ZN(new_n630));
  XNOR2_X1  g429(.A(KEYINPUT102), .B(G85gat), .ZN(new_n631));
  INV_X1    g430(.A(G92gat), .ZN(new_n632));
  NAND2_X1  g431(.A1(new_n631), .A2(new_n632), .ZN(new_n633));
  NAND2_X1  g432(.A1(G85gat), .A2(G92gat), .ZN(new_n634));
  XNOR2_X1  g433(.A(new_n634), .B(KEYINPUT7), .ZN(new_n635));
  INV_X1    g434(.A(G99gat), .ZN(new_n636));
  INV_X1    g435(.A(G106gat), .ZN(new_n637));
  OAI21_X1  g436(.A(KEYINPUT8), .B1(new_n636), .B2(new_n637), .ZN(new_n638));
  NAND3_X1  g437(.A1(new_n633), .A2(new_n635), .A3(new_n638), .ZN(new_n639));
  XOR2_X1   g438(.A(G99gat), .B(G106gat), .Z(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n640), .ZN(new_n642));
  NAND4_X1  g441(.A1(new_n642), .A2(new_n633), .A3(new_n635), .A4(new_n638), .ZN(new_n643));
  NAND3_X1  g442(.A1(new_n641), .A2(KEYINPUT103), .A3(new_n643), .ZN(new_n644));
  OR3_X1    g443(.A1(new_n639), .A2(KEYINPUT103), .A3(new_n640), .ZN(new_n645));
  AND2_X1   g444(.A1(new_n644), .A2(new_n645), .ZN(new_n646));
  OAI21_X1  g445(.A(new_n630), .B1(new_n646), .B2(new_n260), .ZN(new_n647));
  INV_X1    g446(.A(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n644), .A2(new_n645), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n649), .B1(KEYINPUT17), .B2(new_n253), .ZN(new_n650));
  NAND2_X1  g449(.A1(new_n650), .A2(new_n257), .ZN(new_n651));
  XNOR2_X1  g450(.A(G134gat), .B(G162gat), .ZN(new_n652));
  INV_X1    g451(.A(new_n652), .ZN(new_n653));
  NAND3_X1  g452(.A1(new_n648), .A2(new_n651), .A3(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(new_n654), .ZN(new_n655));
  AOI21_X1  g454(.A(new_n653), .B1(new_n648), .B2(new_n651), .ZN(new_n656));
  OAI21_X1  g455(.A(new_n629), .B1(new_n655), .B2(new_n656), .ZN(new_n657));
  INV_X1    g456(.A(new_n656), .ZN(new_n658));
  NAND3_X1  g457(.A1(new_n658), .A2(new_n628), .A3(new_n654), .ZN(new_n659));
  NAND2_X1  g458(.A1(new_n657), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(new_n660), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n624), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(KEYINPUT105), .ZN(new_n663));
  XNOR2_X1  g462(.A(new_n662), .B(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(G230gat), .A2(G233gat), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n644), .A2(new_n645), .A3(new_n609), .ZN(new_n667));
  INV_X1    g466(.A(new_n609), .ZN(new_n668));
  NAND3_X1  g467(.A1(new_n668), .A2(new_n643), .A3(new_n641), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT10), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n667), .A2(new_n669), .A3(new_n670), .ZN(new_n671));
  NAND3_X1  g470(.A1(new_n649), .A2(KEYINPUT10), .A3(new_n668), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n666), .B1(new_n671), .B2(new_n672), .ZN(new_n673));
  INV_X1    g472(.A(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n667), .A2(new_n669), .ZN(new_n675));
  NAND2_X1  g474(.A1(new_n675), .A2(new_n666), .ZN(new_n676));
  XOR2_X1   g475(.A(G120gat), .B(G148gat), .Z(new_n677));
  XNOR2_X1  g476(.A(new_n677), .B(KEYINPUT106), .ZN(new_n678));
  XNOR2_X1  g477(.A(G176gat), .B(G204gat), .ZN(new_n679));
  XNOR2_X1  g478(.A(new_n678), .B(new_n679), .ZN(new_n680));
  AND3_X1   g479(.A1(new_n674), .A2(new_n676), .A3(new_n680), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n680), .B1(new_n674), .B2(new_n676), .ZN(new_n682));
  NOR2_X1   g481(.A1(new_n681), .A2(new_n682), .ZN(new_n683));
  AND2_X1   g482(.A1(new_n664), .A2(new_n683), .ZN(new_n684));
  NAND2_X1  g483(.A1(new_n596), .A2(new_n684), .ZN(new_n685));
  NAND2_X1  g484(.A1(new_n685), .A2(KEYINPUT107), .ZN(new_n686));
  INV_X1    g485(.A(KEYINPUT107), .ZN(new_n687));
  NAND3_X1  g486(.A1(new_n596), .A2(new_n687), .A3(new_n684), .ZN(new_n688));
  NAND2_X1  g487(.A1(new_n686), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n574), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n689), .A2(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G1gat), .ZN(G1324gat));
  AOI21_X1  g491(.A(new_n239), .B1(new_n689), .B2(new_n487), .ZN(new_n693));
  XNOR2_X1  g492(.A(KEYINPUT16), .B(G8gat), .ZN(new_n694));
  AOI211_X1 g493(.A(new_n486), .B(new_n694), .C1(new_n686), .C2(new_n688), .ZN(new_n695));
  OAI21_X1  g494(.A(KEYINPUT42), .B1(new_n693), .B2(new_n695), .ZN(new_n696));
  OAI21_X1  g495(.A(new_n696), .B1(KEYINPUT42), .B2(new_n695), .ZN(G1325gat));
  INV_X1    g496(.A(G15gat), .ZN(new_n698));
  NAND3_X1  g497(.A1(new_n689), .A2(new_n698), .A3(new_n581), .ZN(new_n699));
  INV_X1    g498(.A(new_n699), .ZN(new_n700));
  AOI21_X1  g499(.A(new_n698), .B1(new_n689), .B2(new_n572), .ZN(new_n701));
  OAI21_X1  g500(.A(KEYINPUT108), .B1(new_n700), .B2(new_n701), .ZN(new_n702));
  INV_X1    g501(.A(new_n701), .ZN(new_n703));
  INV_X1    g502(.A(KEYINPUT108), .ZN(new_n704));
  NAND3_X1  g503(.A1(new_n703), .A2(new_n704), .A3(new_n699), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n702), .A2(new_n705), .ZN(G1326gat));
  INV_X1    g505(.A(new_n688), .ZN(new_n707));
  AOI21_X1  g506(.A(new_n687), .B1(new_n596), .B2(new_n684), .ZN(new_n708));
  OAI21_X1  g507(.A(new_n573), .B1(new_n707), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n709), .A2(KEYINPUT109), .ZN(new_n710));
  INV_X1    g509(.A(KEYINPUT109), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n689), .A2(new_n711), .A3(new_n573), .ZN(new_n712));
  XNOR2_X1  g511(.A(KEYINPUT43), .B(G22gat), .ZN(new_n713));
  AND3_X1   g512(.A1(new_n710), .A2(new_n712), .A3(new_n713), .ZN(new_n714));
  AOI21_X1  g513(.A(new_n713), .B1(new_n710), .B2(new_n712), .ZN(new_n715));
  NOR2_X1   g514(.A1(new_n714), .A2(new_n715), .ZN(G1327gat));
  INV_X1    g515(.A(new_n624), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n717), .A2(new_n660), .A3(new_n683), .ZN(new_n718));
  INV_X1    g517(.A(new_n718), .ZN(new_n719));
  NAND2_X1  g518(.A1(new_n596), .A2(new_n719), .ZN(new_n720));
  NOR3_X1   g519(.A1(new_n720), .A2(G29gat), .A3(new_n574), .ZN(new_n721));
  XNOR2_X1  g520(.A(KEYINPUT110), .B(KEYINPUT45), .ZN(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  XNOR2_X1  g522(.A(new_n624), .B(KEYINPUT111), .ZN(new_n724));
  INV_X1    g523(.A(new_n724), .ZN(new_n725));
  INV_X1    g524(.A(new_n683), .ZN(new_n726));
  NOR3_X1   g525(.A1(new_n725), .A2(new_n281), .A3(new_n726), .ZN(new_n727));
  XNOR2_X1  g526(.A(new_n727), .B(KEYINPUT112), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT113), .ZN(new_n729));
  AOI221_X4 g528(.A(new_n729), .B1(new_n593), .B2(KEYINPUT35), .C1(new_n584), .C2(new_n587), .ZN(new_n730));
  AOI21_X1  g529(.A(KEYINPUT113), .B1(new_n588), .B2(new_n594), .ZN(new_n731));
  OAI21_X1  g530(.A(new_n577), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g531(.A1(new_n661), .A2(KEYINPUT44), .ZN(new_n733));
  NAND2_X1  g532(.A1(new_n732), .A2(new_n733), .ZN(new_n734));
  INV_X1    g533(.A(new_n576), .ZN(new_n735));
  NOR2_X1   g534(.A1(new_n488), .A2(KEYINPUT40), .ZN(new_n736));
  NOR3_X1   g535(.A1(new_n736), .A2(new_n364), .A3(new_n381), .ZN(new_n737));
  AOI21_X1  g536(.A(new_n573), .B1(new_n737), .B2(new_n487), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n735), .B1(new_n738), .B2(new_n513), .ZN(new_n739));
  AOI22_X1  g538(.A1(new_n584), .A2(new_n587), .B1(KEYINPUT35), .B2(new_n593), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n660), .B1(new_n739), .B2(new_n740), .ZN(new_n741));
  NAND2_X1  g540(.A1(new_n741), .A2(KEYINPUT44), .ZN(new_n742));
  AOI21_X1  g541(.A(new_n728), .B1(new_n734), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(G29gat), .B1(new_n744), .B2(new_n574), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n723), .A2(new_n745), .ZN(G1328gat));
  NOR3_X1   g545(.A1(new_n720), .A2(G36gat), .A3(new_n486), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n747), .B(KEYINPUT46), .ZN(new_n748));
  OAI21_X1  g547(.A(G36gat), .B1(new_n744), .B2(new_n486), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(G1329gat));
  XNOR2_X1  g549(.A(KEYINPUT114), .B(KEYINPUT47), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n743), .A2(new_n572), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n752), .A2(G43gat), .ZN(new_n753));
  NAND4_X1  g552(.A1(new_n596), .A2(new_n223), .A3(new_n581), .A4(new_n719), .ZN(new_n754));
  AOI21_X1  g553(.A(new_n751), .B1(new_n753), .B2(new_n754), .ZN(new_n755));
  INV_X1    g554(.A(new_n754), .ZN(new_n756));
  INV_X1    g555(.A(new_n751), .ZN(new_n757));
  AOI211_X1 g556(.A(new_n756), .B(new_n757), .C1(new_n752), .C2(G43gat), .ZN(new_n758));
  NOR2_X1   g557(.A1(new_n755), .A2(new_n758), .ZN(G1330gat));
  INV_X1    g558(.A(new_n728), .ZN(new_n760));
  INV_X1    g559(.A(new_n733), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n595), .A2(new_n729), .ZN(new_n762));
  NAND2_X1  g561(.A1(new_n740), .A2(KEYINPUT113), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n761), .B1(new_n764), .B2(new_n577), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT44), .ZN(new_n766));
  NAND2_X1  g565(.A1(new_n577), .A2(new_n595), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n766), .B1(new_n767), .B2(new_n660), .ZN(new_n768));
  OAI211_X1 g567(.A(new_n573), .B(new_n760), .C1(new_n765), .C2(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT115), .ZN(new_n770));
  NAND2_X1  g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  NAND3_X1  g570(.A1(new_n743), .A2(KEYINPUT115), .A3(new_n573), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n771), .A2(new_n235), .A3(new_n772), .ZN(new_n773));
  NOR3_X1   g572(.A1(new_n720), .A2(new_n533), .A3(new_n235), .ZN(new_n774));
  INV_X1    g573(.A(KEYINPUT48), .ZN(new_n775));
  NOR2_X1   g574(.A1(new_n774), .A2(new_n775), .ZN(new_n776));
  NAND2_X1  g575(.A1(new_n773), .A2(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n222), .B1(new_n743), .B2(new_n573), .ZN(new_n778));
  OAI21_X1  g577(.A(new_n775), .B1(new_n778), .B2(new_n774), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n777), .A2(new_n779), .ZN(G1331gat));
  AOI21_X1  g579(.A(new_n739), .B1(new_n762), .B2(new_n763), .ZN(new_n781));
  NAND3_X1  g580(.A1(new_n664), .A2(new_n281), .A3(new_n726), .ZN(new_n782));
  NOR2_X1   g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND2_X1  g582(.A1(new_n783), .A2(new_n690), .ZN(new_n784));
  XNOR2_X1  g583(.A(new_n784), .B(G57gat), .ZN(G1332gat));
  INV_X1    g584(.A(new_n783), .ZN(new_n786));
  NOR2_X1   g585(.A1(new_n786), .A2(new_n486), .ZN(new_n787));
  NOR2_X1   g586(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n788));
  AND2_X1   g587(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n789));
  OAI21_X1  g588(.A(new_n787), .B1(new_n788), .B2(new_n789), .ZN(new_n790));
  OAI21_X1  g589(.A(new_n790), .B1(new_n787), .B2(new_n788), .ZN(G1333gat));
  INV_X1    g590(.A(G71gat), .ZN(new_n792));
  NAND3_X1  g591(.A1(new_n783), .A2(new_n792), .A3(new_n581), .ZN(new_n793));
  INV_X1    g592(.A(new_n572), .ZN(new_n794));
  NOR2_X1   g593(.A1(new_n786), .A2(new_n794), .ZN(new_n795));
  OAI21_X1  g594(.A(new_n793), .B1(new_n795), .B2(new_n792), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT50), .ZN(new_n797));
  NAND2_X1  g596(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  OAI211_X1 g597(.A(KEYINPUT50), .B(new_n793), .C1(new_n795), .C2(new_n792), .ZN(new_n799));
  NAND2_X1  g598(.A1(new_n798), .A2(new_n799), .ZN(G1334gat));
  NAND2_X1  g599(.A1(new_n783), .A2(new_n573), .ZN(new_n801));
  XNOR2_X1  g600(.A(new_n801), .B(G78gat), .ZN(G1335gat));
  INV_X1    g601(.A(KEYINPUT51), .ZN(new_n803));
  NOR2_X1   g602(.A1(new_n280), .A2(new_n624), .ZN(new_n804));
  INV_X1    g603(.A(new_n804), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n805), .A2(new_n661), .ZN(new_n806));
  INV_X1    g605(.A(new_n806), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n803), .B1(new_n781), .B2(new_n807), .ZN(new_n808));
  NAND3_X1  g607(.A1(new_n732), .A2(KEYINPUT51), .A3(new_n806), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND4_X1  g609(.A1(new_n810), .A2(new_n690), .A3(new_n631), .A4(new_n726), .ZN(new_n811));
  NOR2_X1   g610(.A1(new_n805), .A2(new_n683), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  AOI21_X1  g612(.A(new_n813), .B1(new_n734), .B2(new_n742), .ZN(new_n814));
  INV_X1    g613(.A(new_n814), .ZN(new_n815));
  NOR2_X1   g614(.A1(new_n815), .A2(new_n574), .ZN(new_n816));
  OAI21_X1  g615(.A(new_n811), .B1(new_n816), .B2(new_n631), .ZN(G1336gat));
  AOI21_X1  g616(.A(new_n632), .B1(new_n814), .B2(new_n487), .ZN(new_n818));
  NAND3_X1  g617(.A1(new_n487), .A2(new_n632), .A3(new_n726), .ZN(new_n819));
  AOI21_X1  g618(.A(new_n819), .B1(new_n808), .B2(new_n809), .ZN(new_n820));
  OR3_X1    g619(.A1(new_n818), .A2(KEYINPUT52), .A3(new_n820), .ZN(new_n821));
  OAI21_X1  g620(.A(KEYINPUT52), .B1(new_n818), .B2(new_n820), .ZN(new_n822));
  NAND2_X1  g621(.A1(new_n821), .A2(new_n822), .ZN(G1337gat));
  OAI21_X1  g622(.A(G99gat), .B1(new_n815), .B2(new_n794), .ZN(new_n824));
  NAND4_X1  g623(.A1(new_n810), .A2(new_n636), .A3(new_n581), .A4(new_n726), .ZN(new_n825));
  NAND2_X1  g624(.A1(new_n824), .A2(new_n825), .ZN(G1338gat));
  INV_X1    g625(.A(KEYINPUT116), .ZN(new_n827));
  OR2_X1    g626(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n827), .A2(KEYINPUT53), .ZN(new_n829));
  AOI21_X1  g628(.A(new_n637), .B1(new_n814), .B2(new_n573), .ZN(new_n830));
  NOR3_X1   g629(.A1(new_n533), .A2(G106gat), .A3(new_n683), .ZN(new_n831));
  INV_X1    g630(.A(new_n831), .ZN(new_n832));
  AOI21_X1  g631(.A(new_n832), .B1(new_n808), .B2(new_n809), .ZN(new_n833));
  OAI211_X1 g632(.A(new_n828), .B(new_n829), .C1(new_n830), .C2(new_n833), .ZN(new_n834));
  OAI211_X1 g633(.A(new_n573), .B(new_n812), .C1(new_n765), .C2(new_n768), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n835), .A2(G106gat), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n810), .A2(new_n831), .ZN(new_n837));
  NAND4_X1  g636(.A1(new_n836), .A2(new_n837), .A3(new_n827), .A4(KEYINPUT53), .ZN(new_n838));
  AND2_X1   g637(.A1(new_n834), .A2(new_n838), .ZN(G1339gat));
  NAND2_X1  g638(.A1(new_n684), .A2(new_n281), .ZN(new_n840));
  AOI22_X1  g639(.A1(new_n249), .A2(new_n251), .B1(new_n257), .B2(new_n254), .ZN(new_n841));
  INV_X1    g640(.A(KEYINPUT117), .ZN(new_n842));
  OR3_X1    g641(.A1(new_n841), .A2(new_n842), .A3(new_n264), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n263), .A2(new_n265), .ZN(new_n844));
  OAI21_X1  g643(.A(new_n842), .B1(new_n841), .B2(new_n264), .ZN(new_n845));
  NAND3_X1  g644(.A1(new_n843), .A2(new_n844), .A3(new_n845), .ZN(new_n846));
  AOI22_X1  g645(.A1(new_n846), .A2(new_n205), .B1(new_n657), .B2(new_n659), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n671), .A2(new_n666), .A3(new_n672), .ZN(new_n848));
  NAND3_X1  g647(.A1(new_n674), .A2(KEYINPUT54), .A3(new_n848), .ZN(new_n849));
  INV_X1    g648(.A(KEYINPUT54), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n680), .B1(new_n673), .B2(new_n850), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n849), .A2(KEYINPUT55), .A3(new_n851), .ZN(new_n852));
  AOI21_X1  g651(.A(KEYINPUT55), .B1(new_n849), .B2(new_n851), .ZN(new_n853));
  NOR3_X1   g652(.A1(new_n852), .A2(new_n853), .A3(new_n681), .ZN(new_n854));
  OAI211_X1 g653(.A(new_n847), .B(new_n854), .C1(new_n273), .C2(new_n279), .ZN(new_n855));
  NAND2_X1  g654(.A1(new_n855), .A2(KEYINPUT118), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n272), .B1(new_n269), .B2(new_n271), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n275), .A2(KEYINPUT99), .A3(new_n278), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n857), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT118), .ZN(new_n860));
  NAND4_X1  g659(.A1(new_n859), .A2(new_n860), .A3(new_n854), .A4(new_n847), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n856), .A2(new_n861), .ZN(new_n862));
  NAND2_X1  g661(.A1(new_n846), .A2(new_n205), .ZN(new_n863));
  OAI211_X1 g662(.A(new_n726), .B(new_n863), .C1(new_n273), .C2(new_n279), .ZN(new_n864));
  NAND2_X1  g663(.A1(new_n864), .A2(KEYINPUT119), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT119), .ZN(new_n866));
  NAND4_X1  g665(.A1(new_n859), .A2(new_n866), .A3(new_n726), .A4(new_n863), .ZN(new_n867));
  NAND2_X1  g666(.A1(new_n280), .A2(new_n854), .ZN(new_n868));
  NAND3_X1  g667(.A1(new_n865), .A2(new_n867), .A3(new_n868), .ZN(new_n869));
  AOI21_X1  g668(.A(new_n862), .B1(new_n869), .B2(new_n661), .ZN(new_n870));
  OAI21_X1  g669(.A(new_n724), .B1(new_n870), .B2(KEYINPUT120), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT120), .ZN(new_n872));
  AOI211_X1 g671(.A(new_n872), .B(new_n862), .C1(new_n661), .C2(new_n869), .ZN(new_n873));
  OAI21_X1  g672(.A(new_n840), .B1(new_n871), .B2(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n690), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n590), .A2(new_n486), .A3(new_n592), .ZN(new_n876));
  AND2_X1   g675(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  AOI21_X1  g676(.A(G113gat), .B1(new_n877), .B2(new_n280), .ZN(new_n878));
  AND2_X1   g677(.A1(new_n874), .A2(new_n533), .ZN(new_n879));
  NOR2_X1   g678(.A1(new_n487), .A2(new_n574), .ZN(new_n880));
  AND3_X1   g679(.A1(new_n879), .A2(new_n581), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g680(.A1(new_n281), .A2(new_n287), .ZN(new_n882));
  AOI21_X1  g681(.A(new_n878), .B1(new_n881), .B2(new_n882), .ZN(G1340gat));
  AOI21_X1  g682(.A(G120gat), .B1(new_n877), .B2(new_n726), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n683), .A2(new_n289), .ZN(new_n885));
  AOI21_X1  g684(.A(new_n884), .B1(new_n881), .B2(new_n885), .ZN(G1341gat));
  NAND3_X1  g685(.A1(new_n877), .A2(new_n292), .A3(new_n624), .ZN(new_n887));
  AND2_X1   g686(.A1(new_n881), .A2(new_n725), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n887), .B1(new_n888), .B2(new_n292), .ZN(G1342gat));
  NAND3_X1  g688(.A1(new_n877), .A2(new_n294), .A3(new_n660), .ZN(new_n890));
  NAND2_X1  g689(.A1(new_n890), .A2(KEYINPUT56), .ZN(new_n891));
  INV_X1    g690(.A(KEYINPUT56), .ZN(new_n892));
  NAND4_X1  g691(.A1(new_n877), .A2(new_n892), .A3(new_n294), .A4(new_n660), .ZN(new_n893));
  AND2_X1   g692(.A1(new_n881), .A2(new_n660), .ZN(new_n894));
  OAI211_X1 g693(.A(new_n891), .B(new_n893), .C1(new_n294), .C2(new_n894), .ZN(G1343gat));
  NOR3_X1   g694(.A1(new_n572), .A2(new_n574), .A3(new_n487), .ZN(new_n896));
  XOR2_X1   g695(.A(KEYINPUT121), .B(KEYINPUT57), .Z(new_n897));
  INV_X1    g696(.A(new_n897), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n898), .B1(new_n874), .B2(new_n573), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT57), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n660), .B1(new_n868), .B2(new_n864), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n717), .B1(new_n901), .B2(new_n862), .ZN(new_n902));
  AOI211_X1 g701(.A(new_n900), .B(new_n533), .C1(new_n840), .C2(new_n902), .ZN(new_n903));
  OAI211_X1 g702(.A(new_n280), .B(new_n896), .C1(new_n899), .C2(new_n903), .ZN(new_n904));
  NAND2_X1  g703(.A1(new_n904), .A2(G141gat), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n794), .A2(new_n573), .ZN(new_n906));
  NOR2_X1   g705(.A1(new_n906), .A2(new_n487), .ZN(new_n907));
  NOR2_X1   g706(.A1(new_n281), .A2(G141gat), .ZN(new_n908));
  NAND3_X1  g707(.A1(new_n875), .A2(new_n907), .A3(new_n908), .ZN(new_n909));
  NAND2_X1  g708(.A1(new_n905), .A2(new_n909), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n910), .A2(KEYINPUT58), .ZN(new_n911));
  INV_X1    g710(.A(KEYINPUT58), .ZN(new_n912));
  NAND3_X1  g711(.A1(new_n905), .A2(new_n912), .A3(new_n909), .ZN(new_n913));
  NAND2_X1  g712(.A1(new_n911), .A2(new_n913), .ZN(G1344gat));
  AND2_X1   g713(.A1(new_n875), .A2(new_n907), .ZN(new_n915));
  INV_X1    g714(.A(G148gat), .ZN(new_n916));
  NAND3_X1  g715(.A1(new_n915), .A2(new_n916), .A3(new_n726), .ZN(new_n917));
  OAI211_X1 g716(.A(new_n726), .B(new_n896), .C1(new_n899), .C2(new_n903), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT59), .ZN(new_n919));
  AND3_X1   g718(.A1(new_n918), .A2(new_n919), .A3(G148gat), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n874), .A2(new_n573), .A3(new_n898), .ZN(new_n921));
  INV_X1    g720(.A(new_n855), .ZN(new_n922));
  OR2_X1    g721(.A1(new_n901), .A2(new_n922), .ZN(new_n923));
  AOI22_X1  g722(.A1(new_n684), .A2(new_n281), .B1(new_n923), .B2(new_n717), .ZN(new_n924));
  OAI21_X1  g723(.A(new_n900), .B1(new_n924), .B2(new_n533), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n921), .A2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n726), .A3(new_n896), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n919), .B1(new_n927), .B2(G148gat), .ZN(new_n928));
  OAI21_X1  g727(.A(new_n917), .B1(new_n920), .B2(new_n928), .ZN(G1345gat));
  OAI21_X1  g728(.A(new_n896), .B1(new_n899), .B2(new_n903), .ZN(new_n930));
  OAI21_X1  g729(.A(G155gat), .B1(new_n930), .B2(new_n724), .ZN(new_n931));
  INV_X1    g730(.A(G155gat), .ZN(new_n932));
  NAND3_X1  g731(.A1(new_n915), .A2(new_n932), .A3(new_n624), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n931), .A2(new_n933), .ZN(G1346gat));
  OAI21_X1  g733(.A(G162gat), .B1(new_n930), .B2(new_n661), .ZN(new_n935));
  INV_X1    g734(.A(G162gat), .ZN(new_n936));
  NAND3_X1  g735(.A1(new_n915), .A2(new_n936), .A3(new_n660), .ZN(new_n937));
  NAND2_X1  g736(.A1(new_n935), .A2(new_n937), .ZN(G1347gat));
  AND2_X1   g737(.A1(new_n874), .A2(new_n574), .ZN(new_n939));
  NAND3_X1  g738(.A1(new_n590), .A2(new_n487), .A3(new_n592), .ZN(new_n940));
  XNOR2_X1  g739(.A(new_n940), .B(KEYINPUT122), .ZN(new_n941));
  NAND3_X1  g740(.A1(new_n939), .A2(KEYINPUT123), .A3(new_n941), .ZN(new_n942));
  NAND3_X1  g741(.A1(new_n874), .A2(new_n574), .A3(new_n941), .ZN(new_n943));
  INV_X1    g742(.A(KEYINPUT123), .ZN(new_n944));
  NAND2_X1  g743(.A1(new_n943), .A2(new_n944), .ZN(new_n945));
  NOR2_X1   g744(.A1(new_n281), .A2(G169gat), .ZN(new_n946));
  NAND3_X1  g745(.A1(new_n942), .A2(new_n945), .A3(new_n946), .ZN(new_n947));
  INV_X1    g746(.A(KEYINPUT124), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n947), .A2(new_n948), .ZN(new_n949));
  NOR2_X1   g748(.A1(new_n690), .A2(new_n486), .ZN(new_n950));
  NAND2_X1  g749(.A1(new_n950), .A2(new_n581), .ZN(new_n951));
  XOR2_X1   g750(.A(new_n951), .B(KEYINPUT125), .Z(new_n952));
  NAND3_X1  g751(.A1(new_n879), .A2(new_n280), .A3(new_n952), .ZN(new_n953));
  AOI21_X1  g752(.A(KEYINPUT124), .B1(new_n953), .B2(G169gat), .ZN(new_n954));
  AOI21_X1  g753(.A(new_n949), .B1(new_n954), .B2(new_n947), .ZN(G1348gat));
  NAND4_X1  g754(.A1(new_n942), .A2(new_n400), .A3(new_n726), .A4(new_n945), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n879), .A2(new_n952), .ZN(new_n957));
  OAI21_X1  g756(.A(G176gat), .B1(new_n957), .B2(new_n683), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n956), .A2(new_n958), .ZN(G1349gat));
  OAI21_X1  g758(.A(G183gat), .B1(new_n957), .B2(new_n724), .ZN(new_n960));
  NAND4_X1  g759(.A1(new_n939), .A2(new_n429), .A3(new_n624), .A4(new_n941), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n960), .A2(new_n961), .ZN(new_n962));
  NAND2_X1  g761(.A1(new_n962), .A2(KEYINPUT60), .ZN(new_n963));
  INV_X1    g762(.A(KEYINPUT60), .ZN(new_n964));
  NAND3_X1  g763(.A1(new_n960), .A2(new_n964), .A3(new_n961), .ZN(new_n965));
  NAND2_X1  g764(.A1(new_n963), .A2(new_n965), .ZN(G1350gat));
  NAND4_X1  g765(.A1(new_n942), .A2(new_n431), .A3(new_n660), .A4(new_n945), .ZN(new_n967));
  OAI21_X1  g766(.A(G190gat), .B1(new_n957), .B2(new_n661), .ZN(new_n968));
  AND2_X1   g767(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n969));
  NOR2_X1   g768(.A1(new_n968), .A2(KEYINPUT61), .ZN(new_n970));
  OAI21_X1  g769(.A(new_n967), .B1(new_n969), .B2(new_n970), .ZN(G1351gat));
  NOR2_X1   g770(.A1(new_n906), .A2(new_n486), .ZN(new_n972));
  AND2_X1   g771(.A1(new_n939), .A2(new_n972), .ZN(new_n973));
  AOI21_X1  g772(.A(G197gat), .B1(new_n973), .B2(new_n280), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n950), .A2(new_n794), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n975), .B1(new_n921), .B2(new_n925), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n280), .A2(G197gat), .ZN(new_n977));
  AOI21_X1  g776(.A(new_n974), .B1(new_n976), .B2(new_n977), .ZN(G1352gat));
  NAND2_X1  g777(.A1(new_n939), .A2(new_n972), .ZN(new_n979));
  NOR3_X1   g778(.A1(new_n979), .A2(G204gat), .A3(new_n683), .ZN(new_n980));
  NAND2_X1  g779(.A1(KEYINPUT126), .A2(KEYINPUT62), .ZN(new_n981));
  NAND2_X1  g780(.A1(new_n980), .A2(new_n981), .ZN(new_n982));
  NAND2_X1  g781(.A1(new_n976), .A2(new_n726), .ZN(new_n983));
  NAND2_X1  g782(.A1(new_n983), .A2(G204gat), .ZN(new_n984));
  XOR2_X1   g783(.A(KEYINPUT126), .B(KEYINPUT62), .Z(new_n985));
  OAI211_X1 g784(.A(new_n982), .B(new_n984), .C1(new_n980), .C2(new_n985), .ZN(G1353gat));
  NAND3_X1  g785(.A1(new_n973), .A2(new_n388), .A3(new_n624), .ZN(new_n987));
  NAND2_X1  g786(.A1(new_n976), .A2(new_n624), .ZN(new_n988));
  AOI21_X1  g787(.A(KEYINPUT63), .B1(new_n988), .B2(G211gat), .ZN(new_n989));
  INV_X1    g788(.A(KEYINPUT63), .ZN(new_n990));
  AOI211_X1 g789(.A(new_n990), .B(new_n388), .C1(new_n976), .C2(new_n624), .ZN(new_n991));
  OAI21_X1  g790(.A(new_n987), .B1(new_n989), .B2(new_n991), .ZN(G1354gat));
  NAND3_X1  g791(.A1(new_n973), .A2(new_n389), .A3(new_n660), .ZN(new_n993));
  AND2_X1   g792(.A1(new_n976), .A2(new_n660), .ZN(new_n994));
  OAI211_X1 g793(.A(new_n993), .B(KEYINPUT127), .C1(new_n994), .C2(new_n389), .ZN(new_n995));
  INV_X1    g794(.A(KEYINPUT127), .ZN(new_n996));
  NOR3_X1   g795(.A1(new_n979), .A2(G218gat), .A3(new_n661), .ZN(new_n997));
  AOI21_X1  g796(.A(new_n389), .B1(new_n976), .B2(new_n660), .ZN(new_n998));
  OAI21_X1  g797(.A(new_n996), .B1(new_n997), .B2(new_n998), .ZN(new_n999));
  NAND2_X1  g798(.A1(new_n995), .A2(new_n999), .ZN(G1355gat));
endmodule


