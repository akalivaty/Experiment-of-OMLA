//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 0 0 0 1 1 0 0 1 0 1 0 0 0 0 0 0 1 1 0 1 0 1 0 1 1 0 1 0 1 1 1 0 0 0 1 0 0 0 1 1 1 0 1 1 0 1 0 1 1 0 0 0 0 0 1 0 1 1 0 1 0 0 1 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:58 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n667, new_n668, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n679, new_n680, new_n681,
    new_n682, new_n683, new_n684, new_n685, new_n686, new_n687, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n703,
    new_n704, new_n705, new_n706, new_n708, new_n709, new_n710, new_n711,
    new_n712, new_n713, new_n714, new_n715, new_n716, new_n717, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n728, new_n729, new_n730, new_n732, new_n733, new_n734, new_n735,
    new_n736, new_n737, new_n738, new_n740, new_n741, new_n742, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n754, new_n755, new_n756, new_n758,
    new_n759, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n767, new_n768, new_n769, new_n770, new_n771, new_n772, new_n773,
    new_n774, new_n775, new_n776, new_n777, new_n778, new_n779, new_n780,
    new_n781, new_n782, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n790, new_n791, new_n792, new_n793, new_n794, new_n795,
    new_n796, new_n797, new_n799, new_n800, new_n801, new_n802, new_n803,
    new_n804, new_n805, new_n806, new_n807, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n836, new_n837, new_n838, new_n839, new_n840,
    new_n841, new_n842, new_n843, new_n844, new_n845, new_n846, new_n847,
    new_n848, new_n849, new_n850, new_n851, new_n852, new_n853, new_n854,
    new_n855, new_n856, new_n858, new_n859, new_n861, new_n862, new_n863,
    new_n864, new_n865, new_n867, new_n868, new_n869, new_n870, new_n871,
    new_n872, new_n873, new_n874, new_n875, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n882, new_n883, new_n884, new_n885, new_n886,
    new_n887, new_n888, new_n889, new_n890, new_n891, new_n892, new_n893,
    new_n894, new_n895, new_n896, new_n897, new_n898, new_n899, new_n900,
    new_n901, new_n902, new_n903, new_n904, new_n905, new_n906, new_n907,
    new_n908, new_n909, new_n910, new_n911, new_n912, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n928, new_n929, new_n931,
    new_n932, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n943, new_n944, new_n946, new_n947, new_n948,
    new_n950, new_n951, new_n952, new_n953, new_n955, new_n956, new_n957,
    new_n958, new_n959, new_n960, new_n961, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n969, new_n970, new_n971, new_n972, new_n974,
    new_n975, new_n976;
  NAND2_X1  g000(.A1(G227gat), .A2(G233gat), .ZN(new_n202));
  INV_X1    g001(.A(G169gat), .ZN(new_n203));
  INV_X1    g002(.A(G176gat), .ZN(new_n204));
  NAND3_X1  g003(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT26), .ZN(new_n205));
  INV_X1    g004(.A(KEYINPUT26), .ZN(new_n206));
  OAI21_X1  g005(.A(new_n206), .B1(G169gat), .B2(G176gat), .ZN(new_n207));
  AOI22_X1  g006(.A1(new_n205), .A2(new_n207), .B1(G169gat), .B2(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(G183gat), .A2(G190gat), .ZN(new_n209));
  INV_X1    g008(.A(new_n209), .ZN(new_n210));
  XNOR2_X1  g009(.A(KEYINPUT27), .B(G183gat), .ZN(new_n211));
  INV_X1    g010(.A(G190gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n211), .A2(new_n212), .ZN(new_n213));
  INV_X1    g012(.A(KEYINPUT28), .ZN(new_n214));
  NAND2_X1  g013(.A1(new_n213), .A2(new_n214), .ZN(new_n215));
  NAND3_X1  g014(.A1(new_n211), .A2(KEYINPUT28), .A3(new_n212), .ZN(new_n216));
  AOI211_X1 g015(.A(new_n208), .B(new_n210), .C1(new_n215), .C2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(new_n217), .ZN(new_n218));
  INV_X1    g017(.A(KEYINPUT66), .ZN(new_n219));
  INV_X1    g018(.A(KEYINPUT24), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n209), .A2(new_n220), .ZN(new_n221));
  OR2_X1    g020(.A1(G183gat), .A2(G190gat), .ZN(new_n222));
  NAND3_X1  g021(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n223));
  NAND3_X1  g022(.A1(new_n221), .A2(new_n222), .A3(new_n223), .ZN(new_n224));
  NAND3_X1  g023(.A1(new_n203), .A2(new_n204), .A3(KEYINPUT23), .ZN(new_n225));
  INV_X1    g024(.A(KEYINPUT23), .ZN(new_n226));
  OAI21_X1  g025(.A(new_n226), .B1(G169gat), .B2(G176gat), .ZN(new_n227));
  NAND2_X1  g026(.A1(G169gat), .A2(G176gat), .ZN(new_n228));
  AND4_X1   g027(.A1(KEYINPUT25), .A2(new_n225), .A3(new_n227), .A4(new_n228), .ZN(new_n229));
  OAI21_X1  g028(.A(new_n223), .B1(G183gat), .B2(G190gat), .ZN(new_n230));
  AOI21_X1  g029(.A(KEYINPUT24), .B1(G183gat), .B2(G190gat), .ZN(new_n231));
  OAI21_X1  g030(.A(KEYINPUT65), .B1(new_n230), .B2(new_n231), .ZN(new_n232));
  INV_X1    g031(.A(KEYINPUT65), .ZN(new_n233));
  NAND4_X1  g032(.A1(new_n221), .A2(new_n222), .A3(new_n233), .A4(new_n223), .ZN(new_n234));
  AND3_X1   g033(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n235));
  NAND3_X1  g034(.A1(new_n232), .A2(new_n234), .A3(new_n235), .ZN(new_n236));
  XOR2_X1   g035(.A(KEYINPUT64), .B(KEYINPUT25), .Z(new_n237));
  INV_X1    g036(.A(new_n237), .ZN(new_n238));
  AOI221_X4 g037(.A(new_n219), .B1(new_n224), .B2(new_n229), .C1(new_n236), .C2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n236), .A2(new_n238), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n229), .A2(new_n224), .ZN(new_n241));
  AOI21_X1  g040(.A(KEYINPUT66), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  OAI21_X1  g041(.A(new_n218), .B1(new_n239), .B2(new_n242), .ZN(new_n243));
  INV_X1    g042(.A(G134gat), .ZN(new_n244));
  NAND2_X1  g043(.A1(new_n244), .A2(G127gat), .ZN(new_n245));
  INV_X1    g044(.A(KEYINPUT67), .ZN(new_n246));
  NAND2_X1  g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  NAND3_X1  g046(.A1(new_n244), .A2(KEYINPUT67), .A3(G127gat), .ZN(new_n248));
  INV_X1    g047(.A(G127gat), .ZN(new_n249));
  NAND2_X1  g048(.A1(new_n249), .A2(G134gat), .ZN(new_n250));
  NAND3_X1  g049(.A1(new_n247), .A2(new_n248), .A3(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT1), .ZN(new_n252));
  XNOR2_X1  g051(.A(G113gat), .B(G120gat), .ZN(new_n253));
  OAI21_X1  g052(.A(new_n252), .B1(new_n253), .B2(KEYINPUT68), .ZN(new_n254));
  INV_X1    g053(.A(G120gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G113gat), .ZN(new_n256));
  INV_X1    g055(.A(G113gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G120gat), .ZN(new_n258));
  NAND3_X1  g057(.A1(new_n256), .A2(new_n258), .A3(KEYINPUT68), .ZN(new_n259));
  INV_X1    g058(.A(new_n259), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n251), .B1(new_n254), .B2(new_n260), .ZN(new_n261));
  NAND3_X1  g060(.A1(new_n245), .A2(new_n250), .A3(new_n252), .ZN(new_n262));
  NOR2_X1   g061(.A1(new_n262), .A2(new_n253), .ZN(new_n263));
  INV_X1    g062(.A(new_n263), .ZN(new_n264));
  NAND2_X1  g063(.A1(new_n261), .A2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n243), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n225), .A2(new_n227), .A3(new_n228), .ZN(new_n267));
  AOI21_X1  g066(.A(new_n267), .B1(KEYINPUT65), .B2(new_n224), .ZN(new_n268));
  AOI21_X1  g067(.A(new_n237), .B1(new_n268), .B2(new_n234), .ZN(new_n269));
  NOR2_X1   g068(.A1(new_n230), .A2(new_n231), .ZN(new_n270));
  INV_X1    g069(.A(KEYINPUT25), .ZN(new_n271));
  NOR3_X1   g070(.A1(new_n270), .A2(new_n271), .A3(new_n267), .ZN(new_n272));
  OAI21_X1  g071(.A(new_n219), .B1(new_n269), .B2(new_n272), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n240), .A2(KEYINPUT66), .A3(new_n241), .ZN(new_n274));
  NAND2_X1  g073(.A1(new_n273), .A2(new_n274), .ZN(new_n275));
  INV_X1    g074(.A(KEYINPUT68), .ZN(new_n276));
  NOR2_X1   g075(.A1(new_n257), .A2(G120gat), .ZN(new_n277));
  NOR2_X1   g076(.A1(new_n255), .A2(G113gat), .ZN(new_n278));
  OAI21_X1  g077(.A(new_n276), .B1(new_n277), .B2(new_n278), .ZN(new_n279));
  NAND3_X1  g078(.A1(new_n279), .A2(new_n252), .A3(new_n259), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n263), .B1(new_n280), .B2(new_n251), .ZN(new_n281));
  NAND3_X1  g080(.A1(new_n275), .A2(new_n281), .A3(new_n218), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n202), .B1(new_n266), .B2(new_n282), .ZN(new_n283));
  XNOR2_X1  g082(.A(G15gat), .B(G43gat), .ZN(new_n284));
  XNOR2_X1  g083(.A(G71gat), .B(G99gat), .ZN(new_n285));
  XOR2_X1   g084(.A(new_n284), .B(new_n285), .Z(new_n286));
  XOR2_X1   g085(.A(KEYINPUT69), .B(KEYINPUT33), .Z(new_n287));
  NAND2_X1  g086(.A1(new_n286), .A2(new_n287), .ZN(new_n288));
  NAND2_X1  g087(.A1(new_n288), .A2(KEYINPUT32), .ZN(new_n289));
  NOR2_X1   g088(.A1(new_n283), .A2(new_n289), .ZN(new_n290));
  INV_X1    g089(.A(new_n290), .ZN(new_n291));
  INV_X1    g090(.A(new_n202), .ZN(new_n292));
  AOI21_X1  g091(.A(new_n281), .B1(new_n275), .B2(new_n218), .ZN(new_n293));
  AOI211_X1 g092(.A(new_n265), .B(new_n217), .C1(new_n273), .C2(new_n274), .ZN(new_n294));
  OAI21_X1  g093(.A(new_n292), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  INV_X1    g094(.A(new_n287), .ZN(new_n296));
  NOR2_X1   g095(.A1(new_n296), .A2(KEYINPUT32), .ZN(new_n297));
  INV_X1    g096(.A(new_n297), .ZN(new_n298));
  NAND2_X1  g097(.A1(new_n295), .A2(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(KEYINPUT70), .B1(new_n299), .B2(new_n286), .ZN(new_n300));
  INV_X1    g099(.A(KEYINPUT70), .ZN(new_n301));
  INV_X1    g100(.A(new_n286), .ZN(new_n302));
  AOI211_X1 g101(.A(new_n301), .B(new_n302), .C1(new_n295), .C2(new_n298), .ZN(new_n303));
  OAI21_X1  g102(.A(new_n291), .B1(new_n300), .B2(new_n303), .ZN(new_n304));
  INV_X1    g103(.A(KEYINPUT71), .ZN(new_n305));
  AOI21_X1  g104(.A(new_n292), .B1(new_n305), .B2(KEYINPUT34), .ZN(new_n306));
  NAND3_X1  g105(.A1(new_n266), .A2(new_n282), .A3(new_n306), .ZN(new_n307));
  NOR2_X1   g106(.A1(new_n305), .A2(KEYINPUT34), .ZN(new_n308));
  NAND2_X1  g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g108(.A(new_n308), .ZN(new_n310));
  NAND4_X1  g109(.A1(new_n266), .A2(new_n282), .A3(new_n306), .A4(new_n310), .ZN(new_n311));
  NAND2_X1  g110(.A1(new_n309), .A2(new_n311), .ZN(new_n312));
  NAND2_X1  g111(.A1(new_n304), .A2(new_n312), .ZN(new_n313));
  OAI21_X1  g112(.A(new_n286), .B1(new_n283), .B2(new_n297), .ZN(new_n314));
  NAND2_X1  g113(.A1(new_n314), .A2(new_n301), .ZN(new_n315));
  OAI211_X1 g114(.A(KEYINPUT70), .B(new_n286), .C1(new_n283), .C2(new_n297), .ZN(new_n316));
  NAND2_X1  g115(.A1(new_n315), .A2(new_n316), .ZN(new_n317));
  INV_X1    g116(.A(new_n312), .ZN(new_n318));
  NAND3_X1  g117(.A1(new_n317), .A2(new_n291), .A3(new_n318), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n313), .A2(KEYINPUT36), .A3(new_n319), .ZN(new_n320));
  XNOR2_X1  g119(.A(G8gat), .B(G36gat), .ZN(new_n321));
  XNOR2_X1  g120(.A(G64gat), .B(G92gat), .ZN(new_n322));
  XNOR2_X1  g121(.A(new_n321), .B(new_n322), .ZN(new_n323));
  AND2_X1   g122(.A1(G211gat), .A2(G218gat), .ZN(new_n324));
  AND2_X1   g123(.A1(G197gat), .A2(G204gat), .ZN(new_n325));
  NOR2_X1   g124(.A1(G197gat), .A2(G204gat), .ZN(new_n326));
  OAI22_X1  g125(.A1(KEYINPUT22), .A2(new_n324), .B1(new_n325), .B2(new_n326), .ZN(new_n327));
  XOR2_X1   g126(.A(G211gat), .B(G218gat), .Z(new_n328));
  XNOR2_X1  g127(.A(new_n327), .B(new_n328), .ZN(new_n329));
  AOI21_X1  g128(.A(new_n272), .B1(new_n236), .B2(new_n238), .ZN(new_n330));
  INV_X1    g129(.A(G226gat), .ZN(new_n331));
  INV_X1    g130(.A(G233gat), .ZN(new_n332));
  NOR2_X1   g131(.A1(new_n331), .A2(new_n332), .ZN(new_n333));
  INV_X1    g132(.A(new_n333), .ZN(new_n334));
  NOR3_X1   g133(.A1(new_n330), .A2(new_n217), .A3(new_n334), .ZN(new_n335));
  NOR2_X1   g134(.A1(new_n333), .A2(KEYINPUT29), .ZN(new_n336));
  AOI211_X1 g135(.A(new_n329), .B(new_n335), .C1(new_n243), .C2(new_n336), .ZN(new_n337));
  INV_X1    g136(.A(new_n329), .ZN(new_n338));
  INV_X1    g137(.A(new_n330), .ZN(new_n339));
  NAND2_X1  g138(.A1(new_n339), .A2(new_n218), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n336), .ZN(new_n341));
  OAI211_X1 g140(.A(new_n218), .B(new_n333), .C1(new_n239), .C2(new_n242), .ZN(new_n342));
  AOI21_X1  g141(.A(new_n338), .B1(new_n341), .B2(new_n342), .ZN(new_n343));
  OAI21_X1  g142(.A(new_n323), .B1(new_n337), .B2(new_n343), .ZN(new_n344));
  INV_X1    g143(.A(new_n335), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n217), .B1(new_n273), .B2(new_n274), .ZN(new_n346));
  INV_X1    g145(.A(new_n336), .ZN(new_n347));
  OAI211_X1 g146(.A(new_n345), .B(new_n338), .C1(new_n346), .C2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(new_n323), .ZN(new_n349));
  AOI22_X1  g148(.A1(new_n346), .A2(new_n333), .B1(new_n340), .B2(new_n336), .ZN(new_n350));
  OAI211_X1 g149(.A(new_n348), .B(new_n349), .C1(new_n350), .C2(new_n338), .ZN(new_n351));
  NAND3_X1  g150(.A1(new_n344), .A2(KEYINPUT30), .A3(new_n351), .ZN(new_n352));
  INV_X1    g151(.A(new_n343), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND4_X1  g153(.A1(new_n353), .A2(new_n354), .A3(new_n348), .A4(new_n349), .ZN(new_n355));
  AND2_X1   g154(.A1(new_n352), .A2(new_n355), .ZN(new_n356));
  AND2_X1   g155(.A1(G155gat), .A2(G162gat), .ZN(new_n357));
  NOR2_X1   g156(.A1(G155gat), .A2(G162gat), .ZN(new_n358));
  NOR2_X1   g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  XNOR2_X1  g158(.A(G141gat), .B(G148gat), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT2), .ZN(new_n361));
  AOI21_X1  g160(.A(new_n361), .B1(G155gat), .B2(G162gat), .ZN(new_n362));
  OAI21_X1  g161(.A(new_n359), .B1(new_n360), .B2(new_n362), .ZN(new_n363));
  INV_X1    g162(.A(G141gat), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n364), .A2(G148gat), .ZN(new_n365));
  INV_X1    g164(.A(G148gat), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n366), .A2(G141gat), .ZN(new_n367));
  NAND2_X1  g166(.A1(new_n365), .A2(new_n367), .ZN(new_n368));
  XNOR2_X1  g167(.A(G155gat), .B(G162gat), .ZN(new_n369));
  INV_X1    g168(.A(G155gat), .ZN(new_n370));
  INV_X1    g169(.A(G162gat), .ZN(new_n371));
  OAI21_X1  g170(.A(KEYINPUT2), .B1(new_n370), .B2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n368), .A2(new_n369), .A3(new_n372), .ZN(new_n373));
  AND2_X1   g172(.A1(new_n363), .A2(new_n373), .ZN(new_n374));
  NAND3_X1  g173(.A1(new_n374), .A2(new_n261), .A3(new_n264), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT4), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  NAND3_X1  g176(.A1(new_n281), .A2(new_n377), .A3(new_n374), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT3), .ZN(new_n379));
  AND3_X1   g178(.A1(new_n363), .A2(new_n373), .A3(new_n379), .ZN(new_n380));
  AOI21_X1  g179(.A(new_n379), .B1(new_n363), .B2(new_n373), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n380), .A2(new_n381), .ZN(new_n382));
  AOI22_X1  g181(.A1(new_n376), .A2(new_n378), .B1(new_n265), .B2(new_n382), .ZN(new_n383));
  NAND2_X1  g182(.A1(G225gat), .A2(G233gat), .ZN(new_n384));
  XNOR2_X1  g183(.A(new_n384), .B(KEYINPUT72), .ZN(new_n385));
  INV_X1    g184(.A(new_n385), .ZN(new_n386));
  OR3_X1    g185(.A1(new_n383), .A2(KEYINPUT39), .A3(new_n386), .ZN(new_n387));
  XOR2_X1   g186(.A(KEYINPUT73), .B(KEYINPUT0), .Z(new_n388));
  XNOR2_X1  g187(.A(G1gat), .B(G29gat), .ZN(new_n389));
  XNOR2_X1  g188(.A(new_n388), .B(new_n389), .ZN(new_n390));
  XNOR2_X1  g189(.A(G57gat), .B(G85gat), .ZN(new_n391));
  XNOR2_X1  g190(.A(new_n390), .B(new_n391), .ZN(new_n392));
  NOR2_X1   g191(.A1(new_n383), .A2(new_n386), .ZN(new_n393));
  INV_X1    g192(.A(new_n374), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n265), .A2(new_n394), .ZN(new_n395));
  NAND2_X1  g194(.A1(new_n395), .A2(new_n375), .ZN(new_n396));
  OAI21_X1  g195(.A(KEYINPUT39), .B1(new_n396), .B2(new_n385), .ZN(new_n397));
  OAI211_X1 g196(.A(new_n387), .B(new_n392), .C1(new_n393), .C2(new_n397), .ZN(new_n398));
  OR2_X1    g197(.A1(KEYINPUT78), .A2(KEYINPUT40), .ZN(new_n399));
  XNOR2_X1  g198(.A(new_n398), .B(new_n399), .ZN(new_n400));
  NAND2_X1  g199(.A1(new_n382), .A2(new_n265), .ZN(new_n401));
  AND3_X1   g200(.A1(new_n281), .A2(new_n377), .A3(new_n374), .ZN(new_n402));
  AOI21_X1  g201(.A(new_n377), .B1(new_n281), .B2(new_n374), .ZN(new_n403));
  OAI211_X1 g202(.A(new_n401), .B(new_n386), .C1(new_n402), .C2(new_n403), .ZN(new_n404));
  INV_X1    g203(.A(KEYINPUT5), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n404), .A2(new_n405), .ZN(new_n406));
  AOI21_X1  g205(.A(new_n386), .B1(new_n395), .B2(new_n375), .ZN(new_n407));
  AOI21_X1  g206(.A(new_n407), .B1(new_n383), .B2(new_n386), .ZN(new_n408));
  OAI211_X1 g207(.A(KEYINPUT79), .B(new_n406), .C1(new_n408), .C2(new_n405), .ZN(new_n409));
  INV_X1    g208(.A(KEYINPUT79), .ZN(new_n410));
  NAND2_X1  g209(.A1(new_n396), .A2(new_n385), .ZN(new_n411));
  AOI21_X1  g210(.A(new_n405), .B1(new_n404), .B2(new_n411), .ZN(new_n412));
  AOI21_X1  g211(.A(KEYINPUT5), .B1(new_n383), .B2(new_n386), .ZN(new_n413));
  OAI21_X1  g212(.A(new_n410), .B1(new_n412), .B2(new_n413), .ZN(new_n414));
  INV_X1    g213(.A(new_n392), .ZN(new_n415));
  NAND3_X1  g214(.A1(new_n409), .A2(new_n414), .A3(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n356), .A2(new_n400), .A3(new_n416), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT37), .ZN(new_n418));
  NAND3_X1  g217(.A1(new_n353), .A2(new_n418), .A3(new_n348), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(new_n323), .ZN(new_n420));
  AOI21_X1  g219(.A(new_n418), .B1(new_n353), .B2(new_n348), .ZN(new_n421));
  OAI21_X1  g220(.A(KEYINPUT38), .B1(new_n420), .B2(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT6), .ZN(new_n423));
  NOR4_X1   g222(.A1(new_n412), .A2(new_n413), .A3(new_n423), .A4(new_n392), .ZN(new_n424));
  OAI21_X1  g223(.A(new_n406), .B1(new_n408), .B2(new_n405), .ZN(new_n425));
  AOI21_X1  g224(.A(KEYINPUT6), .B1(new_n425), .B2(new_n392), .ZN(new_n426));
  AOI21_X1  g225(.A(new_n424), .B1(new_n416), .B2(new_n426), .ZN(new_n427));
  OAI211_X1 g226(.A(new_n345), .B(new_n329), .C1(new_n346), .C2(new_n347), .ZN(new_n428));
  OAI211_X1 g227(.A(new_n428), .B(KEYINPUT37), .C1(new_n350), .C2(new_n329), .ZN(new_n429));
  NOR2_X1   g228(.A1(new_n349), .A2(KEYINPUT38), .ZN(new_n430));
  NAND3_X1  g229(.A1(new_n419), .A2(new_n429), .A3(new_n430), .ZN(new_n431));
  NAND4_X1  g230(.A1(new_n422), .A2(new_n427), .A3(new_n351), .A4(new_n431), .ZN(new_n432));
  OR3_X1    g231(.A1(new_n380), .A2(KEYINPUT75), .A3(KEYINPUT29), .ZN(new_n433));
  OAI21_X1  g232(.A(KEYINPUT75), .B1(new_n380), .B2(KEYINPUT29), .ZN(new_n434));
  NAND3_X1  g233(.A1(new_n433), .A2(new_n338), .A3(new_n434), .ZN(new_n435));
  AND2_X1   g234(.A1(G228gat), .A2(G233gat), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT29), .ZN(new_n437));
  AOI21_X1  g236(.A(KEYINPUT3), .B1(new_n329), .B2(new_n437), .ZN(new_n438));
  OAI211_X1 g237(.A(new_n435), .B(new_n436), .C1(new_n374), .C2(new_n438), .ZN(new_n439));
  INV_X1    g238(.A(new_n436), .ZN(new_n440));
  NAND3_X1  g239(.A1(new_n327), .A2(KEYINPUT74), .A3(new_n328), .ZN(new_n441));
  OAI211_X1 g240(.A(new_n437), .B(new_n441), .C1(new_n329), .C2(KEYINPUT74), .ZN(new_n442));
  AOI21_X1  g241(.A(new_n374), .B1(new_n442), .B2(new_n379), .ZN(new_n443));
  NOR2_X1   g242(.A1(new_n380), .A2(KEYINPUT29), .ZN(new_n444));
  NOR2_X1   g243(.A1(new_n444), .A2(new_n329), .ZN(new_n445));
  OAI21_X1  g244(.A(new_n440), .B1(new_n443), .B2(new_n445), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n439), .A2(new_n446), .ZN(new_n447));
  OAI21_X1  g246(.A(KEYINPUT76), .B1(new_n447), .B2(G22gat), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT76), .ZN(new_n449));
  INV_X1    g248(.A(G22gat), .ZN(new_n450));
  NAND4_X1  g249(.A1(new_n439), .A2(new_n446), .A3(new_n449), .A4(new_n450), .ZN(new_n451));
  INV_X1    g250(.A(new_n447), .ZN(new_n452));
  OAI211_X1 g251(.A(new_n448), .B(new_n451), .C1(new_n450), .C2(new_n452), .ZN(new_n453));
  XOR2_X1   g252(.A(KEYINPUT31), .B(G50gat), .Z(new_n454));
  XNOR2_X1  g253(.A(G78gat), .B(G106gat), .ZN(new_n455));
  XNOR2_X1  g254(.A(new_n454), .B(new_n455), .ZN(new_n456));
  NAND2_X1  g255(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g256(.A(KEYINPUT77), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n458), .A2(G22gat), .ZN(new_n459));
  AOI21_X1  g258(.A(new_n456), .B1(new_n452), .B2(new_n459), .ZN(new_n460));
  NAND3_X1  g259(.A1(new_n447), .A2(new_n458), .A3(G22gat), .ZN(new_n461));
  NAND2_X1  g260(.A1(new_n460), .A2(new_n461), .ZN(new_n462));
  NAND2_X1  g261(.A1(new_n457), .A2(new_n462), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n417), .A2(new_n432), .A3(new_n463), .ZN(new_n464));
  AOI22_X1  g263(.A1(new_n453), .A2(new_n456), .B1(new_n461), .B2(new_n460), .ZN(new_n465));
  OAI21_X1  g264(.A(new_n426), .B1(new_n392), .B2(new_n425), .ZN(new_n466));
  INV_X1    g265(.A(new_n424), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  INV_X1    g267(.A(new_n468), .ZN(new_n469));
  OAI21_X1  g268(.A(new_n465), .B1(new_n469), .B2(new_n356), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT36), .ZN(new_n471));
  AOI21_X1  g270(.A(new_n318), .B1(new_n317), .B2(new_n291), .ZN(new_n472));
  AOI211_X1 g271(.A(new_n290), .B(new_n312), .C1(new_n315), .C2(new_n316), .ZN(new_n473));
  OAI21_X1  g272(.A(new_n471), .B1(new_n472), .B2(new_n473), .ZN(new_n474));
  AND4_X1   g273(.A1(new_n320), .A2(new_n464), .A3(new_n470), .A4(new_n474), .ZN(new_n475));
  INV_X1    g274(.A(KEYINPUT80), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n476), .B1(new_n356), .B2(new_n427), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n416), .A2(new_n426), .ZN(new_n478));
  NAND2_X1  g277(.A1(new_n478), .A2(new_n467), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n352), .A2(new_n355), .ZN(new_n480));
  NAND3_X1  g279(.A1(new_n479), .A2(KEYINPUT80), .A3(new_n480), .ZN(new_n481));
  NAND2_X1  g280(.A1(new_n477), .A2(new_n481), .ZN(new_n482));
  AOI21_X1  g281(.A(new_n465), .B1(new_n313), .B2(new_n319), .ZN(new_n483));
  XOR2_X1   g282(.A(KEYINPUT81), .B(KEYINPUT35), .Z(new_n484));
  NAND3_X1  g283(.A1(new_n482), .A2(new_n483), .A3(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n313), .A2(new_n319), .ZN(new_n486));
  AND2_X1   g285(.A1(new_n468), .A2(new_n480), .ZN(new_n487));
  NAND3_X1  g286(.A1(new_n486), .A2(new_n487), .A3(new_n463), .ZN(new_n488));
  AOI22_X1  g287(.A1(new_n485), .A2(KEYINPUT82), .B1(KEYINPUT35), .B2(new_n488), .ZN(new_n489));
  INV_X1    g288(.A(KEYINPUT82), .ZN(new_n490));
  NAND4_X1  g289(.A1(new_n482), .A2(new_n483), .A3(new_n490), .A4(new_n484), .ZN(new_n491));
  AOI21_X1  g290(.A(new_n475), .B1(new_n489), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(KEYINPUT93), .ZN(new_n493));
  NAND2_X1  g292(.A1(G229gat), .A2(G233gat), .ZN(new_n494));
  XOR2_X1   g293(.A(new_n494), .B(KEYINPUT13), .Z(new_n495));
  XNOR2_X1  g294(.A(G15gat), .B(G22gat), .ZN(new_n496));
  INV_X1    g295(.A(G1gat), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT16), .ZN(new_n498));
  NAND2_X1  g297(.A1(new_n496), .A2(new_n498), .ZN(new_n499));
  OAI21_X1  g298(.A(new_n499), .B1(G1gat), .B2(new_n496), .ZN(new_n500));
  INV_X1    g299(.A(G8gat), .ZN(new_n501));
  XNOR2_X1  g300(.A(new_n500), .B(new_n501), .ZN(new_n502));
  OR2_X1    g301(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n503));
  NAND2_X1  g302(.A1(new_n502), .A2(KEYINPUT90), .ZN(new_n504));
  AND2_X1   g303(.A1(new_n503), .A2(new_n504), .ZN(new_n505));
  OAI21_X1  g304(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n506));
  XNOR2_X1  g305(.A(new_n506), .B(KEYINPUT85), .ZN(new_n507));
  OR3_X1    g306(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n508));
  AND3_X1   g307(.A1(new_n507), .A2(KEYINPUT88), .A3(new_n508), .ZN(new_n509));
  AOI21_X1  g308(.A(KEYINPUT88), .B1(new_n507), .B2(new_n508), .ZN(new_n510));
  XNOR2_X1  g309(.A(G43gat), .B(G50gat), .ZN(new_n511));
  OR2_X1    g310(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n511), .A2(KEYINPUT15), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT87), .B(G29gat), .ZN(new_n514));
  NAND2_X1  g313(.A1(new_n514), .A2(G36gat), .ZN(new_n515));
  NAND3_X1  g314(.A1(new_n512), .A2(new_n513), .A3(new_n515), .ZN(new_n516));
  OR3_X1    g315(.A1(new_n509), .A2(new_n510), .A3(new_n516), .ZN(new_n517));
  XNOR2_X1  g316(.A(new_n508), .B(KEYINPUT86), .ZN(new_n518));
  INV_X1    g317(.A(new_n507), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NAND3_X1  g319(.A1(new_n520), .A2(KEYINPUT15), .A3(new_n511), .ZN(new_n521));
  NAND2_X1  g320(.A1(new_n517), .A2(new_n521), .ZN(new_n522));
  OAI21_X1  g321(.A(KEYINPUT91), .B1(new_n505), .B2(new_n522), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n505), .A2(new_n522), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n503), .A2(new_n504), .ZN(new_n525));
  INV_X1    g324(.A(KEYINPUT91), .ZN(new_n526));
  AND2_X1   g325(.A1(new_n517), .A2(new_n521), .ZN(new_n527));
  NAND3_X1  g326(.A1(new_n525), .A2(new_n526), .A3(new_n527), .ZN(new_n528));
  NAND3_X1  g327(.A1(new_n523), .A2(new_n524), .A3(new_n528), .ZN(new_n529));
  NAND2_X1  g328(.A1(new_n527), .A2(KEYINPUT17), .ZN(new_n530));
  XOR2_X1   g329(.A(new_n502), .B(KEYINPUT89), .Z(new_n531));
  INV_X1    g330(.A(KEYINPUT17), .ZN(new_n532));
  NAND2_X1  g331(.A1(new_n522), .A2(new_n532), .ZN(new_n533));
  NAND3_X1  g332(.A1(new_n530), .A2(new_n531), .A3(new_n533), .ZN(new_n534));
  NAND3_X1  g333(.A1(new_n534), .A2(new_n494), .A3(new_n524), .ZN(new_n535));
  INV_X1    g334(.A(KEYINPUT18), .ZN(new_n536));
  AOI22_X1  g335(.A1(new_n495), .A2(new_n529), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  OR2_X1    g336(.A1(new_n535), .A2(new_n536), .ZN(new_n538));
  XNOR2_X1  g337(.A(G169gat), .B(G197gat), .ZN(new_n539));
  XNOR2_X1  g338(.A(new_n539), .B(new_n364), .ZN(new_n540));
  XOR2_X1   g339(.A(KEYINPUT83), .B(KEYINPUT11), .Z(new_n541));
  XNOR2_X1  g340(.A(new_n540), .B(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(KEYINPUT84), .B(G113gat), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(new_n544), .B(KEYINPUT12), .ZN(new_n545));
  NAND3_X1  g344(.A1(new_n537), .A2(new_n538), .A3(new_n545), .ZN(new_n546));
  NAND2_X1  g345(.A1(new_n546), .A2(KEYINPUT92), .ZN(new_n547));
  AOI21_X1  g346(.A(new_n545), .B1(new_n537), .B2(new_n538), .ZN(new_n548));
  NOR2_X1   g347(.A1(new_n547), .A2(new_n548), .ZN(new_n549));
  NAND2_X1  g348(.A1(new_n537), .A2(new_n538), .ZN(new_n550));
  INV_X1    g349(.A(KEYINPUT92), .ZN(new_n551));
  INV_X1    g350(.A(new_n545), .ZN(new_n552));
  NAND3_X1  g351(.A1(new_n550), .A2(new_n551), .A3(new_n552), .ZN(new_n553));
  INV_X1    g352(.A(new_n553), .ZN(new_n554));
  OAI21_X1  g353(.A(new_n493), .B1(new_n549), .B2(new_n554), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n550), .A2(new_n552), .ZN(new_n556));
  NAND3_X1  g355(.A1(new_n556), .A2(KEYINPUT92), .A3(new_n546), .ZN(new_n557));
  NAND3_X1  g356(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  INV_X1    g358(.A(new_n559), .ZN(new_n560));
  XNOR2_X1  g359(.A(KEYINPUT94), .B(KEYINPUT19), .ZN(new_n561));
  XNOR2_X1  g360(.A(G57gat), .B(G64gat), .ZN(new_n562));
  AOI21_X1  g361(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n563));
  NOR2_X1   g362(.A1(new_n562), .A2(new_n563), .ZN(new_n564));
  XNOR2_X1  g363(.A(G71gat), .B(G78gat), .ZN(new_n565));
  OR2_X1    g364(.A1(new_n564), .A2(new_n565), .ZN(new_n566));
  NAND2_X1  g365(.A1(new_n564), .A2(new_n565), .ZN(new_n567));
  NAND2_X1  g366(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  INV_X1    g367(.A(new_n568), .ZN(new_n569));
  AOI22_X1  g368(.A1(new_n503), .A2(new_n504), .B1(KEYINPUT21), .B2(new_n569), .ZN(new_n570));
  INV_X1    g369(.A(KEYINPUT21), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  XNOR2_X1  g371(.A(new_n572), .B(KEYINPUT95), .ZN(new_n573));
  NOR2_X1   g372(.A1(new_n570), .A2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n574), .ZN(new_n575));
  NAND2_X1  g374(.A1(new_n570), .A2(new_n573), .ZN(new_n576));
  NAND4_X1  g375(.A1(new_n575), .A2(G231gat), .A3(G233gat), .A4(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  AOI22_X1  g377(.A1(new_n575), .A2(new_n576), .B1(G231gat), .B2(G233gat), .ZN(new_n579));
  OAI21_X1  g378(.A(new_n561), .B1(new_n578), .B2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n579), .ZN(new_n581));
  INV_X1    g380(.A(new_n561), .ZN(new_n582));
  NAND3_X1  g381(.A1(new_n581), .A2(new_n582), .A3(new_n577), .ZN(new_n583));
  NAND2_X1  g382(.A1(new_n580), .A2(new_n583), .ZN(new_n584));
  XOR2_X1   g383(.A(G183gat), .B(G211gat), .Z(new_n585));
  XNOR2_X1  g384(.A(KEYINPUT96), .B(G155gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XOR2_X1   g386(.A(KEYINPUT20), .B(G127gat), .Z(new_n588));
  XOR2_X1   g387(.A(new_n587), .B(new_n588), .Z(new_n589));
  INV_X1    g388(.A(new_n589), .ZN(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  NAND3_X1  g390(.A1(new_n580), .A2(new_n583), .A3(new_n589), .ZN(new_n592));
  NAND2_X1  g391(.A1(new_n591), .A2(new_n592), .ZN(new_n593));
  INV_X1    g392(.A(KEYINPUT7), .ZN(new_n594));
  INV_X1    g393(.A(G85gat), .ZN(new_n595));
  INV_X1    g394(.A(G92gat), .ZN(new_n596));
  OAI21_X1  g395(.A(new_n594), .B1(new_n595), .B2(new_n596), .ZN(new_n597));
  NAND3_X1  g396(.A1(KEYINPUT7), .A2(G85gat), .A3(G92gat), .ZN(new_n598));
  OAI211_X1 g397(.A(new_n597), .B(new_n598), .C1(G85gat), .C2(G92gat), .ZN(new_n599));
  NAND3_X1  g398(.A1(KEYINPUT98), .A2(G99gat), .A3(G106gat), .ZN(new_n600));
  AOI21_X1  g399(.A(KEYINPUT98), .B1(G99gat), .B2(G106gat), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT8), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI21_X1  g402(.A(new_n599), .B1(new_n600), .B2(new_n603), .ZN(new_n604));
  XOR2_X1   g403(.A(G99gat), .B(G106gat), .Z(new_n605));
  INV_X1    g404(.A(new_n605), .ZN(new_n606));
  XNOR2_X1  g405(.A(new_n604), .B(new_n606), .ZN(new_n607));
  NAND3_X1  g406(.A1(new_n530), .A2(new_n533), .A3(new_n607), .ZN(new_n608));
  XNOR2_X1  g407(.A(new_n604), .B(new_n605), .ZN(new_n609));
  AND2_X1   g408(.A1(G232gat), .A2(G233gat), .ZN(new_n610));
  AOI22_X1  g409(.A1(new_n522), .A2(new_n609), .B1(KEYINPUT41), .B2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n608), .A2(new_n611), .ZN(new_n612));
  XNOR2_X1  g411(.A(G190gat), .B(G218gat), .ZN(new_n613));
  XNOR2_X1  g412(.A(new_n613), .B(KEYINPUT99), .ZN(new_n614));
  INV_X1    g413(.A(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(new_n612), .B(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n610), .A2(KEYINPUT41), .ZN(new_n617));
  XNOR2_X1  g416(.A(new_n617), .B(KEYINPUT97), .ZN(new_n618));
  XNOR2_X1  g417(.A(G134gat), .B(G162gat), .ZN(new_n619));
  XNOR2_X1  g418(.A(new_n618), .B(new_n619), .ZN(new_n620));
  XNOR2_X1  g419(.A(new_n616), .B(new_n620), .ZN(new_n621));
  INV_X1    g420(.A(new_n621), .ZN(new_n622));
  NAND2_X1  g421(.A1(new_n607), .A2(new_n568), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n609), .A2(new_n569), .ZN(new_n624));
  INV_X1    g423(.A(KEYINPUT10), .ZN(new_n625));
  NAND3_X1  g424(.A1(new_n623), .A2(new_n624), .A3(new_n625), .ZN(new_n626));
  NAND3_X1  g425(.A1(new_n609), .A2(KEYINPUT10), .A3(new_n569), .ZN(new_n627));
  NAND2_X1  g426(.A1(new_n626), .A2(new_n627), .ZN(new_n628));
  NAND2_X1  g427(.A1(G230gat), .A2(G233gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(KEYINPUT100), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  NAND2_X1  g430(.A1(new_n628), .A2(new_n631), .ZN(new_n632));
  AOI21_X1  g431(.A(new_n631), .B1(new_n623), .B2(new_n624), .ZN(new_n633));
  INV_X1    g432(.A(new_n633), .ZN(new_n634));
  XNOR2_X1  g433(.A(G176gat), .B(G204gat), .ZN(new_n635));
  XNOR2_X1  g434(.A(new_n635), .B(KEYINPUT101), .ZN(new_n636));
  XNOR2_X1  g435(.A(G120gat), .B(G148gat), .ZN(new_n637));
  XOR2_X1   g436(.A(new_n636), .B(new_n637), .Z(new_n638));
  INV_X1    g437(.A(new_n638), .ZN(new_n639));
  NAND3_X1  g438(.A1(new_n632), .A2(new_n634), .A3(new_n639), .ZN(new_n640));
  XOR2_X1   g439(.A(new_n630), .B(KEYINPUT102), .Z(new_n641));
  INV_X1    g440(.A(new_n641), .ZN(new_n642));
  AOI21_X1  g441(.A(new_n642), .B1(new_n626), .B2(new_n627), .ZN(new_n643));
  OAI21_X1  g442(.A(new_n638), .B1(new_n643), .B2(new_n633), .ZN(new_n644));
  NAND2_X1  g443(.A1(new_n640), .A2(new_n644), .ZN(new_n645));
  INV_X1    g444(.A(new_n645), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n593), .A2(new_n622), .A3(new_n646), .ZN(new_n647));
  NOR3_X1   g446(.A1(new_n492), .A2(new_n560), .A3(new_n647), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n648), .A2(new_n469), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n649), .B(G1gat), .ZN(G1324gat));
  AND2_X1   g449(.A1(new_n648), .A2(new_n356), .ZN(new_n651));
  OAI21_X1  g450(.A(KEYINPUT42), .B1(new_n651), .B2(new_n501), .ZN(new_n652));
  XNOR2_X1  g451(.A(KEYINPUT103), .B(KEYINPUT16), .ZN(new_n653));
  XNOR2_X1  g452(.A(new_n653), .B(new_n501), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n651), .A2(new_n654), .ZN(new_n655));
  MUX2_X1   g454(.A(KEYINPUT42), .B(new_n652), .S(new_n655), .Z(G1325gat));
  AOI21_X1  g455(.A(G15gat), .B1(new_n648), .B2(new_n486), .ZN(new_n657));
  INV_X1    g456(.A(new_n320), .ZN(new_n658));
  AOI21_X1  g457(.A(KEYINPUT36), .B1(new_n313), .B2(new_n319), .ZN(new_n659));
  NOR2_X1   g458(.A1(new_n658), .A2(new_n659), .ZN(new_n660));
  INV_X1    g459(.A(KEYINPUT104), .ZN(new_n661));
  NAND2_X1  g460(.A1(new_n660), .A2(new_n661), .ZN(new_n662));
  OAI21_X1  g461(.A(KEYINPUT104), .B1(new_n658), .B2(new_n659), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n662), .A2(new_n663), .ZN(new_n664));
  AND2_X1   g463(.A1(new_n664), .A2(G15gat), .ZN(new_n665));
  AOI21_X1  g464(.A(new_n657), .B1(new_n648), .B2(new_n665), .ZN(G1326gat));
  NAND2_X1  g465(.A1(new_n648), .A2(new_n465), .ZN(new_n667));
  XNOR2_X1  g466(.A(KEYINPUT43), .B(G22gat), .ZN(new_n668));
  XNOR2_X1  g467(.A(new_n667), .B(new_n668), .ZN(G1327gat));
  NOR3_X1   g468(.A1(new_n356), .A2(new_n476), .A3(new_n427), .ZN(new_n670));
  AOI21_X1  g469(.A(KEYINPUT80), .B1(new_n479), .B2(new_n480), .ZN(new_n671));
  NOR2_X1   g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  OAI211_X1 g471(.A(new_n463), .B(new_n484), .C1(new_n472), .C2(new_n473), .ZN(new_n673));
  OAI21_X1  g472(.A(KEYINPUT82), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  NAND2_X1  g473(.A1(new_n488), .A2(KEYINPUT35), .ZN(new_n675));
  NAND3_X1  g474(.A1(new_n674), .A2(new_n675), .A3(new_n491), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n660), .A2(new_n464), .A3(new_n470), .ZN(new_n677));
  AOI21_X1  g476(.A(new_n622), .B1(new_n676), .B2(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n593), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n679), .A2(new_n646), .ZN(new_n680));
  NOR2_X1   g479(.A1(new_n560), .A2(new_n680), .ZN(new_n681));
  NAND2_X1  g480(.A1(new_n678), .A2(new_n681), .ZN(new_n682));
  INV_X1    g481(.A(new_n682), .ZN(new_n683));
  INV_X1    g482(.A(new_n514), .ZN(new_n684));
  NAND3_X1  g483(.A1(new_n683), .A2(new_n469), .A3(new_n684), .ZN(new_n685));
  XNOR2_X1  g484(.A(new_n685), .B(KEYINPUT45), .ZN(new_n686));
  NOR2_X1   g485(.A1(new_n549), .A2(new_n554), .ZN(new_n687));
  INV_X1    g486(.A(new_n687), .ZN(new_n688));
  NOR2_X1   g487(.A1(new_n680), .A2(new_n688), .ZN(new_n689));
  INV_X1    g488(.A(new_n689), .ZN(new_n690));
  NAND2_X1  g489(.A1(new_n676), .A2(new_n677), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n691), .A2(new_n621), .ZN(new_n692));
  INV_X1    g491(.A(KEYINPUT44), .ZN(new_n693));
  NOR2_X1   g492(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n694));
  NAND2_X1  g493(.A1(new_n692), .A2(new_n694), .ZN(new_n695));
  INV_X1    g494(.A(new_n694), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n693), .A2(KEYINPUT105), .ZN(new_n697));
  INV_X1    g496(.A(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n696), .B1(new_n678), .B2(new_n698), .ZN(new_n699));
  AOI21_X1  g498(.A(new_n690), .B1(new_n695), .B2(new_n699), .ZN(new_n700));
  AND2_X1   g499(.A1(new_n700), .A2(new_n469), .ZN(new_n701));
  OAI21_X1  g500(.A(new_n686), .B1(new_n701), .B2(new_n684), .ZN(G1328gat));
  NOR3_X1   g501(.A1(new_n682), .A2(G36gat), .A3(new_n480), .ZN(new_n703));
  XNOR2_X1  g502(.A(new_n703), .B(KEYINPUT46), .ZN(new_n704));
  AND2_X1   g503(.A1(new_n700), .A2(new_n356), .ZN(new_n705));
  INV_X1    g504(.A(G36gat), .ZN(new_n706));
  OAI21_X1  g505(.A(new_n704), .B1(new_n705), .B2(new_n706), .ZN(G1329gat));
  AOI21_X1  g506(.A(G43gat), .B1(new_n313), .B2(new_n319), .ZN(new_n708));
  NAND3_X1  g507(.A1(new_n678), .A2(new_n681), .A3(new_n708), .ZN(new_n709));
  OR2_X1    g508(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n709), .A2(KEYINPUT106), .ZN(new_n711));
  NAND2_X1  g510(.A1(new_n710), .A2(new_n711), .ZN(new_n712));
  AOI211_X1 g511(.A(new_n660), .B(new_n690), .C1(new_n695), .C2(new_n699), .ZN(new_n713));
  INV_X1    g512(.A(G43gat), .ZN(new_n714));
  OAI211_X1 g513(.A(KEYINPUT47), .B(new_n712), .C1(new_n713), .C2(new_n714), .ZN(new_n715));
  NAND2_X1  g514(.A1(new_n700), .A2(new_n664), .ZN(new_n716));
  AOI22_X1  g515(.A1(new_n716), .A2(G43gat), .B1(new_n711), .B2(new_n710), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n715), .B1(new_n717), .B2(KEYINPUT47), .ZN(G1330gat));
  NAND2_X1  g517(.A1(new_n683), .A2(new_n465), .ZN(new_n719));
  INV_X1    g518(.A(G50gat), .ZN(new_n720));
  INV_X1    g519(.A(KEYINPUT107), .ZN(new_n721));
  AOI22_X1  g520(.A1(new_n719), .A2(new_n720), .B1(new_n721), .B2(KEYINPUT48), .ZN(new_n722));
  NAND3_X1  g521(.A1(new_n700), .A2(G50gat), .A3(new_n465), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n721), .A2(KEYINPUT48), .ZN(new_n724));
  AND3_X1   g523(.A1(new_n722), .A2(new_n723), .A3(new_n724), .ZN(new_n725));
  AOI21_X1  g524(.A(new_n724), .B1(new_n722), .B2(new_n723), .ZN(new_n726));
  NOR2_X1   g525(.A1(new_n725), .A2(new_n726), .ZN(G1331gat));
  NAND3_X1  g526(.A1(new_n688), .A2(new_n593), .A3(new_n622), .ZN(new_n728));
  NOR3_X1   g527(.A1(new_n492), .A2(new_n646), .A3(new_n728), .ZN(new_n729));
  NAND2_X1  g528(.A1(new_n729), .A2(new_n469), .ZN(new_n730));
  XNOR2_X1  g529(.A(new_n730), .B(G57gat), .ZN(G1332gat));
  NOR2_X1   g530(.A1(new_n492), .A2(new_n728), .ZN(new_n732));
  XNOR2_X1  g531(.A(new_n480), .B(KEYINPUT108), .ZN(new_n733));
  INV_X1    g532(.A(new_n733), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n734), .A2(new_n646), .ZN(new_n735));
  NAND2_X1  g534(.A1(new_n732), .A2(new_n735), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n736), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n737));
  XOR2_X1   g536(.A(KEYINPUT49), .B(G64gat), .Z(new_n738));
  OAI21_X1  g537(.A(new_n737), .B1(new_n736), .B2(new_n738), .ZN(G1333gat));
  NAND2_X1  g538(.A1(new_n729), .A2(new_n486), .ZN(new_n740));
  NAND2_X1  g539(.A1(new_n740), .A2(KEYINPUT110), .ZN(new_n741));
  INV_X1    g540(.A(G71gat), .ZN(new_n742));
  INV_X1    g541(.A(KEYINPUT110), .ZN(new_n743));
  NAND3_X1  g542(.A1(new_n729), .A2(new_n743), .A3(new_n486), .ZN(new_n744));
  NAND3_X1  g543(.A1(new_n741), .A2(new_n742), .A3(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(new_n664), .ZN(new_n746));
  NOR2_X1   g545(.A1(new_n746), .A2(new_n742), .ZN(new_n747));
  NAND2_X1  g546(.A1(new_n729), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n748), .A2(KEYINPUT109), .ZN(new_n749));
  INV_X1    g548(.A(KEYINPUT109), .ZN(new_n750));
  NAND3_X1  g549(.A1(new_n729), .A2(new_n750), .A3(new_n747), .ZN(new_n751));
  NAND2_X1  g550(.A1(new_n749), .A2(new_n751), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n745), .A2(new_n752), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n753), .A2(KEYINPUT50), .ZN(new_n754));
  INV_X1    g553(.A(KEYINPUT50), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n745), .A2(new_n752), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g555(.A1(new_n754), .A2(new_n756), .ZN(G1334gat));
  NAND2_X1  g556(.A1(new_n729), .A2(new_n465), .ZN(new_n758));
  XNOR2_X1  g557(.A(KEYINPUT111), .B(G78gat), .ZN(new_n759));
  XNOR2_X1  g558(.A(new_n758), .B(new_n759), .ZN(G1335gat));
  NOR2_X1   g559(.A1(new_n687), .A2(new_n593), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n761), .A2(new_n645), .ZN(new_n762));
  XNOR2_X1  g561(.A(new_n762), .B(KEYINPUT112), .ZN(new_n763));
  AOI21_X1  g562(.A(new_n763), .B1(new_n695), .B2(new_n699), .ZN(new_n764));
  AOI21_X1  g563(.A(new_n595), .B1(new_n764), .B2(new_n469), .ZN(new_n765));
  INV_X1    g564(.A(new_n765), .ZN(new_n766));
  NAND3_X1  g565(.A1(new_n469), .A2(new_n595), .A3(new_n645), .ZN(new_n767));
  XNOR2_X1  g566(.A(new_n767), .B(KEYINPUT114), .ZN(new_n768));
  INV_X1    g567(.A(new_n768), .ZN(new_n769));
  INV_X1    g568(.A(KEYINPUT51), .ZN(new_n770));
  OAI21_X1  g569(.A(new_n761), .B1(new_n678), .B2(KEYINPUT113), .ZN(new_n771));
  INV_X1    g570(.A(KEYINPUT113), .ZN(new_n772));
  AOI211_X1 g571(.A(new_n772), .B(new_n622), .C1(new_n676), .C2(new_n677), .ZN(new_n773));
  OAI21_X1  g572(.A(new_n770), .B1(new_n771), .B2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(new_n772), .B1(new_n492), .B2(new_n622), .ZN(new_n775));
  NAND3_X1  g574(.A1(new_n691), .A2(KEYINPUT113), .A3(new_n621), .ZN(new_n776));
  NAND4_X1  g575(.A1(new_n775), .A2(KEYINPUT51), .A3(new_n761), .A4(new_n776), .ZN(new_n777));
  AOI21_X1  g576(.A(new_n769), .B1(new_n774), .B2(new_n777), .ZN(new_n778));
  INV_X1    g577(.A(new_n778), .ZN(new_n779));
  NAND3_X1  g578(.A1(new_n766), .A2(new_n779), .A3(KEYINPUT115), .ZN(new_n780));
  INV_X1    g579(.A(KEYINPUT115), .ZN(new_n781));
  OAI21_X1  g580(.A(new_n781), .B1(new_n765), .B2(new_n778), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n780), .A2(new_n782), .ZN(G1336gat));
  NAND2_X1  g582(.A1(new_n735), .A2(new_n596), .ZN(new_n784));
  AOI21_X1  g583(.A(new_n784), .B1(new_n774), .B2(new_n777), .ZN(new_n785));
  INV_X1    g584(.A(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n695), .A2(new_n699), .ZN(new_n787));
  INV_X1    g586(.A(new_n763), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n787), .A2(new_n733), .A3(new_n788), .ZN(new_n789));
  NOR2_X1   g588(.A1(new_n596), .A2(KEYINPUT52), .ZN(new_n790));
  NAND2_X1  g589(.A1(new_n789), .A2(new_n790), .ZN(new_n791));
  INV_X1    g590(.A(KEYINPUT116), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n792), .A2(KEYINPUT52), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n786), .A2(new_n791), .A3(new_n793), .ZN(new_n794));
  NAND2_X1  g593(.A1(new_n764), .A2(new_n356), .ZN(new_n795));
  AOI22_X1  g594(.A1(new_n785), .A2(new_n792), .B1(new_n795), .B2(G92gat), .ZN(new_n796));
  INV_X1    g595(.A(KEYINPUT52), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n796), .B2(new_n797), .ZN(G1337gat));
  XOR2_X1   g597(.A(KEYINPUT117), .B(G99gat), .Z(new_n799));
  AOI21_X1  g598(.A(new_n799), .B1(new_n313), .B2(new_n319), .ZN(new_n800));
  INV_X1    g599(.A(new_n761), .ZN(new_n801));
  AOI21_X1  g600(.A(new_n801), .B1(new_n692), .B2(new_n772), .ZN(new_n802));
  AOI21_X1  g601(.A(KEYINPUT51), .B1(new_n802), .B2(new_n776), .ZN(new_n803));
  NOR3_X1   g602(.A1(new_n771), .A2(new_n770), .A3(new_n773), .ZN(new_n804));
  OAI211_X1 g603(.A(new_n645), .B(new_n800), .C1(new_n803), .C2(new_n804), .ZN(new_n805));
  NAND2_X1  g604(.A1(new_n787), .A2(new_n788), .ZN(new_n806));
  OAI21_X1  g605(.A(new_n799), .B1(new_n806), .B2(new_n746), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n805), .A2(new_n807), .ZN(G1338gat));
  NOR2_X1   g607(.A1(new_n463), .A2(G106gat), .ZN(new_n809));
  INV_X1    g608(.A(new_n809), .ZN(new_n810));
  AOI211_X1 g609(.A(new_n646), .B(new_n810), .C1(new_n774), .C2(new_n777), .ZN(new_n811));
  INV_X1    g610(.A(G106gat), .ZN(new_n812));
  AOI21_X1  g611(.A(new_n812), .B1(new_n764), .B2(new_n465), .ZN(new_n813));
  OAI21_X1  g612(.A(KEYINPUT53), .B1(new_n811), .B2(new_n813), .ZN(new_n814));
  OAI211_X1 g613(.A(new_n645), .B(new_n809), .C1(new_n803), .C2(new_n804), .ZN(new_n815));
  OAI21_X1  g614(.A(G106gat), .B1(new_n806), .B2(new_n463), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT53), .ZN(new_n817));
  NAND3_X1  g616(.A1(new_n815), .A2(new_n816), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n814), .A2(new_n818), .ZN(G1339gat));
  INV_X1    g618(.A(new_n483), .ZN(new_n820));
  OAI211_X1 g619(.A(new_n632), .B(KEYINPUT54), .C1(new_n628), .C2(new_n641), .ZN(new_n821));
  INV_X1    g620(.A(KEYINPUT54), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n639), .B1(new_n643), .B2(new_n822), .ZN(new_n823));
  NAND2_X1  g622(.A1(new_n821), .A2(new_n823), .ZN(new_n824));
  INV_X1    g623(.A(KEYINPUT55), .ZN(new_n825));
  NAND3_X1  g624(.A1(new_n824), .A2(KEYINPUT118), .A3(new_n825), .ZN(new_n826));
  OAI21_X1  g625(.A(new_n640), .B1(new_n824), .B2(new_n825), .ZN(new_n827));
  AOI21_X1  g626(.A(KEYINPUT118), .B1(new_n824), .B2(new_n825), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n827), .A2(new_n828), .ZN(new_n829));
  NAND4_X1  g628(.A1(new_n557), .A2(new_n826), .A3(new_n829), .A4(new_n553), .ZN(new_n830));
  AOI21_X1  g629(.A(new_n494), .B1(new_n534), .B2(new_n524), .ZN(new_n831));
  INV_X1    g630(.A(KEYINPUT119), .ZN(new_n832));
  NAND2_X1  g631(.A1(new_n831), .A2(new_n832), .ZN(new_n833));
  OAI21_X1  g632(.A(new_n833), .B1(new_n495), .B2(new_n529), .ZN(new_n834));
  NOR2_X1   g633(.A1(new_n831), .A2(new_n832), .ZN(new_n835));
  OAI21_X1  g634(.A(new_n544), .B1(new_n834), .B2(new_n835), .ZN(new_n836));
  NAND3_X1  g635(.A1(new_n836), .A2(new_n546), .A3(new_n645), .ZN(new_n837));
  AOI21_X1  g636(.A(new_n621), .B1(new_n830), .B2(new_n837), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n829), .A2(new_n621), .A3(new_n826), .ZN(new_n839));
  NAND2_X1  g638(.A1(new_n836), .A2(new_n546), .ZN(new_n840));
  NOR2_X1   g639(.A1(new_n839), .A2(new_n840), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n679), .B1(new_n838), .B2(new_n841), .ZN(new_n842));
  NOR2_X1   g641(.A1(new_n647), .A2(new_n687), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  AOI21_X1  g643(.A(new_n820), .B1(new_n842), .B2(new_n844), .ZN(new_n845));
  NOR2_X1   g644(.A1(new_n733), .A2(new_n468), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n845), .A2(new_n846), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n847), .A2(KEYINPUT120), .ZN(new_n848));
  INV_X1    g647(.A(KEYINPUT120), .ZN(new_n849));
  NAND3_X1  g648(.A1(new_n845), .A2(new_n849), .A3(new_n846), .ZN(new_n850));
  NAND4_X1  g649(.A1(new_n848), .A2(new_n257), .A3(new_n687), .A4(new_n850), .ZN(new_n851));
  OAI21_X1  g650(.A(G113gat), .B1(new_n847), .B2(new_n560), .ZN(new_n852));
  NAND2_X1  g651(.A1(new_n851), .A2(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n853), .A2(KEYINPUT121), .ZN(new_n854));
  INV_X1    g653(.A(KEYINPUT121), .ZN(new_n855));
  NAND3_X1  g654(.A1(new_n851), .A2(new_n855), .A3(new_n852), .ZN(new_n856));
  NAND2_X1  g655(.A1(new_n854), .A2(new_n856), .ZN(G1340gat));
  NAND4_X1  g656(.A1(new_n848), .A2(new_n255), .A3(new_n645), .A4(new_n850), .ZN(new_n858));
  OAI21_X1  g657(.A(G120gat), .B1(new_n847), .B2(new_n646), .ZN(new_n859));
  NAND2_X1  g658(.A1(new_n858), .A2(new_n859), .ZN(G1341gat));
  NAND3_X1  g659(.A1(new_n845), .A2(new_n593), .A3(new_n846), .ZN(new_n861));
  OR2_X1    g660(.A1(new_n861), .A2(new_n249), .ZN(new_n862));
  AND2_X1   g661(.A1(new_n862), .A2(KEYINPUT122), .ZN(new_n863));
  NOR2_X1   g662(.A1(new_n862), .A2(KEYINPUT122), .ZN(new_n864));
  AND2_X1   g663(.A1(new_n861), .A2(new_n249), .ZN(new_n865));
  NOR3_X1   g664(.A1(new_n863), .A2(new_n864), .A3(new_n865), .ZN(G1342gat));
  OAI21_X1  g665(.A(G134gat), .B1(new_n847), .B2(new_n622), .ZN(new_n867));
  OR2_X1    g666(.A1(new_n867), .A2(KEYINPUT124), .ZN(new_n868));
  AOI21_X1  g667(.A(new_n468), .B1(new_n842), .B2(new_n844), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n621), .A2(new_n480), .ZN(new_n870));
  XNOR2_X1  g669(.A(new_n870), .B(KEYINPUT123), .ZN(new_n871));
  NOR3_X1   g670(.A1(new_n871), .A2(G134gat), .A3(new_n820), .ZN(new_n872));
  NAND2_X1  g671(.A1(new_n869), .A2(new_n872), .ZN(new_n873));
  XOR2_X1   g672(.A(new_n873), .B(KEYINPUT56), .Z(new_n874));
  NAND2_X1  g673(.A1(new_n867), .A2(KEYINPUT124), .ZN(new_n875));
  NAND3_X1  g674(.A1(new_n868), .A2(new_n874), .A3(new_n875), .ZN(G1343gat));
  NOR2_X1   g675(.A1(new_n664), .A2(new_n463), .ZN(new_n877));
  NAND2_X1  g676(.A1(new_n869), .A2(new_n877), .ZN(new_n878));
  NOR4_X1   g677(.A1(new_n878), .A2(G141gat), .A3(new_n560), .A4(new_n733), .ZN(new_n879));
  NAND2_X1  g678(.A1(new_n660), .A2(new_n846), .ZN(new_n880));
  INV_X1    g679(.A(new_n880), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT57), .ZN(new_n882));
  NOR2_X1   g681(.A1(new_n463), .A2(new_n882), .ZN(new_n883));
  INV_X1    g682(.A(new_n883), .ZN(new_n884));
  OR2_X1    g683(.A1(new_n824), .A2(KEYINPUT125), .ZN(new_n885));
  AOI21_X1  g684(.A(KEYINPUT55), .B1(new_n824), .B2(KEYINPUT125), .ZN(new_n886));
  AOI21_X1  g685(.A(new_n827), .B1(new_n885), .B2(new_n886), .ZN(new_n887));
  AND3_X1   g686(.A1(new_n557), .A2(KEYINPUT93), .A3(new_n553), .ZN(new_n888));
  AOI21_X1  g687(.A(KEYINPUT93), .B1(new_n557), .B2(new_n553), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n888), .B2(new_n889), .ZN(new_n890));
  AOI21_X1  g689(.A(new_n621), .B1(new_n890), .B2(new_n837), .ZN(new_n891));
  OAI21_X1  g690(.A(new_n679), .B1(new_n891), .B2(new_n841), .ZN(new_n892));
  AOI21_X1  g691(.A(new_n884), .B1(new_n892), .B2(new_n844), .ZN(new_n893));
  NAND2_X1  g692(.A1(new_n842), .A2(new_n844), .ZN(new_n894));
  AOI21_X1  g693(.A(KEYINPUT57), .B1(new_n894), .B2(new_n465), .ZN(new_n895));
  OAI211_X1 g694(.A(new_n687), .B(new_n881), .C1(new_n893), .C2(new_n895), .ZN(new_n896));
  AOI21_X1  g695(.A(new_n879), .B1(new_n896), .B2(G141gat), .ZN(new_n897));
  INV_X1    g696(.A(KEYINPUT58), .ZN(new_n898));
  INV_X1    g697(.A(new_n887), .ZN(new_n899));
  AOI21_X1  g698(.A(new_n899), .B1(new_n555), .B2(new_n558), .ZN(new_n900));
  INV_X1    g699(.A(new_n837), .ZN(new_n901));
  OAI21_X1  g700(.A(new_n622), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  INV_X1    g701(.A(new_n841), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n593), .B1(new_n902), .B2(new_n903), .ZN(new_n904));
  OAI21_X1  g703(.A(new_n883), .B1(new_n904), .B2(new_n843), .ZN(new_n905));
  NAND2_X1  g704(.A1(new_n894), .A2(new_n465), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n906), .A2(new_n882), .ZN(new_n907));
  AOI21_X1  g706(.A(new_n880), .B1(new_n905), .B2(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(new_n364), .B1(new_n908), .B2(new_n559), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n878), .A2(new_n733), .ZN(new_n910));
  NAND3_X1  g709(.A1(new_n910), .A2(new_n364), .A3(new_n559), .ZN(new_n911));
  NAND2_X1  g710(.A1(new_n911), .A2(new_n898), .ZN(new_n912));
  OAI22_X1  g711(.A1(new_n897), .A2(new_n898), .B1(new_n909), .B2(new_n912), .ZN(G1344gat));
  NAND3_X1  g712(.A1(new_n910), .A2(new_n366), .A3(new_n645), .ZN(new_n914));
  INV_X1    g713(.A(KEYINPUT59), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(G148gat), .ZN(new_n916));
  AOI21_X1  g715(.A(new_n916), .B1(new_n908), .B2(new_n645), .ZN(new_n917));
  NOR2_X1   g716(.A1(new_n463), .A2(KEYINPUT57), .ZN(new_n918));
  INV_X1    g717(.A(KEYINPUT126), .ZN(new_n919));
  OR3_X1    g718(.A1(new_n559), .A2(new_n919), .A3(new_n647), .ZN(new_n920));
  OAI21_X1  g719(.A(new_n919), .B1(new_n559), .B2(new_n647), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(new_n922));
  OAI21_X1  g721(.A(new_n918), .B1(new_n904), .B2(new_n922), .ZN(new_n923));
  NAND2_X1  g722(.A1(new_n906), .A2(KEYINPUT57), .ZN(new_n924));
  NAND4_X1  g723(.A1(new_n923), .A2(new_n924), .A3(new_n645), .A4(new_n881), .ZN(new_n925));
  AOI21_X1  g724(.A(new_n915), .B1(new_n925), .B2(G148gat), .ZN(new_n926));
  OAI21_X1  g725(.A(new_n914), .B1(new_n917), .B2(new_n926), .ZN(G1345gat));
  AOI21_X1  g726(.A(G155gat), .B1(new_n910), .B2(new_n593), .ZN(new_n928));
  NOR2_X1   g727(.A1(new_n679), .A2(new_n370), .ZN(new_n929));
  AOI21_X1  g728(.A(new_n928), .B1(new_n908), .B2(new_n929), .ZN(G1346gat));
  AOI21_X1  g729(.A(new_n371), .B1(new_n908), .B2(new_n621), .ZN(new_n931));
  NOR3_X1   g730(.A1(new_n878), .A2(G162gat), .A3(new_n871), .ZN(new_n932));
  OR2_X1    g731(.A1(new_n931), .A2(new_n932), .ZN(G1347gat));
  NOR2_X1   g732(.A1(new_n734), .A2(new_n469), .ZN(new_n934));
  AND2_X1   g733(.A1(new_n845), .A2(new_n934), .ZN(new_n935));
  NAND3_X1  g734(.A1(new_n935), .A2(new_n203), .A3(new_n687), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n469), .A2(new_n480), .ZN(new_n937));
  XOR2_X1   g736(.A(new_n937), .B(KEYINPUT127), .Z(new_n938));
  INV_X1    g737(.A(new_n938), .ZN(new_n939));
  NAND2_X1  g738(.A1(new_n845), .A2(new_n939), .ZN(new_n940));
  OAI21_X1  g739(.A(G169gat), .B1(new_n940), .B2(new_n560), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n936), .A2(new_n941), .ZN(G1348gat));
  AOI21_X1  g741(.A(G176gat), .B1(new_n935), .B2(new_n645), .ZN(new_n943));
  NOR3_X1   g742(.A1(new_n940), .A2(new_n204), .A3(new_n646), .ZN(new_n944));
  NOR2_X1   g743(.A1(new_n943), .A2(new_n944), .ZN(G1349gat));
  NAND3_X1  g744(.A1(new_n935), .A2(new_n211), .A3(new_n593), .ZN(new_n946));
  OAI21_X1  g745(.A(G183gat), .B1(new_n940), .B2(new_n679), .ZN(new_n947));
  NAND2_X1  g746(.A1(new_n946), .A2(new_n947), .ZN(new_n948));
  XNOR2_X1  g747(.A(new_n948), .B(KEYINPUT60), .ZN(G1350gat));
  NAND3_X1  g748(.A1(new_n935), .A2(new_n212), .A3(new_n621), .ZN(new_n950));
  OAI21_X1  g749(.A(G190gat), .B1(new_n940), .B2(new_n622), .ZN(new_n951));
  AND2_X1   g750(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n952));
  NOR2_X1   g751(.A1(new_n951), .A2(KEYINPUT61), .ZN(new_n953));
  OAI21_X1  g752(.A(new_n950), .B1(new_n952), .B2(new_n953), .ZN(G1351gat));
  NOR2_X1   g753(.A1(new_n664), .A2(new_n938), .ZN(new_n955));
  AND3_X1   g754(.A1(new_n923), .A2(new_n924), .A3(new_n955), .ZN(new_n956));
  NAND2_X1  g755(.A1(new_n956), .A2(new_n559), .ZN(new_n957));
  NAND2_X1  g756(.A1(new_n957), .A2(G197gat), .ZN(new_n958));
  AND2_X1   g757(.A1(new_n894), .A2(new_n934), .ZN(new_n959));
  NAND2_X1  g758(.A1(new_n959), .A2(new_n877), .ZN(new_n960));
  OR3_X1    g759(.A1(new_n960), .A2(G197gat), .A3(new_n688), .ZN(new_n961));
  NAND2_X1  g760(.A1(new_n958), .A2(new_n961), .ZN(G1352gat));
  NOR2_X1   g761(.A1(new_n646), .A2(G204gat), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n959), .A2(new_n877), .A3(new_n963), .ZN(new_n964));
  XOR2_X1   g763(.A(new_n964), .B(KEYINPUT62), .Z(new_n965));
  NAND4_X1  g764(.A1(new_n923), .A2(new_n924), .A3(new_n645), .A4(new_n955), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n966), .A2(G204gat), .ZN(new_n967));
  NAND2_X1  g766(.A1(new_n965), .A2(new_n967), .ZN(G1353gat));
  OR3_X1    g767(.A1(new_n960), .A2(G211gat), .A3(new_n679), .ZN(new_n969));
  NAND4_X1  g768(.A1(new_n923), .A2(new_n924), .A3(new_n593), .A4(new_n955), .ZN(new_n970));
  AND3_X1   g769(.A1(new_n970), .A2(KEYINPUT63), .A3(G211gat), .ZN(new_n971));
  AOI21_X1  g770(.A(KEYINPUT63), .B1(new_n970), .B2(G211gat), .ZN(new_n972));
  OAI21_X1  g771(.A(new_n969), .B1(new_n971), .B2(new_n972), .ZN(G1354gat));
  NAND3_X1  g772(.A1(new_n956), .A2(G218gat), .A3(new_n621), .ZN(new_n974));
  INV_X1    g773(.A(G218gat), .ZN(new_n975));
  OAI21_X1  g774(.A(new_n975), .B1(new_n960), .B2(new_n622), .ZN(new_n976));
  AND2_X1   g775(.A1(new_n974), .A2(new_n976), .ZN(G1355gat));
endmodule


