//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 0 0 0 1 1 1 0 0 1 1 0 1 1 0 0 0 1 0 0 0 1 1 1 1 0 1 0 1 1 0 1 1 0 0 1 1 1 0 0 1 0 1 0 1 0 1 0 0 1 1 1 0 0 1 1 0 0 0 0 0 0 0 0 1' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:29:08 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n459, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n472,
    new_n473, new_n474, new_n475, new_n476, new_n477, new_n478, new_n479,
    new_n480, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n515, new_n516, new_n517,
    new_n518, new_n519, new_n520, new_n521, new_n522, new_n523, new_n524,
    new_n525, new_n526, new_n527, new_n528, new_n529, new_n530, new_n531,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n539, new_n540,
    new_n541, new_n542, new_n543, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n563, new_n564, new_n566, new_n567,
    new_n568, new_n569, new_n570, new_n571, new_n572, new_n574, new_n575,
    new_n577, new_n578, new_n579, new_n580, new_n582, new_n583, new_n584,
    new_n585, new_n586, new_n587, new_n588, new_n589, new_n590, new_n591,
    new_n593, new_n594, new_n595, new_n596, new_n597, new_n598, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n619, new_n620, new_n623, new_n625, new_n626,
    new_n627, new_n628, new_n629, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n653, new_n654, new_n655, new_n656, new_n657,
    new_n658, new_n659, new_n660, new_n661, new_n662, new_n663, new_n664,
    new_n665, new_n666, new_n667, new_n668, new_n669, new_n670, new_n671,
    new_n672, new_n673, new_n674, new_n675, new_n677, new_n678, new_n679,
    new_n680, new_n681, new_n682, new_n683, new_n684, new_n685, new_n686,
    new_n687, new_n688, new_n689, new_n690, new_n691, new_n692, new_n693,
    new_n694, new_n695, new_n696, new_n697, new_n698, new_n699, new_n701,
    new_n702, new_n703, new_n704, new_n705, new_n706, new_n707, new_n708,
    new_n709, new_n710, new_n711, new_n712, new_n713, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n822, new_n823, new_n824, new_n825, new_n826, new_n827, new_n828,
    new_n829, new_n830, new_n831, new_n832, new_n833, new_n834, new_n835,
    new_n836, new_n837, new_n838, new_n839, new_n840, new_n841, new_n842,
    new_n843, new_n844, new_n845, new_n846, new_n847, new_n848, new_n849,
    new_n850, new_n851, new_n852, new_n853, new_n854, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n880, new_n881, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n914, new_n915,
    new_n916, new_n917, new_n918, new_n919, new_n920, new_n921, new_n922,
    new_n923, new_n924, new_n925, new_n926, new_n927, new_n928, new_n929,
    new_n930, new_n931, new_n932, new_n933, new_n935, new_n936, new_n937,
    new_n938, new_n939, new_n940, new_n941, new_n942, new_n943, new_n944,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n976, new_n977, new_n978, new_n979, new_n980, new_n981,
    new_n982, new_n983, new_n984, new_n985, new_n986, new_n987, new_n988,
    new_n989, new_n990, new_n991, new_n992, new_n993, new_n994, new_n995,
    new_n996, new_n997, new_n998, new_n999, new_n1000, new_n1001,
    new_n1002, new_n1003, new_n1004, new_n1005, new_n1006, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1185, new_n1186, new_n1187, new_n1188,
    new_n1189, new_n1190, new_n1191, new_n1192, new_n1193, new_n1194,
    new_n1195, new_n1196, new_n1197, new_n1198, new_n1199, new_n1200,
    new_n1201, new_n1202, new_n1203, new_n1204, new_n1205, new_n1206,
    new_n1207, new_n1208, new_n1211, new_n1212, new_n1213, new_n1214,
    new_n1215, new_n1216, new_n1217, new_n1218, new_n1219;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  XOR2_X1   g002(.A(KEYINPUT64), .B(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  XOR2_X1   g007(.A(KEYINPUT65), .B(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  XNOR2_X1  g015(.A(KEYINPUT66), .B(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  XNOR2_X1  g018(.A(KEYINPUT67), .B(G452), .ZN(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XNOR2_X1  g025(.A(new_n450), .B(KEYINPUT2), .ZN(new_n451));
  NOR4_X1   g026(.A1(G238), .A2(G237), .A3(G235), .A4(G236), .ZN(new_n452));
  NAND2_X1  g027(.A1(new_n451), .A2(new_n452), .ZN(G261));
  INV_X1    g028(.A(G261), .ZN(G325));
  INV_X1    g029(.A(G567), .ZN(new_n455));
  NOR2_X1   g030(.A1(new_n452), .A2(new_n455), .ZN(new_n456));
  INV_X1    g031(.A(new_n451), .ZN(new_n457));
  AOI21_X1  g032(.A(new_n456), .B1(new_n457), .B2(G2106), .ZN(G319));
  INV_X1    g033(.A(G2105), .ZN(new_n459));
  AND2_X1   g034(.A1(G113), .A2(G2104), .ZN(new_n460));
  AND2_X1   g035(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n461));
  NOR2_X1   g036(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n462));
  OAI21_X1  g037(.A(G125), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g038(.A(KEYINPUT68), .ZN(new_n464));
  AOI21_X1  g039(.A(new_n460), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  OR2_X1    g040(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n466));
  NAND2_X1  g041(.A1(KEYINPUT3), .A2(G2104), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n466), .A2(new_n467), .ZN(new_n468));
  NAND3_X1  g043(.A1(new_n468), .A2(KEYINPUT68), .A3(G125), .ZN(new_n469));
  AOI21_X1  g044(.A(new_n459), .B1(new_n465), .B2(new_n469), .ZN(new_n470));
  INV_X1    g045(.A(G2104), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n471), .A2(G2105), .ZN(new_n472));
  INV_X1    g047(.A(KEYINPUT69), .ZN(new_n473));
  AND3_X1   g048(.A1(new_n472), .A2(new_n473), .A3(G101), .ZN(new_n474));
  AOI21_X1  g049(.A(new_n473), .B1(new_n472), .B2(G101), .ZN(new_n475));
  INV_X1    g050(.A(G137), .ZN(new_n476));
  OAI21_X1  g051(.A(new_n459), .B1(new_n461), .B2(new_n462), .ZN(new_n477));
  OAI22_X1  g052(.A1(new_n474), .A2(new_n475), .B1(new_n476), .B2(new_n477), .ZN(new_n478));
  NOR2_X1   g053(.A1(new_n470), .A2(new_n478), .ZN(new_n479));
  INV_X1    g054(.A(KEYINPUT70), .ZN(new_n480));
  XNOR2_X1  g055(.A(new_n479), .B(new_n480), .ZN(G160));
  INV_X1    g056(.A(KEYINPUT71), .ZN(new_n482));
  NAND2_X1  g057(.A1(new_n468), .A2(new_n482), .ZN(new_n483));
  NOR2_X1   g058(.A1(new_n461), .A2(new_n462), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(KEYINPUT71), .ZN(new_n485));
  AOI21_X1  g060(.A(G2105), .B1(new_n483), .B2(new_n485), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n486), .A2(G136), .ZN(new_n487));
  AOI21_X1  g062(.A(new_n459), .B1(new_n483), .B2(new_n485), .ZN(new_n488));
  NAND2_X1  g063(.A1(new_n488), .A2(G124), .ZN(new_n489));
  NOR2_X1   g064(.A1(G100), .A2(G2105), .ZN(new_n490));
  OAI21_X1  g065(.A(G2104), .B1(new_n459), .B2(G112), .ZN(new_n491));
  OAI211_X1 g066(.A(new_n487), .B(new_n489), .C1(new_n490), .C2(new_n491), .ZN(new_n492));
  XOR2_X1   g067(.A(new_n492), .B(KEYINPUT72), .Z(G162));
  NAND2_X1  g068(.A1(G126), .A2(G2105), .ZN(new_n494));
  NAND2_X1  g069(.A1(KEYINPUT75), .A2(G138), .ZN(new_n495));
  OAI21_X1  g070(.A(new_n494), .B1(new_n495), .B2(G2105), .ZN(new_n496));
  INV_X1    g071(.A(KEYINPUT4), .ZN(new_n497));
  NOR2_X1   g072(.A1(new_n497), .A2(KEYINPUT74), .ZN(new_n498));
  NAND3_X1  g073(.A1(new_n468), .A2(new_n496), .A3(new_n498), .ZN(new_n499));
  INV_X1    g074(.A(KEYINPUT73), .ZN(new_n500));
  OAI21_X1  g075(.A(new_n500), .B1(new_n459), .B2(G114), .ZN(new_n501));
  INV_X1    g076(.A(G114), .ZN(new_n502));
  NAND3_X1  g077(.A1(new_n502), .A2(KEYINPUT73), .A3(G2105), .ZN(new_n503));
  OR2_X1    g078(.A1(G102), .A2(G2105), .ZN(new_n504));
  NAND4_X1  g079(.A1(new_n501), .A2(new_n503), .A3(new_n504), .A4(G2104), .ZN(new_n505));
  OAI21_X1  g080(.A(G138), .B1(KEYINPUT75), .B2(KEYINPUT4), .ZN(new_n506));
  NOR2_X1   g081(.A1(new_n477), .A2(new_n506), .ZN(new_n507));
  OAI211_X1 g082(.A(new_n499), .B(new_n505), .C1(new_n507), .C2(new_n498), .ZN(new_n508));
  INV_X1    g083(.A(new_n508), .ZN(G164));
  INV_X1    g084(.A(KEYINPUT77), .ZN(new_n510));
  NAND2_X1  g085(.A1(KEYINPUT76), .A2(G543), .ZN(new_n511));
  NAND2_X1  g086(.A1(new_n511), .A2(KEYINPUT5), .ZN(new_n512));
  INV_X1    g087(.A(KEYINPUT5), .ZN(new_n513));
  NAND3_X1  g088(.A1(new_n513), .A2(KEYINPUT76), .A3(G543), .ZN(new_n514));
  NAND2_X1  g089(.A1(new_n512), .A2(new_n514), .ZN(new_n515));
  INV_X1    g090(.A(G651), .ZN(new_n516));
  NAND2_X1  g091(.A1(new_n516), .A2(KEYINPUT6), .ZN(new_n517));
  INV_X1    g092(.A(KEYINPUT6), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(G651), .ZN(new_n519));
  NAND2_X1  g094(.A1(new_n517), .A2(new_n519), .ZN(new_n520));
  OAI21_X1  g095(.A(new_n510), .B1(new_n515), .B2(new_n520), .ZN(new_n521));
  XNOR2_X1  g096(.A(KEYINPUT6), .B(G651), .ZN(new_n522));
  NAND4_X1  g097(.A1(new_n522), .A2(KEYINPUT77), .A3(new_n512), .A4(new_n514), .ZN(new_n523));
  AND2_X1   g098(.A1(new_n521), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g099(.A1(new_n524), .A2(G88), .ZN(new_n525));
  NAND2_X1  g100(.A1(G75), .A2(G543), .ZN(new_n526));
  INV_X1    g101(.A(G62), .ZN(new_n527));
  OAI21_X1  g102(.A(new_n526), .B1(new_n515), .B2(new_n527), .ZN(new_n528));
  INV_X1    g103(.A(G543), .ZN(new_n529));
  NOR2_X1   g104(.A1(new_n520), .A2(new_n529), .ZN(new_n530));
  AOI22_X1  g105(.A1(new_n528), .A2(G651), .B1(new_n530), .B2(G50), .ZN(new_n531));
  NAND2_X1  g106(.A1(new_n525), .A2(new_n531), .ZN(G303));
  INV_X1    g107(.A(G303), .ZN(G166));
  NAND3_X1  g108(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n534));
  NAND2_X1  g109(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n535));
  OR2_X1    g110(.A1(new_n534), .A2(KEYINPUT7), .ZN(new_n536));
  AOI22_X1  g111(.A1(new_n530), .A2(G51), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n538));
  NAND2_X1  g113(.A1(new_n515), .A2(new_n538), .ZN(new_n539));
  NAND3_X1  g114(.A1(new_n512), .A2(new_n514), .A3(KEYINPUT78), .ZN(new_n540));
  NAND4_X1  g115(.A1(new_n539), .A2(G63), .A3(G651), .A4(new_n540), .ZN(new_n541));
  NAND2_X1  g116(.A1(new_n521), .A2(new_n523), .ZN(new_n542));
  INV_X1    g117(.A(G89), .ZN(new_n543));
  OAI211_X1 g118(.A(new_n537), .B(new_n541), .C1(new_n542), .C2(new_n543), .ZN(G286));
  INV_X1    g119(.A(G286), .ZN(G168));
  NAND2_X1  g120(.A1(new_n530), .A2(G52), .ZN(new_n546));
  INV_X1    g121(.A(G90), .ZN(new_n547));
  OAI21_X1  g122(.A(new_n546), .B1(new_n542), .B2(new_n547), .ZN(new_n548));
  NAND3_X1  g123(.A1(new_n539), .A2(G64), .A3(new_n540), .ZN(new_n549));
  NAND2_X1  g124(.A1(G77), .A2(G543), .ZN(new_n550));
  AOI21_X1  g125(.A(new_n516), .B1(new_n549), .B2(new_n550), .ZN(new_n551));
  NOR2_X1   g126(.A1(new_n548), .A2(new_n551), .ZN(G171));
  NAND2_X1  g127(.A1(new_n530), .A2(G43), .ZN(new_n553));
  INV_X1    g128(.A(G81), .ZN(new_n554));
  OAI21_X1  g129(.A(new_n553), .B1(new_n542), .B2(new_n554), .ZN(new_n555));
  NAND3_X1  g130(.A1(new_n539), .A2(G56), .A3(new_n540), .ZN(new_n556));
  NAND2_X1  g131(.A1(G68), .A2(G543), .ZN(new_n557));
  AOI21_X1  g132(.A(new_n516), .B1(new_n556), .B2(new_n557), .ZN(new_n558));
  NOR2_X1   g133(.A1(new_n555), .A2(new_n558), .ZN(new_n559));
  NAND2_X1  g134(.A1(new_n559), .A2(G860), .ZN(new_n560));
  XOR2_X1   g135(.A(new_n560), .B(KEYINPUT79), .Z(G153));
  NAND4_X1  g136(.A1(G319), .A2(G36), .A3(G483), .A4(G661), .ZN(G176));
  NAND2_X1  g137(.A1(G1), .A2(G3), .ZN(new_n563));
  XNOR2_X1  g138(.A(new_n563), .B(KEYINPUT8), .ZN(new_n564));
  NAND4_X1  g139(.A1(G319), .A2(G483), .A3(G661), .A4(new_n564), .ZN(G188));
  NAND4_X1  g140(.A1(new_n517), .A2(new_n519), .A3(G53), .A4(G543), .ZN(new_n566));
  XNOR2_X1  g141(.A(new_n566), .B(KEYINPUT9), .ZN(new_n567));
  NAND2_X1  g142(.A1(G78), .A2(G543), .ZN(new_n568));
  INV_X1    g143(.A(G65), .ZN(new_n569));
  OAI21_X1  g144(.A(new_n568), .B1(new_n515), .B2(new_n569), .ZN(new_n570));
  NAND2_X1  g145(.A1(new_n570), .A2(G651), .ZN(new_n571));
  INV_X1    g146(.A(G91), .ZN(new_n572));
  OAI211_X1 g147(.A(new_n567), .B(new_n571), .C1(new_n572), .C2(new_n542), .ZN(G299));
  AOI22_X1  g148(.A1(new_n524), .A2(G90), .B1(G52), .B2(new_n530), .ZN(new_n574));
  INV_X1    g149(.A(new_n551), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n574), .A2(new_n575), .ZN(G301));
  AND2_X1   g151(.A1(new_n539), .A2(new_n540), .ZN(new_n577));
  OAI21_X1  g152(.A(G651), .B1(new_n577), .B2(G74), .ZN(new_n578));
  NAND2_X1  g153(.A1(new_n524), .A2(G87), .ZN(new_n579));
  NAND2_X1  g154(.A1(new_n530), .A2(G49), .ZN(new_n580));
  NAND3_X1  g155(.A1(new_n578), .A2(new_n579), .A3(new_n580), .ZN(G288));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  INV_X1    g157(.A(G61), .ZN(new_n583));
  OAI21_X1  g158(.A(new_n582), .B1(new_n515), .B2(new_n583), .ZN(new_n584));
  AND3_X1   g159(.A1(new_n584), .A2(KEYINPUT80), .A3(G651), .ZN(new_n585));
  AOI21_X1  g160(.A(KEYINPUT80), .B1(new_n584), .B2(G651), .ZN(new_n586));
  NOR2_X1   g161(.A1(new_n585), .A2(new_n586), .ZN(new_n587));
  NAND3_X1  g162(.A1(new_n521), .A2(G86), .A3(new_n523), .ZN(new_n588));
  NAND2_X1  g163(.A1(new_n530), .A2(G48), .ZN(new_n589));
  NAND2_X1  g164(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  INV_X1    g165(.A(new_n590), .ZN(new_n591));
  NAND2_X1  g166(.A1(new_n587), .A2(new_n591), .ZN(G305));
  AOI22_X1  g167(.A1(new_n577), .A2(G60), .B1(G72), .B2(G543), .ZN(new_n593));
  NOR2_X1   g168(.A1(new_n593), .A2(new_n516), .ZN(new_n594));
  NAND2_X1  g169(.A1(new_n530), .A2(G47), .ZN(new_n595));
  INV_X1    g170(.A(G85), .ZN(new_n596));
  OAI21_X1  g171(.A(new_n595), .B1(new_n542), .B2(new_n596), .ZN(new_n597));
  NOR2_X1   g172(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g173(.A(new_n598), .ZN(G290));
  NAND2_X1  g174(.A1(G301), .A2(G868), .ZN(new_n600));
  NAND2_X1  g175(.A1(G79), .A2(G543), .ZN(new_n601));
  INV_X1    g176(.A(G66), .ZN(new_n602));
  OAI21_X1  g177(.A(new_n601), .B1(new_n515), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g178(.A1(new_n603), .A2(G651), .ZN(new_n604));
  NAND2_X1  g179(.A1(new_n530), .A2(G54), .ZN(new_n605));
  AND2_X1   g180(.A1(new_n604), .A2(new_n605), .ZN(new_n606));
  INV_X1    g181(.A(new_n606), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n521), .A2(G92), .A3(new_n523), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n608), .A2(KEYINPUT81), .ZN(new_n609));
  INV_X1    g184(.A(KEYINPUT81), .ZN(new_n610));
  NAND4_X1  g185(.A1(new_n521), .A2(new_n610), .A3(G92), .A4(new_n523), .ZN(new_n611));
  NAND2_X1  g186(.A1(new_n609), .A2(new_n611), .ZN(new_n612));
  NAND2_X1  g187(.A1(new_n612), .A2(KEYINPUT10), .ZN(new_n613));
  INV_X1    g188(.A(KEYINPUT10), .ZN(new_n614));
  NAND3_X1  g189(.A1(new_n609), .A2(new_n614), .A3(new_n611), .ZN(new_n615));
  AOI21_X1  g190(.A(new_n607), .B1(new_n613), .B2(new_n615), .ZN(new_n616));
  OAI21_X1  g191(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G284));
  OAI21_X1  g192(.A(new_n600), .B1(new_n616), .B2(G868), .ZN(G321));
  NAND2_X1  g193(.A1(G286), .A2(G868), .ZN(new_n619));
  INV_X1    g194(.A(G299), .ZN(new_n620));
  OAI21_X1  g195(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G297));
  OAI21_X1  g196(.A(new_n619), .B1(new_n620), .B2(G868), .ZN(G280));
  INV_X1    g197(.A(G559), .ZN(new_n623));
  OAI21_X1  g198(.A(new_n616), .B1(new_n623), .B2(G860), .ZN(G148));
  NAND2_X1  g199(.A1(new_n616), .A2(new_n623), .ZN(new_n625));
  NAND2_X1  g200(.A1(new_n625), .A2(G868), .ZN(new_n626));
  INV_X1    g201(.A(G868), .ZN(new_n627));
  INV_X1    g202(.A(new_n559), .ZN(new_n628));
  AOI22_X1  g203(.A1(new_n626), .A2(KEYINPUT82), .B1(new_n627), .B2(new_n628), .ZN(new_n629));
  OAI21_X1  g204(.A(new_n629), .B1(KEYINPUT82), .B2(new_n626), .ZN(G323));
  XNOR2_X1  g205(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g206(.A1(new_n486), .A2(G135), .ZN(new_n632));
  NAND2_X1  g207(.A1(new_n488), .A2(G123), .ZN(new_n633));
  NOR2_X1   g208(.A1(G99), .A2(G2105), .ZN(new_n634));
  OAI21_X1  g209(.A(G2104), .B1(new_n459), .B2(G111), .ZN(new_n635));
  OAI211_X1 g210(.A(new_n632), .B(new_n633), .C1(new_n634), .C2(new_n635), .ZN(new_n636));
  XNOR2_X1  g211(.A(new_n636), .B(KEYINPUT84), .ZN(new_n637));
  XOR2_X1   g212(.A(new_n637), .B(G2096), .Z(new_n638));
  NAND2_X1  g213(.A1(new_n468), .A2(new_n472), .ZN(new_n639));
  XOR2_X1   g214(.A(KEYINPUT83), .B(KEYINPUT12), .Z(new_n640));
  XNOR2_X1  g215(.A(new_n639), .B(new_n640), .ZN(new_n641));
  XNOR2_X1  g216(.A(KEYINPUT13), .B(G2100), .ZN(new_n642));
  XNOR2_X1  g217(.A(new_n641), .B(new_n642), .ZN(new_n643));
  NAND2_X1  g218(.A1(new_n638), .A2(new_n643), .ZN(G156));
  XNOR2_X1  g219(.A(G2451), .B(G2454), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n645), .B(KEYINPUT16), .ZN(new_n646));
  INV_X1    g221(.A(new_n646), .ZN(new_n647));
  XNOR2_X1  g222(.A(G2443), .B(G2446), .ZN(new_n648));
  INV_X1    g223(.A(new_n648), .ZN(new_n649));
  XNOR2_X1  g224(.A(G1341), .B(G1348), .ZN(new_n650));
  XOR2_X1   g225(.A(new_n650), .B(KEYINPUT87), .Z(new_n651));
  INV_X1    g226(.A(new_n651), .ZN(new_n652));
  XNOR2_X1  g227(.A(KEYINPUT85), .B(KEYINPUT14), .ZN(new_n653));
  XNOR2_X1  g228(.A(KEYINPUT15), .B(G2435), .ZN(new_n654));
  XNOR2_X1  g229(.A(new_n654), .B(G2438), .ZN(new_n655));
  INV_X1    g230(.A(new_n655), .ZN(new_n656));
  XNOR2_X1  g231(.A(G2427), .B(G2430), .ZN(new_n657));
  INV_X1    g232(.A(new_n657), .ZN(new_n658));
  OAI21_X1  g233(.A(new_n653), .B1(new_n656), .B2(new_n658), .ZN(new_n659));
  XOR2_X1   g234(.A(new_n659), .B(KEYINPUT86), .Z(new_n660));
  NAND2_X1  g235(.A1(new_n656), .A2(new_n658), .ZN(new_n661));
  AOI21_X1  g236(.A(new_n652), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  INV_X1    g237(.A(new_n662), .ZN(new_n663));
  NAND3_X1  g238(.A1(new_n660), .A2(new_n652), .A3(new_n661), .ZN(new_n664));
  AOI21_X1  g239(.A(new_n649), .B1(new_n663), .B2(new_n664), .ZN(new_n665));
  INV_X1    g240(.A(new_n664), .ZN(new_n666));
  NOR3_X1   g241(.A1(new_n666), .A2(new_n648), .A3(new_n662), .ZN(new_n667));
  OAI21_X1  g242(.A(new_n647), .B1(new_n665), .B2(new_n667), .ZN(new_n668));
  OAI21_X1  g243(.A(new_n648), .B1(new_n666), .B2(new_n662), .ZN(new_n669));
  NAND3_X1  g244(.A1(new_n663), .A2(new_n649), .A3(new_n664), .ZN(new_n670));
  NAND3_X1  g245(.A1(new_n669), .A2(new_n670), .A3(new_n646), .ZN(new_n671));
  NAND3_X1  g246(.A1(new_n668), .A2(G14), .A3(new_n671), .ZN(new_n672));
  INV_X1    g247(.A(KEYINPUT88), .ZN(new_n673));
  NAND2_X1  g248(.A1(new_n672), .A2(new_n673), .ZN(new_n674));
  NAND4_X1  g249(.A1(new_n668), .A2(KEYINPUT88), .A3(G14), .A4(new_n671), .ZN(new_n675));
  AND2_X1   g250(.A1(new_n674), .A2(new_n675), .ZN(G401));
  INV_X1    g251(.A(G2100), .ZN(new_n677));
  XOR2_X1   g252(.A(G2072), .B(G2078), .Z(new_n678));
  XNOR2_X1  g253(.A(new_n678), .B(KEYINPUT17), .ZN(new_n679));
  XNOR2_X1  g254(.A(G2067), .B(G2678), .ZN(new_n680));
  XNOR2_X1  g255(.A(new_n680), .B(KEYINPUT90), .ZN(new_n681));
  XOR2_X1   g256(.A(G2084), .B(G2090), .Z(new_n682));
  NAND3_X1  g257(.A1(new_n679), .A2(new_n681), .A3(new_n682), .ZN(new_n683));
  NAND2_X1  g258(.A1(new_n682), .A2(new_n680), .ZN(new_n684));
  NOR2_X1   g259(.A1(new_n684), .A2(new_n678), .ZN(new_n685));
  XNOR2_X1  g260(.A(KEYINPUT89), .B(KEYINPUT18), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n685), .B(new_n686), .ZN(new_n687));
  AOI21_X1  g262(.A(new_n682), .B1(new_n681), .B2(new_n678), .ZN(new_n688));
  OAI21_X1  g263(.A(new_n688), .B1(new_n681), .B2(new_n679), .ZN(new_n689));
  AND2_X1   g264(.A1(new_n689), .A2(KEYINPUT91), .ZN(new_n690));
  NOR2_X1   g265(.A1(new_n689), .A2(KEYINPUT91), .ZN(new_n691));
  OAI211_X1 g266(.A(new_n683), .B(new_n687), .C1(new_n690), .C2(new_n691), .ZN(new_n692));
  NAND2_X1  g267(.A1(new_n692), .A2(G2096), .ZN(new_n693));
  INV_X1    g268(.A(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(new_n692), .A2(G2096), .ZN(new_n695));
  OAI21_X1  g270(.A(new_n677), .B1(new_n694), .B2(new_n695), .ZN(new_n696));
  INV_X1    g271(.A(new_n695), .ZN(new_n697));
  NAND3_X1  g272(.A1(new_n697), .A2(G2100), .A3(new_n693), .ZN(new_n698));
  AND2_X1   g273(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(new_n699), .ZN(G227));
  XNOR2_X1  g275(.A(G1971), .B(G1976), .ZN(new_n701));
  INV_X1    g276(.A(KEYINPUT19), .ZN(new_n702));
  XNOR2_X1  g277(.A(new_n701), .B(new_n702), .ZN(new_n703));
  XOR2_X1   g278(.A(G1956), .B(G2474), .Z(new_n704));
  XOR2_X1   g279(.A(G1961), .B(G1966), .Z(new_n705));
  AND2_X1   g280(.A1(new_n704), .A2(new_n705), .ZN(new_n706));
  NAND2_X1  g281(.A1(new_n703), .A2(new_n706), .ZN(new_n707));
  XNOR2_X1  g282(.A(new_n707), .B(KEYINPUT20), .ZN(new_n708));
  NOR2_X1   g283(.A1(new_n704), .A2(new_n705), .ZN(new_n709));
  NOR3_X1   g284(.A1(new_n703), .A2(new_n706), .A3(new_n709), .ZN(new_n710));
  AOI21_X1  g285(.A(new_n710), .B1(new_n703), .B2(new_n709), .ZN(new_n711));
  AND2_X1   g286(.A1(new_n708), .A2(new_n711), .ZN(new_n712));
  XNOR2_X1  g287(.A(new_n712), .B(G1986), .ZN(new_n713));
  XOR2_X1   g288(.A(KEYINPUT21), .B(KEYINPUT22), .Z(new_n714));
  INV_X1    g289(.A(new_n714), .ZN(new_n715));
  NAND2_X1  g290(.A1(new_n713), .A2(new_n715), .ZN(new_n716));
  INV_X1    g291(.A(G1986), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n712), .B(new_n717), .ZN(new_n718));
  NAND2_X1  g293(.A1(new_n718), .A2(new_n714), .ZN(new_n719));
  XNOR2_X1  g294(.A(G1991), .B(G1996), .ZN(new_n720));
  INV_X1    g295(.A(G1981), .ZN(new_n721));
  XNOR2_X1  g296(.A(new_n720), .B(new_n721), .ZN(new_n722));
  AND3_X1   g297(.A1(new_n716), .A2(new_n719), .A3(new_n722), .ZN(new_n723));
  AOI21_X1  g298(.A(new_n722), .B1(new_n716), .B2(new_n719), .ZN(new_n724));
  NOR2_X1   g299(.A1(new_n723), .A2(new_n724), .ZN(G229));
  INV_X1    g300(.A(G16), .ZN(new_n726));
  NAND2_X1  g301(.A1(new_n726), .A2(G4), .ZN(new_n727));
  OAI21_X1  g302(.A(new_n727), .B1(new_n616), .B2(new_n726), .ZN(new_n728));
  XNOR2_X1  g303(.A(new_n728), .B(KEYINPUT95), .ZN(new_n729));
  INV_X1    g304(.A(G1348), .ZN(new_n730));
  XNOR2_X1  g305(.A(new_n729), .B(new_n730), .ZN(new_n731));
  INV_X1    g306(.A(G29), .ZN(new_n732));
  NAND2_X1  g307(.A1(new_n732), .A2(G35), .ZN(new_n733));
  XOR2_X1   g308(.A(new_n733), .B(KEYINPUT101), .Z(new_n734));
  OAI21_X1  g309(.A(new_n734), .B1(G162), .B2(new_n732), .ZN(new_n735));
  XOR2_X1   g310(.A(KEYINPUT29), .B(G2090), .Z(new_n736));
  XNOR2_X1  g311(.A(new_n735), .B(new_n736), .ZN(new_n737));
  NAND2_X1  g312(.A1(new_n726), .A2(G19), .ZN(new_n738));
  OAI21_X1  g313(.A(new_n738), .B1(new_n559), .B2(new_n726), .ZN(new_n739));
  XOR2_X1   g314(.A(new_n739), .B(G1341), .Z(new_n740));
  NAND2_X1  g315(.A1(new_n726), .A2(G20), .ZN(new_n741));
  XOR2_X1   g316(.A(new_n741), .B(KEYINPUT23), .Z(new_n742));
  AOI21_X1  g317(.A(new_n742), .B1(G299), .B2(G16), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(G1956), .ZN(new_n744));
  INV_X1    g319(.A(G28), .ZN(new_n745));
  OR2_X1    g320(.A1(new_n745), .A2(KEYINPUT30), .ZN(new_n746));
  AOI21_X1  g321(.A(G29), .B1(new_n745), .B2(KEYINPUT30), .ZN(new_n747));
  OR2_X1    g322(.A1(KEYINPUT31), .A2(G11), .ZN(new_n748));
  NAND2_X1  g323(.A1(KEYINPUT31), .A2(G11), .ZN(new_n749));
  AOI22_X1  g324(.A1(new_n746), .A2(new_n747), .B1(new_n748), .B2(new_n749), .ZN(new_n750));
  OAI21_X1  g325(.A(new_n750), .B1(new_n636), .B2(new_n732), .ZN(new_n751));
  XOR2_X1   g326(.A(new_n751), .B(KEYINPUT98), .Z(new_n752));
  NAND4_X1  g327(.A1(new_n737), .A2(new_n740), .A3(new_n744), .A4(new_n752), .ZN(new_n753));
  NAND2_X1  g328(.A1(new_n486), .A2(G141), .ZN(new_n754));
  NAND2_X1  g329(.A1(new_n488), .A2(G129), .ZN(new_n755));
  NAND3_X1  g330(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n756));
  INV_X1    g331(.A(KEYINPUT26), .ZN(new_n757));
  OR2_X1    g332(.A1(new_n756), .A2(new_n757), .ZN(new_n758));
  NAND2_X1  g333(.A1(new_n756), .A2(new_n757), .ZN(new_n759));
  AOI22_X1  g334(.A1(new_n758), .A2(new_n759), .B1(G105), .B2(new_n472), .ZN(new_n760));
  NAND3_X1  g335(.A1(new_n754), .A2(new_n755), .A3(new_n760), .ZN(new_n761));
  INV_X1    g336(.A(new_n761), .ZN(new_n762));
  NOR2_X1   g337(.A1(new_n762), .A2(new_n732), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n732), .B2(G32), .ZN(new_n764));
  XNOR2_X1  g339(.A(KEYINPUT27), .B(G1996), .ZN(new_n765));
  AND2_X1   g340(.A1(new_n764), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g341(.A1(new_n764), .A2(new_n765), .ZN(new_n767));
  NAND2_X1  g342(.A1(new_n732), .A2(G33), .ZN(new_n768));
  NAND3_X1  g343(.A1(new_n459), .A2(G103), .A3(G2104), .ZN(new_n769));
  XOR2_X1   g344(.A(new_n769), .B(KEYINPUT25), .Z(new_n770));
  AOI22_X1  g345(.A1(new_n468), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n771));
  OAI21_X1  g346(.A(new_n770), .B1(new_n771), .B2(new_n459), .ZN(new_n772));
  AOI21_X1  g347(.A(new_n772), .B1(G139), .B2(new_n486), .ZN(new_n773));
  OAI21_X1  g348(.A(new_n768), .B1(new_n773), .B2(new_n732), .ZN(new_n774));
  XNOR2_X1  g349(.A(new_n774), .B(G2072), .ZN(new_n775));
  NOR3_X1   g350(.A1(new_n766), .A2(new_n767), .A3(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n732), .A2(G27), .ZN(new_n777));
  OAI21_X1  g352(.A(new_n777), .B1(G164), .B2(new_n732), .ZN(new_n778));
  XNOR2_X1  g353(.A(new_n778), .B(G2078), .ZN(new_n779));
  XNOR2_X1  g354(.A(new_n779), .B(KEYINPUT100), .ZN(new_n780));
  NAND2_X1  g355(.A1(new_n726), .A2(G21), .ZN(new_n781));
  OAI21_X1  g356(.A(new_n781), .B1(G168), .B2(new_n726), .ZN(new_n782));
  XNOR2_X1  g357(.A(new_n782), .B(G1966), .ZN(new_n783));
  NOR2_X1   g358(.A1(new_n780), .A2(new_n783), .ZN(new_n784));
  NAND2_X1  g359(.A1(new_n726), .A2(G5), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n785), .B1(G171), .B2(new_n726), .ZN(new_n786));
  XOR2_X1   g361(.A(KEYINPUT99), .B(G1961), .Z(new_n787));
  XNOR2_X1  g362(.A(new_n786), .B(new_n787), .ZN(new_n788));
  NAND2_X1  g363(.A1(new_n732), .A2(G26), .ZN(new_n789));
  XOR2_X1   g364(.A(new_n789), .B(KEYINPUT28), .Z(new_n790));
  OAI21_X1  g365(.A(G2104), .B1(new_n459), .B2(G116), .ZN(new_n791));
  INV_X1    g366(.A(G104), .ZN(new_n792));
  AOI21_X1  g367(.A(new_n791), .B1(new_n792), .B2(new_n459), .ZN(new_n793));
  OR2_X1    g368(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n794));
  NAND2_X1  g369(.A1(new_n793), .A2(KEYINPUT97), .ZN(new_n795));
  AOI22_X1  g370(.A1(new_n794), .A2(new_n795), .B1(new_n486), .B2(G140), .ZN(new_n796));
  NAND3_X1  g371(.A1(new_n488), .A2(KEYINPUT96), .A3(G128), .ZN(new_n797));
  INV_X1    g372(.A(new_n797), .ZN(new_n798));
  AOI21_X1  g373(.A(KEYINPUT96), .B1(new_n488), .B2(G128), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n796), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  AOI21_X1  g375(.A(new_n790), .B1(new_n800), .B2(G29), .ZN(new_n801));
  XNOR2_X1  g376(.A(new_n801), .B(G2067), .ZN(new_n802));
  NAND4_X1  g377(.A1(new_n776), .A2(new_n784), .A3(new_n788), .A4(new_n802), .ZN(new_n803));
  INV_X1    g378(.A(G34), .ZN(new_n804));
  AND2_X1   g379(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n805));
  NOR2_X1   g380(.A1(new_n804), .A2(KEYINPUT24), .ZN(new_n806));
  OAI21_X1  g381(.A(new_n732), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  OAI21_X1  g382(.A(new_n807), .B1(G160), .B2(new_n732), .ZN(new_n808));
  XNOR2_X1  g383(.A(new_n808), .B(G2084), .ZN(new_n809));
  NOR3_X1   g384(.A1(new_n753), .A2(new_n803), .A3(new_n809), .ZN(new_n810));
  MUX2_X1   g385(.A(G6), .B(G305), .S(G16), .Z(new_n811));
  XNOR2_X1  g386(.A(KEYINPUT32), .B(G1981), .ZN(new_n812));
  XNOR2_X1  g387(.A(new_n811), .B(new_n812), .ZN(new_n813));
  INV_X1    g388(.A(KEYINPUT93), .ZN(new_n814));
  NAND2_X1  g389(.A1(new_n813), .A2(new_n814), .ZN(new_n815));
  OR2_X1    g390(.A1(new_n811), .A2(new_n812), .ZN(new_n816));
  NAND2_X1  g391(.A1(new_n811), .A2(new_n812), .ZN(new_n817));
  NAND3_X1  g392(.A1(new_n816), .A2(KEYINPUT93), .A3(new_n817), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n726), .A2(G23), .ZN(new_n819));
  INV_X1    g394(.A(G288), .ZN(new_n820));
  OAI21_X1  g395(.A(new_n819), .B1(new_n820), .B2(new_n726), .ZN(new_n821));
  XOR2_X1   g396(.A(KEYINPUT33), .B(G1976), .Z(new_n822));
  NAND2_X1  g397(.A1(new_n821), .A2(new_n822), .ZN(new_n823));
  NAND2_X1  g398(.A1(new_n726), .A2(G22), .ZN(new_n824));
  OAI21_X1  g399(.A(new_n824), .B1(G166), .B2(new_n726), .ZN(new_n825));
  XNOR2_X1  g400(.A(new_n825), .B(G1971), .ZN(new_n826));
  NOR2_X1   g401(.A1(new_n821), .A2(new_n822), .ZN(new_n827));
  NOR2_X1   g402(.A1(new_n826), .A2(new_n827), .ZN(new_n828));
  NAND4_X1  g403(.A1(new_n815), .A2(new_n818), .A3(new_n823), .A4(new_n828), .ZN(new_n829));
  OR2_X1    g404(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n830));
  NAND2_X1  g405(.A1(new_n829), .A2(KEYINPUT34), .ZN(new_n831));
  NAND2_X1  g406(.A1(new_n732), .A2(G25), .ZN(new_n832));
  OAI21_X1  g407(.A(G2104), .B1(new_n459), .B2(G107), .ZN(new_n833));
  INV_X1    g408(.A(G95), .ZN(new_n834));
  AOI21_X1  g409(.A(new_n833), .B1(new_n834), .B2(new_n459), .ZN(new_n835));
  AOI21_X1  g410(.A(new_n835), .B1(new_n488), .B2(G119), .ZN(new_n836));
  NAND2_X1  g411(.A1(new_n486), .A2(G131), .ZN(new_n837));
  NAND2_X1  g412(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  INV_X1    g413(.A(new_n838), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n832), .B1(new_n839), .B2(new_n732), .ZN(new_n840));
  XOR2_X1   g415(.A(KEYINPUT35), .B(G1991), .Z(new_n841));
  XNOR2_X1  g416(.A(new_n840), .B(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n843));
  NAND2_X1  g418(.A1(new_n598), .A2(KEYINPUT92), .ZN(new_n844));
  NAND3_X1  g419(.A1(new_n843), .A2(G16), .A3(new_n844), .ZN(new_n845));
  INV_X1    g420(.A(G24), .ZN(new_n846));
  OAI21_X1  g421(.A(new_n845), .B1(G16), .B2(new_n846), .ZN(new_n847));
  OAI21_X1  g422(.A(new_n842), .B1(new_n847), .B2(G1986), .ZN(new_n848));
  AOI21_X1  g423(.A(new_n848), .B1(G1986), .B2(new_n847), .ZN(new_n849));
  NAND3_X1  g424(.A1(new_n830), .A2(new_n831), .A3(new_n849), .ZN(new_n850));
  NAND2_X1  g425(.A1(KEYINPUT94), .A2(KEYINPUT36), .ZN(new_n851));
  OAI211_X1 g426(.A(new_n731), .B(new_n810), .C1(new_n850), .C2(new_n851), .ZN(new_n852));
  XOR2_X1   g427(.A(KEYINPUT94), .B(KEYINPUT36), .Z(new_n853));
  AND2_X1   g428(.A1(new_n850), .A2(new_n853), .ZN(new_n854));
  NOR2_X1   g429(.A1(new_n852), .A2(new_n854), .ZN(G311));
  OR2_X1    g430(.A1(new_n852), .A2(new_n854), .ZN(G150));
  NAND3_X1  g431(.A1(new_n539), .A2(G67), .A3(new_n540), .ZN(new_n857));
  INV_X1    g432(.A(KEYINPUT102), .ZN(new_n858));
  AND2_X1   g433(.A1(G80), .A2(G543), .ZN(new_n859));
  INV_X1    g434(.A(new_n859), .ZN(new_n860));
  NAND3_X1  g435(.A1(new_n857), .A2(new_n858), .A3(new_n860), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  AOI21_X1  g437(.A(new_n858), .B1(new_n857), .B2(new_n860), .ZN(new_n863));
  NOR3_X1   g438(.A1(new_n862), .A2(new_n863), .A3(new_n516), .ZN(new_n864));
  AOI22_X1  g439(.A1(new_n524), .A2(G93), .B1(G55), .B2(new_n530), .ZN(new_n865));
  INV_X1    g440(.A(new_n865), .ZN(new_n866));
  OAI21_X1  g441(.A(new_n628), .B1(new_n864), .B2(new_n866), .ZN(new_n867));
  NAND2_X1  g442(.A1(new_n857), .A2(new_n860), .ZN(new_n868));
  NAND2_X1  g443(.A1(new_n868), .A2(KEYINPUT102), .ZN(new_n869));
  NAND3_X1  g444(.A1(new_n869), .A2(G651), .A3(new_n861), .ZN(new_n870));
  NAND3_X1  g445(.A1(new_n870), .A2(new_n559), .A3(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  NAND2_X1  g447(.A1(new_n616), .A2(G559), .ZN(new_n873));
  XNOR2_X1  g448(.A(new_n872), .B(new_n873), .ZN(new_n874));
  XNOR2_X1  g449(.A(KEYINPUT103), .B(KEYINPUT38), .ZN(new_n875));
  XNOR2_X1  g450(.A(new_n874), .B(new_n875), .ZN(new_n876));
  INV_X1    g451(.A(KEYINPUT39), .ZN(new_n877));
  AOI21_X1  g452(.A(G860), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  OAI21_X1  g453(.A(new_n878), .B1(new_n877), .B2(new_n876), .ZN(new_n879));
  OAI21_X1  g454(.A(G860), .B1(new_n864), .B2(new_n866), .ZN(new_n880));
  XOR2_X1   g455(.A(new_n880), .B(KEYINPUT37), .Z(new_n881));
  NAND2_X1  g456(.A1(new_n879), .A2(new_n881), .ZN(G145));
  XNOR2_X1  g457(.A(KEYINPUT106), .B(G37), .ZN(new_n883));
  INV_X1    g458(.A(new_n883), .ZN(new_n884));
  NAND2_X1  g459(.A1(new_n486), .A2(G142), .ZN(new_n885));
  NAND2_X1  g460(.A1(new_n488), .A2(G130), .ZN(new_n886));
  NOR3_X1   g461(.A1(new_n459), .A2(KEYINPUT104), .A3(G118), .ZN(new_n887));
  OAI21_X1  g462(.A(KEYINPUT104), .B1(new_n459), .B2(G118), .ZN(new_n888));
  OR2_X1    g463(.A1(G106), .A2(G2105), .ZN(new_n889));
  NAND3_X1  g464(.A1(new_n888), .A2(G2104), .A3(new_n889), .ZN(new_n890));
  OAI211_X1 g465(.A(new_n885), .B(new_n886), .C1(new_n887), .C2(new_n890), .ZN(new_n891));
  XNOR2_X1  g466(.A(new_n891), .B(new_n838), .ZN(new_n892));
  AND2_X1   g467(.A1(new_n892), .A2(new_n641), .ZN(new_n893));
  NOR2_X1   g468(.A1(new_n892), .A2(new_n641), .ZN(new_n894));
  NOR2_X1   g469(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  INV_X1    g470(.A(new_n773), .ZN(new_n896));
  NAND2_X1  g471(.A1(new_n800), .A2(G164), .ZN(new_n897));
  INV_X1    g472(.A(KEYINPUT96), .ZN(new_n898));
  NAND2_X1  g473(.A1(new_n483), .A2(new_n485), .ZN(new_n899));
  NAND2_X1  g474(.A1(new_n899), .A2(G2105), .ZN(new_n900));
  INV_X1    g475(.A(G128), .ZN(new_n901));
  OAI21_X1  g476(.A(new_n898), .B1(new_n900), .B2(new_n901), .ZN(new_n902));
  NAND2_X1  g477(.A1(new_n902), .A2(new_n797), .ZN(new_n903));
  NAND3_X1  g478(.A1(new_n903), .A2(new_n508), .A3(new_n796), .ZN(new_n904));
  AND3_X1   g479(.A1(new_n897), .A2(new_n761), .A3(new_n904), .ZN(new_n905));
  AOI21_X1  g480(.A(new_n761), .B1(new_n897), .B2(new_n904), .ZN(new_n906));
  OAI21_X1  g481(.A(new_n896), .B1(new_n905), .B2(new_n906), .ZN(new_n907));
  NAND2_X1  g482(.A1(new_n897), .A2(new_n904), .ZN(new_n908));
  NAND2_X1  g483(.A1(new_n908), .A2(new_n762), .ZN(new_n909));
  NAND3_X1  g484(.A1(new_n897), .A2(new_n761), .A3(new_n904), .ZN(new_n910));
  NAND3_X1  g485(.A1(new_n909), .A2(new_n773), .A3(new_n910), .ZN(new_n911));
  NAND3_X1  g486(.A1(new_n895), .A2(new_n907), .A3(new_n911), .ZN(new_n912));
  NAND2_X1  g487(.A1(new_n907), .A2(new_n911), .ZN(new_n913));
  INV_X1    g488(.A(new_n895), .ZN(new_n914));
  INV_X1    g489(.A(KEYINPUT105), .ZN(new_n915));
  NAND3_X1  g490(.A1(new_n913), .A2(new_n914), .A3(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(new_n916), .ZN(new_n917));
  AOI21_X1  g492(.A(new_n915), .B1(new_n913), .B2(new_n914), .ZN(new_n918));
  OAI21_X1  g493(.A(new_n912), .B1(new_n917), .B2(new_n918), .ZN(new_n919));
  XNOR2_X1  g494(.A(G160), .B(new_n636), .ZN(new_n920));
  AND2_X1   g495(.A1(new_n920), .A2(G162), .ZN(new_n921));
  NOR2_X1   g496(.A1(new_n920), .A2(G162), .ZN(new_n922));
  NOR2_X1   g497(.A1(new_n921), .A2(new_n922), .ZN(new_n923));
  INV_X1    g498(.A(new_n923), .ZN(new_n924));
  AOI21_X1  g499(.A(new_n884), .B1(new_n919), .B2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n913), .A2(new_n914), .ZN(new_n926));
  NAND3_X1  g501(.A1(new_n926), .A2(new_n923), .A3(new_n912), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(KEYINPUT107), .ZN(new_n928));
  INV_X1    g503(.A(KEYINPUT107), .ZN(new_n929));
  NAND4_X1  g504(.A1(new_n926), .A2(new_n923), .A3(new_n929), .A4(new_n912), .ZN(new_n930));
  NAND2_X1  g505(.A1(new_n928), .A2(new_n930), .ZN(new_n931));
  AND3_X1   g506(.A1(new_n925), .A2(KEYINPUT40), .A3(new_n931), .ZN(new_n932));
  AOI21_X1  g507(.A(KEYINPUT40), .B1(new_n925), .B2(new_n931), .ZN(new_n933));
  NOR2_X1   g508(.A1(new_n932), .A2(new_n933), .ZN(G395));
  XNOR2_X1  g509(.A(new_n598), .B(G305), .ZN(new_n935));
  XNOR2_X1  g510(.A(G166), .B(G288), .ZN(new_n936));
  XNOR2_X1  g511(.A(new_n935), .B(new_n936), .ZN(new_n937));
  INV_X1    g512(.A(new_n937), .ZN(new_n938));
  NAND2_X1  g513(.A1(new_n938), .A2(KEYINPUT42), .ZN(new_n939));
  INV_X1    g514(.A(KEYINPUT42), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n937), .A2(new_n940), .ZN(new_n941));
  NAND2_X1  g516(.A1(new_n939), .A2(new_n941), .ZN(new_n942));
  XOR2_X1   g517(.A(new_n872), .B(new_n625), .Z(new_n943));
  NAND2_X1  g518(.A1(new_n616), .A2(G299), .ZN(new_n944));
  AND3_X1   g519(.A1(new_n609), .A2(new_n614), .A3(new_n611), .ZN(new_n945));
  AOI21_X1  g520(.A(new_n614), .B1(new_n609), .B2(new_n611), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n606), .B1(new_n945), .B2(new_n946), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(new_n620), .ZN(new_n948));
  NAND2_X1  g523(.A1(new_n944), .A2(new_n948), .ZN(new_n949));
  OR2_X1    g524(.A1(new_n943), .A2(new_n949), .ZN(new_n950));
  OAI21_X1  g525(.A(KEYINPUT108), .B1(new_n616), .B2(G299), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT108), .ZN(new_n952));
  NAND3_X1  g527(.A1(new_n947), .A2(new_n952), .A3(new_n620), .ZN(new_n953));
  NAND3_X1  g528(.A1(new_n951), .A2(new_n944), .A3(new_n953), .ZN(new_n954));
  INV_X1    g529(.A(KEYINPUT41), .ZN(new_n955));
  AOI21_X1  g530(.A(new_n955), .B1(new_n616), .B2(G299), .ZN(new_n956));
  AOI22_X1  g531(.A1(new_n954), .A2(new_n955), .B1(new_n948), .B2(new_n956), .ZN(new_n957));
  NAND2_X1  g532(.A1(new_n957), .A2(new_n943), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n950), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n942), .A2(new_n959), .ZN(new_n960));
  NAND4_X1  g535(.A1(new_n939), .A2(new_n950), .A3(new_n941), .A4(new_n958), .ZN(new_n961));
  NAND3_X1  g536(.A1(new_n960), .A2(G868), .A3(new_n961), .ZN(new_n962));
  INV_X1    g537(.A(KEYINPUT109), .ZN(new_n963));
  NAND2_X1  g538(.A1(new_n962), .A2(new_n963), .ZN(new_n964));
  NAND4_X1  g539(.A1(new_n960), .A2(KEYINPUT109), .A3(G868), .A4(new_n961), .ZN(new_n965));
  OAI21_X1  g540(.A(new_n627), .B1(new_n864), .B2(new_n866), .ZN(new_n966));
  NAND3_X1  g541(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G295));
  NAND3_X1  g542(.A1(new_n964), .A2(new_n965), .A3(new_n966), .ZN(G331));
  NOR2_X1   g543(.A1(G171), .A2(KEYINPUT110), .ZN(new_n969));
  INV_X1    g544(.A(new_n969), .ZN(new_n970));
  AND3_X1   g545(.A1(new_n870), .A2(new_n559), .A3(new_n865), .ZN(new_n971));
  AOI21_X1  g546(.A(new_n559), .B1(new_n870), .B2(new_n865), .ZN(new_n972));
  AOI21_X1  g547(.A(G286), .B1(G171), .B2(KEYINPUT110), .ZN(new_n973));
  NOR3_X1   g548(.A1(new_n971), .A2(new_n972), .A3(new_n973), .ZN(new_n974));
  INV_X1    g549(.A(KEYINPUT110), .ZN(new_n975));
  OAI21_X1  g550(.A(G168), .B1(G301), .B2(new_n975), .ZN(new_n976));
  AOI21_X1  g551(.A(new_n976), .B1(new_n867), .B2(new_n871), .ZN(new_n977));
  OAI21_X1  g552(.A(new_n970), .B1(new_n974), .B2(new_n977), .ZN(new_n978));
  OAI21_X1  g553(.A(new_n973), .B1(new_n971), .B2(new_n972), .ZN(new_n979));
  NAND3_X1  g554(.A1(new_n867), .A2(new_n976), .A3(new_n871), .ZN(new_n980));
  NAND3_X1  g555(.A1(new_n979), .A2(new_n980), .A3(new_n969), .ZN(new_n981));
  NAND3_X1  g556(.A1(new_n978), .A2(new_n949), .A3(new_n981), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n978), .A2(new_n981), .ZN(new_n983));
  NAND3_X1  g558(.A1(new_n951), .A2(new_n956), .A3(new_n953), .ZN(new_n984));
  NAND2_X1  g559(.A1(new_n949), .A2(new_n955), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n984), .A2(new_n985), .ZN(new_n986));
  AOI22_X1  g561(.A1(new_n982), .A2(KEYINPUT111), .B1(new_n983), .B2(new_n986), .ZN(new_n987));
  OR2_X1    g562(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n988));
  AOI21_X1  g563(.A(new_n937), .B1(new_n987), .B2(new_n988), .ZN(new_n989));
  INV_X1    g564(.A(KEYINPUT43), .ZN(new_n990));
  AND3_X1   g565(.A1(new_n979), .A2(new_n980), .A3(new_n969), .ZN(new_n991));
  AOI21_X1  g566(.A(new_n969), .B1(new_n979), .B2(new_n980), .ZN(new_n992));
  NOR2_X1   g567(.A1(new_n991), .A2(new_n992), .ZN(new_n993));
  OAI211_X1 g568(.A(new_n982), .B(new_n937), .C1(new_n993), .C2(new_n957), .ZN(new_n994));
  NAND2_X1  g569(.A1(new_n994), .A2(new_n883), .ZN(new_n995));
  NOR3_X1   g570(.A1(new_n989), .A2(new_n990), .A3(new_n995), .ZN(new_n996));
  INV_X1    g571(.A(G37), .ZN(new_n997));
  AND2_X1   g572(.A1(new_n994), .A2(new_n997), .ZN(new_n998));
  OAI21_X1  g573(.A(new_n982), .B1(new_n993), .B2(new_n957), .ZN(new_n999));
  NAND2_X1  g574(.A1(new_n999), .A2(new_n938), .ZN(new_n1000));
  AOI21_X1  g575(.A(KEYINPUT43), .B1(new_n998), .B2(new_n1000), .ZN(new_n1001));
  OAI21_X1  g576(.A(KEYINPUT44), .B1(new_n996), .B2(new_n1001), .ZN(new_n1002));
  INV_X1    g577(.A(KEYINPUT44), .ZN(new_n1003));
  NOR3_X1   g578(.A1(new_n989), .A2(KEYINPUT43), .A3(new_n995), .ZN(new_n1004));
  AOI21_X1  g579(.A(new_n990), .B1(new_n998), .B2(new_n1000), .ZN(new_n1005));
  OAI21_X1  g580(.A(new_n1003), .B1(new_n1004), .B2(new_n1005), .ZN(new_n1006));
  NAND2_X1  g581(.A1(new_n1002), .A2(new_n1006), .ZN(G397));
  INV_X1    g582(.A(G40), .ZN(new_n1008));
  NOR3_X1   g583(.A1(new_n470), .A2(new_n1008), .A3(new_n478), .ZN(new_n1009));
  INV_X1    g584(.A(G1384), .ZN(new_n1010));
  AOI21_X1  g585(.A(KEYINPUT45), .B1(new_n508), .B2(new_n1010), .ZN(new_n1011));
  NAND2_X1  g586(.A1(new_n1009), .A2(new_n1011), .ZN(new_n1012));
  XOR2_X1   g587(.A(new_n1012), .B(KEYINPUT112), .Z(new_n1013));
  NAND2_X1  g588(.A1(new_n800), .A2(G2067), .ZN(new_n1014));
  INV_X1    g589(.A(G2067), .ZN(new_n1015));
  NAND3_X1  g590(.A1(new_n903), .A2(new_n1015), .A3(new_n796), .ZN(new_n1016));
  NAND2_X1  g591(.A1(new_n1014), .A2(new_n1016), .ZN(new_n1017));
  INV_X1    g592(.A(new_n1017), .ZN(new_n1018));
  INV_X1    g593(.A(G1996), .ZN(new_n1019));
  XNOR2_X1  g594(.A(new_n761), .B(new_n1019), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n839), .A2(new_n841), .ZN(new_n1021));
  OR2_X1    g596(.A1(new_n839), .A2(new_n841), .ZN(new_n1022));
  NAND4_X1  g597(.A1(new_n1018), .A2(new_n1020), .A3(new_n1021), .A4(new_n1022), .ZN(new_n1023));
  XNOR2_X1  g598(.A(new_n598), .B(new_n717), .ZN(new_n1024));
  OAI21_X1  g599(.A(new_n1013), .B1(new_n1023), .B2(new_n1024), .ZN(new_n1025));
  INV_X1    g600(.A(KEYINPUT127), .ZN(new_n1026));
  NAND2_X1  g601(.A1(new_n499), .A2(new_n505), .ZN(new_n1027));
  AOI21_X1  g602(.A(G2105), .B1(new_n466), .B2(new_n467), .ZN(new_n1028));
  INV_X1    g603(.A(new_n506), .ZN(new_n1029));
  AOI21_X1  g604(.A(new_n498), .B1(new_n1028), .B2(new_n1029), .ZN(new_n1030));
  OAI21_X1  g605(.A(new_n1010), .B1(new_n1027), .B2(new_n1030), .ZN(new_n1031));
  NAND2_X1  g606(.A1(new_n1031), .A2(KEYINPUT50), .ZN(new_n1032));
  INV_X1    g607(.A(KEYINPUT50), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n508), .A2(new_n1033), .A3(new_n1010), .ZN(new_n1034));
  AND3_X1   g609(.A1(new_n1009), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1035));
  INV_X1    g610(.A(G2090), .ZN(new_n1036));
  INV_X1    g611(.A(KEYINPUT45), .ZN(new_n1037));
  NAND2_X1  g612(.A1(new_n1031), .A2(new_n1037), .ZN(new_n1038));
  OAI211_X1 g613(.A(KEYINPUT45), .B(new_n1010), .C1(new_n1027), .C2(new_n1030), .ZN(new_n1039));
  NAND3_X1  g614(.A1(new_n1009), .A2(new_n1038), .A3(new_n1039), .ZN(new_n1040));
  INV_X1    g615(.A(G1971), .ZN(new_n1041));
  AOI22_X1  g616(.A1(new_n1035), .A2(new_n1036), .B1(new_n1040), .B2(new_n1041), .ZN(new_n1042));
  INV_X1    g617(.A(G8), .ZN(new_n1043));
  NOR2_X1   g618(.A1(new_n1042), .A2(new_n1043), .ZN(new_n1044));
  NAND2_X1  g619(.A1(G303), .A2(G8), .ZN(new_n1045));
  XOR2_X1   g620(.A(new_n1045), .B(KEYINPUT55), .Z(new_n1046));
  NAND2_X1  g621(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1047));
  INV_X1    g622(.A(G2078), .ZN(new_n1048));
  NAND4_X1  g623(.A1(new_n1009), .A2(new_n1038), .A3(new_n1048), .A4(new_n1039), .ZN(new_n1049));
  INV_X1    g624(.A(KEYINPUT53), .ZN(new_n1050));
  NAND3_X1  g625(.A1(new_n1009), .A2(new_n1032), .A3(new_n1034), .ZN(new_n1051));
  XNOR2_X1  g626(.A(KEYINPUT125), .B(G1961), .ZN(new_n1052));
  AOI22_X1  g627(.A1(new_n1049), .A2(new_n1050), .B1(new_n1051), .B2(new_n1052), .ZN(new_n1053));
  OR2_X1    g628(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1054));
  AOI21_X1  g629(.A(G301), .B1(new_n1053), .B2(new_n1054), .ZN(new_n1055));
  AND2_X1   g630(.A1(new_n1047), .A2(new_n1055), .ZN(new_n1056));
  XOR2_X1   g631(.A(KEYINPUT122), .B(KEYINPUT51), .Z(new_n1057));
  INV_X1    g632(.A(G1966), .ZN(new_n1058));
  NAND2_X1  g633(.A1(new_n1040), .A2(new_n1058), .ZN(new_n1059));
  INV_X1    g634(.A(G2084), .ZN(new_n1060));
  NAND4_X1  g635(.A1(new_n1009), .A2(new_n1032), .A3(new_n1060), .A4(new_n1034), .ZN(new_n1061));
  AOI21_X1  g636(.A(new_n1043), .B1(new_n1059), .B2(new_n1061), .ZN(new_n1062));
  NAND2_X1  g637(.A1(G286), .A2(G8), .ZN(new_n1063));
  NAND2_X1  g638(.A1(new_n1063), .A2(KEYINPUT121), .ZN(new_n1064));
  INV_X1    g639(.A(KEYINPUT121), .ZN(new_n1065));
  NAND3_X1  g640(.A1(G286), .A2(new_n1065), .A3(G8), .ZN(new_n1066));
  NAND2_X1  g641(.A1(new_n1064), .A2(new_n1066), .ZN(new_n1067));
  OAI21_X1  g642(.A(new_n1057), .B1(new_n1062), .B2(new_n1067), .ZN(new_n1068));
  INV_X1    g643(.A(KEYINPUT51), .ZN(new_n1069));
  NAND3_X1  g644(.A1(new_n1064), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1070));
  OAI21_X1  g645(.A(KEYINPUT123), .B1(new_n1062), .B2(new_n1070), .ZN(new_n1071));
  INV_X1    g646(.A(KEYINPUT123), .ZN(new_n1072));
  AND3_X1   g647(.A1(new_n1064), .A2(new_n1069), .A3(new_n1066), .ZN(new_n1073));
  AOI22_X1  g648(.A1(new_n1035), .A2(new_n1060), .B1(new_n1040), .B2(new_n1058), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1072), .B(new_n1073), .C1(new_n1074), .C2(new_n1043), .ZN(new_n1075));
  NAND3_X1  g650(.A1(new_n1068), .A2(new_n1071), .A3(new_n1075), .ZN(new_n1076));
  INV_X1    g651(.A(new_n1074), .ZN(new_n1077));
  NAND2_X1  g652(.A1(new_n1077), .A2(new_n1067), .ZN(new_n1078));
  AND3_X1   g653(.A1(new_n1076), .A2(KEYINPUT62), .A3(new_n1078), .ZN(new_n1079));
  AOI21_X1  g654(.A(KEYINPUT62), .B1(new_n1076), .B2(new_n1078), .ZN(new_n1080));
  OAI21_X1  g655(.A(new_n1056), .B1(new_n1079), .B2(new_n1080), .ZN(new_n1081));
  NOR4_X1   g656(.A1(new_n1031), .A2(new_n470), .A3(new_n1008), .A4(new_n478), .ZN(new_n1082));
  NOR2_X1   g657(.A1(new_n1082), .A2(new_n1043), .ZN(new_n1083));
  NAND3_X1  g658(.A1(new_n587), .A2(new_n591), .A3(new_n721), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT114), .ZN(new_n1085));
  AND3_X1   g660(.A1(new_n588), .A2(new_n1085), .A3(new_n589), .ZN(new_n1086));
  AOI21_X1  g661(.A(new_n1085), .B1(new_n588), .B2(new_n589), .ZN(new_n1087));
  AND2_X1   g662(.A1(new_n584), .A2(G651), .ZN(new_n1088));
  NOR3_X1   g663(.A1(new_n1086), .A2(new_n1087), .A3(new_n1088), .ZN(new_n1089));
  OAI21_X1  g664(.A(new_n1084), .B1(new_n1089), .B2(new_n721), .ZN(new_n1090));
  INV_X1    g665(.A(KEYINPUT49), .ZN(new_n1091));
  OAI21_X1  g666(.A(new_n1083), .B1(new_n1090), .B2(new_n1091), .ZN(new_n1092));
  AOI21_X1  g667(.A(new_n1088), .B1(new_n590), .B2(KEYINPUT114), .ZN(new_n1093));
  NAND3_X1  g668(.A1(new_n588), .A2(new_n1085), .A3(new_n589), .ZN(new_n1094));
  AOI21_X1  g669(.A(new_n721), .B1(new_n1093), .B2(new_n1094), .ZN(new_n1095));
  NOR4_X1   g670(.A1(new_n590), .A2(new_n585), .A3(new_n586), .A4(G1981), .ZN(new_n1096));
  OAI21_X1  g671(.A(KEYINPUT115), .B1(new_n1095), .B2(new_n1096), .ZN(new_n1097));
  INV_X1    g672(.A(KEYINPUT115), .ZN(new_n1098));
  OAI211_X1 g673(.A(new_n1098), .B(new_n1084), .C1(new_n1089), .C2(new_n721), .ZN(new_n1099));
  NAND3_X1  g674(.A1(new_n1097), .A2(new_n1099), .A3(new_n1091), .ZN(new_n1100));
  INV_X1    g675(.A(KEYINPUT116), .ZN(new_n1101));
  NAND2_X1  g676(.A1(new_n1100), .A2(new_n1101), .ZN(new_n1102));
  NAND4_X1  g677(.A1(new_n1097), .A2(new_n1099), .A3(KEYINPUT116), .A4(new_n1091), .ZN(new_n1103));
  AOI21_X1  g678(.A(new_n1092), .B1(new_n1102), .B2(new_n1103), .ZN(new_n1104));
  INV_X1    g679(.A(G1976), .ZN(new_n1105));
  OAI21_X1  g680(.A(new_n1083), .B1(new_n1105), .B2(G288), .ZN(new_n1106));
  NAND2_X1  g681(.A1(new_n1106), .A2(KEYINPUT52), .ZN(new_n1107));
  XOR2_X1   g682(.A(KEYINPUT113), .B(G1976), .Z(new_n1108));
  AOI21_X1  g683(.A(KEYINPUT52), .B1(G288), .B2(new_n1108), .ZN(new_n1109));
  OAI211_X1 g684(.A(new_n1109), .B(new_n1083), .C1(new_n1105), .C2(G288), .ZN(new_n1110));
  NAND2_X1  g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  NOR2_X1   g686(.A1(new_n1044), .A2(new_n1046), .ZN(new_n1112));
  NOR3_X1   g687(.A1(new_n1104), .A2(new_n1111), .A3(new_n1112), .ZN(new_n1113));
  INV_X1    g688(.A(new_n1113), .ZN(new_n1114));
  OAI21_X1  g689(.A(new_n1026), .B1(new_n1081), .B2(new_n1114), .ZN(new_n1115));
  NAND2_X1  g690(.A1(new_n1076), .A2(new_n1078), .ZN(new_n1116));
  INV_X1    g691(.A(KEYINPUT62), .ZN(new_n1117));
  NAND2_X1  g692(.A1(new_n1116), .A2(new_n1117), .ZN(new_n1118));
  NAND3_X1  g693(.A1(new_n1076), .A2(KEYINPUT62), .A3(new_n1078), .ZN(new_n1119));
  NAND2_X1  g694(.A1(new_n1118), .A2(new_n1119), .ZN(new_n1120));
  NAND4_X1  g695(.A1(new_n1120), .A2(KEYINPUT127), .A3(new_n1113), .A4(new_n1056), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1115), .A2(new_n1121), .ZN(new_n1122));
  INV_X1    g697(.A(new_n1111), .ZN(new_n1123));
  NAND2_X1  g698(.A1(new_n1062), .A2(G168), .ZN(new_n1124));
  NOR2_X1   g699(.A1(new_n1112), .A2(new_n1124), .ZN(new_n1125));
  AND2_X1   g700(.A1(new_n1102), .A2(new_n1103), .ZN(new_n1126));
  OAI211_X1 g701(.A(new_n1123), .B(new_n1125), .C1(new_n1126), .C2(new_n1092), .ZN(new_n1127));
  NAND2_X1  g702(.A1(new_n820), .A2(new_n1105), .ZN(new_n1128));
  OAI21_X1  g703(.A(new_n1084), .B1(new_n1104), .B2(new_n1128), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1127), .A2(KEYINPUT63), .B1(new_n1129), .B2(new_n1083), .ZN(new_n1130));
  OAI21_X1  g705(.A(new_n1047), .B1(KEYINPUT63), .B2(new_n1124), .ZN(new_n1131));
  XNOR2_X1  g706(.A(KEYINPUT124), .B(KEYINPUT54), .ZN(new_n1132));
  NAND2_X1  g707(.A1(new_n1049), .A2(new_n1050), .ZN(new_n1133));
  NAND2_X1  g708(.A1(new_n1051), .A2(new_n1052), .ZN(new_n1134));
  OR2_X1    g709(.A1(KEYINPUT126), .A2(G2078), .ZN(new_n1135));
  NAND2_X1  g710(.A1(KEYINPUT126), .A2(G2078), .ZN(new_n1136));
  AOI21_X1  g711(.A(new_n1050), .B1(new_n1135), .B2(new_n1136), .ZN(new_n1137));
  NAND4_X1  g712(.A1(new_n1009), .A2(new_n1038), .A3(new_n1039), .A4(new_n1137), .ZN(new_n1138));
  AND4_X1   g713(.A1(G301), .A2(new_n1133), .A3(new_n1134), .A4(new_n1138), .ZN(new_n1139));
  OAI21_X1  g714(.A(new_n1132), .B1(new_n1055), .B2(new_n1139), .ZN(new_n1140));
  NAND3_X1  g715(.A1(new_n1133), .A2(new_n1134), .A3(new_n1138), .ZN(new_n1141));
  NAND2_X1  g716(.A1(new_n1141), .A2(G171), .ZN(new_n1142));
  NAND3_X1  g717(.A1(new_n1053), .A2(new_n1054), .A3(G301), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1142), .A2(new_n1143), .A3(KEYINPUT54), .ZN(new_n1144));
  NAND2_X1  g719(.A1(new_n1140), .A2(new_n1144), .ZN(new_n1145));
  AOI21_X1  g720(.A(new_n1145), .B1(new_n1078), .B2(new_n1076), .ZN(new_n1146));
  INV_X1    g721(.A(new_n1039), .ZN(new_n1147));
  NOR2_X1   g722(.A1(new_n1147), .A2(new_n1011), .ZN(new_n1148));
  XNOR2_X1  g723(.A(KEYINPUT117), .B(KEYINPUT56), .ZN(new_n1149));
  XNOR2_X1  g724(.A(new_n1149), .B(G2072), .ZN(new_n1150));
  NAND4_X1  g725(.A1(new_n1148), .A2(KEYINPUT118), .A3(new_n1009), .A4(new_n1150), .ZN(new_n1151));
  NAND4_X1  g726(.A1(new_n1009), .A2(new_n1038), .A3(new_n1039), .A4(new_n1150), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT118), .ZN(new_n1153));
  NAND2_X1  g728(.A1(new_n1152), .A2(new_n1153), .ZN(new_n1154));
  INV_X1    g729(.A(KEYINPUT57), .ZN(new_n1155));
  XNOR2_X1  g730(.A(G299), .B(new_n1155), .ZN(new_n1156));
  INV_X1    g731(.A(G1956), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1051), .A2(new_n1157), .ZN(new_n1158));
  NAND4_X1  g733(.A1(new_n1151), .A2(new_n1154), .A3(new_n1156), .A4(new_n1158), .ZN(new_n1159));
  INV_X1    g734(.A(KEYINPUT119), .ZN(new_n1160));
  NAND2_X1  g735(.A1(new_n1159), .A2(new_n1160), .ZN(new_n1161));
  INV_X1    g736(.A(KEYINPUT61), .ZN(new_n1162));
  AOI22_X1  g737(.A1(new_n1152), .A2(new_n1153), .B1(new_n1051), .B2(new_n1157), .ZN(new_n1163));
  NAND4_X1  g738(.A1(new_n1163), .A2(KEYINPUT119), .A3(new_n1156), .A4(new_n1151), .ZN(new_n1164));
  NAND3_X1  g739(.A1(new_n1161), .A2(new_n1162), .A3(new_n1164), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n1051), .A2(new_n730), .ZN(new_n1166));
  NAND2_X1  g741(.A1(new_n1082), .A2(new_n1015), .ZN(new_n1167));
  AND4_X1   g742(.A1(KEYINPUT60), .A2(new_n947), .A3(new_n1166), .A4(new_n1167), .ZN(new_n1168));
  AOI22_X1  g743(.A1(new_n1051), .A2(new_n730), .B1(new_n1082), .B2(new_n1015), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1169), .A2(KEYINPUT60), .ZN(new_n1170));
  AOI21_X1  g745(.A(new_n947), .B1(new_n1169), .B2(KEYINPUT60), .ZN(new_n1171));
  AOI21_X1  g746(.A(new_n1168), .B1(new_n1170), .B2(new_n1171), .ZN(new_n1172));
  NAND3_X1  g747(.A1(new_n1151), .A2(new_n1154), .A3(new_n1158), .ZN(new_n1173));
  INV_X1    g748(.A(new_n1156), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n1173), .A2(new_n1174), .ZN(new_n1175));
  NAND3_X1  g750(.A1(new_n1175), .A2(KEYINPUT61), .A3(new_n1159), .ZN(new_n1176));
  XNOR2_X1  g751(.A(KEYINPUT58), .B(G1341), .ZN(new_n1177));
  OAI22_X1  g752(.A1(new_n1040), .A2(G1996), .B1(new_n1082), .B2(new_n1177), .ZN(new_n1178));
  INV_X1    g753(.A(KEYINPUT120), .ZN(new_n1179));
  NAND3_X1  g754(.A1(new_n1178), .A2(new_n1179), .A3(new_n559), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1180), .A2(KEYINPUT59), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT59), .ZN(new_n1182));
  NAND4_X1  g757(.A1(new_n1178), .A2(new_n1179), .A3(new_n1182), .A4(new_n559), .ZN(new_n1183));
  NAND2_X1  g758(.A1(new_n1181), .A2(new_n1183), .ZN(new_n1184));
  NAND4_X1  g759(.A1(new_n1165), .A2(new_n1172), .A3(new_n1176), .A4(new_n1184), .ZN(new_n1185));
  OAI21_X1  g760(.A(new_n1175), .B1(new_n947), .B2(new_n1169), .ZN(new_n1186));
  NAND2_X1  g761(.A1(new_n1161), .A2(new_n1164), .ZN(new_n1187));
  NAND2_X1  g762(.A1(new_n1186), .A2(new_n1187), .ZN(new_n1188));
  NAND2_X1  g763(.A1(new_n1185), .A2(new_n1188), .ZN(new_n1189));
  AOI21_X1  g764(.A(new_n1131), .B1(new_n1146), .B2(new_n1189), .ZN(new_n1190));
  OAI21_X1  g765(.A(new_n1130), .B1(new_n1190), .B2(new_n1114), .ZN(new_n1191));
  OAI21_X1  g766(.A(new_n1025), .B1(new_n1122), .B2(new_n1191), .ZN(new_n1192));
  AND2_X1   g767(.A1(new_n1013), .A2(new_n1019), .ZN(new_n1193));
  OR2_X1    g768(.A1(new_n1193), .A2(KEYINPUT46), .ZN(new_n1194));
  NAND2_X1  g769(.A1(new_n1193), .A2(KEYINPUT46), .ZN(new_n1195));
  OAI21_X1  g770(.A(new_n1013), .B1(new_n761), .B2(new_n1017), .ZN(new_n1196));
  NAND3_X1  g771(.A1(new_n1194), .A2(new_n1195), .A3(new_n1196), .ZN(new_n1197));
  XNOR2_X1  g772(.A(new_n1197), .B(KEYINPUT47), .ZN(new_n1198));
  NAND3_X1  g773(.A1(new_n1013), .A2(new_n717), .A3(new_n598), .ZN(new_n1199));
  INV_X1    g774(.A(KEYINPUT48), .ZN(new_n1200));
  OR2_X1    g775(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1201));
  NAND2_X1  g776(.A1(new_n1023), .A2(new_n1013), .ZN(new_n1202));
  NAND2_X1  g777(.A1(new_n1199), .A2(new_n1200), .ZN(new_n1203));
  NAND3_X1  g778(.A1(new_n1201), .A2(new_n1202), .A3(new_n1203), .ZN(new_n1204));
  NAND2_X1  g779(.A1(new_n1018), .A2(new_n1020), .ZN(new_n1205));
  OAI21_X1  g780(.A(new_n1016), .B1(new_n1205), .B2(new_n1021), .ZN(new_n1206));
  NAND2_X1  g781(.A1(new_n1206), .A2(new_n1013), .ZN(new_n1207));
  AND3_X1   g782(.A1(new_n1198), .A2(new_n1204), .A3(new_n1207), .ZN(new_n1208));
  NAND2_X1  g783(.A1(new_n1192), .A2(new_n1208), .ZN(G329));
  assign    G231 = 1'b0;
  NOR2_X1   g784(.A1(new_n1004), .A2(new_n1005), .ZN(new_n1211));
  OAI211_X1 g785(.A(new_n699), .B(G319), .C1(new_n723), .C2(new_n724), .ZN(new_n1212));
  AOI21_X1  g786(.A(new_n1212), .B1(new_n674), .B2(new_n675), .ZN(new_n1213));
  INV_X1    g787(.A(new_n912), .ZN(new_n1214));
  NAND2_X1  g788(.A1(new_n926), .A2(KEYINPUT105), .ZN(new_n1215));
  AOI21_X1  g789(.A(new_n1214), .B1(new_n1215), .B2(new_n916), .ZN(new_n1216));
  OAI21_X1  g790(.A(new_n883), .B1(new_n1216), .B2(new_n923), .ZN(new_n1217));
  INV_X1    g791(.A(new_n931), .ZN(new_n1218));
  OAI21_X1  g792(.A(new_n1213), .B1(new_n1217), .B2(new_n1218), .ZN(new_n1219));
  NOR2_X1   g793(.A1(new_n1211), .A2(new_n1219), .ZN(G308));
  OAI221_X1 g794(.A(new_n1213), .B1(new_n1218), .B2(new_n1217), .C1(new_n1004), .C2(new_n1005), .ZN(G225));
endmodule


