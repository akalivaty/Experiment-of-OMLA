//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 0 0 1 0 1 0 0 1 1 1 1 0 1 0 0 0 0 1 1 0 1 1 0 0 0 0 0 0 1 1 1 1 0 1 1 0 0 1 1 0 0 1 1 1 1 1 1 0 0 0 1 1 1 1 1 1 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:49 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n582, new_n583, new_n584, new_n585,
    new_n586, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n612, new_n613, new_n614, new_n615,
    new_n616, new_n617, new_n619, new_n620, new_n621, new_n622, new_n623,
    new_n624, new_n625, new_n626, new_n627, new_n629, new_n630, new_n631,
    new_n632, new_n633, new_n634, new_n635, new_n636, new_n637, new_n638,
    new_n639, new_n640, new_n642, new_n643, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n664, new_n665, new_n667, new_n668, new_n669,
    new_n670, new_n671, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n680, new_n681, new_n683, new_n685,
    new_n686, new_n687, new_n688, new_n689, new_n690, new_n691, new_n692,
    new_n693, new_n695, new_n696, new_n697, new_n698, new_n699, new_n700,
    new_n701, new_n702, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n710, new_n711, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n726, new_n728, new_n729, new_n730, new_n731, new_n732,
    new_n733, new_n734, new_n735, new_n736, new_n737, new_n738, new_n739,
    new_n740, new_n741, new_n742, new_n743, new_n744, new_n745, new_n746,
    new_n748, new_n749, new_n750, new_n751, new_n752, new_n753, new_n754,
    new_n756, new_n757, new_n758, new_n759, new_n760, new_n761, new_n762,
    new_n763, new_n764, new_n765, new_n766, new_n767, new_n768, new_n769,
    new_n770, new_n771, new_n772, new_n773, new_n774, new_n775, new_n776,
    new_n777, new_n778, new_n779, new_n780, new_n781, new_n782, new_n783,
    new_n784, new_n785, new_n786, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n891, new_n892, new_n893, new_n894, new_n895, new_n896, new_n897,
    new_n899, new_n900, new_n901, new_n902, new_n904, new_n905, new_n906,
    new_n907, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n942, new_n943,
    new_n945, new_n946, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n969, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980,
    new_n981, new_n982, new_n983, new_n984;
  INV_X1    g000(.A(G143), .ZN(new_n187));
  NOR2_X1   g001(.A1(new_n187), .A2(G146), .ZN(new_n188));
  INV_X1    g002(.A(new_n188), .ZN(new_n189));
  INV_X1    g003(.A(KEYINPUT64), .ZN(new_n190));
  AOI21_X1  g004(.A(new_n190), .B1(new_n187), .B2(G146), .ZN(new_n191));
  INV_X1    g005(.A(G146), .ZN(new_n192));
  NOR3_X1   g006(.A1(new_n192), .A2(KEYINPUT64), .A3(G143), .ZN(new_n193));
  OAI21_X1  g007(.A(new_n189), .B1(new_n191), .B2(new_n193), .ZN(new_n194));
  OR2_X1    g008(.A1(KEYINPUT0), .A2(G128), .ZN(new_n195));
  NAND2_X1  g009(.A1(KEYINPUT0), .A2(G128), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n194), .A2(new_n195), .A3(new_n196), .ZN(new_n197));
  NAND2_X1  g011(.A1(new_n197), .A2(KEYINPUT65), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT65), .ZN(new_n199));
  NAND4_X1  g013(.A1(new_n194), .A2(new_n199), .A3(new_n195), .A4(new_n196), .ZN(new_n200));
  INV_X1    g014(.A(KEYINPUT66), .ZN(new_n201));
  OAI21_X1  g015(.A(new_n201), .B1(new_n187), .B2(G146), .ZN(new_n202));
  NAND3_X1  g016(.A1(new_n192), .A2(KEYINPUT66), .A3(G143), .ZN(new_n203));
  AOI22_X1  g017(.A1(new_n202), .A2(new_n203), .B1(new_n187), .B2(G146), .ZN(new_n204));
  NAND3_X1  g018(.A1(new_n204), .A2(KEYINPUT0), .A3(G128), .ZN(new_n205));
  NAND3_X1  g019(.A1(new_n198), .A2(new_n200), .A3(new_n205), .ZN(new_n206));
  NAND2_X1  g020(.A1(new_n206), .A2(G125), .ZN(new_n207));
  NAND2_X1  g021(.A1(new_n202), .A2(new_n203), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n187), .A2(G146), .ZN(new_n209));
  XNOR2_X1  g023(.A(KEYINPUT68), .B(KEYINPUT1), .ZN(new_n210));
  NAND4_X1  g024(.A1(new_n208), .A2(G128), .A3(new_n209), .A4(new_n210), .ZN(new_n211));
  NAND2_X1  g025(.A1(new_n211), .A2(KEYINPUT69), .ZN(new_n212));
  INV_X1    g026(.A(KEYINPUT69), .ZN(new_n213));
  NAND4_X1  g027(.A1(new_n204), .A2(new_n213), .A3(G128), .A4(new_n210), .ZN(new_n214));
  OAI21_X1  g028(.A(G128), .B1(new_n210), .B2(new_n188), .ZN(new_n215));
  AOI22_X1  g029(.A1(new_n212), .A2(new_n214), .B1(new_n194), .B2(new_n215), .ZN(new_n216));
  INV_X1    g030(.A(G125), .ZN(new_n217));
  NAND2_X1  g031(.A1(new_n216), .A2(new_n217), .ZN(new_n218));
  NAND2_X1  g032(.A1(new_n207), .A2(new_n218), .ZN(new_n219));
  INV_X1    g033(.A(G953), .ZN(new_n220));
  AND2_X1   g034(.A1(new_n220), .A2(G224), .ZN(new_n221));
  INV_X1    g035(.A(KEYINPUT7), .ZN(new_n222));
  NOR2_X1   g036(.A1(new_n221), .A2(new_n222), .ZN(new_n223));
  XNOR2_X1  g037(.A(new_n219), .B(new_n223), .ZN(new_n224));
  INV_X1    g038(.A(G119), .ZN(new_n225));
  NAND2_X1  g039(.A1(new_n225), .A2(G116), .ZN(new_n226));
  INV_X1    g040(.A(G116), .ZN(new_n227));
  AND3_X1   g041(.A1(new_n227), .A2(KEYINPUT70), .A3(G119), .ZN(new_n228));
  AOI21_X1  g042(.A(KEYINPUT70), .B1(new_n227), .B2(G119), .ZN(new_n229));
  OAI211_X1 g043(.A(KEYINPUT5), .B(new_n226), .C1(new_n228), .C2(new_n229), .ZN(new_n230));
  NOR2_X1   g044(.A1(new_n226), .A2(KEYINPUT5), .ZN(new_n231));
  INV_X1    g045(.A(new_n231), .ZN(new_n232));
  NAND3_X1  g046(.A1(new_n230), .A2(G113), .A3(new_n232), .ZN(new_n233));
  NOR2_X1   g047(.A1(new_n227), .A2(G119), .ZN(new_n234));
  INV_X1    g048(.A(KEYINPUT70), .ZN(new_n235));
  OAI21_X1  g049(.A(new_n235), .B1(new_n225), .B2(G116), .ZN(new_n236));
  NAND3_X1  g050(.A1(new_n227), .A2(KEYINPUT70), .A3(G119), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n234), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  XOR2_X1   g052(.A(KEYINPUT2), .B(G113), .Z(new_n239));
  AND3_X1   g053(.A1(new_n238), .A2(KEYINPUT71), .A3(new_n239), .ZN(new_n240));
  AOI21_X1  g054(.A(KEYINPUT71), .B1(new_n238), .B2(new_n239), .ZN(new_n241));
  OAI21_X1  g055(.A(new_n233), .B1(new_n240), .B2(new_n241), .ZN(new_n242));
  INV_X1    g056(.A(G107), .ZN(new_n243));
  NAND3_X1  g057(.A1(new_n243), .A2(KEYINPUT83), .A3(G104), .ZN(new_n244));
  NAND2_X1  g058(.A1(new_n244), .A2(KEYINPUT3), .ZN(new_n245));
  NOR2_X1   g059(.A1(new_n243), .A2(G104), .ZN(new_n246));
  INV_X1    g060(.A(new_n246), .ZN(new_n247));
  INV_X1    g061(.A(G101), .ZN(new_n248));
  INV_X1    g062(.A(KEYINPUT3), .ZN(new_n249));
  NAND4_X1  g063(.A1(new_n249), .A2(new_n243), .A3(KEYINPUT83), .A4(G104), .ZN(new_n250));
  NAND4_X1  g064(.A1(new_n245), .A2(new_n247), .A3(new_n248), .A4(new_n250), .ZN(new_n251));
  INV_X1    g065(.A(G104), .ZN(new_n252));
  NOR2_X1   g066(.A1(new_n252), .A2(G107), .ZN(new_n253));
  OAI21_X1  g067(.A(G101), .B1(new_n253), .B2(new_n246), .ZN(new_n254));
  NAND2_X1  g068(.A1(new_n251), .A2(new_n254), .ZN(new_n255));
  NOR2_X1   g069(.A1(new_n242), .A2(new_n255), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n238), .A2(new_n239), .ZN(new_n257));
  INV_X1    g071(.A(KEYINPUT71), .ZN(new_n258));
  NAND2_X1  g072(.A1(new_n257), .A2(new_n258), .ZN(new_n259));
  NAND3_X1  g073(.A1(new_n238), .A2(KEYINPUT71), .A3(new_n239), .ZN(new_n260));
  AOI21_X1  g074(.A(new_n231), .B1(new_n238), .B2(KEYINPUT5), .ZN(new_n261));
  AOI22_X1  g075(.A1(new_n259), .A2(new_n260), .B1(new_n261), .B2(G113), .ZN(new_n262));
  INV_X1    g076(.A(new_n255), .ZN(new_n263));
  OAI21_X1  g077(.A(KEYINPUT86), .B1(new_n262), .B2(new_n263), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT86), .ZN(new_n265));
  NAND3_X1  g079(.A1(new_n242), .A2(new_n265), .A3(new_n255), .ZN(new_n266));
  AOI21_X1  g080(.A(new_n256), .B1(new_n264), .B2(new_n266), .ZN(new_n267));
  INV_X1    g081(.A(KEYINPUT87), .ZN(new_n268));
  XOR2_X1   g082(.A(G110), .B(G122), .Z(new_n269));
  XNOR2_X1  g083(.A(new_n269), .B(KEYINPUT8), .ZN(new_n270));
  NOR3_X1   g084(.A1(new_n267), .A2(new_n268), .A3(new_n270), .ZN(new_n271));
  NAND2_X1  g085(.A1(new_n262), .A2(new_n263), .ZN(new_n272));
  AND3_X1   g086(.A1(new_n242), .A2(new_n265), .A3(new_n255), .ZN(new_n273));
  AOI21_X1  g087(.A(new_n265), .B1(new_n242), .B2(new_n255), .ZN(new_n274));
  OAI21_X1  g088(.A(new_n272), .B1(new_n273), .B2(new_n274), .ZN(new_n275));
  INV_X1    g089(.A(new_n270), .ZN(new_n276));
  AOI21_X1  g090(.A(KEYINPUT87), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  OAI21_X1  g091(.A(new_n224), .B1(new_n271), .B2(new_n277), .ZN(new_n278));
  INV_X1    g092(.A(KEYINPUT88), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n278), .A2(new_n279), .ZN(new_n280));
  NAND3_X1  g094(.A1(new_n245), .A2(new_n247), .A3(new_n250), .ZN(new_n281));
  NAND2_X1  g095(.A1(new_n281), .A2(G101), .ZN(new_n282));
  NAND3_X1  g096(.A1(new_n282), .A2(KEYINPUT4), .A3(new_n251), .ZN(new_n283));
  INV_X1    g097(.A(KEYINPUT4), .ZN(new_n284));
  NAND3_X1  g098(.A1(new_n281), .A2(new_n284), .A3(G101), .ZN(new_n285));
  AND2_X1   g099(.A1(new_n283), .A2(new_n285), .ZN(new_n286));
  NOR2_X1   g100(.A1(new_n238), .A2(new_n239), .ZN(new_n287));
  AOI21_X1  g101(.A(new_n287), .B1(new_n259), .B2(new_n260), .ZN(new_n288));
  INV_X1    g102(.A(new_n288), .ZN(new_n289));
  NAND2_X1  g103(.A1(new_n286), .A2(new_n289), .ZN(new_n290));
  INV_X1    g104(.A(new_n269), .ZN(new_n291));
  NAND3_X1  g105(.A1(new_n290), .A2(new_n291), .A3(new_n272), .ZN(new_n292));
  OAI211_X1 g106(.A(new_n224), .B(KEYINPUT88), .C1(new_n271), .C2(new_n277), .ZN(new_n293));
  NAND3_X1  g107(.A1(new_n280), .A2(new_n292), .A3(new_n293), .ZN(new_n294));
  NAND2_X1  g108(.A1(new_n290), .A2(new_n272), .ZN(new_n295));
  NAND2_X1  g109(.A1(new_n295), .A2(new_n269), .ZN(new_n296));
  NAND3_X1  g110(.A1(new_n296), .A2(KEYINPUT6), .A3(new_n292), .ZN(new_n297));
  INV_X1    g111(.A(KEYINPUT6), .ZN(new_n298));
  NAND3_X1  g112(.A1(new_n295), .A2(new_n298), .A3(new_n269), .ZN(new_n299));
  NAND2_X1  g113(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  INV_X1    g114(.A(new_n300), .ZN(new_n301));
  XNOR2_X1  g115(.A(new_n219), .B(new_n221), .ZN(new_n302));
  AOI21_X1  g116(.A(G902), .B1(new_n301), .B2(new_n302), .ZN(new_n303));
  NAND2_X1  g117(.A1(new_n294), .A2(new_n303), .ZN(new_n304));
  OAI21_X1  g118(.A(G210), .B1(G237), .B2(G902), .ZN(new_n305));
  INV_X1    g119(.A(new_n305), .ZN(new_n306));
  NAND2_X1  g120(.A1(new_n304), .A2(new_n306), .ZN(new_n307));
  NAND3_X1  g121(.A1(new_n294), .A2(new_n303), .A3(new_n305), .ZN(new_n308));
  NAND2_X1  g122(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  INV_X1    g123(.A(G475), .ZN(new_n310));
  INV_X1    g124(.A(G902), .ZN(new_n311));
  AND2_X1   g125(.A1(KEYINPUT79), .A2(G140), .ZN(new_n312));
  NOR2_X1   g126(.A1(KEYINPUT79), .A2(G140), .ZN(new_n313));
  OAI21_X1  g127(.A(G125), .B1(new_n312), .B2(new_n313), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n314), .A2(KEYINPUT80), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n217), .A2(G140), .ZN(new_n316));
  INV_X1    g130(.A(KEYINPUT80), .ZN(new_n317));
  OAI211_X1 g131(.A(new_n317), .B(G125), .C1(new_n312), .C2(new_n313), .ZN(new_n318));
  NAND3_X1  g132(.A1(new_n315), .A2(new_n316), .A3(new_n318), .ZN(new_n319));
  AND2_X1   g133(.A1(new_n319), .A2(KEYINPUT16), .ZN(new_n320));
  INV_X1    g134(.A(G140), .ZN(new_n321));
  AOI21_X1  g135(.A(KEYINPUT16), .B1(new_n321), .B2(G125), .ZN(new_n322));
  OAI21_X1  g136(.A(G146), .B1(new_n320), .B2(new_n322), .ZN(new_n323));
  NAND2_X1  g137(.A1(new_n220), .A2(KEYINPUT72), .ZN(new_n324));
  INV_X1    g138(.A(KEYINPUT72), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G953), .ZN(new_n326));
  NAND2_X1  g140(.A1(new_n324), .A2(new_n326), .ZN(new_n327));
  INV_X1    g141(.A(G237), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n327), .A2(G214), .A3(new_n328), .ZN(new_n329));
  XOR2_X1   g143(.A(KEYINPUT89), .B(G143), .Z(new_n330));
  NAND2_X1  g144(.A1(new_n329), .A2(new_n330), .ZN(new_n331));
  AOI21_X1  g145(.A(G237), .B1(new_n324), .B2(new_n326), .ZN(new_n332));
  NOR2_X1   g146(.A1(KEYINPUT89), .A2(G143), .ZN(new_n333));
  NAND3_X1  g147(.A1(new_n332), .A2(G214), .A3(new_n333), .ZN(new_n334));
  NAND2_X1  g148(.A1(new_n331), .A2(new_n334), .ZN(new_n335));
  INV_X1    g149(.A(G131), .ZN(new_n336));
  NAND2_X1  g150(.A1(new_n335), .A2(new_n336), .ZN(new_n337));
  INV_X1    g151(.A(KEYINPUT17), .ZN(new_n338));
  NAND3_X1  g152(.A1(new_n331), .A2(G131), .A3(new_n334), .ZN(new_n339));
  NAND3_X1  g153(.A1(new_n337), .A2(new_n338), .A3(new_n339), .ZN(new_n340));
  AOI21_X1  g154(.A(new_n322), .B1(new_n319), .B2(KEYINPUT16), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(new_n192), .ZN(new_n342));
  OR2_X1    g156(.A1(new_n339), .A2(new_n338), .ZN(new_n343));
  NAND4_X1  g157(.A1(new_n323), .A2(new_n340), .A3(new_n342), .A4(new_n343), .ZN(new_n344));
  XNOR2_X1  g158(.A(G113), .B(G122), .ZN(new_n345));
  XNOR2_X1  g159(.A(new_n345), .B(new_n252), .ZN(new_n346));
  INV_X1    g160(.A(KEYINPUT18), .ZN(new_n347));
  OAI21_X1  g161(.A(new_n335), .B1(new_n347), .B2(new_n336), .ZN(new_n348));
  NAND2_X1  g162(.A1(new_n319), .A2(G146), .ZN(new_n349));
  NAND2_X1  g163(.A1(new_n321), .A2(G125), .ZN(new_n350));
  NAND3_X1  g164(.A1(new_n316), .A2(new_n350), .A3(new_n192), .ZN(new_n351));
  NAND2_X1  g165(.A1(new_n349), .A2(new_n351), .ZN(new_n352));
  OAI211_X1 g166(.A(new_n348), .B(new_n352), .C1(new_n347), .C2(new_n339), .ZN(new_n353));
  AND3_X1   g167(.A1(new_n344), .A2(new_n346), .A3(new_n353), .ZN(new_n354));
  NAND2_X1  g168(.A1(new_n337), .A2(new_n339), .ZN(new_n355));
  NAND2_X1  g169(.A1(new_n319), .A2(KEYINPUT19), .ZN(new_n356));
  NAND2_X1  g170(.A1(new_n316), .A2(new_n350), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n356), .B1(KEYINPUT19), .B2(new_n357), .ZN(new_n358));
  OAI211_X1 g172(.A(new_n323), .B(new_n355), .C1(G146), .C2(new_n358), .ZN(new_n359));
  AOI21_X1  g173(.A(new_n346), .B1(new_n359), .B2(new_n353), .ZN(new_n360));
  OAI211_X1 g174(.A(new_n310), .B(new_n311), .C1(new_n354), .C2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT20), .ZN(new_n362));
  NAND2_X1  g176(.A1(new_n361), .A2(new_n362), .ZN(new_n363));
  NAND2_X1  g177(.A1(new_n323), .A2(new_n355), .ZN(new_n364));
  NOR2_X1   g178(.A1(new_n358), .A2(G146), .ZN(new_n365));
  OAI21_X1  g179(.A(new_n353), .B1(new_n364), .B2(new_n365), .ZN(new_n366));
  INV_X1    g180(.A(new_n346), .ZN(new_n367));
  NAND2_X1  g181(.A1(new_n366), .A2(new_n367), .ZN(new_n368));
  NAND3_X1  g182(.A1(new_n344), .A2(new_n346), .A3(new_n353), .ZN(new_n369));
  NAND2_X1  g183(.A1(new_n368), .A2(new_n369), .ZN(new_n370));
  NAND4_X1  g184(.A1(new_n370), .A2(KEYINPUT20), .A3(new_n310), .A4(new_n311), .ZN(new_n371));
  AOI21_X1  g185(.A(new_n346), .B1(new_n344), .B2(new_n353), .ZN(new_n372));
  OAI21_X1  g186(.A(new_n311), .B1(new_n354), .B2(new_n372), .ZN(new_n373));
  NAND2_X1  g187(.A1(new_n373), .A2(G475), .ZN(new_n374));
  NAND3_X1  g188(.A1(new_n363), .A2(new_n371), .A3(new_n374), .ZN(new_n375));
  INV_X1    g189(.A(G478), .ZN(new_n376));
  NOR2_X1   g190(.A1(new_n376), .A2(KEYINPUT15), .ZN(new_n377));
  NAND2_X1  g191(.A1(new_n187), .A2(G128), .ZN(new_n378));
  INV_X1    g192(.A(G128), .ZN(new_n379));
  NAND2_X1  g193(.A1(new_n379), .A2(G143), .ZN(new_n380));
  AND2_X1   g194(.A1(new_n378), .A2(new_n380), .ZN(new_n381));
  INV_X1    g195(.A(G134), .ZN(new_n382));
  XNOR2_X1  g196(.A(new_n381), .B(new_n382), .ZN(new_n383));
  NAND2_X1  g197(.A1(new_n227), .A2(G122), .ZN(new_n384));
  NAND2_X1  g198(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n385));
  INV_X1    g199(.A(G122), .ZN(new_n386));
  NAND2_X1  g200(.A1(new_n386), .A2(G116), .ZN(new_n387));
  NAND2_X1  g201(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NOR2_X1   g202(.A1(new_n384), .A2(KEYINPUT14), .ZN(new_n389));
  OAI21_X1  g203(.A(G107), .B1(new_n388), .B2(new_n389), .ZN(new_n390));
  AND3_X1   g204(.A1(new_n387), .A2(new_n384), .A3(new_n243), .ZN(new_n391));
  INV_X1    g205(.A(KEYINPUT91), .ZN(new_n392));
  OR2_X1    g206(.A1(new_n391), .A2(new_n392), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n391), .A2(new_n392), .ZN(new_n394));
  NAND4_X1  g208(.A1(new_n383), .A2(new_n390), .A3(new_n393), .A4(new_n394), .ZN(new_n395));
  INV_X1    g209(.A(KEYINPUT13), .ZN(new_n396));
  OAI21_X1  g210(.A(KEYINPUT90), .B1(new_n378), .B2(new_n396), .ZN(new_n397));
  NAND2_X1  g211(.A1(new_n378), .A2(new_n396), .ZN(new_n398));
  INV_X1    g212(.A(KEYINPUT90), .ZN(new_n399));
  NAND4_X1  g213(.A1(new_n399), .A2(new_n187), .A3(KEYINPUT13), .A4(G128), .ZN(new_n400));
  NAND4_X1  g214(.A1(new_n397), .A2(new_n398), .A3(new_n400), .A4(new_n380), .ZN(new_n401));
  NAND2_X1  g215(.A1(new_n401), .A2(G134), .ZN(new_n402));
  NAND2_X1  g216(.A1(new_n381), .A2(new_n382), .ZN(new_n403));
  AND2_X1   g217(.A1(new_n387), .A2(new_n384), .ZN(new_n404));
  NOR2_X1   g218(.A1(new_n404), .A2(new_n243), .ZN(new_n405));
  OAI211_X1 g219(.A(new_n402), .B(new_n403), .C1(new_n405), .C2(new_n391), .ZN(new_n406));
  NAND2_X1  g220(.A1(new_n395), .A2(new_n406), .ZN(new_n407));
  XOR2_X1   g221(.A(KEYINPUT76), .B(G217), .Z(new_n408));
  XOR2_X1   g222(.A(KEYINPUT9), .B(G234), .Z(new_n409));
  NAND3_X1  g223(.A1(new_n408), .A2(new_n409), .A3(new_n220), .ZN(new_n410));
  AND2_X1   g224(.A1(new_n407), .A2(new_n410), .ZN(new_n411));
  NOR2_X1   g225(.A1(new_n407), .A2(new_n410), .ZN(new_n412));
  OAI21_X1  g226(.A(new_n311), .B1(new_n411), .B2(new_n412), .ZN(new_n413));
  INV_X1    g227(.A(KEYINPUT92), .ZN(new_n414));
  NOR2_X1   g228(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  XNOR2_X1  g229(.A(new_n407), .B(new_n410), .ZN(new_n416));
  AOI21_X1  g230(.A(KEYINPUT92), .B1(new_n416), .B2(new_n311), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n377), .B1(new_n415), .B2(new_n417), .ZN(new_n418));
  OAI21_X1  g232(.A(new_n418), .B1(new_n377), .B2(new_n417), .ZN(new_n419));
  INV_X1    g233(.A(G234), .ZN(new_n420));
  OAI211_X1 g234(.A(G952), .B(new_n220), .C1(new_n420), .C2(new_n328), .ZN(new_n421));
  XNOR2_X1  g235(.A(new_n421), .B(KEYINPUT93), .ZN(new_n422));
  INV_X1    g236(.A(new_n327), .ZN(new_n423));
  OAI211_X1 g237(.A(new_n423), .B(G902), .C1(new_n420), .C2(new_n328), .ZN(new_n424));
  XOR2_X1   g238(.A(KEYINPUT21), .B(G898), .Z(new_n425));
  OAI21_X1  g239(.A(new_n422), .B1(new_n424), .B2(new_n425), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NOR3_X1   g241(.A1(new_n375), .A2(new_n419), .A3(new_n427), .ZN(new_n428));
  INV_X1    g242(.A(G221), .ZN(new_n429));
  AOI21_X1  g243(.A(new_n429), .B1(new_n409), .B2(new_n311), .ZN(new_n430));
  INV_X1    g244(.A(G469), .ZN(new_n431));
  NAND2_X1  g245(.A1(new_n327), .A2(G227), .ZN(new_n432));
  XNOR2_X1  g246(.A(G110), .B(G140), .ZN(new_n433));
  XNOR2_X1  g247(.A(new_n432), .B(new_n433), .ZN(new_n434));
  AND3_X1   g248(.A1(new_n198), .A2(new_n200), .A3(new_n205), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n286), .A3(KEYINPUT84), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT84), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n283), .A2(new_n285), .ZN(new_n438));
  OAI21_X1  g252(.A(new_n437), .B1(new_n206), .B2(new_n438), .ZN(new_n439));
  NAND2_X1  g253(.A1(new_n436), .A2(new_n439), .ZN(new_n440));
  NAND2_X1  g254(.A1(new_n212), .A2(new_n214), .ZN(new_n441));
  AOI21_X1  g255(.A(new_n379), .B1(new_n189), .B2(KEYINPUT1), .ZN(new_n442));
  OR2_X1    g256(.A1(new_n442), .A2(new_n204), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n441), .A2(new_n443), .ZN(new_n444));
  INV_X1    g258(.A(KEYINPUT10), .ZN(new_n445));
  NAND3_X1  g259(.A1(new_n444), .A2(new_n445), .A3(new_n263), .ZN(new_n446));
  OAI21_X1  g260(.A(KEYINPUT10), .B1(new_n216), .B2(new_n255), .ZN(new_n447));
  NAND2_X1  g261(.A1(new_n446), .A2(new_n447), .ZN(new_n448));
  NAND2_X1  g262(.A1(new_n440), .A2(new_n448), .ZN(new_n449));
  INV_X1    g263(.A(KEYINPUT85), .ZN(new_n450));
  INV_X1    g264(.A(KEYINPUT11), .ZN(new_n451));
  OAI21_X1  g265(.A(new_n451), .B1(new_n382), .B2(G137), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n382), .A2(G137), .ZN(new_n453));
  INV_X1    g267(.A(G137), .ZN(new_n454));
  NAND3_X1  g268(.A1(new_n454), .A2(KEYINPUT11), .A3(G134), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n452), .A2(new_n453), .A3(new_n455), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n456), .A2(G131), .ZN(new_n457));
  NAND4_X1  g271(.A1(new_n452), .A2(new_n455), .A3(new_n336), .A4(new_n453), .ZN(new_n458));
  NAND2_X1  g272(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  NAND3_X1  g273(.A1(new_n449), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  AOI22_X1  g274(.A1(new_n436), .A2(new_n439), .B1(new_n446), .B2(new_n447), .ZN(new_n461));
  INV_X1    g275(.A(new_n459), .ZN(new_n462));
  OAI21_X1  g276(.A(KEYINPUT85), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  NAND2_X1  g277(.A1(new_n460), .A2(new_n463), .ZN(new_n464));
  NAND3_X1  g278(.A1(new_n440), .A2(new_n462), .A3(new_n448), .ZN(new_n465));
  AOI21_X1  g279(.A(new_n434), .B1(new_n464), .B2(new_n465), .ZN(new_n466));
  NAND2_X1  g280(.A1(new_n215), .A2(new_n194), .ZN(new_n467));
  AND3_X1   g281(.A1(new_n441), .A2(new_n467), .A3(new_n255), .ZN(new_n468));
  AOI21_X1  g282(.A(new_n255), .B1(new_n441), .B2(new_n443), .ZN(new_n469));
  OAI21_X1  g283(.A(new_n459), .B1(new_n468), .B2(new_n469), .ZN(new_n470));
  INV_X1    g284(.A(KEYINPUT12), .ZN(new_n471));
  NAND2_X1  g285(.A1(new_n470), .A2(new_n471), .ZN(new_n472));
  OAI211_X1 g286(.A(KEYINPUT12), .B(new_n459), .C1(new_n468), .C2(new_n469), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n472), .A2(new_n473), .ZN(new_n474));
  INV_X1    g288(.A(new_n474), .ZN(new_n475));
  NAND2_X1  g289(.A1(new_n465), .A2(new_n434), .ZN(new_n476));
  NOR2_X1   g290(.A1(new_n475), .A2(new_n476), .ZN(new_n477));
  OAI211_X1 g291(.A(new_n431), .B(new_n311), .C1(new_n466), .C2(new_n477), .ZN(new_n478));
  AOI21_X1  g292(.A(new_n434), .B1(new_n474), .B2(new_n465), .ZN(new_n479));
  INV_X1    g293(.A(new_n476), .ZN(new_n480));
  AOI21_X1  g294(.A(new_n479), .B1(new_n464), .B2(new_n480), .ZN(new_n481));
  OAI21_X1  g295(.A(G469), .B1(new_n481), .B2(G902), .ZN(new_n482));
  AOI21_X1  g296(.A(new_n430), .B1(new_n478), .B2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(G214), .B1(G237), .B2(G902), .ZN(new_n484));
  NAND4_X1  g298(.A1(new_n309), .A2(new_n428), .A3(new_n483), .A4(new_n484), .ZN(new_n485));
  INV_X1    g299(.A(new_n485), .ZN(new_n486));
  INV_X1    g300(.A(KEYINPUT23), .ZN(new_n487));
  OAI21_X1  g301(.A(new_n487), .B1(new_n225), .B2(G128), .ZN(new_n488));
  NAND3_X1  g302(.A1(new_n379), .A2(KEYINPUT23), .A3(G119), .ZN(new_n489));
  OAI211_X1 g303(.A(new_n488), .B(new_n489), .C1(G119), .C2(new_n379), .ZN(new_n490));
  NAND2_X1  g304(.A1(new_n490), .A2(G110), .ZN(new_n491));
  XNOR2_X1  g305(.A(KEYINPUT24), .B(G110), .ZN(new_n492));
  XNOR2_X1  g306(.A(new_n492), .B(KEYINPUT78), .ZN(new_n493));
  XNOR2_X1  g307(.A(G119), .B(G128), .ZN(new_n494));
  NAND2_X1  g308(.A1(new_n493), .A2(new_n494), .ZN(new_n495));
  NOR2_X1   g309(.A1(new_n341), .A2(new_n192), .ZN(new_n496));
  AOI211_X1 g310(.A(G146), .B(new_n322), .C1(new_n319), .C2(KEYINPUT16), .ZN(new_n497));
  OAI211_X1 g311(.A(new_n491), .B(new_n495), .C1(new_n496), .C2(new_n497), .ZN(new_n498));
  OAI22_X1  g312(.A1(new_n493), .A2(new_n494), .B1(G110), .B2(new_n490), .ZN(new_n499));
  NAND3_X1  g313(.A1(new_n323), .A2(new_n351), .A3(new_n499), .ZN(new_n500));
  NAND2_X1  g314(.A1(new_n498), .A2(new_n500), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n327), .A2(G221), .A3(G234), .ZN(new_n502));
  XOR2_X1   g316(.A(new_n502), .B(KEYINPUT22), .Z(new_n503));
  XNOR2_X1  g317(.A(new_n503), .B(new_n454), .ZN(new_n504));
  INV_X1    g318(.A(new_n504), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n501), .A2(new_n505), .ZN(new_n506));
  NAND3_X1  g320(.A1(new_n498), .A2(new_n504), .A3(new_n500), .ZN(new_n507));
  NAND3_X1  g321(.A1(new_n506), .A2(new_n311), .A3(new_n507), .ZN(new_n508));
  AOI21_X1  g322(.A(KEYINPUT81), .B1(KEYINPUT82), .B2(KEYINPUT25), .ZN(new_n509));
  INV_X1    g323(.A(new_n509), .ZN(new_n510));
  NAND2_X1  g324(.A1(new_n508), .A2(new_n510), .ZN(new_n511));
  OAI21_X1  g325(.A(new_n408), .B1(new_n420), .B2(G902), .ZN(new_n512));
  XNOR2_X1  g326(.A(new_n512), .B(KEYINPUT77), .ZN(new_n513));
  INV_X1    g327(.A(new_n513), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n511), .A2(new_n514), .ZN(new_n515));
  INV_X1    g329(.A(KEYINPUT81), .ZN(new_n516));
  NAND4_X1  g330(.A1(new_n506), .A2(new_n516), .A3(new_n311), .A4(new_n507), .ZN(new_n517));
  AOI21_X1  g331(.A(KEYINPUT25), .B1(new_n517), .B2(KEYINPUT82), .ZN(new_n518));
  NOR2_X1   g332(.A1(new_n515), .A2(new_n518), .ZN(new_n519));
  INV_X1    g333(.A(new_n519), .ZN(new_n520));
  AND2_X1   g334(.A1(new_n506), .A2(new_n507), .ZN(new_n521));
  AOI21_X1  g335(.A(G902), .B1(new_n408), .B2(new_n420), .ZN(new_n522));
  NAND2_X1  g336(.A1(new_n521), .A2(new_n522), .ZN(new_n523));
  NAND2_X1  g337(.A1(new_n520), .A2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(KEYINPUT75), .ZN(new_n525));
  INV_X1    g339(.A(KEYINPUT28), .ZN(new_n526));
  NAND4_X1  g340(.A1(new_n198), .A2(new_n459), .A3(new_n200), .A4(new_n205), .ZN(new_n527));
  INV_X1    g341(.A(new_n527), .ZN(new_n528));
  INV_X1    g342(.A(KEYINPUT67), .ZN(new_n529));
  OAI21_X1  g343(.A(new_n529), .B1(new_n382), .B2(G137), .ZN(new_n530));
  NAND3_X1  g344(.A1(new_n454), .A2(KEYINPUT67), .A3(G134), .ZN(new_n531));
  AND3_X1   g345(.A1(new_n530), .A2(new_n453), .A3(new_n531), .ZN(new_n532));
  OAI21_X1  g346(.A(new_n458), .B1(new_n532), .B2(new_n336), .ZN(new_n533));
  AOI21_X1  g347(.A(new_n533), .B1(new_n441), .B2(new_n467), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n289), .B1(new_n528), .B2(new_n534), .ZN(new_n535));
  OAI211_X1 g349(.A(new_n527), .B(new_n288), .C1(new_n216), .C2(new_n533), .ZN(new_n536));
  AOI21_X1  g350(.A(new_n526), .B1(new_n535), .B2(new_n536), .ZN(new_n537));
  AND3_X1   g351(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n526), .ZN(new_n538));
  AOI21_X1  g352(.A(KEYINPUT74), .B1(new_n536), .B2(new_n526), .ZN(new_n539));
  NOR3_X1   g353(.A1(new_n537), .A2(new_n538), .A3(new_n539), .ZN(new_n540));
  INV_X1    g354(.A(KEYINPUT27), .ZN(new_n541));
  NAND3_X1  g355(.A1(new_n332), .A2(new_n541), .A3(G210), .ZN(new_n542));
  INV_X1    g356(.A(new_n542), .ZN(new_n543));
  AOI21_X1  g357(.A(new_n541), .B1(new_n332), .B2(G210), .ZN(new_n544));
  OAI21_X1  g358(.A(KEYINPUT26), .B1(new_n543), .B2(new_n544), .ZN(new_n545));
  INV_X1    g359(.A(new_n544), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT26), .ZN(new_n547));
  NAND3_X1  g361(.A1(new_n546), .A2(new_n547), .A3(new_n542), .ZN(new_n548));
  AND3_X1   g362(.A1(new_n545), .A2(new_n548), .A3(G101), .ZN(new_n549));
  AOI21_X1  g363(.A(G101), .B1(new_n545), .B2(new_n548), .ZN(new_n550));
  NOR2_X1   g364(.A1(new_n549), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g365(.A(new_n525), .B1(new_n540), .B2(new_n551), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n536), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n553), .A2(KEYINPUT73), .ZN(new_n554));
  INV_X1    g368(.A(KEYINPUT31), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT30), .ZN(new_n556));
  OAI21_X1  g370(.A(new_n556), .B1(new_n528), .B2(new_n534), .ZN(new_n557));
  OAI211_X1 g371(.A(new_n527), .B(KEYINPUT30), .C1(new_n216), .C2(new_n533), .ZN(new_n558));
  NAND3_X1  g372(.A1(new_n557), .A2(new_n289), .A3(new_n558), .ZN(new_n559));
  INV_X1    g373(.A(KEYINPUT73), .ZN(new_n560));
  NAND3_X1  g374(.A1(new_n551), .A2(new_n560), .A3(new_n536), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n554), .A2(new_n555), .A3(new_n559), .A4(new_n561), .ZN(new_n562));
  NAND3_X1  g376(.A1(new_n554), .A2(new_n559), .A3(new_n561), .ZN(new_n563));
  NAND2_X1  g377(.A1(new_n563), .A2(KEYINPUT31), .ZN(new_n564));
  INV_X1    g378(.A(new_n551), .ZN(new_n565));
  NAND2_X1  g379(.A1(new_n536), .A2(new_n526), .ZN(new_n566));
  INV_X1    g380(.A(KEYINPUT74), .ZN(new_n567));
  NAND2_X1  g381(.A1(new_n566), .A2(new_n567), .ZN(new_n568));
  NAND3_X1  g382(.A1(new_n536), .A2(KEYINPUT74), .A3(new_n526), .ZN(new_n569));
  NAND2_X1  g383(.A1(new_n568), .A2(new_n569), .ZN(new_n570));
  OAI211_X1 g384(.A(KEYINPUT75), .B(new_n565), .C1(new_n570), .C2(new_n537), .ZN(new_n571));
  NAND4_X1  g385(.A1(new_n552), .A2(new_n562), .A3(new_n564), .A4(new_n571), .ZN(new_n572));
  NOR2_X1   g386(.A1(G472), .A2(G902), .ZN(new_n573));
  AND3_X1   g387(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n574));
  AOI21_X1  g388(.A(KEYINPUT32), .B1(new_n572), .B2(new_n573), .ZN(new_n575));
  NOR2_X1   g389(.A1(new_n574), .A2(new_n575), .ZN(new_n576));
  NAND2_X1  g390(.A1(new_n540), .A2(new_n551), .ZN(new_n577));
  INV_X1    g391(.A(KEYINPUT29), .ZN(new_n578));
  NAND2_X1  g392(.A1(new_n559), .A2(new_n536), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n579), .A2(new_n565), .ZN(new_n580));
  NAND3_X1  g394(.A1(new_n577), .A2(new_n578), .A3(new_n580), .ZN(new_n581));
  NAND2_X1  g395(.A1(new_n581), .A2(new_n311), .ZN(new_n582));
  NOR2_X1   g396(.A1(new_n577), .A2(new_n578), .ZN(new_n583));
  OAI21_X1  g397(.A(G472), .B1(new_n582), .B2(new_n583), .ZN(new_n584));
  AOI21_X1  g398(.A(new_n524), .B1(new_n576), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g399(.A1(new_n486), .A2(new_n585), .ZN(new_n586));
  XNOR2_X1  g400(.A(new_n586), .B(G101), .ZN(G3));
  INV_X1    g401(.A(new_n430), .ZN(new_n588));
  OAI211_X1 g402(.A(new_n523), .B(new_n588), .C1(new_n515), .C2(new_n518), .ZN(new_n589));
  AOI21_X1  g403(.A(new_n589), .B1(new_n478), .B2(new_n482), .ZN(new_n590));
  NAND2_X1  g404(.A1(new_n572), .A2(new_n573), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n572), .A2(new_n311), .ZN(new_n592));
  NAND2_X1  g406(.A1(new_n592), .A2(G472), .ZN(new_n593));
  NAND3_X1  g407(.A1(new_n590), .A2(new_n591), .A3(new_n593), .ZN(new_n594));
  AND3_X1   g408(.A1(new_n294), .A2(new_n305), .A3(new_n303), .ZN(new_n595));
  AOI21_X1  g409(.A(new_n305), .B1(new_n294), .B2(new_n303), .ZN(new_n596));
  OAI211_X1 g410(.A(new_n426), .B(new_n484), .C1(new_n595), .C2(new_n596), .ZN(new_n597));
  NOR2_X1   g411(.A1(new_n594), .A2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(KEYINPUT33), .ZN(new_n599));
  INV_X1    g413(.A(KEYINPUT94), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n599), .B1(new_n410), .B2(new_n600), .ZN(new_n601));
  XNOR2_X1  g415(.A(new_n416), .B(new_n601), .ZN(new_n602));
  NAND3_X1  g416(.A1(new_n602), .A2(G478), .A3(new_n311), .ZN(new_n603));
  XOR2_X1   g417(.A(KEYINPUT95), .B(G478), .Z(new_n604));
  NAND2_X1  g418(.A1(new_n413), .A2(new_n604), .ZN(new_n605));
  NAND2_X1  g419(.A1(new_n603), .A2(new_n605), .ZN(new_n606));
  NAND2_X1  g420(.A1(new_n606), .A2(new_n375), .ZN(new_n607));
  XOR2_X1   g421(.A(new_n607), .B(KEYINPUT96), .Z(new_n608));
  NAND2_X1  g422(.A1(new_n598), .A2(new_n608), .ZN(new_n609));
  XOR2_X1   g423(.A(KEYINPUT34), .B(G104), .Z(new_n610));
  XNOR2_X1  g424(.A(new_n609), .B(new_n610), .ZN(G6));
  INV_X1    g425(.A(new_n375), .ZN(new_n612));
  NAND2_X1  g426(.A1(new_n612), .A2(new_n419), .ZN(new_n613));
  INV_X1    g427(.A(new_n613), .ZN(new_n614));
  NAND2_X1  g428(.A1(new_n598), .A2(new_n614), .ZN(new_n615));
  XNOR2_X1  g429(.A(KEYINPUT35), .B(G107), .ZN(new_n616));
  XNOR2_X1  g430(.A(new_n616), .B(KEYINPUT97), .ZN(new_n617));
  XNOR2_X1  g431(.A(new_n615), .B(new_n617), .ZN(G9));
  NOR2_X1   g432(.A1(new_n505), .A2(KEYINPUT36), .ZN(new_n619));
  XNOR2_X1  g433(.A(new_n619), .B(new_n501), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n620), .A2(new_n522), .ZN(new_n621));
  NAND2_X1  g435(.A1(new_n520), .A2(new_n621), .ZN(new_n622));
  NAND3_X1  g436(.A1(new_n593), .A2(new_n591), .A3(new_n622), .ZN(new_n623));
  INV_X1    g437(.A(new_n623), .ZN(new_n624));
  NAND2_X1  g438(.A1(new_n486), .A2(new_n624), .ZN(new_n625));
  XNOR2_X1  g439(.A(new_n625), .B(KEYINPUT98), .ZN(new_n626));
  XOR2_X1   g440(.A(KEYINPUT37), .B(G110), .Z(new_n627));
  XNOR2_X1  g441(.A(new_n626), .B(new_n627), .ZN(G12));
  OAI21_X1  g442(.A(new_n484), .B1(new_n595), .B2(new_n596), .ZN(new_n629));
  NAND2_X1  g443(.A1(new_n478), .A2(new_n482), .ZN(new_n630));
  NAND2_X1  g444(.A1(new_n630), .A2(new_n588), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n629), .A2(new_n631), .ZN(new_n632));
  INV_X1    g446(.A(KEYINPUT32), .ZN(new_n633));
  NAND2_X1  g447(.A1(new_n591), .A2(new_n633), .ZN(new_n634));
  NAND3_X1  g448(.A1(new_n572), .A2(KEYINPUT32), .A3(new_n573), .ZN(new_n635));
  NAND3_X1  g449(.A1(new_n634), .A2(new_n635), .A3(new_n584), .ZN(new_n636));
  OAI21_X1  g450(.A(new_n422), .B1(new_n424), .B2(G900), .ZN(new_n637));
  INV_X1    g451(.A(new_n637), .ZN(new_n638));
  NOR2_X1   g452(.A1(new_n613), .A2(new_n638), .ZN(new_n639));
  NAND4_X1  g453(.A1(new_n632), .A2(new_n636), .A3(new_n622), .A4(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(new_n640), .B(G128), .ZN(G30));
  XNOR2_X1  g455(.A(new_n637), .B(KEYINPUT101), .ZN(new_n642));
  XNOR2_X1  g456(.A(new_n642), .B(KEYINPUT39), .ZN(new_n643));
  OR2_X1    g457(.A1(new_n631), .A2(new_n643), .ZN(new_n644));
  OR2_X1    g458(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n645));
  NAND2_X1  g459(.A1(new_n644), .A2(KEYINPUT102), .ZN(new_n646));
  NAND2_X1  g460(.A1(new_n645), .A2(new_n646), .ZN(new_n647));
  NAND2_X1  g461(.A1(new_n647), .A2(KEYINPUT40), .ZN(new_n648));
  NAND2_X1  g462(.A1(new_n535), .A2(new_n536), .ZN(new_n649));
  NAND2_X1  g463(.A1(new_n649), .A2(new_n565), .ZN(new_n650));
  AND2_X1   g464(.A1(new_n563), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g465(.A(G472), .B1(new_n651), .B2(G902), .ZN(new_n652));
  NAND2_X1  g466(.A1(new_n576), .A2(new_n652), .ZN(new_n653));
  AND3_X1   g467(.A1(new_n375), .A2(new_n419), .A3(new_n484), .ZN(new_n654));
  AND2_X1   g468(.A1(new_n653), .A2(new_n654), .ZN(new_n655));
  INV_X1    g469(.A(KEYINPUT40), .ZN(new_n656));
  NAND3_X1  g470(.A1(new_n645), .A2(new_n656), .A3(new_n646), .ZN(new_n657));
  XNOR2_X1  g471(.A(KEYINPUT99), .B(KEYINPUT38), .ZN(new_n658));
  XNOR2_X1  g472(.A(new_n658), .B(KEYINPUT100), .ZN(new_n659));
  XNOR2_X1  g473(.A(new_n309), .B(new_n659), .ZN(new_n660));
  NOR2_X1   g474(.A1(new_n660), .A2(new_n622), .ZN(new_n661));
  NAND4_X1  g475(.A1(new_n648), .A2(new_n655), .A3(new_n657), .A4(new_n661), .ZN(new_n662));
  XNOR2_X1  g476(.A(new_n662), .B(G143), .ZN(G45));
  NOR2_X1   g477(.A1(new_n607), .A2(new_n638), .ZN(new_n664));
  NAND4_X1  g478(.A1(new_n632), .A2(new_n636), .A3(new_n622), .A4(new_n664), .ZN(new_n665));
  XNOR2_X1  g479(.A(new_n665), .B(G146), .ZN(G48));
  AOI22_X1  g480(.A1(new_n460), .A2(new_n463), .B1(new_n462), .B2(new_n461), .ZN(new_n667));
  OAI22_X1  g481(.A1(new_n667), .A2(new_n434), .B1(new_n475), .B2(new_n476), .ZN(new_n668));
  NAND2_X1  g482(.A1(new_n668), .A2(new_n311), .ZN(new_n669));
  NAND2_X1  g483(.A1(new_n669), .A2(G469), .ZN(new_n670));
  NAND3_X1  g484(.A1(new_n670), .A2(new_n588), .A3(new_n478), .ZN(new_n671));
  INV_X1    g485(.A(KEYINPUT103), .ZN(new_n672));
  NAND2_X1  g486(.A1(new_n671), .A2(new_n672), .ZN(new_n673));
  INV_X1    g487(.A(new_n478), .ZN(new_n674));
  AOI21_X1  g488(.A(new_n431), .B1(new_n668), .B2(new_n311), .ZN(new_n675));
  NOR2_X1   g489(.A1(new_n674), .A2(new_n675), .ZN(new_n676));
  NAND3_X1  g490(.A1(new_n676), .A2(KEYINPUT103), .A3(new_n588), .ZN(new_n677));
  NAND2_X1  g491(.A1(new_n673), .A2(new_n677), .ZN(new_n678));
  INV_X1    g492(.A(new_n597), .ZN(new_n679));
  NAND4_X1  g493(.A1(new_n678), .A2(new_n585), .A3(new_n608), .A4(new_n679), .ZN(new_n680));
  XNOR2_X1  g494(.A(KEYINPUT41), .B(G113), .ZN(new_n681));
  XNOR2_X1  g495(.A(new_n680), .B(new_n681), .ZN(G15));
  NAND4_X1  g496(.A1(new_n678), .A2(new_n585), .A3(new_n679), .A4(new_n614), .ZN(new_n683));
  XNOR2_X1  g497(.A(new_n683), .B(G116), .ZN(G18));
  AOI21_X1  g498(.A(new_n519), .B1(new_n522), .B2(new_n620), .ZN(new_n685));
  AOI21_X1  g499(.A(new_n685), .B1(new_n576), .B2(new_n584), .ZN(new_n686));
  NOR2_X1   g500(.A1(new_n671), .A2(new_n629), .ZN(new_n687));
  NAND4_X1  g501(.A1(new_n686), .A2(KEYINPUT104), .A3(new_n687), .A4(new_n428), .ZN(new_n688));
  INV_X1    g502(.A(KEYINPUT104), .ZN(new_n689));
  NAND3_X1  g503(.A1(new_n636), .A2(new_n428), .A3(new_n622), .ZN(new_n690));
  NAND4_X1  g504(.A1(new_n676), .A2(new_n309), .A3(new_n484), .A4(new_n588), .ZN(new_n691));
  OAI21_X1  g505(.A(new_n689), .B1(new_n690), .B2(new_n691), .ZN(new_n692));
  NAND2_X1  g506(.A1(new_n688), .A2(new_n692), .ZN(new_n693));
  XNOR2_X1  g507(.A(new_n693), .B(G119), .ZN(G21));
  OAI21_X1  g508(.A(new_n654), .B1(new_n595), .B2(new_n596), .ZN(new_n695));
  NAND2_X1  g509(.A1(new_n695), .A2(KEYINPUT105), .ZN(new_n696));
  INV_X1    g510(.A(KEYINPUT105), .ZN(new_n697));
  OAI211_X1 g511(.A(new_n654), .B(new_n697), .C1(new_n595), .C2(new_n596), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n696), .A2(new_n698), .ZN(new_n699));
  AND2_X1   g513(.A1(new_n564), .A2(new_n562), .ZN(new_n700));
  OAI21_X1  g514(.A(new_n565), .B1(new_n570), .B2(new_n537), .ZN(new_n701));
  NAND2_X1  g515(.A1(new_n700), .A2(new_n701), .ZN(new_n702));
  NAND2_X1  g516(.A1(new_n702), .A2(new_n573), .ZN(new_n703));
  INV_X1    g517(.A(new_n703), .ZN(new_n704));
  INV_X1    g518(.A(G472), .ZN(new_n705));
  AOI21_X1  g519(.A(new_n705), .B1(new_n572), .B2(new_n311), .ZN(new_n706));
  NOR3_X1   g520(.A1(new_n704), .A2(new_n706), .A3(new_n524), .ZN(new_n707));
  NAND4_X1  g521(.A1(new_n678), .A2(new_n699), .A3(new_n426), .A4(new_n707), .ZN(new_n708));
  XNOR2_X1  g522(.A(new_n708), .B(G122), .ZN(G24));
  NOR3_X1   g523(.A1(new_n704), .A2(new_n685), .A3(new_n706), .ZN(new_n710));
  NAND3_X1  g524(.A1(new_n687), .A2(new_n664), .A3(new_n710), .ZN(new_n711));
  XNOR2_X1  g525(.A(new_n711), .B(G125), .ZN(G27));
  INV_X1    g526(.A(new_n589), .ZN(new_n713));
  NAND2_X1  g527(.A1(new_n630), .A2(new_n713), .ZN(new_n714));
  AOI21_X1  g528(.A(new_n714), .B1(new_n576), .B2(new_n584), .ZN(new_n715));
  INV_X1    g529(.A(new_n484), .ZN(new_n716));
  NOR3_X1   g530(.A1(new_n595), .A2(new_n596), .A3(new_n716), .ZN(new_n717));
  XOR2_X1   g531(.A(KEYINPUT106), .B(KEYINPUT42), .Z(new_n718));
  INV_X1    g532(.A(new_n718), .ZN(new_n719));
  NAND4_X1  g533(.A1(new_n715), .A2(new_n664), .A3(new_n717), .A4(new_n719), .ZN(new_n720));
  NAND4_X1  g534(.A1(new_n636), .A2(new_n717), .A3(new_n590), .A4(new_n664), .ZN(new_n721));
  NAND2_X1  g535(.A1(KEYINPUT106), .A2(KEYINPUT42), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n721), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n720), .A2(new_n723), .ZN(new_n724));
  XNOR2_X1  g538(.A(new_n724), .B(G131), .ZN(G33));
  AND4_X1   g539(.A1(new_n636), .A2(new_n590), .A3(new_n717), .A4(new_n639), .ZN(new_n726));
  XNOR2_X1  g540(.A(new_n726), .B(new_n382), .ZN(G36));
  OR2_X1    g541(.A1(new_n481), .A2(KEYINPUT45), .ZN(new_n728));
  NAND2_X1  g542(.A1(new_n481), .A2(KEYINPUT45), .ZN(new_n729));
  NAND3_X1  g543(.A1(new_n728), .A2(G469), .A3(new_n729), .ZN(new_n730));
  NAND2_X1  g544(.A1(G469), .A2(G902), .ZN(new_n731));
  AOI21_X1  g545(.A(KEYINPUT46), .B1(new_n730), .B2(new_n731), .ZN(new_n732));
  NOR2_X1   g546(.A1(new_n732), .A2(new_n674), .ZN(new_n733));
  NAND3_X1  g547(.A1(new_n730), .A2(KEYINPUT46), .A3(new_n731), .ZN(new_n734));
  NAND2_X1  g548(.A1(new_n733), .A2(new_n734), .ZN(new_n735));
  NAND2_X1  g549(.A1(new_n735), .A2(new_n588), .ZN(new_n736));
  NOR2_X1   g550(.A1(new_n736), .A2(new_n643), .ZN(new_n737));
  NAND3_X1  g551(.A1(new_n307), .A2(new_n484), .A3(new_n308), .ZN(new_n738));
  AOI21_X1  g552(.A(new_n685), .B1(new_n593), .B2(new_n591), .ZN(new_n739));
  NAND2_X1  g553(.A1(new_n612), .A2(new_n606), .ZN(new_n740));
  XOR2_X1   g554(.A(new_n740), .B(KEYINPUT43), .Z(new_n741));
  NAND2_X1  g555(.A1(new_n739), .A2(new_n741), .ZN(new_n742));
  INV_X1    g556(.A(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n738), .B1(new_n743), .B2(KEYINPUT44), .ZN(new_n744));
  OAI211_X1 g558(.A(new_n737), .B(new_n744), .C1(KEYINPUT44), .C2(new_n743), .ZN(new_n745));
  XNOR2_X1  g559(.A(new_n745), .B(KEYINPUT107), .ZN(new_n746));
  XNOR2_X1  g560(.A(new_n746), .B(G137), .ZN(G39));
  NAND2_X1  g561(.A1(new_n736), .A2(KEYINPUT47), .ZN(new_n748));
  INV_X1    g562(.A(new_n524), .ZN(new_n749));
  NOR2_X1   g563(.A1(new_n636), .A2(new_n749), .ZN(new_n750));
  INV_X1    g564(.A(KEYINPUT47), .ZN(new_n751));
  NAND3_X1  g565(.A1(new_n735), .A2(new_n751), .A3(new_n588), .ZN(new_n752));
  NOR3_X1   g566(.A1(new_n738), .A2(new_n607), .A3(new_n638), .ZN(new_n753));
  NAND4_X1  g567(.A1(new_n748), .A2(new_n750), .A3(new_n752), .A4(new_n753), .ZN(new_n754));
  XNOR2_X1  g568(.A(new_n754), .B(G140), .ZN(G42));
  INV_X1    g569(.A(KEYINPUT117), .ZN(new_n756));
  AOI22_X1  g570(.A1(new_n748), .A2(new_n752), .B1(new_n430), .B2(new_n676), .ZN(new_n757));
  OR3_X1    g571(.A1(new_n671), .A2(KEYINPUT116), .A3(new_n484), .ZN(new_n758));
  OAI21_X1  g572(.A(KEYINPUT116), .B1(new_n671), .B2(new_n484), .ZN(new_n759));
  NAND3_X1  g573(.A1(new_n758), .A2(new_n660), .A3(new_n759), .ZN(new_n760));
  OAI22_X1  g574(.A1(new_n757), .A2(new_n738), .B1(KEYINPUT50), .B2(new_n760), .ZN(new_n761));
  INV_X1    g575(.A(new_n422), .ZN(new_n762));
  AND2_X1   g576(.A1(new_n741), .A2(new_n762), .ZN(new_n763));
  NAND2_X1  g577(.A1(new_n763), .A2(new_n707), .ZN(new_n764));
  INV_X1    g578(.A(new_n764), .ZN(new_n765));
  NAND2_X1  g579(.A1(new_n761), .A2(new_n765), .ZN(new_n766));
  NOR2_X1   g580(.A1(new_n671), .A2(new_n738), .ZN(new_n767));
  NAND3_X1  g581(.A1(new_n763), .A2(new_n710), .A3(new_n767), .ZN(new_n768));
  OR2_X1    g582(.A1(new_n764), .A2(new_n760), .ZN(new_n769));
  NAND2_X1  g583(.A1(new_n769), .A2(KEYINPUT50), .ZN(new_n770));
  INV_X1    g584(.A(new_n653), .ZN(new_n771));
  NAND4_X1  g585(.A1(new_n771), .A2(new_n749), .A3(new_n762), .A4(new_n767), .ZN(new_n772));
  NOR2_X1   g586(.A1(new_n772), .A2(new_n606), .ZN(new_n773));
  NAND2_X1  g587(.A1(new_n773), .A2(new_n612), .ZN(new_n774));
  NAND2_X1  g588(.A1(new_n770), .A2(new_n774), .ZN(new_n775));
  INV_X1    g589(.A(new_n775), .ZN(new_n776));
  NAND3_X1  g590(.A1(new_n766), .A2(new_n768), .A3(new_n776), .ZN(new_n777));
  INV_X1    g591(.A(KEYINPUT51), .ZN(new_n778));
  OAI21_X1  g592(.A(new_n756), .B1(new_n777), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n220), .A2(G952), .ZN(new_n780));
  INV_X1    g594(.A(new_n772), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n780), .B1(new_n781), .B2(new_n608), .ZN(new_n782));
  NAND3_X1  g596(.A1(new_n763), .A2(new_n585), .A3(new_n767), .ZN(new_n783));
  INV_X1    g597(.A(KEYINPUT118), .ZN(new_n784));
  NOR2_X1   g598(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n785));
  XOR2_X1   g599(.A(new_n783), .B(new_n785), .Z(new_n786));
  AND2_X1   g600(.A1(new_n784), .A2(KEYINPUT48), .ZN(new_n787));
  OAI21_X1  g601(.A(new_n782), .B1(new_n786), .B2(new_n787), .ZN(new_n788));
  AOI21_X1  g602(.A(new_n788), .B1(new_n777), .B2(new_n778), .ZN(new_n789));
  AOI21_X1  g603(.A(new_n775), .B1(new_n761), .B2(new_n765), .ZN(new_n790));
  NAND4_X1  g604(.A1(new_n790), .A2(KEYINPUT117), .A3(KEYINPUT51), .A4(new_n768), .ZN(new_n791));
  AND3_X1   g605(.A1(new_n779), .A2(new_n789), .A3(new_n791), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n636), .A2(new_n428), .A3(new_n622), .ZN(new_n793));
  AOI21_X1  g607(.A(KEYINPUT104), .B1(new_n793), .B2(new_n687), .ZN(new_n794));
  NOR3_X1   g608(.A1(new_n690), .A2(new_n691), .A3(new_n689), .ZN(new_n795));
  OAI21_X1  g609(.A(new_n683), .B1(new_n794), .B2(new_n795), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n708), .A2(new_n680), .ZN(new_n797));
  NOR2_X1   g611(.A1(new_n796), .A2(new_n797), .ZN(new_n798));
  INV_X1    g612(.A(new_n726), .ZN(new_n799));
  AND2_X1   g613(.A1(new_n721), .A2(new_n722), .ZN(new_n800));
  NOR2_X1   g614(.A1(new_n721), .A2(new_n718), .ZN(new_n801));
  OAI21_X1  g615(.A(new_n799), .B1(new_n800), .B2(new_n801), .ZN(new_n802));
  INV_X1    g616(.A(KEYINPUT110), .ZN(new_n803));
  NOR2_X1   g617(.A1(new_n375), .A2(new_n419), .ZN(new_n804));
  NAND4_X1  g618(.A1(new_n717), .A2(new_n803), .A3(new_n804), .A4(new_n637), .ZN(new_n805));
  NAND4_X1  g619(.A1(new_n307), .A2(new_n804), .A3(new_n484), .A4(new_n308), .ZN(new_n806));
  OAI21_X1  g620(.A(KEYINPUT110), .B1(new_n806), .B2(new_n638), .ZN(new_n807));
  NAND4_X1  g621(.A1(new_n686), .A2(new_n805), .A3(new_n807), .A4(new_n483), .ZN(new_n808));
  OAI21_X1  g622(.A(new_n486), .B1(new_n585), .B2(new_n624), .ZN(new_n809));
  NAND2_X1  g623(.A1(new_n613), .A2(new_n607), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n598), .A2(new_n810), .ZN(new_n811));
  NAND4_X1  g625(.A1(new_n710), .A2(new_n483), .A3(new_n664), .A4(new_n717), .ZN(new_n812));
  NAND4_X1  g626(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n813));
  NOR2_X1   g627(.A1(new_n802), .A2(new_n813), .ZN(new_n814));
  INV_X1    g628(.A(KEYINPUT111), .ZN(new_n815));
  NAND3_X1  g629(.A1(new_n798), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  AOI21_X1  g630(.A(new_n726), .B1(new_n720), .B2(new_n723), .ZN(new_n817));
  NAND2_X1  g631(.A1(new_n636), .A2(new_n749), .ZN(new_n818));
  AOI21_X1  g632(.A(new_n485), .B1(new_n818), .B2(new_n623), .ZN(new_n819));
  INV_X1    g633(.A(new_n810), .ZN(new_n820));
  NOR3_X1   g634(.A1(new_n594), .A2(new_n597), .A3(new_n820), .ZN(new_n821));
  NAND4_X1  g635(.A1(new_n593), .A2(new_n664), .A3(new_n622), .A4(new_n703), .ZN(new_n822));
  NOR3_X1   g636(.A1(new_n822), .A2(new_n631), .A3(new_n738), .ZN(new_n823));
  NOR3_X1   g637(.A1(new_n819), .A2(new_n821), .A3(new_n823), .ZN(new_n824));
  NAND3_X1  g638(.A1(new_n817), .A2(new_n824), .A3(new_n808), .ZN(new_n825));
  NAND4_X1  g639(.A1(new_n693), .A2(new_n680), .A3(new_n683), .A4(new_n708), .ZN(new_n826));
  OAI21_X1  g640(.A(KEYINPUT111), .B1(new_n825), .B2(new_n826), .ZN(new_n827));
  NAND4_X1  g641(.A1(new_n520), .A2(KEYINPUT113), .A3(new_n621), .A4(new_n637), .ZN(new_n828));
  OAI211_X1 g642(.A(new_n621), .B(new_n637), .C1(new_n515), .C2(new_n518), .ZN(new_n829));
  INV_X1    g643(.A(KEYINPUT113), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n829), .A2(new_n830), .ZN(new_n831));
  AND3_X1   g645(.A1(new_n828), .A2(new_n483), .A3(new_n831), .ZN(new_n832));
  AOI21_X1  g646(.A(new_n697), .B1(new_n309), .B2(new_n654), .ZN(new_n833));
  INV_X1    g647(.A(new_n698), .ZN(new_n834));
  OAI211_X1 g648(.A(new_n653), .B(new_n832), .C1(new_n833), .C2(new_n834), .ZN(new_n835));
  NAND4_X1  g649(.A1(new_n835), .A2(new_n640), .A3(new_n665), .A4(new_n711), .ZN(new_n836));
  INV_X1    g650(.A(KEYINPUT52), .ZN(new_n837));
  NAND2_X1  g651(.A1(new_n836), .A2(new_n837), .ZN(new_n838));
  OAI211_X1 g652(.A(new_n686), .B(new_n632), .C1(new_n639), .C2(new_n664), .ZN(new_n839));
  NAND4_X1  g653(.A1(new_n839), .A2(KEYINPUT52), .A3(new_n711), .A4(new_n835), .ZN(new_n840));
  NAND2_X1  g654(.A1(new_n838), .A2(new_n840), .ZN(new_n841));
  NAND3_X1  g655(.A1(new_n816), .A2(new_n827), .A3(new_n841), .ZN(new_n842));
  INV_X1    g656(.A(KEYINPUT53), .ZN(new_n843));
  NAND2_X1  g657(.A1(new_n842), .A2(new_n843), .ZN(new_n844));
  XOR2_X1   g658(.A(KEYINPUT114), .B(KEYINPUT54), .Z(new_n845));
  INV_X1    g659(.A(new_n845), .ZN(new_n846));
  NAND2_X1  g660(.A1(new_n841), .A2(KEYINPUT53), .ZN(new_n847));
  AND3_X1   g661(.A1(new_n678), .A2(new_n585), .A3(new_n679), .ZN(new_n848));
  AOI22_X1  g662(.A1(new_n848), .A2(new_n614), .B1(new_n692), .B2(new_n688), .ZN(new_n849));
  INV_X1    g663(.A(new_n797), .ZN(new_n850));
  AND4_X1   g664(.A1(new_n808), .A2(new_n809), .A3(new_n811), .A4(new_n812), .ZN(new_n851));
  NAND4_X1  g665(.A1(new_n849), .A2(new_n850), .A3(new_n851), .A4(new_n817), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n847), .A2(new_n852), .ZN(new_n853));
  INV_X1    g667(.A(new_n853), .ZN(new_n854));
  AND4_X1   g668(.A1(KEYINPUT115), .A2(new_n844), .A3(new_n846), .A4(new_n854), .ZN(new_n855));
  AOI21_X1  g669(.A(new_n853), .B1(new_n842), .B2(new_n843), .ZN(new_n856));
  AOI21_X1  g670(.A(KEYINPUT115), .B1(new_n856), .B2(new_n846), .ZN(new_n857));
  NOR2_X1   g671(.A1(new_n855), .A2(new_n857), .ZN(new_n858));
  AOI21_X1  g672(.A(KEYINPUT53), .B1(new_n841), .B2(KEYINPUT112), .ZN(new_n859));
  NAND2_X1  g673(.A1(new_n842), .A2(new_n859), .ZN(new_n860));
  NAND2_X1  g674(.A1(new_n841), .A2(KEYINPUT112), .ZN(new_n861));
  NAND2_X1  g675(.A1(new_n861), .A2(new_n843), .ZN(new_n862));
  NAND4_X1  g676(.A1(new_n862), .A2(new_n841), .A3(new_n816), .A4(new_n827), .ZN(new_n863));
  NAND2_X1  g677(.A1(new_n860), .A2(new_n863), .ZN(new_n864));
  NAND2_X1  g678(.A1(new_n864), .A2(KEYINPUT54), .ZN(new_n865));
  NAND3_X1  g679(.A1(new_n792), .A2(new_n858), .A3(new_n865), .ZN(new_n866));
  NOR2_X1   g680(.A1(new_n764), .A2(new_n691), .ZN(new_n867));
  OAI22_X1  g681(.A1(new_n866), .A2(new_n867), .B1(G952), .B2(G953), .ZN(new_n868));
  NOR2_X1   g682(.A1(new_n589), .A2(new_n716), .ZN(new_n869));
  XNOR2_X1  g683(.A(new_n869), .B(KEYINPUT108), .ZN(new_n870));
  AND3_X1   g684(.A1(new_n870), .A2(new_n612), .A3(new_n606), .ZN(new_n871));
  XNOR2_X1  g685(.A(new_n676), .B(KEYINPUT49), .ZN(new_n872));
  NAND4_X1  g686(.A1(new_n871), .A2(new_n771), .A3(new_n660), .A4(new_n872), .ZN(new_n873));
  XNOR2_X1  g687(.A(new_n873), .B(KEYINPUT109), .ZN(new_n874));
  NAND2_X1  g688(.A1(new_n868), .A2(new_n874), .ZN(G75));
  XOR2_X1   g689(.A(new_n300), .B(new_n302), .Z(new_n876));
  XNOR2_X1  g690(.A(new_n876), .B(KEYINPUT55), .ZN(new_n877));
  INV_X1    g691(.A(new_n877), .ZN(new_n878));
  INV_X1    g692(.A(KEYINPUT56), .ZN(new_n879));
  NAND2_X1  g693(.A1(new_n844), .A2(new_n854), .ZN(new_n880));
  NAND2_X1  g694(.A1(new_n880), .A2(G902), .ZN(new_n881));
  INV_X1    g695(.A(G210), .ZN(new_n882));
  OAI21_X1  g696(.A(new_n879), .B1(new_n881), .B2(new_n882), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n883), .A2(KEYINPUT119), .ZN(new_n884));
  INV_X1    g698(.A(KEYINPUT119), .ZN(new_n885));
  OAI211_X1 g699(.A(new_n885), .B(new_n879), .C1(new_n881), .C2(new_n882), .ZN(new_n886));
  AOI21_X1  g700(.A(new_n878), .B1(new_n884), .B2(new_n886), .ZN(new_n887));
  NOR2_X1   g701(.A1(new_n327), .A2(G952), .ZN(new_n888));
  AOI21_X1  g702(.A(new_n877), .B1(new_n883), .B2(KEYINPUT119), .ZN(new_n889));
  NOR3_X1   g703(.A1(new_n887), .A2(new_n888), .A3(new_n889), .ZN(G51));
  XOR2_X1   g704(.A(new_n731), .B(KEYINPUT57), .Z(new_n891));
  NAND3_X1  g705(.A1(new_n844), .A2(new_n846), .A3(new_n854), .ZN(new_n892));
  INV_X1    g706(.A(new_n892), .ZN(new_n893));
  NOR2_X1   g707(.A1(new_n856), .A2(new_n846), .ZN(new_n894));
  OAI21_X1  g708(.A(new_n891), .B1(new_n893), .B2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n895), .A2(new_n668), .ZN(new_n896));
  OR2_X1    g710(.A1(new_n881), .A2(new_n730), .ZN(new_n897));
  AOI21_X1  g711(.A(new_n888), .B1(new_n896), .B2(new_n897), .ZN(G54));
  NAND4_X1  g712(.A1(new_n880), .A2(KEYINPUT58), .A3(G475), .A4(G902), .ZN(new_n899));
  INV_X1    g713(.A(new_n370), .ZN(new_n900));
  AND2_X1   g714(.A1(new_n899), .A2(new_n900), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n899), .A2(new_n900), .ZN(new_n902));
  NOR3_X1   g716(.A1(new_n901), .A2(new_n902), .A3(new_n888), .ZN(G60));
  NAND2_X1  g717(.A1(G478), .A2(G902), .ZN(new_n904));
  XOR2_X1   g718(.A(new_n904), .B(KEYINPUT59), .Z(new_n905));
  NAND2_X1  g719(.A1(new_n880), .A2(new_n845), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n905), .B1(new_n906), .B2(new_n892), .ZN(new_n907));
  AOI21_X1  g721(.A(new_n888), .B1(new_n907), .B2(new_n602), .ZN(new_n908));
  AOI21_X1  g722(.A(new_n905), .B1(new_n858), .B2(new_n865), .ZN(new_n909));
  OAI211_X1 g723(.A(KEYINPUT120), .B(new_n908), .C1(new_n909), .C2(new_n602), .ZN(new_n910));
  INV_X1    g724(.A(KEYINPUT120), .ZN(new_n911));
  INV_X1    g725(.A(KEYINPUT115), .ZN(new_n912));
  NAND2_X1  g726(.A1(new_n892), .A2(new_n912), .ZN(new_n913));
  NAND3_X1  g727(.A1(new_n856), .A2(KEYINPUT115), .A3(new_n846), .ZN(new_n914));
  NAND3_X1  g728(.A1(new_n913), .A2(new_n865), .A3(new_n914), .ZN(new_n915));
  INV_X1    g729(.A(new_n905), .ZN(new_n916));
  AOI21_X1  g730(.A(new_n602), .B1(new_n915), .B2(new_n916), .ZN(new_n917));
  OAI211_X1 g731(.A(new_n602), .B(new_n916), .C1(new_n893), .C2(new_n894), .ZN(new_n918));
  INV_X1    g732(.A(new_n888), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n918), .A2(new_n919), .ZN(new_n920));
  OAI21_X1  g734(.A(new_n911), .B1(new_n917), .B2(new_n920), .ZN(new_n921));
  NAND2_X1  g735(.A1(new_n910), .A2(new_n921), .ZN(G63));
  NAND2_X1  g736(.A1(G217), .A2(G902), .ZN(new_n923));
  XNOR2_X1  g737(.A(new_n923), .B(KEYINPUT121), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  NAND2_X1  g739(.A1(new_n880), .A2(new_n925), .ZN(new_n926));
  INV_X1    g740(.A(new_n521), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n888), .B1(new_n926), .B2(new_n927), .ZN(new_n928));
  NAND3_X1  g742(.A1(new_n880), .A2(new_n620), .A3(new_n925), .ZN(new_n929));
  AOI22_X1  g743(.A1(new_n928), .A2(new_n929), .B1(KEYINPUT122), .B2(KEYINPUT61), .ZN(new_n930));
  INV_X1    g744(.A(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT61), .ZN(new_n932));
  NAND2_X1  g746(.A1(new_n931), .A2(new_n932), .ZN(new_n933));
  NAND2_X1  g747(.A1(new_n930), .A2(new_n933), .ZN(new_n934));
  NAND4_X1  g748(.A1(new_n928), .A2(new_n931), .A3(new_n932), .A4(new_n929), .ZN(new_n935));
  AND2_X1   g749(.A1(new_n934), .A2(new_n935), .ZN(G66));
  NAND2_X1  g750(.A1(new_n809), .A2(new_n811), .ZN(new_n937));
  NOR2_X1   g751(.A1(new_n826), .A2(new_n937), .ZN(new_n938));
  NOR2_X1   g752(.A1(new_n938), .A2(new_n423), .ZN(new_n939));
  XNOR2_X1  g753(.A(new_n939), .B(KEYINPUT123), .ZN(new_n940));
  AOI21_X1  g754(.A(new_n220), .B1(new_n425), .B2(G224), .ZN(new_n941));
  NOR2_X1   g755(.A1(new_n940), .A2(new_n941), .ZN(new_n942));
  OAI21_X1  g756(.A(new_n300), .B1(G898), .B2(new_n327), .ZN(new_n943));
  XOR2_X1   g757(.A(new_n942), .B(new_n943), .Z(G69));
  NAND2_X1  g758(.A1(new_n557), .A2(new_n558), .ZN(new_n945));
  XNOR2_X1  g759(.A(new_n945), .B(new_n358), .ZN(new_n946));
  XNOR2_X1  g760(.A(KEYINPUT124), .B(KEYINPUT125), .ZN(new_n947));
  XOR2_X1   g761(.A(new_n946), .B(new_n947), .Z(new_n948));
  INV_X1    g762(.A(new_n948), .ZN(new_n949));
  NAND3_X1  g763(.A1(new_n737), .A2(new_n585), .A3(new_n699), .ZN(new_n950));
  NAND3_X1  g764(.A1(new_n745), .A2(new_n950), .A3(new_n754), .ZN(new_n951));
  INV_X1    g765(.A(KEYINPUT126), .ZN(new_n952));
  AND2_X1   g766(.A1(new_n839), .A2(new_n711), .ZN(new_n953));
  NAND2_X1  g767(.A1(new_n953), .A2(new_n817), .ZN(new_n954));
  OR3_X1    g768(.A1(new_n951), .A2(new_n952), .A3(new_n954), .ZN(new_n955));
  OAI21_X1  g769(.A(new_n952), .B1(new_n951), .B2(new_n954), .ZN(new_n956));
  NAND2_X1  g770(.A1(new_n955), .A2(new_n956), .ZN(new_n957));
  AOI21_X1  g771(.A(new_n949), .B1(new_n957), .B2(new_n327), .ZN(new_n958));
  INV_X1    g772(.A(G900), .ZN(new_n959));
  NAND2_X1  g773(.A1(new_n423), .A2(new_n959), .ZN(new_n960));
  AND2_X1   g774(.A1(new_n745), .A2(new_n754), .ZN(new_n961));
  OR4_X1    g775(.A1(new_n818), .A2(new_n647), .A3(new_n738), .A4(new_n820), .ZN(new_n962));
  AND3_X1   g776(.A1(new_n662), .A2(KEYINPUT62), .A3(new_n953), .ZN(new_n963));
  AOI21_X1  g777(.A(KEYINPUT62), .B1(new_n662), .B2(new_n953), .ZN(new_n964));
  OAI211_X1 g778(.A(new_n961), .B(new_n962), .C1(new_n963), .C2(new_n964), .ZN(new_n965));
  NOR2_X1   g779(.A1(new_n948), .A2(new_n423), .ZN(new_n966));
  AOI22_X1  g780(.A1(new_n958), .A2(new_n960), .B1(new_n965), .B2(new_n966), .ZN(new_n967));
  INV_X1    g781(.A(G227), .ZN(new_n968));
  OAI21_X1  g782(.A(new_n423), .B1(new_n968), .B2(new_n959), .ZN(new_n969));
  XOR2_X1   g783(.A(new_n967), .B(new_n969), .Z(G72));
  NAND3_X1  g784(.A1(new_n955), .A2(new_n956), .A3(new_n938), .ZN(new_n971));
  NAND2_X1  g785(.A1(G472), .A2(G902), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n972), .B(KEYINPUT63), .Z(new_n973));
  AOI21_X1  g787(.A(new_n579), .B1(new_n971), .B2(new_n973), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n888), .B1(new_n974), .B2(new_n565), .ZN(new_n975));
  INV_X1    g789(.A(new_n938), .ZN(new_n976));
  OAI21_X1  g790(.A(new_n973), .B1(new_n965), .B2(new_n976), .ZN(new_n977));
  NAND3_X1  g791(.A1(new_n977), .A2(new_n551), .A3(new_n579), .ZN(new_n978));
  NAND2_X1  g792(.A1(new_n580), .A2(new_n563), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n864), .A2(new_n973), .A3(new_n979), .ZN(new_n980));
  NAND3_X1  g794(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(new_n981));
  INV_X1    g795(.A(KEYINPUT127), .ZN(new_n982));
  NAND2_X1  g796(.A1(new_n981), .A2(new_n982), .ZN(new_n983));
  NAND4_X1  g797(.A1(new_n975), .A2(KEYINPUT127), .A3(new_n978), .A4(new_n980), .ZN(new_n984));
  NAND2_X1  g798(.A1(new_n983), .A2(new_n984), .ZN(G57));
endmodule


