//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 1 0 1 0 0 1 0 0 0 0 1 0 1 1 0 1 0 1 0 0 0 0 0 1 1 0 1 0 0 1 1 0 0 1 1 1 1 1 0 0 0 1 1 1 0 0 1 1 0 1 0 1 1 1 1 0 0 0 1 0 0 0 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:19:35 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n674, new_n675, new_n676, new_n677, new_n678,
    new_n679, new_n680, new_n682, new_n683, new_n684, new_n686, new_n687,
    new_n688, new_n689, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n719, new_n720, new_n721, new_n722, new_n724, new_n725,
    new_n726, new_n728, new_n729, new_n730, new_n731, new_n732, new_n733,
    new_n734, new_n736, new_n737, new_n738, new_n740, new_n741, new_n742,
    new_n744, new_n745, new_n746, new_n747, new_n748, new_n749, new_n750,
    new_n751, new_n752, new_n753, new_n755, new_n757, new_n758, new_n759,
    new_n760, new_n761, new_n762, new_n763, new_n764, new_n765, new_n766,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n777, new_n778, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n786, new_n787, new_n788, new_n789,
    new_n790, new_n791, new_n792, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n810, new_n811, new_n812,
    new_n813, new_n814, new_n815, new_n816, new_n817, new_n818, new_n819,
    new_n820, new_n821, new_n822, new_n823, new_n824, new_n825, new_n826,
    new_n827, new_n828, new_n829, new_n830, new_n831, new_n832, new_n833,
    new_n834, new_n835, new_n837, new_n838, new_n840, new_n841, new_n843,
    new_n844, new_n845, new_n846, new_n847, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n854, new_n855, new_n856, new_n857, new_n858,
    new_n859, new_n860, new_n861, new_n862, new_n863, new_n864, new_n865,
    new_n866, new_n867, new_n868, new_n869, new_n870, new_n871, new_n872,
    new_n873, new_n874, new_n875, new_n876, new_n877, new_n878, new_n879,
    new_n881, new_n882, new_n883, new_n884, new_n885, new_n886, new_n887,
    new_n888, new_n889, new_n890, new_n891, new_n892, new_n893, new_n894,
    new_n895, new_n896, new_n897, new_n898, new_n899, new_n900, new_n901,
    new_n902, new_n903, new_n904, new_n905, new_n907, new_n908, new_n909,
    new_n910, new_n912, new_n913, new_n915, new_n916, new_n917, new_n918,
    new_n920, new_n921, new_n923, new_n924, new_n925, new_n926, new_n927,
    new_n929, new_n930, new_n931, new_n933, new_n934, new_n935, new_n936,
    new_n937, new_n938, new_n939, new_n940, new_n941, new_n943, new_n944,
    new_n945, new_n946, new_n948, new_n949, new_n950, new_n951, new_n952,
    new_n953, new_n954, new_n956, new_n957;
  XOR2_X1   g000(.A(G15gat), .B(G43gat), .Z(new_n202));
  XNOR2_X1  g001(.A(G71gat), .B(G99gat), .ZN(new_n203));
  XNOR2_X1  g002(.A(new_n202), .B(new_n203), .ZN(new_n204));
  INV_X1    g003(.A(new_n204), .ZN(new_n205));
  NAND2_X1  g004(.A1(G183gat), .A2(G190gat), .ZN(new_n206));
  INV_X1    g005(.A(G169gat), .ZN(new_n207));
  INV_X1    g006(.A(G176gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(new_n208), .ZN(new_n209));
  NOR2_X1   g008(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n210));
  XNOR2_X1  g009(.A(new_n210), .B(KEYINPUT68), .ZN(new_n211));
  NAND2_X1  g010(.A1(G169gat), .A2(G176gat), .ZN(new_n212));
  NAND2_X1  g011(.A1(new_n209), .A2(KEYINPUT26), .ZN(new_n213));
  NAND3_X1  g012(.A1(new_n211), .A2(new_n212), .A3(new_n213), .ZN(new_n214));
  XNOR2_X1  g013(.A(KEYINPUT27), .B(G183gat), .ZN(new_n215));
  INV_X1    g014(.A(G190gat), .ZN(new_n216));
  NAND2_X1  g015(.A1(new_n215), .A2(new_n216), .ZN(new_n217));
  INV_X1    g016(.A(KEYINPUT28), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(new_n219), .B(KEYINPUT67), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n217), .A2(new_n218), .ZN(new_n221));
  XNOR2_X1  g020(.A(new_n221), .B(KEYINPUT66), .ZN(new_n222));
  OAI211_X1 g021(.A(new_n206), .B(new_n214), .C1(new_n220), .C2(new_n222), .ZN(new_n223));
  NOR2_X1   g022(.A1(G169gat), .A2(G176gat), .ZN(new_n224));
  NAND2_X1  g023(.A1(new_n224), .A2(KEYINPUT23), .ZN(new_n225));
  NAND2_X1  g024(.A1(new_n225), .A2(new_n212), .ZN(new_n226));
  XOR2_X1   g025(.A(new_n226), .B(KEYINPUT65), .Z(new_n227));
  INV_X1    g026(.A(KEYINPUT23), .ZN(new_n228));
  NAND2_X1  g027(.A1(new_n209), .A2(new_n228), .ZN(new_n229));
  NOR2_X1   g028(.A1(new_n206), .A2(KEYINPUT24), .ZN(new_n230));
  XOR2_X1   g029(.A(G183gat), .B(G190gat), .Z(new_n231));
  AOI21_X1  g030(.A(new_n230), .B1(new_n231), .B2(KEYINPUT24), .ZN(new_n232));
  NAND4_X1  g031(.A1(new_n227), .A2(KEYINPUT25), .A3(new_n229), .A4(new_n232), .ZN(new_n233));
  INV_X1    g032(.A(KEYINPUT25), .ZN(new_n234));
  NAND3_X1  g033(.A1(new_n229), .A2(new_n212), .A3(new_n225), .ZN(new_n235));
  NAND2_X1  g034(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n236), .A2(new_n232), .ZN(new_n237));
  NOR2_X1   g036(.A1(new_n235), .A2(KEYINPUT64), .ZN(new_n238));
  OAI21_X1  g037(.A(new_n234), .B1(new_n237), .B2(new_n238), .ZN(new_n239));
  NAND2_X1  g038(.A1(new_n233), .A2(new_n239), .ZN(new_n240));
  NAND2_X1  g039(.A1(new_n223), .A2(new_n240), .ZN(new_n241));
  XNOR2_X1  g040(.A(G127gat), .B(G134gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(G113gat), .A2(G120gat), .ZN(new_n243));
  INV_X1    g042(.A(G113gat), .ZN(new_n244));
  INV_X1    g043(.A(G120gat), .ZN(new_n245));
  AOI21_X1  g044(.A(KEYINPUT1), .B1(new_n244), .B2(new_n245), .ZN(new_n246));
  AOI21_X1  g045(.A(new_n242), .B1(new_n243), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT69), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n248), .A2(G120gat), .ZN(new_n249));
  NOR2_X1   g048(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n250));
  OAI21_X1  g049(.A(G113gat), .B1(new_n249), .B2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(KEYINPUT70), .ZN(new_n252));
  NAND4_X1  g051(.A1(new_n251), .A2(new_n252), .A3(new_n246), .A4(new_n242), .ZN(new_n253));
  NAND2_X1  g052(.A1(new_n244), .A2(new_n245), .ZN(new_n254));
  INV_X1    g053(.A(G134gat), .ZN(new_n255));
  NAND2_X1  g054(.A1(new_n255), .A2(G127gat), .ZN(new_n256));
  INV_X1    g055(.A(G127gat), .ZN(new_n257));
  NAND2_X1  g056(.A1(new_n257), .A2(G134gat), .ZN(new_n258));
  INV_X1    g057(.A(KEYINPUT1), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n254), .A2(new_n256), .A3(new_n258), .A4(new_n259), .ZN(new_n260));
  NAND2_X1  g059(.A1(new_n245), .A2(KEYINPUT69), .ZN(new_n261));
  NAND2_X1  g060(.A1(new_n248), .A2(G120gat), .ZN(new_n262));
  AOI21_X1  g061(.A(new_n244), .B1(new_n261), .B2(new_n262), .ZN(new_n263));
  OAI21_X1  g062(.A(KEYINPUT70), .B1(new_n260), .B2(new_n263), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n247), .B1(new_n253), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n241), .A2(new_n265), .ZN(new_n266));
  INV_X1    g065(.A(G227gat), .ZN(new_n267));
  INV_X1    g066(.A(G233gat), .ZN(new_n268));
  NOR2_X1   g067(.A1(new_n267), .A2(new_n268), .ZN(new_n269));
  NAND2_X1  g068(.A1(new_n253), .A2(new_n264), .ZN(new_n270));
  INV_X1    g069(.A(new_n247), .ZN(new_n271));
  NAND2_X1  g070(.A1(new_n270), .A2(new_n271), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n223), .A2(new_n272), .A3(new_n240), .ZN(new_n273));
  NAND3_X1  g072(.A1(new_n266), .A2(new_n269), .A3(new_n273), .ZN(new_n274));
  INV_X1    g073(.A(KEYINPUT33), .ZN(new_n275));
  AOI21_X1  g074(.A(new_n205), .B1(new_n274), .B2(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(KEYINPUT34), .ZN(new_n277));
  NAND2_X1  g076(.A1(new_n266), .A2(new_n273), .ZN(new_n278));
  INV_X1    g077(.A(new_n269), .ZN(new_n279));
  AOI21_X1  g078(.A(new_n277), .B1(new_n278), .B2(new_n279), .ZN(new_n280));
  AOI211_X1 g079(.A(KEYINPUT34), .B(new_n269), .C1(new_n266), .C2(new_n273), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n276), .A2(new_n280), .A3(new_n281), .ZN(new_n282));
  INV_X1    g081(.A(new_n282), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n274), .A2(KEYINPUT32), .ZN(new_n284));
  INV_X1    g083(.A(new_n284), .ZN(new_n285));
  OAI21_X1  g084(.A(new_n276), .B1(new_n280), .B2(new_n281), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n283), .A2(new_n285), .A3(new_n286), .ZN(new_n287));
  INV_X1    g086(.A(new_n286), .ZN(new_n288));
  OAI21_X1  g087(.A(new_n284), .B1(new_n288), .B2(new_n282), .ZN(new_n289));
  NAND2_X1  g088(.A1(new_n287), .A2(new_n289), .ZN(new_n290));
  NAND2_X1  g089(.A1(G228gat), .A2(G233gat), .ZN(new_n291));
  INV_X1    g090(.A(new_n291), .ZN(new_n292));
  AND2_X1   g091(.A1(G141gat), .A2(G148gat), .ZN(new_n293));
  NOR2_X1   g092(.A1(G141gat), .A2(G148gat), .ZN(new_n294));
  NOR2_X1   g093(.A1(new_n293), .A2(new_n294), .ZN(new_n295));
  NAND2_X1  g094(.A1(G155gat), .A2(G162gat), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT2), .ZN(new_n297));
  NAND2_X1  g096(.A1(new_n295), .A2(new_n297), .ZN(new_n298));
  INV_X1    g097(.A(new_n296), .ZN(new_n299));
  NOR2_X1   g098(.A1(G155gat), .A2(G162gat), .ZN(new_n300));
  OAI21_X1  g099(.A(KEYINPUT74), .B1(new_n299), .B2(new_n300), .ZN(new_n301));
  INV_X1    g100(.A(new_n300), .ZN(new_n302));
  INV_X1    g101(.A(KEYINPUT74), .ZN(new_n303));
  NAND3_X1  g102(.A1(new_n302), .A2(new_n303), .A3(new_n296), .ZN(new_n304));
  NAND3_X1  g103(.A1(new_n298), .A2(new_n301), .A3(new_n304), .ZN(new_n305));
  NOR2_X1   g104(.A1(new_n299), .A2(new_n300), .ZN(new_n306));
  NAND4_X1  g105(.A1(new_n306), .A2(new_n295), .A3(new_n303), .A4(new_n297), .ZN(new_n307));
  NAND2_X1  g106(.A1(new_n305), .A2(new_n307), .ZN(new_n308));
  XNOR2_X1  g107(.A(G197gat), .B(G204gat), .ZN(new_n309));
  INV_X1    g108(.A(G211gat), .ZN(new_n310));
  INV_X1    g109(.A(G218gat), .ZN(new_n311));
  NOR2_X1   g110(.A1(new_n310), .A2(new_n311), .ZN(new_n312));
  OAI21_X1  g111(.A(new_n309), .B1(KEYINPUT22), .B2(new_n312), .ZN(new_n313));
  XOR2_X1   g112(.A(G211gat), .B(G218gat), .Z(new_n314));
  XOR2_X1   g113(.A(new_n313), .B(new_n314), .Z(new_n315));
  OR2_X1    g114(.A1(new_n315), .A2(KEYINPUT29), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT3), .ZN(new_n317));
  AOI21_X1  g116(.A(new_n308), .B1(new_n316), .B2(new_n317), .ZN(new_n318));
  INV_X1    g117(.A(KEYINPUT71), .ZN(new_n319));
  NAND2_X1  g118(.A1(new_n315), .A2(new_n319), .ZN(new_n320));
  NAND3_X1  g119(.A1(new_n313), .A2(KEYINPUT71), .A3(new_n314), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n320), .A2(new_n321), .ZN(new_n322));
  NAND2_X1  g121(.A1(new_n308), .A2(new_n317), .ZN(new_n323));
  INV_X1    g122(.A(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n322), .B1(new_n324), .B2(KEYINPUT29), .ZN(new_n325));
  AOI21_X1  g124(.A(new_n318), .B1(new_n325), .B2(KEYINPUT85), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT85), .ZN(new_n327));
  OAI211_X1 g126(.A(new_n322), .B(new_n327), .C1(KEYINPUT29), .C2(new_n324), .ZN(new_n328));
  AOI21_X1  g127(.A(new_n292), .B1(new_n326), .B2(new_n328), .ZN(new_n329));
  OAI21_X1  g128(.A(new_n317), .B1(new_n322), .B2(KEYINPUT29), .ZN(new_n330));
  INV_X1    g129(.A(new_n308), .ZN(new_n331));
  NAND2_X1  g130(.A1(new_n330), .A2(new_n331), .ZN(new_n332));
  AND3_X1   g131(.A1(new_n332), .A2(new_n292), .A3(new_n325), .ZN(new_n333));
  OAI21_X1  g132(.A(G22gat), .B1(new_n329), .B2(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n325), .A2(KEYINPUT85), .ZN(new_n335));
  INV_X1    g134(.A(new_n318), .ZN(new_n336));
  NAND3_X1  g135(.A1(new_n335), .A2(new_n328), .A3(new_n336), .ZN(new_n337));
  NAND2_X1  g136(.A1(new_n337), .A2(new_n291), .ZN(new_n338));
  INV_X1    g137(.A(G22gat), .ZN(new_n339));
  AND2_X1   g138(.A1(new_n325), .A2(new_n292), .ZN(new_n340));
  NAND2_X1  g139(.A1(new_n340), .A2(new_n332), .ZN(new_n341));
  NAND3_X1  g140(.A1(new_n338), .A2(new_n339), .A3(new_n341), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n334), .A2(new_n342), .ZN(new_n343));
  INV_X1    g142(.A(KEYINPUT86), .ZN(new_n344));
  AOI22_X1  g143(.A1(new_n337), .A2(new_n291), .B1(new_n340), .B2(new_n332), .ZN(new_n345));
  AOI21_X1  g144(.A(new_n344), .B1(new_n345), .B2(new_n339), .ZN(new_n346));
  XOR2_X1   g145(.A(G78gat), .B(G106gat), .Z(new_n347));
  XNOR2_X1  g146(.A(KEYINPUT84), .B(G50gat), .ZN(new_n348));
  XNOR2_X1  g147(.A(new_n347), .B(new_n348), .ZN(new_n349));
  XOR2_X1   g148(.A(KEYINPUT83), .B(KEYINPUT31), .Z(new_n350));
  XOR2_X1   g149(.A(new_n349), .B(new_n350), .Z(new_n351));
  INV_X1    g150(.A(new_n351), .ZN(new_n352));
  OAI21_X1  g151(.A(new_n343), .B1(new_n346), .B2(new_n352), .ZN(new_n353));
  NAND4_X1  g152(.A1(new_n334), .A2(new_n342), .A3(new_n344), .A4(new_n351), .ZN(new_n354));
  NAND2_X1  g153(.A1(new_n353), .A2(new_n354), .ZN(new_n355));
  NOR2_X1   g154(.A1(new_n290), .A2(new_n355), .ZN(new_n356));
  XOR2_X1   g155(.A(G1gat), .B(G29gat), .Z(new_n357));
  XNOR2_X1  g156(.A(new_n357), .B(KEYINPUT81), .ZN(new_n358));
  XOR2_X1   g157(.A(G57gat), .B(G85gat), .Z(new_n359));
  XNOR2_X1  g158(.A(new_n358), .B(new_n359), .ZN(new_n360));
  XNOR2_X1  g159(.A(KEYINPUT80), .B(KEYINPUT0), .ZN(new_n361));
  XOR2_X1   g160(.A(new_n360), .B(new_n361), .Z(new_n362));
  NAND2_X1  g161(.A1(G225gat), .A2(G233gat), .ZN(new_n363));
  INV_X1    g162(.A(new_n363), .ZN(new_n364));
  NAND2_X1  g163(.A1(new_n272), .A2(KEYINPUT76), .ZN(new_n365));
  INV_X1    g164(.A(KEYINPUT76), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n265), .A2(new_n366), .ZN(new_n367));
  NAND4_X1  g166(.A1(new_n365), .A2(KEYINPUT79), .A3(new_n331), .A4(new_n367), .ZN(new_n368));
  NOR2_X1   g167(.A1(new_n265), .A2(new_n366), .ZN(new_n369));
  AOI211_X1 g168(.A(KEYINPUT76), .B(new_n247), .C1(new_n253), .C2(new_n264), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n369), .A2(new_n370), .A3(new_n308), .ZN(new_n371));
  NAND2_X1  g170(.A1(new_n265), .A2(new_n308), .ZN(new_n372));
  INV_X1    g171(.A(KEYINPUT79), .ZN(new_n373));
  NAND2_X1  g172(.A1(new_n372), .A2(new_n373), .ZN(new_n374));
  OAI211_X1 g173(.A(new_n364), .B(new_n368), .C1(new_n371), .C2(new_n374), .ZN(new_n375));
  NAND2_X1  g174(.A1(new_n375), .A2(KEYINPUT5), .ZN(new_n376));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n377), .B1(new_n265), .B2(new_n308), .ZN(new_n378));
  NAND3_X1  g177(.A1(new_n265), .A2(new_n377), .A3(new_n308), .ZN(new_n379));
  AOI21_X1  g178(.A(new_n378), .B1(KEYINPUT77), .B2(new_n379), .ZN(new_n380));
  NAND3_X1  g179(.A1(new_n372), .A2(KEYINPUT77), .A3(KEYINPUT4), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(new_n382), .ZN(new_n383));
  NAND3_X1  g182(.A1(new_n305), .A2(KEYINPUT3), .A3(new_n307), .ZN(new_n384));
  NAND2_X1  g183(.A1(new_n384), .A2(KEYINPUT75), .ZN(new_n385));
  INV_X1    g184(.A(KEYINPUT75), .ZN(new_n386));
  NAND4_X1  g185(.A1(new_n305), .A2(new_n307), .A3(new_n386), .A4(KEYINPUT3), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n385), .A2(new_n387), .ZN(new_n388));
  NAND4_X1  g187(.A1(new_n388), .A2(new_n365), .A3(new_n367), .A4(new_n323), .ZN(new_n389));
  NAND2_X1  g188(.A1(new_n389), .A2(new_n363), .ZN(new_n390));
  OAI21_X1  g189(.A(KEYINPUT78), .B1(new_n383), .B2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n379), .A2(KEYINPUT77), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n372), .A2(KEYINPUT4), .ZN(new_n393));
  NAND2_X1  g192(.A1(new_n392), .A2(new_n393), .ZN(new_n394));
  NAND2_X1  g193(.A1(new_n394), .A2(new_n381), .ZN(new_n395));
  INV_X1    g194(.A(KEYINPUT78), .ZN(new_n396));
  NAND4_X1  g195(.A1(new_n395), .A2(new_n396), .A3(new_n363), .A4(new_n389), .ZN(new_n397));
  AOI21_X1  g196(.A(new_n376), .B1(new_n391), .B2(new_n397), .ZN(new_n398));
  NAND2_X1  g197(.A1(new_n393), .A2(new_n379), .ZN(new_n399));
  INV_X1    g198(.A(new_n399), .ZN(new_n400));
  NOR3_X1   g199(.A1(new_n390), .A2(new_n400), .A3(KEYINPUT5), .ZN(new_n401));
  OAI21_X1  g200(.A(new_n362), .B1(new_n398), .B2(new_n401), .ZN(new_n402));
  INV_X1    g201(.A(KEYINPUT6), .ZN(new_n403));
  AND2_X1   g202(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  NOR3_X1   g203(.A1(new_n398), .A2(new_n362), .A3(new_n401), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n405), .A2(KEYINPUT82), .ZN(new_n406));
  INV_X1    g205(.A(new_n362), .ZN(new_n407));
  INV_X1    g206(.A(new_n401), .ZN(new_n408));
  AND2_X1   g207(.A1(new_n391), .A2(new_n397), .ZN(new_n409));
  OAI211_X1 g208(.A(new_n407), .B(new_n408), .C1(new_n409), .C2(new_n376), .ZN(new_n410));
  INV_X1    g209(.A(KEYINPUT82), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n410), .A2(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n404), .A2(new_n406), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(new_n402), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n414), .A2(KEYINPUT6), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n413), .A2(new_n415), .ZN(new_n416));
  XNOR2_X1  g215(.A(G8gat), .B(G36gat), .ZN(new_n417));
  XNOR2_X1  g216(.A(G64gat), .B(G92gat), .ZN(new_n418));
  XOR2_X1   g217(.A(new_n417), .B(new_n418), .Z(new_n419));
  NAND2_X1  g218(.A1(G226gat), .A2(G233gat), .ZN(new_n420));
  XNOR2_X1  g219(.A(new_n420), .B(KEYINPUT72), .ZN(new_n421));
  INV_X1    g220(.A(new_n421), .ZN(new_n422));
  INV_X1    g221(.A(KEYINPUT29), .ZN(new_n423));
  NAND2_X1  g222(.A1(new_n422), .A2(new_n423), .ZN(new_n424));
  NAND2_X1  g223(.A1(new_n241), .A2(new_n424), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n223), .A2(new_n422), .A3(new_n240), .ZN(new_n426));
  AND3_X1   g225(.A1(new_n425), .A2(new_n322), .A3(new_n426), .ZN(new_n427));
  AOI21_X1  g226(.A(new_n322), .B1(new_n425), .B2(new_n426), .ZN(new_n428));
  OAI21_X1  g227(.A(new_n419), .B1(new_n427), .B2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT30), .ZN(new_n430));
  OR2_X1    g229(.A1(new_n429), .A2(new_n430), .ZN(new_n431));
  INV_X1    g230(.A(KEYINPUT73), .ZN(new_n432));
  OAI21_X1  g231(.A(new_n432), .B1(new_n427), .B2(new_n428), .ZN(new_n433));
  INV_X1    g232(.A(new_n426), .ZN(new_n434));
  AOI22_X1  g233(.A1(new_n223), .A2(new_n240), .B1(new_n423), .B2(new_n422), .ZN(new_n435));
  OAI211_X1 g234(.A(new_n321), .B(new_n320), .C1(new_n434), .C2(new_n435), .ZN(new_n436));
  NAND3_X1  g235(.A1(new_n425), .A2(new_n322), .A3(new_n426), .ZN(new_n437));
  NAND3_X1  g236(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT73), .ZN(new_n438));
  INV_X1    g237(.A(new_n419), .ZN(new_n439));
  NAND3_X1  g238(.A1(new_n433), .A2(new_n438), .A3(new_n439), .ZN(new_n440));
  NAND2_X1  g239(.A1(new_n429), .A2(new_n430), .ZN(new_n441));
  NAND3_X1  g240(.A1(new_n431), .A2(new_n440), .A3(new_n441), .ZN(new_n442));
  INV_X1    g241(.A(new_n442), .ZN(new_n443));
  NAND3_X1  g242(.A1(new_n356), .A2(new_n416), .A3(new_n443), .ZN(new_n444));
  NOR4_X1   g243(.A1(new_n290), .A2(new_n355), .A3(KEYINPUT35), .A4(new_n442), .ZN(new_n445));
  INV_X1    g244(.A(KEYINPUT88), .ZN(new_n446));
  OAI211_X1 g245(.A(new_n403), .B(new_n402), .C1(new_n405), .C2(KEYINPUT82), .ZN(new_n447));
  NOR2_X1   g246(.A1(new_n410), .A2(new_n411), .ZN(new_n448));
  OAI21_X1  g247(.A(new_n446), .B1(new_n447), .B2(new_n448), .ZN(new_n449));
  NAND4_X1  g248(.A1(new_n404), .A2(new_n412), .A3(KEYINPUT88), .A4(new_n406), .ZN(new_n450));
  NAND3_X1  g249(.A1(new_n449), .A2(new_n415), .A3(new_n450), .ZN(new_n451));
  AOI22_X1  g250(.A1(KEYINPUT35), .A2(new_n444), .B1(new_n445), .B2(new_n451), .ZN(new_n452));
  INV_X1    g251(.A(KEYINPUT37), .ZN(new_n453));
  OAI21_X1  g252(.A(new_n453), .B1(new_n427), .B2(new_n428), .ZN(new_n454));
  NAND3_X1  g253(.A1(new_n436), .A2(new_n437), .A3(KEYINPUT37), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n419), .A2(KEYINPUT38), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n454), .A2(new_n455), .A3(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n457), .A2(new_n429), .ZN(new_n458));
  AOI21_X1  g257(.A(new_n458), .B1(KEYINPUT6), .B2(new_n414), .ZN(new_n459));
  NAND3_X1  g258(.A1(new_n449), .A2(new_n450), .A3(new_n459), .ZN(new_n460));
  NAND2_X1  g259(.A1(new_n460), .A2(KEYINPUT89), .ZN(new_n461));
  INV_X1    g260(.A(KEYINPUT89), .ZN(new_n462));
  NAND4_X1  g261(.A1(new_n449), .A2(new_n459), .A3(new_n462), .A4(new_n450), .ZN(new_n463));
  NAND3_X1  g262(.A1(new_n433), .A2(new_n438), .A3(KEYINPUT37), .ZN(new_n464));
  NAND2_X1  g263(.A1(new_n464), .A2(new_n439), .ZN(new_n465));
  INV_X1    g264(.A(KEYINPUT90), .ZN(new_n466));
  NAND2_X1  g265(.A1(new_n465), .A2(new_n466), .ZN(new_n467));
  NAND3_X1  g266(.A1(new_n464), .A2(KEYINPUT90), .A3(new_n439), .ZN(new_n468));
  NAND3_X1  g267(.A1(new_n467), .A2(new_n454), .A3(new_n468), .ZN(new_n469));
  NAND2_X1  g268(.A1(new_n469), .A2(KEYINPUT38), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n461), .A2(new_n463), .A3(new_n470), .ZN(new_n471));
  INV_X1    g270(.A(new_n355), .ZN(new_n472));
  AOI21_X1  g271(.A(new_n363), .B1(new_n389), .B2(new_n399), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT39), .ZN(new_n474));
  AOI21_X1  g273(.A(new_n362), .B1(new_n473), .B2(new_n474), .ZN(new_n475));
  OR2_X1    g274(.A1(new_n473), .A2(new_n474), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n368), .B1(new_n371), .B2(new_n374), .ZN(new_n477));
  AND2_X1   g276(.A1(new_n477), .A2(new_n363), .ZN(new_n478));
  OAI21_X1  g277(.A(new_n475), .B1(new_n476), .B2(new_n478), .ZN(new_n479));
  NOR2_X1   g278(.A1(KEYINPUT87), .A2(KEYINPUT40), .ZN(new_n480));
  NAND2_X1  g279(.A1(new_n479), .A2(new_n480), .ZN(new_n481));
  OR2_X1    g280(.A1(new_n479), .A2(new_n480), .ZN(new_n482));
  NAND4_X1  g281(.A1(new_n442), .A2(new_n402), .A3(new_n481), .A4(new_n482), .ZN(new_n483));
  NAND2_X1  g282(.A1(new_n472), .A2(new_n483), .ZN(new_n484));
  INV_X1    g283(.A(new_n484), .ZN(new_n485));
  NAND2_X1  g284(.A1(new_n471), .A2(new_n485), .ZN(new_n486));
  XNOR2_X1  g285(.A(new_n290), .B(KEYINPUT36), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n416), .A2(new_n443), .ZN(new_n488));
  AOI21_X1  g287(.A(new_n487), .B1(new_n488), .B2(new_n355), .ZN(new_n489));
  AOI21_X1  g288(.A(new_n452), .B1(new_n486), .B2(new_n489), .ZN(new_n490));
  INV_X1    g289(.A(KEYINPUT100), .ZN(new_n491));
  NAND2_X1  g290(.A1(G229gat), .A2(G233gat), .ZN(new_n492));
  INV_X1    g291(.A(G50gat), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n493), .A2(G43gat), .ZN(new_n494));
  INV_X1    g293(.A(G43gat), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n495), .A2(G50gat), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n494), .A2(new_n496), .A3(KEYINPUT15), .ZN(new_n497));
  NOR3_X1   g296(.A1(KEYINPUT14), .A2(G29gat), .A3(G36gat), .ZN(new_n498));
  OAI21_X1  g297(.A(KEYINPUT14), .B1(G29gat), .B2(G36gat), .ZN(new_n499));
  AOI21_X1  g298(.A(new_n498), .B1(KEYINPUT92), .B2(new_n499), .ZN(new_n500));
  OR2_X1    g299(.A1(new_n499), .A2(KEYINPUT92), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n500), .A2(new_n501), .ZN(new_n502));
  XOR2_X1   g301(.A(KEYINPUT93), .B(G36gat), .Z(new_n503));
  NAND2_X1  g302(.A1(new_n503), .A2(G29gat), .ZN(new_n504));
  AOI21_X1  g303(.A(new_n497), .B1(new_n502), .B2(new_n504), .ZN(new_n505));
  INV_X1    g304(.A(KEYINPUT94), .ZN(new_n506));
  OR2_X1    g305(.A1(new_n505), .A2(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n505), .A2(new_n506), .ZN(new_n508));
  NAND2_X1  g307(.A1(new_n507), .A2(new_n508), .ZN(new_n509));
  INV_X1    g308(.A(KEYINPUT15), .ZN(new_n510));
  AOI21_X1  g309(.A(KEYINPUT95), .B1(new_n493), .B2(G43gat), .ZN(new_n511));
  NAND3_X1  g310(.A1(new_n493), .A2(KEYINPUT95), .A3(G43gat), .ZN(new_n512));
  NAND2_X1  g311(.A1(new_n512), .A2(new_n496), .ZN(new_n513));
  OAI21_X1  g312(.A(new_n510), .B1(new_n511), .B2(new_n513), .ZN(new_n514));
  OR2_X1    g313(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n515));
  OAI21_X1  g314(.A(KEYINPUT96), .B1(new_n515), .B2(G36gat), .ZN(new_n516));
  INV_X1    g315(.A(KEYINPUT96), .ZN(new_n517));
  NAND2_X1  g316(.A1(new_n498), .A2(new_n517), .ZN(new_n518));
  NAND3_X1  g317(.A1(new_n516), .A2(new_n518), .A3(new_n499), .ZN(new_n519));
  NAND4_X1  g318(.A1(new_n514), .A2(new_n519), .A3(new_n504), .A4(new_n497), .ZN(new_n520));
  INV_X1    g319(.A(KEYINPUT97), .ZN(new_n521));
  OR2_X1    g320(.A1(new_n520), .A2(new_n521), .ZN(new_n522));
  NAND2_X1  g321(.A1(new_n520), .A2(new_n521), .ZN(new_n523));
  NAND2_X1  g322(.A1(new_n522), .A2(new_n523), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n509), .A2(new_n524), .ZN(new_n525));
  XNOR2_X1  g324(.A(G15gat), .B(G22gat), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT16), .ZN(new_n527));
  OAI21_X1  g326(.A(new_n526), .B1(new_n527), .B2(G1gat), .ZN(new_n528));
  OAI21_X1  g327(.A(new_n528), .B1(G1gat), .B2(new_n526), .ZN(new_n529));
  XOR2_X1   g328(.A(new_n529), .B(G8gat), .Z(new_n530));
  INV_X1    g329(.A(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n525), .A2(new_n531), .ZN(new_n532));
  AOI22_X1  g331(.A1(new_n507), .A2(new_n508), .B1(new_n522), .B2(new_n523), .ZN(new_n533));
  OAI21_X1  g332(.A(new_n530), .B1(new_n533), .B2(KEYINPUT17), .ZN(new_n534));
  INV_X1    g333(.A(KEYINPUT17), .ZN(new_n535));
  NOR2_X1   g334(.A1(new_n525), .A2(new_n535), .ZN(new_n536));
  OAI211_X1 g335(.A(new_n492), .B(new_n532), .C1(new_n534), .C2(new_n536), .ZN(new_n537));
  INV_X1    g336(.A(KEYINPUT18), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(new_n525), .A2(new_n535), .ZN(new_n540));
  NAND2_X1  g339(.A1(new_n533), .A2(KEYINPUT17), .ZN(new_n541));
  NAND3_X1  g340(.A1(new_n540), .A2(new_n541), .A3(new_n530), .ZN(new_n542));
  NAND4_X1  g341(.A1(new_n542), .A2(KEYINPUT18), .A3(new_n492), .A4(new_n532), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n533), .A2(new_n530), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n532), .A2(new_n544), .A3(KEYINPUT99), .ZN(new_n545));
  OR3_X1    g344(.A1(new_n533), .A2(KEYINPUT99), .A3(new_n530), .ZN(new_n546));
  XOR2_X1   g345(.A(KEYINPUT98), .B(KEYINPUT13), .Z(new_n547));
  XNOR2_X1  g346(.A(new_n547), .B(new_n492), .ZN(new_n548));
  NAND3_X1  g347(.A1(new_n545), .A2(new_n546), .A3(new_n548), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n539), .A2(new_n543), .A3(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(G113gat), .B(G141gat), .ZN(new_n551));
  XNOR2_X1  g350(.A(new_n551), .B(G197gat), .ZN(new_n552));
  XOR2_X1   g351(.A(KEYINPUT11), .B(G169gat), .Z(new_n553));
  XNOR2_X1  g352(.A(new_n552), .B(new_n553), .ZN(new_n554));
  XOR2_X1   g353(.A(new_n554), .B(KEYINPUT12), .Z(new_n555));
  INV_X1    g354(.A(new_n555), .ZN(new_n556));
  AND3_X1   g355(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n557));
  AOI21_X1  g356(.A(new_n556), .B1(new_n550), .B2(KEYINPUT91), .ZN(new_n558));
  OAI21_X1  g357(.A(new_n491), .B1(new_n557), .B2(new_n558), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n550), .A2(KEYINPUT91), .ZN(new_n560));
  NAND2_X1  g359(.A1(new_n560), .A2(new_n555), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n550), .A2(KEYINPUT91), .A3(new_n556), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n561), .A2(KEYINPUT100), .A3(new_n562), .ZN(new_n563));
  NAND2_X1  g362(.A1(new_n559), .A2(new_n563), .ZN(new_n564));
  INV_X1    g363(.A(new_n564), .ZN(new_n565));
  NOR2_X1   g364(.A1(new_n490), .A2(new_n565), .ZN(new_n566));
  XOR2_X1   g365(.A(KEYINPUT106), .B(G92gat), .Z(new_n567));
  INV_X1    g366(.A(G85gat), .ZN(new_n568));
  NAND2_X1  g367(.A1(new_n567), .A2(new_n568), .ZN(new_n569));
  NAND2_X1  g368(.A1(G85gat), .A2(G92gat), .ZN(new_n570));
  XNOR2_X1  g369(.A(new_n570), .B(KEYINPUT7), .ZN(new_n571));
  INV_X1    g370(.A(G99gat), .ZN(new_n572));
  INV_X1    g371(.A(G106gat), .ZN(new_n573));
  OAI21_X1  g372(.A(KEYINPUT8), .B1(new_n572), .B2(new_n573), .ZN(new_n574));
  NAND3_X1  g373(.A1(new_n569), .A2(new_n571), .A3(new_n574), .ZN(new_n575));
  XNOR2_X1  g374(.A(G99gat), .B(G106gat), .ZN(new_n576));
  XNOR2_X1  g375(.A(new_n575), .B(new_n576), .ZN(new_n577));
  INV_X1    g376(.A(new_n577), .ZN(new_n578));
  NAND3_X1  g377(.A1(new_n540), .A2(new_n541), .A3(new_n578), .ZN(new_n579));
  XOR2_X1   g378(.A(G190gat), .B(G218gat), .Z(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  AND2_X1   g380(.A1(G232gat), .A2(G233gat), .ZN(new_n582));
  AOI22_X1  g381(.A1(new_n525), .A2(new_n577), .B1(KEYINPUT41), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n579), .A2(new_n581), .A3(new_n583), .ZN(new_n584));
  INV_X1    g383(.A(new_n584), .ZN(new_n585));
  AOI21_X1  g384(.A(new_n581), .B1(new_n579), .B2(new_n583), .ZN(new_n586));
  INV_X1    g385(.A(KEYINPUT107), .ZN(new_n587));
  NOR2_X1   g386(.A1(new_n582), .A2(KEYINPUT41), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n588), .B(KEYINPUT105), .ZN(new_n589));
  XOR2_X1   g388(.A(G134gat), .B(G162gat), .Z(new_n590));
  XNOR2_X1  g389(.A(new_n589), .B(new_n590), .ZN(new_n591));
  OAI22_X1  g390(.A1(new_n585), .A2(new_n586), .B1(new_n587), .B2(new_n591), .ZN(new_n592));
  INV_X1    g391(.A(new_n586), .ZN(new_n593));
  XNOR2_X1  g392(.A(new_n591), .B(new_n587), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n593), .A2(new_n584), .A3(new_n594), .ZN(new_n595));
  NAND2_X1  g394(.A1(new_n592), .A2(new_n595), .ZN(new_n596));
  INV_X1    g395(.A(new_n596), .ZN(new_n597));
  INV_X1    g396(.A(KEYINPUT108), .ZN(new_n598));
  XOR2_X1   g397(.A(G71gat), .B(G78gat), .Z(new_n599));
  INV_X1    g398(.A(new_n599), .ZN(new_n600));
  XNOR2_X1  g399(.A(G57gat), .B(G64gat), .ZN(new_n601));
  NOR2_X1   g400(.A1(new_n601), .A2(KEYINPUT101), .ZN(new_n602));
  AOI21_X1  g401(.A(KEYINPUT9), .B1(G71gat), .B2(G78gat), .ZN(new_n603));
  NOR2_X1   g402(.A1(new_n602), .A2(new_n603), .ZN(new_n604));
  NAND2_X1  g403(.A1(new_n601), .A2(KEYINPUT101), .ZN(new_n605));
  AOI21_X1  g404(.A(new_n600), .B1(new_n604), .B2(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(G57gat), .ZN(new_n607));
  INV_X1    g406(.A(G64gat), .ZN(new_n608));
  OR2_X1    g407(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n609));
  NAND2_X1  g408(.A1(new_n608), .A2(KEYINPUT102), .ZN(new_n610));
  AOI21_X1  g409(.A(new_n607), .B1(new_n609), .B2(new_n610), .ZN(new_n611));
  INV_X1    g410(.A(KEYINPUT103), .ZN(new_n612));
  AOI22_X1  g411(.A1(new_n611), .A2(new_n612), .B1(new_n607), .B2(G64gat), .ZN(new_n613));
  AND2_X1   g412(.A1(new_n609), .A2(new_n610), .ZN(new_n614));
  OAI21_X1  g413(.A(KEYINPUT103), .B1(new_n614), .B2(new_n607), .ZN(new_n615));
  NAND2_X1  g414(.A1(new_n613), .A2(new_n615), .ZN(new_n616));
  NOR2_X1   g415(.A1(new_n599), .A2(new_n603), .ZN(new_n617));
  AOI21_X1  g416(.A(new_n606), .B1(new_n616), .B2(new_n617), .ZN(new_n618));
  NOR2_X1   g417(.A1(new_n618), .A2(KEYINPUT21), .ZN(new_n619));
  XNOR2_X1  g418(.A(G127gat), .B(G155gat), .ZN(new_n620));
  INV_X1    g419(.A(new_n620), .ZN(new_n621));
  NAND2_X1  g420(.A1(new_n619), .A2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n620), .B1(new_n618), .B2(KEYINPUT21), .ZN(new_n623));
  NAND2_X1  g422(.A1(new_n622), .A2(new_n623), .ZN(new_n624));
  AOI21_X1  g423(.A(new_n531), .B1(new_n618), .B2(KEYINPUT21), .ZN(new_n625));
  OR2_X1    g424(.A1(new_n624), .A2(new_n625), .ZN(new_n626));
  NAND2_X1  g425(.A1(new_n624), .A2(new_n625), .ZN(new_n627));
  NAND2_X1  g426(.A1(G231gat), .A2(G233gat), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(KEYINPUT104), .ZN(new_n629));
  XOR2_X1   g428(.A(KEYINPUT19), .B(KEYINPUT20), .Z(new_n630));
  XNOR2_X1  g429(.A(new_n629), .B(new_n630), .ZN(new_n631));
  XNOR2_X1  g430(.A(G183gat), .B(G211gat), .ZN(new_n632));
  XNOR2_X1  g431(.A(new_n631), .B(new_n632), .ZN(new_n633));
  AND3_X1   g432(.A1(new_n626), .A2(new_n627), .A3(new_n633), .ZN(new_n634));
  AOI21_X1  g433(.A(new_n633), .B1(new_n626), .B2(new_n627), .ZN(new_n635));
  OR2_X1    g434(.A1(new_n634), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  NAND3_X1  g436(.A1(new_n597), .A2(new_n598), .A3(new_n637), .ZN(new_n638));
  OAI21_X1  g437(.A(KEYINPUT108), .B1(new_n596), .B2(new_n636), .ZN(new_n639));
  INV_X1    g438(.A(new_n603), .ZN(new_n640));
  NAND3_X1  g439(.A1(new_n616), .A2(new_n600), .A3(new_n640), .ZN(new_n641));
  INV_X1    g440(.A(new_n606), .ZN(new_n642));
  NAND2_X1  g441(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  NAND2_X1  g442(.A1(new_n643), .A2(new_n578), .ZN(new_n644));
  INV_X1    g443(.A(KEYINPUT10), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n618), .A2(new_n577), .ZN(new_n646));
  NAND3_X1  g445(.A1(new_n644), .A2(new_n645), .A3(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n618), .A2(KEYINPUT10), .A3(new_n577), .ZN(new_n648));
  NAND2_X1  g447(.A1(new_n647), .A2(new_n648), .ZN(new_n649));
  INV_X1    g448(.A(G230gat), .ZN(new_n650));
  NOR2_X1   g449(.A1(new_n650), .A2(new_n268), .ZN(new_n651));
  INV_X1    g450(.A(new_n651), .ZN(new_n652));
  NAND2_X1  g451(.A1(new_n649), .A2(new_n652), .ZN(new_n653));
  NAND2_X1  g452(.A1(new_n644), .A2(new_n646), .ZN(new_n654));
  NAND2_X1  g453(.A1(new_n654), .A2(new_n651), .ZN(new_n655));
  NAND2_X1  g454(.A1(new_n653), .A2(new_n655), .ZN(new_n656));
  XNOR2_X1  g455(.A(G120gat), .B(G148gat), .ZN(new_n657));
  XNOR2_X1  g456(.A(G176gat), .B(G204gat), .ZN(new_n658));
  XOR2_X1   g457(.A(new_n657), .B(new_n658), .Z(new_n659));
  INV_X1    g458(.A(new_n659), .ZN(new_n660));
  NAND2_X1  g459(.A1(new_n656), .A2(new_n660), .ZN(new_n661));
  OR2_X1    g460(.A1(new_n655), .A2(KEYINPUT109), .ZN(new_n662));
  NAND2_X1  g461(.A1(new_n655), .A2(KEYINPUT109), .ZN(new_n663));
  NAND4_X1  g462(.A1(new_n662), .A2(new_n653), .A3(new_n659), .A4(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n661), .A2(new_n664), .ZN(new_n665));
  INV_X1    g464(.A(new_n665), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n638), .A2(new_n639), .A3(new_n666), .ZN(new_n667));
  INV_X1    g466(.A(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n566), .A2(new_n668), .ZN(new_n669));
  INV_X1    g468(.A(new_n669), .ZN(new_n670));
  INV_X1    g469(.A(new_n416), .ZN(new_n671));
  NAND2_X1  g470(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  XNOR2_X1  g471(.A(new_n672), .B(G1gat), .ZN(G1324gat));
  XOR2_X1   g472(.A(KEYINPUT16), .B(G8gat), .Z(new_n674));
  NAND4_X1  g473(.A1(new_n670), .A2(KEYINPUT42), .A3(new_n442), .A4(new_n674), .ZN(new_n675));
  OR3_X1    g474(.A1(new_n669), .A2(KEYINPUT110), .A3(new_n443), .ZN(new_n676));
  OAI21_X1  g475(.A(KEYINPUT110), .B1(new_n669), .B2(new_n443), .ZN(new_n677));
  NAND3_X1  g476(.A1(new_n676), .A2(G8gat), .A3(new_n677), .ZN(new_n678));
  INV_X1    g477(.A(new_n674), .ZN(new_n679));
  AOI21_X1  g478(.A(new_n679), .B1(new_n676), .B2(new_n677), .ZN(new_n680));
  OAI211_X1 g479(.A(new_n675), .B(new_n678), .C1(new_n680), .C2(KEYINPUT42), .ZN(G1325gat));
  INV_X1    g480(.A(new_n487), .ZN(new_n682));
  OAI21_X1  g481(.A(G15gat), .B1(new_n669), .B2(new_n682), .ZN(new_n683));
  OR2_X1    g482(.A1(new_n290), .A2(G15gat), .ZN(new_n684));
  OAI21_X1  g483(.A(new_n683), .B1(new_n669), .B2(new_n684), .ZN(G1326gat));
  OR3_X1    g484(.A1(new_n669), .A2(KEYINPUT111), .A3(new_n472), .ZN(new_n686));
  OAI21_X1  g485(.A(KEYINPUT111), .B1(new_n669), .B2(new_n472), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n686), .A2(new_n687), .ZN(new_n688));
  XNOR2_X1  g487(.A(KEYINPUT43), .B(G22gat), .ZN(new_n689));
  XNOR2_X1  g488(.A(new_n688), .B(new_n689), .ZN(G1327gat));
  OAI21_X1  g489(.A(KEYINPUT44), .B1(new_n490), .B2(new_n597), .ZN(new_n691));
  NAND2_X1  g490(.A1(new_n444), .A2(KEYINPUT35), .ZN(new_n692));
  NAND2_X1  g491(.A1(new_n445), .A2(new_n451), .ZN(new_n693));
  NAND2_X1  g492(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  AOI22_X1  g493(.A1(new_n460), .A2(KEYINPUT89), .B1(KEYINPUT38), .B2(new_n469), .ZN(new_n695));
  AOI21_X1  g494(.A(new_n484), .B1(new_n695), .B2(new_n463), .ZN(new_n696));
  NAND2_X1  g495(.A1(new_n488), .A2(new_n355), .ZN(new_n697));
  NAND2_X1  g496(.A1(new_n682), .A2(new_n697), .ZN(new_n698));
  OAI21_X1  g497(.A(new_n694), .B1(new_n696), .B2(new_n698), .ZN(new_n699));
  XNOR2_X1  g498(.A(KEYINPUT113), .B(KEYINPUT44), .ZN(new_n700));
  XNOR2_X1  g499(.A(new_n596), .B(KEYINPUT114), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n699), .A2(new_n700), .A3(new_n701), .ZN(new_n702));
  NAND2_X1  g501(.A1(new_n691), .A2(new_n702), .ZN(new_n703));
  NOR2_X1   g502(.A1(new_n557), .A2(new_n558), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g504(.A1(new_n666), .A2(new_n636), .ZN(new_n706));
  NOR2_X1   g505(.A1(new_n705), .A2(new_n706), .ZN(new_n707));
  NAND2_X1  g506(.A1(new_n703), .A2(new_n707), .ZN(new_n708));
  OAI21_X1  g507(.A(G29gat), .B1(new_n708), .B2(new_n416), .ZN(new_n709));
  NOR2_X1   g508(.A1(new_n706), .A2(new_n597), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n416), .A2(G29gat), .ZN(new_n711));
  NAND3_X1  g510(.A1(new_n566), .A2(new_n710), .A3(new_n711), .ZN(new_n712));
  OR2_X1    g511(.A1(new_n712), .A2(KEYINPUT112), .ZN(new_n713));
  INV_X1    g512(.A(KEYINPUT45), .ZN(new_n714));
  NAND2_X1  g513(.A1(new_n712), .A2(KEYINPUT112), .ZN(new_n715));
  AND3_X1   g514(.A1(new_n713), .A2(new_n714), .A3(new_n715), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n714), .B1(new_n713), .B2(new_n715), .ZN(new_n717));
  OAI21_X1  g516(.A(new_n709), .B1(new_n716), .B2(new_n717), .ZN(G1328gat));
  NAND3_X1  g517(.A1(new_n699), .A2(new_n564), .A3(new_n710), .ZN(new_n719));
  NOR3_X1   g518(.A1(new_n719), .A2(new_n443), .A3(new_n503), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT46), .ZN(new_n721));
  OAI21_X1  g520(.A(new_n503), .B1(new_n708), .B2(new_n443), .ZN(new_n722));
  NAND2_X1  g521(.A1(new_n721), .A2(new_n722), .ZN(G1329gat));
  OAI21_X1  g522(.A(new_n495), .B1(new_n719), .B2(new_n290), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n487), .A2(G43gat), .ZN(new_n725));
  OAI21_X1  g524(.A(new_n724), .B1(new_n708), .B2(new_n725), .ZN(new_n726));
  XNOR2_X1  g525(.A(new_n726), .B(KEYINPUT47), .ZN(G1330gat));
  OAI21_X1  g526(.A(G50gat), .B1(new_n708), .B2(new_n472), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT115), .ZN(new_n729));
  AOI211_X1 g528(.A(G50gat), .B(new_n472), .C1(new_n719), .C2(new_n729), .ZN(new_n730));
  OAI21_X1  g529(.A(new_n730), .B1(new_n729), .B2(new_n719), .ZN(new_n731));
  INV_X1    g530(.A(KEYINPUT48), .ZN(new_n732));
  AND3_X1   g531(.A1(new_n728), .A2(new_n731), .A3(new_n732), .ZN(new_n733));
  AOI21_X1  g532(.A(new_n732), .B1(new_n728), .B2(new_n731), .ZN(new_n734));
  NOR2_X1   g533(.A1(new_n733), .A2(new_n734), .ZN(G1331gat));
  NAND4_X1  g534(.A1(new_n705), .A2(new_n638), .A3(new_n639), .A4(new_n665), .ZN(new_n736));
  NOR2_X1   g535(.A1(new_n490), .A2(new_n736), .ZN(new_n737));
  NAND2_X1  g536(.A1(new_n737), .A2(new_n671), .ZN(new_n738));
  XNOR2_X1  g537(.A(new_n738), .B(G57gat), .ZN(G1332gat));
  NAND2_X1  g538(.A1(new_n737), .A2(new_n442), .ZN(new_n740));
  OAI21_X1  g539(.A(new_n740), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n741));
  XOR2_X1   g540(.A(KEYINPUT49), .B(G64gat), .Z(new_n742));
  OAI21_X1  g541(.A(new_n741), .B1(new_n740), .B2(new_n742), .ZN(G1333gat));
  INV_X1    g542(.A(new_n290), .ZN(new_n744));
  NAND2_X1  g543(.A1(new_n737), .A2(new_n744), .ZN(new_n745));
  INV_X1    g544(.A(KEYINPUT116), .ZN(new_n746));
  AOI21_X1  g545(.A(G71gat), .B1(new_n745), .B2(new_n746), .ZN(new_n747));
  OAI21_X1  g546(.A(new_n747), .B1(new_n746), .B2(new_n745), .ZN(new_n748));
  NAND3_X1  g547(.A1(new_n737), .A2(G71gat), .A3(new_n487), .ZN(new_n749));
  NAND2_X1  g548(.A1(new_n748), .A2(new_n749), .ZN(new_n750));
  NAND2_X1  g549(.A1(new_n750), .A2(KEYINPUT50), .ZN(new_n751));
  INV_X1    g550(.A(KEYINPUT50), .ZN(new_n752));
  NAND3_X1  g551(.A1(new_n748), .A2(new_n752), .A3(new_n749), .ZN(new_n753));
  NAND2_X1  g552(.A1(new_n751), .A2(new_n753), .ZN(G1334gat));
  NAND2_X1  g553(.A1(new_n737), .A2(new_n355), .ZN(new_n755));
  XNOR2_X1  g554(.A(new_n755), .B(G78gat), .ZN(G1335gat));
  NOR2_X1   g555(.A1(new_n704), .A2(new_n637), .ZN(new_n757));
  NAND2_X1  g556(.A1(new_n757), .A2(new_n665), .ZN(new_n758));
  AOI21_X1  g557(.A(new_n758), .B1(new_n691), .B2(new_n702), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n671), .ZN(new_n760));
  NAND2_X1  g559(.A1(new_n760), .A2(G85gat), .ZN(new_n761));
  NAND3_X1  g560(.A1(new_n699), .A2(new_n596), .A3(new_n757), .ZN(new_n762));
  INV_X1    g561(.A(KEYINPUT51), .ZN(new_n763));
  XNOR2_X1  g562(.A(new_n762), .B(new_n763), .ZN(new_n764));
  INV_X1    g563(.A(new_n764), .ZN(new_n765));
  NAND3_X1  g564(.A1(new_n671), .A2(new_n568), .A3(new_n665), .ZN(new_n766));
  OAI21_X1  g565(.A(new_n761), .B1(new_n765), .B2(new_n766), .ZN(G1336gat));
  NOR2_X1   g566(.A1(new_n666), .A2(G92gat), .ZN(new_n768));
  NAND3_X1  g567(.A1(new_n764), .A2(new_n442), .A3(new_n768), .ZN(new_n769));
  NAND2_X1  g568(.A1(new_n759), .A2(new_n442), .ZN(new_n770));
  INV_X1    g569(.A(new_n770), .ZN(new_n771));
  OAI21_X1  g570(.A(new_n769), .B1(new_n771), .B2(new_n567), .ZN(new_n772));
  NAND2_X1  g571(.A1(new_n772), .A2(KEYINPUT52), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT52), .ZN(new_n774));
  OAI211_X1 g573(.A(new_n769), .B(new_n774), .C1(new_n771), .C2(new_n567), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n773), .A2(new_n775), .ZN(G1337gat));
  INV_X1    g575(.A(new_n758), .ZN(new_n777));
  INV_X1    g576(.A(KEYINPUT44), .ZN(new_n778));
  AOI21_X1  g577(.A(new_n778), .B1(new_n699), .B2(new_n596), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n701), .A2(new_n700), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n486), .A2(new_n489), .ZN(new_n781));
  AOI21_X1  g580(.A(new_n780), .B1(new_n781), .B2(new_n694), .ZN(new_n782));
  OAI211_X1 g581(.A(new_n487), .B(new_n777), .C1(new_n779), .C2(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(KEYINPUT117), .ZN(new_n784));
  NAND2_X1  g583(.A1(new_n783), .A2(new_n784), .ZN(new_n785));
  NAND4_X1  g584(.A1(new_n703), .A2(KEYINPUT117), .A3(new_n487), .A4(new_n777), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n785), .A2(new_n786), .A3(G99gat), .ZN(new_n787));
  NAND4_X1  g586(.A1(new_n764), .A2(new_n572), .A3(new_n744), .A4(new_n665), .ZN(new_n788));
  NAND2_X1  g587(.A1(new_n787), .A2(new_n788), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n789), .A2(KEYINPUT118), .ZN(new_n790));
  INV_X1    g589(.A(KEYINPUT118), .ZN(new_n791));
  NAND3_X1  g590(.A1(new_n787), .A2(new_n788), .A3(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n790), .A2(new_n792), .ZN(G1338gat));
  AOI21_X1  g592(.A(new_n573), .B1(new_n759), .B2(new_n355), .ZN(new_n794));
  NOR3_X1   g593(.A1(new_n472), .A2(G106gat), .A3(new_n666), .ZN(new_n795));
  XNOR2_X1  g594(.A(new_n795), .B(KEYINPUT119), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n794), .B1(new_n764), .B2(new_n796), .ZN(new_n797));
  INV_X1    g596(.A(KEYINPUT53), .ZN(new_n798));
  INV_X1    g597(.A(new_n795), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n798), .B1(new_n765), .B2(new_n799), .ZN(new_n800));
  OAI22_X1  g599(.A1(new_n797), .A2(new_n798), .B1(new_n800), .B2(new_n794), .ZN(G1339gat));
  NOR2_X1   g600(.A1(new_n667), .A2(new_n704), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n647), .A2(new_n651), .A3(new_n648), .ZN(new_n803));
  NAND3_X1  g602(.A1(new_n653), .A2(KEYINPUT54), .A3(new_n803), .ZN(new_n804));
  AOI21_X1  g603(.A(new_n651), .B1(new_n647), .B2(new_n648), .ZN(new_n805));
  INV_X1    g604(.A(KEYINPUT54), .ZN(new_n806));
  AOI21_X1  g605(.A(new_n659), .B1(new_n805), .B2(new_n806), .ZN(new_n807));
  NAND2_X1  g606(.A1(new_n804), .A2(new_n807), .ZN(new_n808));
  INV_X1    g607(.A(KEYINPUT55), .ZN(new_n809));
  NAND2_X1  g608(.A1(new_n808), .A2(new_n809), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n804), .A2(KEYINPUT55), .A3(new_n807), .ZN(new_n811));
  NAND3_X1  g610(.A1(new_n810), .A2(new_n811), .A3(new_n664), .ZN(new_n812));
  INV_X1    g611(.A(new_n812), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n550), .A2(new_n555), .ZN(new_n814));
  AND2_X1   g613(.A1(new_n542), .A2(new_n532), .ZN(new_n815));
  AOI21_X1  g614(.A(new_n548), .B1(new_n545), .B2(new_n546), .ZN(new_n816));
  INV_X1    g615(.A(KEYINPUT120), .ZN(new_n817));
  OAI22_X1  g616(.A1(new_n815), .A2(new_n492), .B1(new_n816), .B2(new_n817), .ZN(new_n818));
  AND2_X1   g617(.A1(new_n816), .A2(new_n817), .ZN(new_n819));
  OAI21_X1  g618(.A(new_n554), .B1(new_n818), .B2(new_n819), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n814), .A2(new_n820), .ZN(new_n821));
  NAND3_X1  g620(.A1(new_n701), .A2(new_n813), .A3(new_n821), .ZN(new_n822));
  AOI22_X1  g621(.A1(new_n821), .A2(new_n665), .B1(new_n704), .B2(new_n813), .ZN(new_n823));
  OAI21_X1  g622(.A(new_n822), .B1(new_n823), .B2(new_n701), .ZN(new_n824));
  AOI21_X1  g623(.A(new_n802), .B1(new_n824), .B2(new_n636), .ZN(new_n825));
  NOR2_X1   g624(.A1(new_n825), .A2(new_n416), .ZN(new_n826));
  INV_X1    g625(.A(new_n356), .ZN(new_n827));
  NOR2_X1   g626(.A1(new_n827), .A2(new_n442), .ZN(new_n828));
  NAND2_X1  g627(.A1(new_n826), .A2(new_n828), .ZN(new_n829));
  INV_X1    g628(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g629(.A(G113gat), .B1(new_n830), .B2(new_n704), .ZN(new_n831));
  NOR2_X1   g630(.A1(new_n825), .A2(new_n355), .ZN(new_n832));
  NOR2_X1   g631(.A1(new_n416), .A2(new_n442), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n832), .A2(new_n744), .A3(new_n833), .ZN(new_n834));
  NOR3_X1   g633(.A1(new_n834), .A2(new_n244), .A3(new_n565), .ZN(new_n835));
  NOR2_X1   g634(.A1(new_n831), .A2(new_n835), .ZN(G1340gat));
  OAI21_X1  g635(.A(G120gat), .B1(new_n834), .B2(new_n666), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n665), .A2(new_n261), .A3(new_n262), .ZN(new_n838));
  OAI21_X1  g637(.A(new_n837), .B1(new_n829), .B2(new_n838), .ZN(G1341gat));
  NAND3_X1  g638(.A1(new_n830), .A2(new_n257), .A3(new_n637), .ZN(new_n840));
  OAI21_X1  g639(.A(G127gat), .B1(new_n834), .B2(new_n636), .ZN(new_n841));
  NAND2_X1  g640(.A1(new_n840), .A2(new_n841), .ZN(G1342gat));
  NOR3_X1   g641(.A1(new_n829), .A2(G134gat), .A3(new_n597), .ZN(new_n843));
  INV_X1    g642(.A(new_n843), .ZN(new_n844));
  OR2_X1    g643(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n845));
  OAI21_X1  g644(.A(G134gat), .B1(new_n834), .B2(new_n597), .ZN(new_n846));
  NAND2_X1  g645(.A1(new_n844), .A2(KEYINPUT56), .ZN(new_n847));
  NAND3_X1  g646(.A1(new_n845), .A2(new_n846), .A3(new_n847), .ZN(G1343gat));
  INV_X1    g647(.A(KEYINPUT121), .ZN(new_n849));
  INV_X1    g648(.A(new_n802), .ZN(new_n850));
  AOI21_X1  g649(.A(new_n812), .B1(new_n559), .B2(new_n563), .ZN(new_n851));
  AND3_X1   g650(.A1(new_n814), .A2(new_n820), .A3(new_n665), .ZN(new_n852));
  OAI21_X1  g651(.A(new_n597), .B1(new_n851), .B2(new_n852), .ZN(new_n853));
  AND2_X1   g652(.A1(new_n853), .A2(new_n822), .ZN(new_n854));
  OAI21_X1  g653(.A(new_n850), .B1(new_n854), .B2(new_n637), .ZN(new_n855));
  INV_X1    g654(.A(KEYINPUT57), .ZN(new_n856));
  NOR2_X1   g655(.A1(new_n472), .A2(new_n856), .ZN(new_n857));
  AOI21_X1  g656(.A(new_n849), .B1(new_n855), .B2(new_n857), .ZN(new_n858));
  AOI21_X1  g657(.A(new_n637), .B1(new_n853), .B2(new_n822), .ZN(new_n859));
  OAI211_X1 g658(.A(new_n849), .B(new_n857), .C1(new_n859), .C2(new_n802), .ZN(new_n860));
  OAI21_X1  g659(.A(new_n856), .B1(new_n825), .B2(new_n472), .ZN(new_n861));
  NAND2_X1  g660(.A1(new_n860), .A2(new_n861), .ZN(new_n862));
  NOR2_X1   g661(.A1(new_n858), .A2(new_n862), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n682), .A2(new_n833), .ZN(new_n864));
  NOR2_X1   g663(.A1(new_n863), .A2(new_n864), .ZN(new_n865));
  NAND2_X1  g664(.A1(new_n865), .A2(new_n564), .ZN(new_n866));
  NAND2_X1  g665(.A1(new_n866), .A2(G141gat), .ZN(new_n867));
  NOR3_X1   g666(.A1(new_n487), .A2(new_n472), .A3(new_n442), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n826), .A2(new_n868), .ZN(new_n869));
  NOR3_X1   g668(.A1(new_n869), .A2(G141gat), .A3(new_n565), .ZN(new_n870));
  NOR2_X1   g669(.A1(new_n870), .A2(KEYINPUT58), .ZN(new_n871));
  NAND2_X1  g670(.A1(new_n867), .A2(new_n871), .ZN(new_n872));
  INV_X1    g671(.A(new_n864), .ZN(new_n873));
  OAI211_X1 g672(.A(new_n704), .B(new_n873), .C1(new_n858), .C2(new_n862), .ZN(new_n874));
  INV_X1    g673(.A(KEYINPUT122), .ZN(new_n875));
  AND3_X1   g674(.A1(new_n874), .A2(new_n875), .A3(G141gat), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n875), .B1(new_n874), .B2(G141gat), .ZN(new_n877));
  NOR3_X1   g676(.A1(new_n876), .A2(new_n877), .A3(new_n870), .ZN(new_n878));
  INV_X1    g677(.A(KEYINPUT58), .ZN(new_n879));
  OAI21_X1  g678(.A(new_n872), .B1(new_n878), .B2(new_n879), .ZN(G1344gat));
  INV_X1    g679(.A(new_n869), .ZN(new_n881));
  INV_X1    g680(.A(G148gat), .ZN(new_n882));
  NAND3_X1  g681(.A1(new_n881), .A2(new_n882), .A3(new_n665), .ZN(new_n883));
  INV_X1    g682(.A(KEYINPUT59), .ZN(new_n884));
  NOR2_X1   g683(.A1(new_n864), .A2(new_n666), .ZN(new_n885));
  INV_X1    g684(.A(new_n885), .ZN(new_n886));
  INV_X1    g685(.A(KEYINPUT123), .ZN(new_n887));
  INV_X1    g686(.A(new_n857), .ZN(new_n888));
  OR3_X1    g687(.A1(new_n825), .A2(new_n887), .A3(new_n888), .ZN(new_n889));
  OAI21_X1  g688(.A(new_n887), .B1(new_n825), .B2(new_n888), .ZN(new_n890));
  AND2_X1   g689(.A1(new_n889), .A2(new_n890), .ZN(new_n891));
  NAND3_X1  g690(.A1(new_n813), .A2(KEYINPUT124), .A3(new_n596), .ZN(new_n892));
  INV_X1    g691(.A(KEYINPUT124), .ZN(new_n893));
  OAI21_X1  g692(.A(new_n893), .B1(new_n597), .B2(new_n812), .ZN(new_n894));
  NAND3_X1  g693(.A1(new_n892), .A2(new_n821), .A3(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n853), .A2(new_n895), .ZN(new_n896));
  AOI22_X1  g695(.A1(new_n896), .A2(new_n636), .B1(new_n565), .B2(new_n668), .ZN(new_n897));
  OAI21_X1  g696(.A(new_n856), .B1(new_n897), .B2(new_n472), .ZN(new_n898));
  AOI21_X1  g697(.A(new_n886), .B1(new_n891), .B2(new_n898), .ZN(new_n899));
  INV_X1    g698(.A(KEYINPUT125), .ZN(new_n900));
  AOI21_X1  g699(.A(new_n882), .B1(new_n899), .B2(new_n900), .ZN(new_n901));
  AND3_X1   g700(.A1(new_n898), .A2(new_n890), .A3(new_n889), .ZN(new_n902));
  OAI21_X1  g701(.A(KEYINPUT125), .B1(new_n902), .B2(new_n886), .ZN(new_n903));
  AOI21_X1  g702(.A(new_n884), .B1(new_n901), .B2(new_n903), .ZN(new_n904));
  AOI211_X1 g703(.A(KEYINPUT59), .B(new_n882), .C1(new_n865), .C2(new_n665), .ZN(new_n905));
  OAI21_X1  g704(.A(new_n883), .B1(new_n904), .B2(new_n905), .ZN(G1345gat));
  INV_X1    g705(.A(G155gat), .ZN(new_n907));
  NAND3_X1  g706(.A1(new_n881), .A2(new_n907), .A3(new_n637), .ZN(new_n908));
  NAND2_X1  g707(.A1(new_n865), .A2(new_n637), .ZN(new_n909));
  INV_X1    g708(.A(new_n909), .ZN(new_n910));
  OAI21_X1  g709(.A(new_n908), .B1(new_n910), .B2(new_n907), .ZN(G1346gat));
  AOI21_X1  g710(.A(G162gat), .B1(new_n881), .B2(new_n596), .ZN(new_n912));
  AND2_X1   g711(.A1(new_n701), .A2(G162gat), .ZN(new_n913));
  AOI21_X1  g712(.A(new_n912), .B1(new_n865), .B2(new_n913), .ZN(G1347gat));
  NAND4_X1  g713(.A1(new_n832), .A2(new_n416), .A3(new_n442), .A4(new_n744), .ZN(new_n915));
  NOR3_X1   g714(.A1(new_n915), .A2(new_n207), .A3(new_n565), .ZN(new_n916));
  NOR4_X1   g715(.A1(new_n825), .A2(new_n671), .A3(new_n443), .A4(new_n827), .ZN(new_n917));
  AOI21_X1  g716(.A(G169gat), .B1(new_n917), .B2(new_n704), .ZN(new_n918));
  NOR2_X1   g717(.A1(new_n916), .A2(new_n918), .ZN(G1348gat));
  OAI21_X1  g718(.A(G176gat), .B1(new_n915), .B2(new_n666), .ZN(new_n920));
  NAND3_X1  g719(.A1(new_n917), .A2(new_n208), .A3(new_n665), .ZN(new_n921));
  NAND2_X1  g720(.A1(new_n920), .A2(new_n921), .ZN(G1349gat));
  OAI21_X1  g721(.A(G183gat), .B1(new_n915), .B2(new_n636), .ZN(new_n923));
  AND2_X1   g722(.A1(new_n637), .A2(new_n215), .ZN(new_n924));
  AOI22_X1  g723(.A1(new_n917), .A2(new_n924), .B1(KEYINPUT126), .B2(KEYINPUT60), .ZN(new_n925));
  NAND2_X1  g724(.A1(new_n923), .A2(new_n925), .ZN(new_n926));
  NOR2_X1   g725(.A1(KEYINPUT126), .A2(KEYINPUT60), .ZN(new_n927));
  XOR2_X1   g726(.A(new_n926), .B(new_n927), .Z(G1350gat));
  OAI21_X1  g727(.A(G190gat), .B1(new_n915), .B2(new_n597), .ZN(new_n929));
  XNOR2_X1  g728(.A(new_n929), .B(KEYINPUT61), .ZN(new_n930));
  NAND3_X1  g729(.A1(new_n917), .A2(new_n216), .A3(new_n701), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(G1351gat));
  NOR2_X1   g731(.A1(new_n825), .A2(new_n671), .ZN(new_n933));
  NOR3_X1   g732(.A1(new_n487), .A2(new_n472), .A3(new_n443), .ZN(new_n934));
  NAND2_X1  g733(.A1(new_n933), .A2(new_n934), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(G197gat), .B1(new_n936), .B2(new_n704), .ZN(new_n937));
  NAND3_X1  g736(.A1(new_n682), .A2(new_n416), .A3(new_n442), .ZN(new_n938));
  XOR2_X1   g737(.A(new_n938), .B(KEYINPUT127), .Z(new_n939));
  NOR2_X1   g738(.A1(new_n902), .A2(new_n939), .ZN(new_n940));
  AND2_X1   g739(.A1(new_n564), .A2(G197gat), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n937), .B1(new_n940), .B2(new_n941), .ZN(G1352gat));
  NOR3_X1   g741(.A1(new_n935), .A2(G204gat), .A3(new_n666), .ZN(new_n943));
  XNOR2_X1  g742(.A(new_n943), .B(KEYINPUT62), .ZN(new_n944));
  NOR3_X1   g743(.A1(new_n902), .A2(new_n666), .A3(new_n939), .ZN(new_n945));
  INV_X1    g744(.A(G204gat), .ZN(new_n946));
  OAI21_X1  g745(.A(new_n944), .B1(new_n945), .B2(new_n946), .ZN(G1353gat));
  NAND3_X1  g746(.A1(new_n936), .A2(new_n310), .A3(new_n637), .ZN(new_n948));
  NOR2_X1   g747(.A1(new_n938), .A2(new_n636), .ZN(new_n949));
  INV_X1    g748(.A(new_n949), .ZN(new_n950));
  OAI21_X1  g749(.A(G211gat), .B1(new_n902), .B2(new_n950), .ZN(new_n951));
  INV_X1    g750(.A(KEYINPUT63), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NOR2_X1   g752(.A1(new_n951), .A2(new_n952), .ZN(new_n954));
  OAI21_X1  g753(.A(new_n948), .B1(new_n953), .B2(new_n954), .ZN(G1354gat));
  NAND3_X1  g754(.A1(new_n936), .A2(new_n311), .A3(new_n701), .ZN(new_n956));
  NOR3_X1   g755(.A1(new_n902), .A2(new_n597), .A3(new_n939), .ZN(new_n957));
  OAI21_X1  g756(.A(new_n956), .B1(new_n957), .B2(new_n311), .ZN(G1355gat));
endmodule


