//Secret key is'1 0 1 0 1 1 1 1 0 0 1 1 0 1 0 0 1 0 1 1 1 0 0 1 1 0 0 1 1 0 1 0 1 1 0 0 0 0 1 1 1 1 0 1 0 0 0 1 1 1 0 0 1 0 1 0 0 1 1 0 1 1 1 1 1 1 1 1 1 1 1 0 1 0 0 0 1 0 1 1 1 1 0 0 0 0 1 0 0 0 1 1 0 0 1 1 0 1 0 0 0 0 1 0 1 1 1 1 0 0 1 1 0 0 1 0 0 1 1 0 0 1 1 1 1 1 1 1' ..
// Benchmark "locked_locked_c1908" written by ABC on Sat Dec 16 05:26:56 2023

module locked_locked_c1908 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G101, G104, G107, G110, G113, G116, G119, G122, G125, G128,
    G131, G134, G137, G140, G143, G146, G210, G214, G217, G221, G224, G227,
    G234, G237, G469, G472, G475, G478, G898, G900, G902, G952, G953,
    G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36, G39,
    G42, G75, G51, G54, G60, G63, G66, G69, G72, G57  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G101, G104, G107, G110, G113, G116,
    G119, G122, G125, G128, G131, G134, G137, G140, G143, G146, G210, G214,
    G217, G221, G224, G227, G234, G237, G469, G472, G475, G478, G898, G900,
    G902, G952, G953;
  output G3, G6, G9, G12, G30, G45, G48, G15, G18, G21, G24, G27, G33, G36,
    G39, G42, G75, G51, G54, G60, G63, G66, G69, G72, G57;
  wire new_n187, new_n188, new_n189, new_n190, new_n191, new_n192, new_n193,
    new_n194, new_n195, new_n196, new_n197, new_n198, new_n199, new_n200,
    new_n201, new_n202, new_n203, new_n204, new_n205, new_n206, new_n207,
    new_n208, new_n209, new_n210, new_n211, new_n212, new_n213, new_n214,
    new_n215, new_n216, new_n217, new_n218, new_n219, new_n220, new_n221,
    new_n222, new_n223, new_n224, new_n225, new_n226, new_n227, new_n228,
    new_n229, new_n230, new_n231, new_n232, new_n233, new_n234, new_n235,
    new_n236, new_n237, new_n238, new_n239, new_n240, new_n241, new_n242,
    new_n243, new_n244, new_n245, new_n246, new_n247, new_n248, new_n249,
    new_n250, new_n251, new_n252, new_n253, new_n254, new_n255, new_n256,
    new_n257, new_n258, new_n259, new_n260, new_n261, new_n262, new_n263,
    new_n264, new_n265, new_n266, new_n267, new_n268, new_n269, new_n270,
    new_n271, new_n272, new_n273, new_n274, new_n275, new_n276, new_n277,
    new_n278, new_n279, new_n280, new_n281, new_n282, new_n283, new_n284,
    new_n285, new_n286, new_n287, new_n288, new_n289, new_n290, new_n291,
    new_n292, new_n293, new_n294, new_n295, new_n296, new_n297, new_n298,
    new_n299, new_n300, new_n301, new_n302, new_n303, new_n304, new_n305,
    new_n306, new_n307, new_n308, new_n309, new_n310, new_n311, new_n312,
    new_n313, new_n314, new_n315, new_n316, new_n317, new_n318, new_n319,
    new_n320, new_n321, new_n322, new_n323, new_n324, new_n325, new_n326,
    new_n327, new_n328, new_n329, new_n330, new_n331, new_n332, new_n333,
    new_n334, new_n335, new_n336, new_n337, new_n338, new_n339, new_n340,
    new_n341, new_n342, new_n343, new_n344, new_n345, new_n346, new_n347,
    new_n348, new_n349, new_n350, new_n351, new_n352, new_n353, new_n354,
    new_n355, new_n356, new_n357, new_n358, new_n359, new_n360, new_n361,
    new_n362, new_n363, new_n364, new_n365, new_n366, new_n367, new_n368,
    new_n369, new_n370, new_n371, new_n372, new_n373, new_n374, new_n375,
    new_n376, new_n377, new_n378, new_n379, new_n380, new_n381, new_n382,
    new_n383, new_n384, new_n385, new_n386, new_n387, new_n388, new_n389,
    new_n390, new_n391, new_n392, new_n393, new_n394, new_n395, new_n396,
    new_n397, new_n398, new_n399, new_n400, new_n401, new_n402, new_n403,
    new_n404, new_n405, new_n406, new_n407, new_n408, new_n409, new_n410,
    new_n411, new_n412, new_n413, new_n414, new_n415, new_n416, new_n417,
    new_n418, new_n419, new_n420, new_n421, new_n422, new_n423, new_n424,
    new_n425, new_n426, new_n427, new_n428, new_n429, new_n430, new_n431,
    new_n432, new_n433, new_n434, new_n435, new_n436, new_n437, new_n438,
    new_n439, new_n440, new_n441, new_n442, new_n443, new_n444, new_n445,
    new_n446, new_n447, new_n448, new_n449, new_n450, new_n451, new_n452,
    new_n453, new_n454, new_n455, new_n456, new_n457, new_n458, new_n459,
    new_n460, new_n461, new_n462, new_n463, new_n464, new_n465, new_n466,
    new_n467, new_n468, new_n469, new_n470, new_n471, new_n472, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n482, new_n483, new_n484, new_n485, new_n486, new_n487,
    new_n488, new_n489, new_n490, new_n491, new_n492, new_n493, new_n494,
    new_n495, new_n496, new_n497, new_n498, new_n499, new_n500, new_n501,
    new_n502, new_n503, new_n504, new_n505, new_n506, new_n507, new_n508,
    new_n509, new_n510, new_n511, new_n512, new_n513, new_n514, new_n515,
    new_n516, new_n517, new_n518, new_n519, new_n520, new_n521, new_n522,
    new_n523, new_n524, new_n525, new_n526, new_n527, new_n528, new_n529,
    new_n530, new_n531, new_n532, new_n533, new_n534, new_n535, new_n536,
    new_n537, new_n538, new_n539, new_n540, new_n541, new_n542, new_n543,
    new_n544, new_n545, new_n546, new_n547, new_n548, new_n549, new_n550,
    new_n551, new_n552, new_n553, new_n554, new_n555, new_n556, new_n557,
    new_n558, new_n559, new_n560, new_n561, new_n562, new_n563, new_n564,
    new_n565, new_n566, new_n567, new_n568, new_n569, new_n570, new_n571,
    new_n572, new_n573, new_n574, new_n575, new_n576, new_n577, new_n578,
    new_n579, new_n580, new_n581, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n614, new_n615,
    new_n616, new_n617, new_n618, new_n619, new_n620, new_n621, new_n622,
    new_n623, new_n625, new_n626, new_n627, new_n628, new_n629, new_n630,
    new_n631, new_n632, new_n633, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n639, new_n640, new_n641, new_n643, new_n644, new_n645,
    new_n646, new_n647, new_n648, new_n649, new_n650, new_n651, new_n652,
    new_n653, new_n654, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n664, new_n665, new_n666, new_n667,
    new_n668, new_n669, new_n670, new_n671, new_n672, new_n673, new_n674,
    new_n675, new_n676, new_n677, new_n678, new_n680, new_n681, new_n682,
    new_n684, new_n685, new_n686, new_n687, new_n688, new_n689, new_n690,
    new_n692, new_n693, new_n694, new_n696, new_n697, new_n698, new_n699,
    new_n700, new_n701, new_n703, new_n704, new_n705, new_n706, new_n707,
    new_n708, new_n709, new_n710, new_n711, new_n712, new_n714, new_n715,
    new_n716, new_n717, new_n718, new_n719, new_n720, new_n721, new_n722,
    new_n723, new_n724, new_n725, new_n726, new_n727, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n747, new_n749, new_n750, new_n751, new_n752, new_n753,
    new_n754, new_n755, new_n756, new_n757, new_n758, new_n759, new_n760,
    new_n761, new_n762, new_n763, new_n764, new_n765, new_n766, new_n767,
    new_n768, new_n769, new_n770, new_n771, new_n772, new_n773, new_n774,
    new_n775, new_n776, new_n777, new_n779, new_n780, new_n781, new_n782,
    new_n783, new_n784, new_n785, new_n787, new_n788, new_n789, new_n790,
    new_n791, new_n792, new_n793, new_n794, new_n795, new_n796, new_n797,
    new_n798, new_n799, new_n800, new_n801, new_n802, new_n803, new_n804,
    new_n805, new_n806, new_n807, new_n808, new_n809, new_n810, new_n811,
    new_n812, new_n813, new_n814, new_n815, new_n816, new_n817, new_n818,
    new_n819, new_n820, new_n821, new_n822, new_n823, new_n824, new_n825,
    new_n826, new_n827, new_n828, new_n829, new_n830, new_n831, new_n832,
    new_n833, new_n834, new_n835, new_n836, new_n837, new_n838, new_n839,
    new_n840, new_n841, new_n842, new_n843, new_n844, new_n845, new_n846,
    new_n847, new_n848, new_n849, new_n850, new_n851, new_n852, new_n853,
    new_n854, new_n855, new_n856, new_n857, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n867,
    new_n868, new_n869, new_n870, new_n871, new_n872, new_n873, new_n874,
    new_n875, new_n876, new_n877, new_n878, new_n879, new_n880, new_n881,
    new_n882, new_n883, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n900, new_n901, new_n902, new_n903, new_n904,
    new_n905, new_n906, new_n908, new_n909, new_n910, new_n911, new_n913,
    new_n914, new_n915, new_n916, new_n917, new_n918, new_n919, new_n920,
    new_n921, new_n922, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n941, new_n942, new_n943,
    new_n944, new_n945, new_n947, new_n948, new_n949, new_n950, new_n951,
    new_n952, new_n953, new_n954, new_n955, new_n956, new_n957, new_n958,
    new_n959, new_n960, new_n961, new_n962, new_n963, new_n964, new_n965,
    new_n966, new_n967, new_n968, new_n970, new_n971, new_n972, new_n973,
    new_n974, new_n975, new_n976, new_n977, new_n978, new_n979, new_n980;
  INV_X1    g000(.A(G475), .ZN(new_n187));
  INV_X1    g001(.A(G140), .ZN(new_n188));
  NAND2_X1  g002(.A1(new_n188), .A2(G125), .ZN(new_n189));
  INV_X1    g003(.A(G125), .ZN(new_n190));
  NAND2_X1  g004(.A1(new_n190), .A2(G140), .ZN(new_n191));
  NAND3_X1  g005(.A1(new_n189), .A2(new_n191), .A3(KEYINPUT16), .ZN(new_n192));
  OR3_X1    g006(.A1(new_n190), .A2(KEYINPUT16), .A3(G140), .ZN(new_n193));
  NAND2_X1  g007(.A1(new_n192), .A2(new_n193), .ZN(new_n194));
  INV_X1    g008(.A(G146), .ZN(new_n195));
  NAND2_X1  g009(.A1(new_n194), .A2(new_n195), .ZN(new_n196));
  NAND3_X1  g010(.A1(new_n192), .A2(new_n193), .A3(G146), .ZN(new_n197));
  NAND3_X1  g011(.A1(new_n196), .A2(KEYINPUT72), .A3(new_n197), .ZN(new_n198));
  INV_X1    g012(.A(KEYINPUT72), .ZN(new_n199));
  NAND3_X1  g013(.A1(new_n194), .A2(new_n199), .A3(new_n195), .ZN(new_n200));
  NAND2_X1  g014(.A1(new_n198), .A2(new_n200), .ZN(new_n201));
  INV_X1    g015(.A(G237), .ZN(new_n202));
  INV_X1    g016(.A(G953), .ZN(new_n203));
  NAND3_X1  g017(.A1(new_n202), .A2(new_n203), .A3(G214), .ZN(new_n204));
  INV_X1    g018(.A(G143), .ZN(new_n205));
  NAND2_X1  g019(.A1(new_n204), .A2(new_n205), .ZN(new_n206));
  NOR2_X1   g020(.A1(G237), .A2(G953), .ZN(new_n207));
  NAND3_X1  g021(.A1(new_n207), .A2(G143), .A3(G214), .ZN(new_n208));
  NAND2_X1  g022(.A1(new_n206), .A2(new_n208), .ZN(new_n209));
  NAND2_X1  g023(.A1(new_n209), .A2(G131), .ZN(new_n210));
  NAND2_X1  g024(.A1(new_n210), .A2(KEYINPUT86), .ZN(new_n211));
  INV_X1    g025(.A(KEYINPUT86), .ZN(new_n212));
  NAND3_X1  g026(.A1(new_n209), .A2(new_n212), .A3(G131), .ZN(new_n213));
  NAND3_X1  g027(.A1(new_n211), .A2(KEYINPUT17), .A3(new_n213), .ZN(new_n214));
  INV_X1    g028(.A(G131), .ZN(new_n215));
  NAND3_X1  g029(.A1(new_n206), .A2(new_n215), .A3(new_n208), .ZN(new_n216));
  AOI21_X1  g030(.A(new_n212), .B1(new_n209), .B2(G131), .ZN(new_n217));
  AOI211_X1 g031(.A(KEYINPUT86), .B(new_n215), .C1(new_n206), .C2(new_n208), .ZN(new_n218));
  OAI21_X1  g032(.A(new_n216), .B1(new_n217), .B2(new_n218), .ZN(new_n219));
  OAI211_X1 g033(.A(new_n201), .B(new_n214), .C1(new_n219), .C2(KEYINPUT17), .ZN(new_n220));
  XNOR2_X1  g034(.A(G113), .B(G122), .ZN(new_n221));
  INV_X1    g035(.A(G104), .ZN(new_n222));
  XNOR2_X1  g036(.A(new_n221), .B(new_n222), .ZN(new_n223));
  AND2_X1   g037(.A1(new_n189), .A2(new_n191), .ZN(new_n224));
  OR3_X1    g038(.A1(new_n224), .A2(KEYINPUT85), .A3(new_n195), .ZN(new_n225));
  XNOR2_X1  g039(.A(KEYINPUT66), .B(G146), .ZN(new_n226));
  INV_X1    g040(.A(new_n226), .ZN(new_n227));
  NAND2_X1  g041(.A1(new_n227), .A2(new_n224), .ZN(new_n228));
  OAI21_X1  g042(.A(KEYINPUT85), .B1(new_n224), .B2(new_n195), .ZN(new_n229));
  NAND3_X1  g043(.A1(new_n225), .A2(new_n228), .A3(new_n229), .ZN(new_n230));
  NAND2_X1  g044(.A1(KEYINPUT18), .A2(G131), .ZN(new_n231));
  XNOR2_X1  g045(.A(new_n209), .B(new_n231), .ZN(new_n232));
  NAND2_X1  g046(.A1(new_n230), .A2(new_n232), .ZN(new_n233));
  AND3_X1   g047(.A1(new_n220), .A2(new_n223), .A3(new_n233), .ZN(new_n234));
  AOI21_X1  g048(.A(new_n223), .B1(new_n220), .B2(new_n233), .ZN(new_n235));
  OR2_X1    g049(.A1(new_n234), .A2(new_n235), .ZN(new_n236));
  INV_X1    g050(.A(G902), .ZN(new_n237));
  AOI21_X1  g051(.A(new_n187), .B1(new_n236), .B2(new_n237), .ZN(new_n238));
  NOR2_X1   g052(.A1(G475), .A2(G902), .ZN(new_n239));
  NAND2_X1  g053(.A1(new_n219), .A2(KEYINPUT87), .ZN(new_n240));
  INV_X1    g054(.A(new_n197), .ZN(new_n241));
  XNOR2_X1  g055(.A(KEYINPUT88), .B(KEYINPUT19), .ZN(new_n242));
  INV_X1    g056(.A(KEYINPUT19), .ZN(new_n243));
  NOR2_X1   g057(.A1(new_n243), .A2(KEYINPUT88), .ZN(new_n244));
  MUX2_X1   g058(.A(new_n242), .B(new_n244), .S(new_n224), .Z(new_n245));
  AOI21_X1  g059(.A(new_n241), .B1(new_n245), .B2(new_n227), .ZN(new_n246));
  INV_X1    g060(.A(KEYINPUT87), .ZN(new_n247));
  OAI211_X1 g061(.A(new_n247), .B(new_n216), .C1(new_n217), .C2(new_n218), .ZN(new_n248));
  NAND3_X1  g062(.A1(new_n240), .A2(new_n246), .A3(new_n248), .ZN(new_n249));
  AOI21_X1  g063(.A(new_n223), .B1(new_n249), .B2(new_n233), .ZN(new_n250));
  OAI21_X1  g064(.A(new_n239), .B1(new_n250), .B2(new_n234), .ZN(new_n251));
  NAND2_X1  g065(.A1(new_n251), .A2(KEYINPUT20), .ZN(new_n252));
  INV_X1    g066(.A(KEYINPUT89), .ZN(new_n253));
  NAND2_X1  g067(.A1(new_n252), .A2(new_n253), .ZN(new_n254));
  INV_X1    g068(.A(KEYINPUT20), .ZN(new_n255));
  OAI211_X1 g069(.A(new_n255), .B(new_n239), .C1(new_n250), .C2(new_n234), .ZN(new_n256));
  NAND2_X1  g070(.A1(new_n254), .A2(new_n256), .ZN(new_n257));
  NOR3_X1   g071(.A1(new_n251), .A2(KEYINPUT89), .A3(KEYINPUT20), .ZN(new_n258));
  INV_X1    g072(.A(new_n258), .ZN(new_n259));
  AOI21_X1  g073(.A(new_n238), .B1(new_n257), .B2(new_n259), .ZN(new_n260));
  XNOR2_X1  g074(.A(G128), .B(G143), .ZN(new_n261));
  INV_X1    g075(.A(G134), .ZN(new_n262));
  XNOR2_X1  g076(.A(new_n261), .B(new_n262), .ZN(new_n263));
  XNOR2_X1  g077(.A(G116), .B(G122), .ZN(new_n264));
  INV_X1    g078(.A(KEYINPUT14), .ZN(new_n265));
  NAND2_X1  g079(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  INV_X1    g080(.A(G116), .ZN(new_n267));
  NAND3_X1  g081(.A1(new_n267), .A2(KEYINPUT14), .A3(G122), .ZN(new_n268));
  NAND3_X1  g082(.A1(new_n266), .A2(G107), .A3(new_n268), .ZN(new_n269));
  INV_X1    g083(.A(G107), .ZN(new_n270));
  NAND2_X1  g084(.A1(new_n264), .A2(new_n270), .ZN(new_n271));
  NAND3_X1  g085(.A1(new_n263), .A2(new_n269), .A3(new_n271), .ZN(new_n272));
  XNOR2_X1  g086(.A(new_n272), .B(KEYINPUT90), .ZN(new_n273));
  NAND2_X1  g087(.A1(new_n261), .A2(KEYINPUT13), .ZN(new_n274));
  NAND2_X1  g088(.A1(new_n205), .A2(G128), .ZN(new_n275));
  OAI211_X1 g089(.A(new_n274), .B(G134), .C1(KEYINPUT13), .C2(new_n275), .ZN(new_n276));
  XNOR2_X1  g090(.A(new_n264), .B(new_n270), .ZN(new_n277));
  NAND2_X1  g091(.A1(new_n261), .A2(new_n262), .ZN(new_n278));
  NAND3_X1  g092(.A1(new_n276), .A2(new_n277), .A3(new_n278), .ZN(new_n279));
  NAND2_X1  g093(.A1(new_n273), .A2(new_n279), .ZN(new_n280));
  XOR2_X1   g094(.A(KEYINPUT9), .B(G234), .Z(new_n281));
  INV_X1    g095(.A(new_n281), .ZN(new_n282));
  INV_X1    g096(.A(G217), .ZN(new_n283));
  NOR3_X1   g097(.A1(new_n282), .A2(new_n283), .A3(G953), .ZN(new_n284));
  INV_X1    g098(.A(new_n284), .ZN(new_n285));
  NAND2_X1  g099(.A1(new_n280), .A2(new_n285), .ZN(new_n286));
  NAND3_X1  g100(.A1(new_n273), .A2(new_n279), .A3(new_n284), .ZN(new_n287));
  AOI21_X1  g101(.A(G902), .B1(new_n286), .B2(new_n287), .ZN(new_n288));
  INV_X1    g102(.A(G478), .ZN(new_n289));
  NOR2_X1   g103(.A1(new_n289), .A2(KEYINPUT15), .ZN(new_n290));
  INV_X1    g104(.A(new_n290), .ZN(new_n291));
  XNOR2_X1  g105(.A(new_n288), .B(new_n291), .ZN(new_n292));
  INV_X1    g106(.A(new_n292), .ZN(new_n293));
  NAND2_X1  g107(.A1(new_n260), .A2(new_n293), .ZN(new_n294));
  INV_X1    g108(.A(new_n294), .ZN(new_n295));
  OAI21_X1  g109(.A(G214), .B1(G237), .B2(G902), .ZN(new_n296));
  INV_X1    g110(.A(new_n296), .ZN(new_n297));
  NAND2_X1  g111(.A1(G234), .A2(G237), .ZN(new_n298));
  AND3_X1   g112(.A1(new_n298), .A2(G952), .A3(new_n203), .ZN(new_n299));
  XNOR2_X1  g113(.A(KEYINPUT21), .B(G898), .ZN(new_n300));
  XOR2_X1   g114(.A(new_n300), .B(KEYINPUT91), .Z(new_n301));
  INV_X1    g115(.A(new_n301), .ZN(new_n302));
  AND3_X1   g116(.A1(new_n298), .A2(G902), .A3(G953), .ZN(new_n303));
  AOI21_X1  g117(.A(new_n299), .B1(new_n302), .B2(new_n303), .ZN(new_n304));
  AND2_X1   g118(.A1(KEYINPUT0), .A2(G128), .ZN(new_n305));
  NOR2_X1   g119(.A1(new_n195), .A2(G143), .ZN(new_n306));
  INV_X1    g120(.A(new_n306), .ZN(new_n307));
  OAI211_X1 g121(.A(new_n305), .B(new_n307), .C1(new_n226), .C2(new_n205), .ZN(new_n308));
  INV_X1    g122(.A(KEYINPUT67), .ZN(new_n309));
  NAND2_X1  g123(.A1(new_n308), .A2(new_n309), .ZN(new_n310));
  NAND2_X1  g124(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n311));
  INV_X1    g125(.A(KEYINPUT66), .ZN(new_n312));
  NAND2_X1  g126(.A1(new_n312), .A2(G146), .ZN(new_n313));
  NAND3_X1  g127(.A1(new_n311), .A2(new_n313), .A3(new_n205), .ZN(new_n314));
  NAND2_X1  g128(.A1(new_n195), .A2(G143), .ZN(new_n315));
  NAND2_X1  g129(.A1(new_n314), .A2(new_n315), .ZN(new_n316));
  NOR2_X1   g130(.A1(KEYINPUT0), .A2(G128), .ZN(new_n317));
  AOI21_X1  g131(.A(new_n305), .B1(KEYINPUT65), .B2(new_n317), .ZN(new_n318));
  OR2_X1    g132(.A1(new_n317), .A2(KEYINPUT65), .ZN(new_n319));
  NAND3_X1  g133(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NOR2_X1   g134(.A1(new_n312), .A2(G146), .ZN(new_n321));
  NOR2_X1   g135(.A1(new_n195), .A2(KEYINPUT66), .ZN(new_n322));
  OAI21_X1  g136(.A(G143), .B1(new_n321), .B2(new_n322), .ZN(new_n323));
  NAND4_X1  g137(.A1(new_n323), .A2(KEYINPUT67), .A3(new_n305), .A4(new_n307), .ZN(new_n324));
  NAND3_X1  g138(.A1(new_n310), .A2(new_n320), .A3(new_n324), .ZN(new_n325));
  NAND2_X1  g139(.A1(new_n325), .A2(G125), .ZN(new_n326));
  INV_X1    g140(.A(G128), .ZN(new_n327));
  NOR2_X1   g141(.A1(new_n327), .A2(KEYINPUT1), .ZN(new_n328));
  NAND3_X1  g142(.A1(new_n323), .A2(new_n307), .A3(new_n328), .ZN(new_n329));
  AOI21_X1  g143(.A(new_n327), .B1(new_n323), .B2(KEYINPUT1), .ZN(new_n330));
  INV_X1    g144(.A(new_n316), .ZN(new_n331));
  OAI211_X1 g145(.A(new_n190), .B(new_n329), .C1(new_n330), .C2(new_n331), .ZN(new_n332));
  NAND2_X1  g146(.A1(new_n326), .A2(new_n332), .ZN(new_n333));
  NAND2_X1  g147(.A1(new_n203), .A2(G224), .ZN(new_n334));
  XOR2_X1   g148(.A(new_n334), .B(KEYINPUT82), .Z(new_n335));
  INV_X1    g149(.A(new_n335), .ZN(new_n336));
  XNOR2_X1  g150(.A(new_n333), .B(new_n336), .ZN(new_n337));
  NAND2_X1  g151(.A1(new_n222), .A2(KEYINPUT78), .ZN(new_n338));
  INV_X1    g152(.A(KEYINPUT78), .ZN(new_n339));
  NAND2_X1  g153(.A1(new_n339), .A2(G104), .ZN(new_n340));
  NAND3_X1  g154(.A1(new_n338), .A2(new_n340), .A3(new_n270), .ZN(new_n341));
  NAND2_X1  g155(.A1(new_n341), .A2(KEYINPUT3), .ZN(new_n342));
  NAND2_X1  g156(.A1(new_n338), .A2(new_n340), .ZN(new_n343));
  NAND2_X1  g157(.A1(new_n343), .A2(G107), .ZN(new_n344));
  OR3_X1    g158(.A1(new_n222), .A2(KEYINPUT3), .A3(G107), .ZN(new_n345));
  NAND3_X1  g159(.A1(new_n342), .A2(new_n344), .A3(new_n345), .ZN(new_n346));
  NAND2_X1  g160(.A1(new_n346), .A2(G101), .ZN(new_n347));
  INV_X1    g161(.A(G101), .ZN(new_n348));
  NAND4_X1  g162(.A1(new_n342), .A2(new_n344), .A3(new_n348), .A4(new_n345), .ZN(new_n349));
  NAND3_X1  g163(.A1(new_n347), .A2(KEYINPUT4), .A3(new_n349), .ZN(new_n350));
  XOR2_X1   g164(.A(KEYINPUT2), .B(G113), .Z(new_n351));
  XNOR2_X1  g165(.A(G116), .B(G119), .ZN(new_n352));
  NAND2_X1  g166(.A1(new_n351), .A2(new_n352), .ZN(new_n353));
  XNOR2_X1  g167(.A(KEYINPUT2), .B(G113), .ZN(new_n354));
  NOR2_X1   g168(.A1(new_n267), .A2(G119), .ZN(new_n355));
  INV_X1    g169(.A(G119), .ZN(new_n356));
  NOR2_X1   g170(.A1(new_n356), .A2(G116), .ZN(new_n357));
  OAI21_X1  g171(.A(new_n354), .B1(new_n355), .B2(new_n357), .ZN(new_n358));
  AND3_X1   g172(.A1(new_n353), .A2(new_n358), .A3(KEYINPUT70), .ZN(new_n359));
  AOI21_X1  g173(.A(KEYINPUT70), .B1(new_n353), .B2(new_n358), .ZN(new_n360));
  NOR2_X1   g174(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g175(.A(KEYINPUT4), .ZN(new_n362));
  NAND3_X1  g176(.A1(new_n346), .A2(new_n362), .A3(G101), .ZN(new_n363));
  NAND3_X1  g177(.A1(new_n350), .A2(new_n361), .A3(new_n363), .ZN(new_n364));
  NAND2_X1  g178(.A1(new_n222), .A2(G107), .ZN(new_n365));
  NAND3_X1  g179(.A1(new_n341), .A2(KEYINPUT79), .A3(new_n365), .ZN(new_n366));
  OR2_X1    g180(.A1(new_n365), .A2(KEYINPUT79), .ZN(new_n367));
  NAND3_X1  g181(.A1(new_n366), .A2(G101), .A3(new_n367), .ZN(new_n368));
  NAND2_X1  g182(.A1(new_n368), .A2(new_n349), .ZN(new_n369));
  INV_X1    g183(.A(new_n369), .ZN(new_n370));
  NAND2_X1  g184(.A1(new_n352), .A2(KEYINPUT5), .ZN(new_n371));
  INV_X1    g185(.A(G113), .ZN(new_n372));
  INV_X1    g186(.A(KEYINPUT5), .ZN(new_n373));
  AOI21_X1  g187(.A(new_n372), .B1(new_n355), .B2(new_n373), .ZN(new_n374));
  AOI22_X1  g188(.A1(new_n371), .A2(new_n374), .B1(new_n351), .B2(new_n352), .ZN(new_n375));
  NAND2_X1  g189(.A1(new_n370), .A2(new_n375), .ZN(new_n376));
  NAND2_X1  g190(.A1(new_n364), .A2(new_n376), .ZN(new_n377));
  XOR2_X1   g191(.A(G110), .B(G122), .Z(new_n378));
  NAND2_X1  g192(.A1(new_n377), .A2(new_n378), .ZN(new_n379));
  INV_X1    g193(.A(new_n378), .ZN(new_n380));
  NAND3_X1  g194(.A1(new_n364), .A2(new_n380), .A3(new_n376), .ZN(new_n381));
  NAND3_X1  g195(.A1(new_n379), .A2(KEYINPUT6), .A3(new_n381), .ZN(new_n382));
  AOI21_X1  g196(.A(new_n380), .B1(new_n364), .B2(new_n376), .ZN(new_n383));
  INV_X1    g197(.A(KEYINPUT81), .ZN(new_n384));
  INV_X1    g198(.A(KEYINPUT6), .ZN(new_n385));
  AND3_X1   g199(.A1(new_n383), .A2(new_n384), .A3(new_n385), .ZN(new_n386));
  AOI21_X1  g200(.A(new_n384), .B1(new_n383), .B2(new_n385), .ZN(new_n387));
  OAI211_X1 g201(.A(new_n337), .B(new_n382), .C1(new_n386), .C2(new_n387), .ZN(new_n388));
  NAND2_X1  g202(.A1(new_n333), .A2(new_n336), .ZN(new_n389));
  INV_X1    g203(.A(KEYINPUT7), .ZN(new_n390));
  NAND2_X1  g204(.A1(new_n333), .A2(new_n390), .ZN(new_n391));
  NAND4_X1  g205(.A1(new_n326), .A2(KEYINPUT7), .A3(new_n335), .A4(new_n332), .ZN(new_n392));
  NAND2_X1  g206(.A1(new_n369), .A2(new_n375), .ZN(new_n393));
  NAND2_X1  g207(.A1(new_n356), .A2(G116), .ZN(new_n394));
  OAI211_X1 g208(.A(KEYINPUT83), .B(G113), .C1(new_n394), .C2(KEYINPUT5), .ZN(new_n395));
  NAND2_X1  g209(.A1(new_n371), .A2(new_n395), .ZN(new_n396));
  NOR2_X1   g210(.A1(new_n374), .A2(KEYINPUT83), .ZN(new_n397));
  OAI21_X1  g211(.A(new_n353), .B1(new_n396), .B2(new_n397), .ZN(new_n398));
  NAND3_X1  g212(.A1(new_n398), .A2(new_n349), .A3(new_n368), .ZN(new_n399));
  XOR2_X1   g213(.A(new_n378), .B(KEYINPUT8), .Z(new_n400));
  NAND3_X1  g214(.A1(new_n393), .A2(new_n399), .A3(new_n400), .ZN(new_n401));
  NAND4_X1  g215(.A1(new_n389), .A2(new_n391), .A3(new_n392), .A4(new_n401), .ZN(new_n402));
  INV_X1    g216(.A(KEYINPUT84), .ZN(new_n403));
  NAND2_X1  g217(.A1(new_n402), .A2(new_n403), .ZN(new_n404));
  AND2_X1   g218(.A1(new_n392), .A2(new_n401), .ZN(new_n405));
  NAND4_X1  g219(.A1(new_n405), .A2(KEYINPUT84), .A3(new_n389), .A4(new_n391), .ZN(new_n406));
  NAND3_X1  g220(.A1(new_n404), .A2(new_n406), .A3(new_n381), .ZN(new_n407));
  NAND3_X1  g221(.A1(new_n388), .A2(new_n407), .A3(new_n237), .ZN(new_n408));
  OAI21_X1  g222(.A(G210), .B1(G237), .B2(G902), .ZN(new_n409));
  INV_X1    g223(.A(new_n409), .ZN(new_n410));
  NAND2_X1  g224(.A1(new_n408), .A2(new_n410), .ZN(new_n411));
  NAND4_X1  g225(.A1(new_n388), .A2(new_n407), .A3(new_n237), .A4(new_n409), .ZN(new_n412));
  AOI211_X1 g226(.A(new_n297), .B(new_n304), .C1(new_n411), .C2(new_n412), .ZN(new_n413));
  OAI21_X1  g227(.A(G221), .B1(new_n282), .B2(G902), .ZN(new_n414));
  INV_X1    g228(.A(new_n414), .ZN(new_n415));
  INV_X1    g229(.A(new_n325), .ZN(new_n416));
  NAND3_X1  g230(.A1(new_n350), .A2(new_n416), .A3(new_n363), .ZN(new_n417));
  OAI21_X1  g231(.A(new_n329), .B1(new_n330), .B2(new_n331), .ZN(new_n418));
  NAND3_X1  g232(.A1(new_n370), .A2(KEYINPUT10), .A3(new_n418), .ZN(new_n419));
  INV_X1    g233(.A(KEYINPUT11), .ZN(new_n420));
  OAI21_X1  g234(.A(new_n420), .B1(new_n262), .B2(G137), .ZN(new_n421));
  INV_X1    g235(.A(G137), .ZN(new_n422));
  NAND3_X1  g236(.A1(new_n422), .A2(KEYINPUT11), .A3(G134), .ZN(new_n423));
  NAND2_X1  g237(.A1(new_n262), .A2(G137), .ZN(new_n424));
  NAND3_X1  g238(.A1(new_n421), .A2(new_n423), .A3(new_n424), .ZN(new_n425));
  NAND2_X1  g239(.A1(KEYINPUT68), .A2(G131), .ZN(new_n426));
  INV_X1    g240(.A(new_n426), .ZN(new_n427));
  NAND2_X1  g241(.A1(new_n425), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g242(.A1(new_n421), .A2(new_n423), .A3(new_n426), .A4(new_n424), .ZN(new_n429));
  NAND2_X1  g243(.A1(new_n428), .A2(new_n429), .ZN(new_n430));
  INV_X1    g244(.A(new_n430), .ZN(new_n431));
  AOI21_X1  g245(.A(new_n205), .B1(new_n311), .B2(new_n313), .ZN(new_n432));
  NOR2_X1   g246(.A1(new_n432), .A2(new_n306), .ZN(new_n433));
  AOI21_X1  g247(.A(new_n327), .B1(new_n315), .B2(KEYINPUT1), .ZN(new_n434));
  OAI21_X1  g248(.A(new_n329), .B1(new_n433), .B2(new_n434), .ZN(new_n435));
  NAND3_X1  g249(.A1(new_n435), .A2(new_n368), .A3(new_n349), .ZN(new_n436));
  INV_X1    g250(.A(KEYINPUT10), .ZN(new_n437));
  NAND2_X1  g251(.A1(new_n436), .A2(new_n437), .ZN(new_n438));
  NAND4_X1  g252(.A1(new_n417), .A2(new_n419), .A3(new_n431), .A4(new_n438), .ZN(new_n439));
  INV_X1    g253(.A(KEYINPUT1), .ZN(new_n440));
  OAI21_X1  g254(.A(G128), .B1(new_n432), .B2(new_n440), .ZN(new_n441));
  AOI22_X1  g255(.A1(new_n441), .A2(new_n316), .B1(new_n433), .B2(new_n328), .ZN(new_n442));
  NAND2_X1  g256(.A1(new_n369), .A2(new_n442), .ZN(new_n443));
  NAND2_X1  g257(.A1(new_n443), .A2(new_n436), .ZN(new_n444));
  AOI21_X1  g258(.A(KEYINPUT12), .B1(new_n444), .B2(new_n430), .ZN(new_n445));
  INV_X1    g259(.A(KEYINPUT12), .ZN(new_n446));
  AOI211_X1 g260(.A(new_n446), .B(new_n431), .C1(new_n443), .C2(new_n436), .ZN(new_n447));
  OAI21_X1  g261(.A(new_n439), .B1(new_n445), .B2(new_n447), .ZN(new_n448));
  XNOR2_X1  g262(.A(G110), .B(G140), .ZN(new_n449));
  NAND2_X1  g263(.A1(new_n203), .A2(G227), .ZN(new_n450));
  XNOR2_X1  g264(.A(new_n449), .B(new_n450), .ZN(new_n451));
  INV_X1    g265(.A(new_n451), .ZN(new_n452));
  NAND2_X1  g266(.A1(new_n448), .A2(new_n452), .ZN(new_n453));
  NAND3_X1  g267(.A1(new_n417), .A2(new_n419), .A3(new_n438), .ZN(new_n454));
  NAND2_X1  g268(.A1(new_n454), .A2(new_n430), .ZN(new_n455));
  NAND3_X1  g269(.A1(new_n455), .A2(new_n439), .A3(new_n451), .ZN(new_n456));
  NAND2_X1  g270(.A1(new_n453), .A2(new_n456), .ZN(new_n457));
  INV_X1    g271(.A(new_n457), .ZN(new_n458));
  INV_X1    g272(.A(KEYINPUT80), .ZN(new_n459));
  NAND2_X1  g273(.A1(new_n458), .A2(new_n459), .ZN(new_n460));
  NAND2_X1  g274(.A1(new_n457), .A2(KEYINPUT80), .ZN(new_n461));
  NAND3_X1  g275(.A1(new_n460), .A2(G469), .A3(new_n461), .ZN(new_n462));
  INV_X1    g276(.A(G469), .ZN(new_n463));
  NOR2_X1   g277(.A1(new_n445), .A2(new_n447), .ZN(new_n464));
  NAND2_X1  g278(.A1(new_n439), .A2(new_n451), .ZN(new_n465));
  NOR2_X1   g279(.A1(new_n464), .A2(new_n465), .ZN(new_n466));
  AOI21_X1  g280(.A(new_n451), .B1(new_n455), .B2(new_n439), .ZN(new_n467));
  OAI211_X1 g281(.A(new_n463), .B(new_n237), .C1(new_n466), .C2(new_n467), .ZN(new_n468));
  NOR2_X1   g282(.A1(new_n463), .A2(new_n237), .ZN(new_n469));
  INV_X1    g283(.A(new_n469), .ZN(new_n470));
  AND2_X1   g284(.A1(new_n468), .A2(new_n470), .ZN(new_n471));
  AOI21_X1  g285(.A(new_n415), .B1(new_n462), .B2(new_n471), .ZN(new_n472));
  NAND3_X1  g286(.A1(new_n295), .A2(new_n413), .A3(new_n472), .ZN(new_n473));
  NAND2_X1  g287(.A1(new_n207), .A2(G210), .ZN(new_n474));
  XNOR2_X1  g288(.A(new_n474), .B(new_n348), .ZN(new_n475));
  XNOR2_X1  g289(.A(KEYINPUT26), .B(KEYINPUT27), .ZN(new_n476));
  XOR2_X1   g290(.A(new_n475), .B(new_n476), .Z(new_n477));
  INV_X1    g291(.A(new_n361), .ZN(new_n478));
  NAND4_X1  g292(.A1(new_n310), .A2(new_n430), .A3(new_n320), .A4(new_n324), .ZN(new_n479));
  NAND2_X1  g293(.A1(new_n425), .A2(new_n215), .ZN(new_n480));
  NAND2_X1  g294(.A1(new_n422), .A2(G134), .ZN(new_n481));
  NAND3_X1  g295(.A1(new_n481), .A2(new_n424), .A3(G131), .ZN(new_n482));
  NAND2_X1  g296(.A1(new_n480), .A2(new_n482), .ZN(new_n483));
  OAI21_X1  g297(.A(KEYINPUT1), .B1(new_n226), .B2(new_n205), .ZN(new_n484));
  AOI22_X1  g298(.A1(new_n484), .A2(G128), .B1(new_n315), .B2(new_n314), .ZN(new_n485));
  AND3_X1   g299(.A1(new_n323), .A2(new_n307), .A3(new_n328), .ZN(new_n486));
  OAI21_X1  g300(.A(new_n483), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND3_X1  g301(.A1(new_n478), .A2(new_n479), .A3(new_n487), .ZN(new_n488));
  NAND2_X1  g302(.A1(new_n488), .A2(KEYINPUT28), .ZN(new_n489));
  AND2_X1   g303(.A1(new_n487), .A2(new_n479), .ZN(new_n490));
  INV_X1    g304(.A(KEYINPUT28), .ZN(new_n491));
  NAND3_X1  g305(.A1(new_n490), .A2(new_n491), .A3(new_n478), .ZN(new_n492));
  NAND2_X1  g306(.A1(new_n489), .A2(new_n492), .ZN(new_n493));
  AND3_X1   g307(.A1(new_n480), .A2(KEYINPUT69), .A3(new_n482), .ZN(new_n494));
  AOI21_X1  g308(.A(KEYINPUT69), .B1(new_n480), .B2(new_n482), .ZN(new_n495));
  NOR3_X1   g309(.A1(new_n442), .A2(new_n494), .A3(new_n495), .ZN(new_n496));
  INV_X1    g310(.A(new_n479), .ZN(new_n497));
  OAI21_X1  g311(.A(new_n361), .B1(new_n496), .B2(new_n497), .ZN(new_n498));
  AOI21_X1  g312(.A(new_n477), .B1(new_n493), .B2(new_n498), .ZN(new_n499));
  XOR2_X1   g313(.A(KEYINPUT64), .B(KEYINPUT30), .Z(new_n500));
  OAI21_X1  g314(.A(new_n500), .B1(new_n496), .B2(new_n497), .ZN(new_n501));
  NAND3_X1  g315(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n479), .ZN(new_n502));
  NAND3_X1  g316(.A1(new_n501), .A2(new_n361), .A3(new_n502), .ZN(new_n503));
  NAND3_X1  g317(.A1(new_n503), .A2(new_n488), .A3(new_n477), .ZN(new_n504));
  INV_X1    g318(.A(KEYINPUT31), .ZN(new_n505));
  NAND2_X1  g319(.A1(new_n504), .A2(new_n505), .ZN(new_n506));
  NAND4_X1  g320(.A1(new_n503), .A2(KEYINPUT31), .A3(new_n488), .A4(new_n477), .ZN(new_n507));
  AOI21_X1  g321(.A(new_n499), .B1(new_n506), .B2(new_n507), .ZN(new_n508));
  NOR3_X1   g322(.A1(new_n508), .A2(G472), .A3(G902), .ZN(new_n509));
  NAND2_X1  g323(.A1(new_n509), .A2(KEYINPUT32), .ZN(new_n510));
  INV_X1    g324(.A(new_n499), .ZN(new_n511));
  INV_X1    g325(.A(new_n488), .ZN(new_n512));
  INV_X1    g326(.A(new_n500), .ZN(new_n513));
  INV_X1    g327(.A(KEYINPUT69), .ZN(new_n514));
  NAND2_X1  g328(.A1(new_n483), .A2(new_n514), .ZN(new_n515));
  NAND3_X1  g329(.A1(new_n480), .A2(KEYINPUT69), .A3(new_n482), .ZN(new_n516));
  NAND3_X1  g330(.A1(new_n418), .A2(new_n515), .A3(new_n516), .ZN(new_n517));
  AOI21_X1  g331(.A(new_n513), .B1(new_n517), .B2(new_n479), .ZN(new_n518));
  AND3_X1   g332(.A1(new_n487), .A2(KEYINPUT30), .A3(new_n479), .ZN(new_n519));
  NOR2_X1   g333(.A1(new_n518), .A2(new_n519), .ZN(new_n520));
  AOI21_X1  g334(.A(new_n512), .B1(new_n520), .B2(new_n361), .ZN(new_n521));
  AOI21_X1  g335(.A(KEYINPUT31), .B1(new_n521), .B2(new_n477), .ZN(new_n522));
  INV_X1    g336(.A(new_n507), .ZN(new_n523));
  OAI21_X1  g337(.A(new_n511), .B1(new_n522), .B2(new_n523), .ZN(new_n524));
  INV_X1    g338(.A(G472), .ZN(new_n525));
  NAND3_X1  g339(.A1(new_n524), .A2(new_n525), .A3(new_n237), .ZN(new_n526));
  INV_X1    g340(.A(KEYINPUT32), .ZN(new_n527));
  NAND2_X1  g341(.A1(new_n526), .A2(new_n527), .ZN(new_n528));
  NOR2_X1   g342(.A1(new_n521), .A2(new_n477), .ZN(new_n529));
  AND3_X1   g343(.A1(new_n493), .A2(new_n498), .A3(new_n477), .ZN(new_n530));
  NOR3_X1   g344(.A1(new_n529), .A2(new_n530), .A3(KEYINPUT29), .ZN(new_n531));
  OR2_X1    g345(.A1(new_n490), .A2(new_n478), .ZN(new_n532));
  NAND2_X1  g346(.A1(new_n493), .A2(new_n532), .ZN(new_n533));
  NAND2_X1  g347(.A1(new_n477), .A2(KEYINPUT29), .ZN(new_n534));
  OAI21_X1  g348(.A(new_n237), .B1(new_n533), .B2(new_n534), .ZN(new_n535));
  OAI21_X1  g349(.A(G472), .B1(new_n531), .B2(new_n535), .ZN(new_n536));
  NAND3_X1  g350(.A1(new_n510), .A2(new_n528), .A3(new_n536), .ZN(new_n537));
  XNOR2_X1  g351(.A(KEYINPUT22), .B(G137), .ZN(new_n538));
  NAND3_X1  g352(.A1(new_n203), .A2(G221), .A3(G234), .ZN(new_n539));
  XNOR2_X1  g353(.A(new_n538), .B(new_n539), .ZN(new_n540));
  XNOR2_X1  g354(.A(new_n540), .B(KEYINPUT75), .ZN(new_n541));
  INV_X1    g355(.A(KEYINPUT71), .ZN(new_n542));
  OAI21_X1  g356(.A(new_n542), .B1(new_n356), .B2(G128), .ZN(new_n543));
  NAND2_X1  g357(.A1(new_n543), .A2(KEYINPUT23), .ZN(new_n544));
  INV_X1    g358(.A(G110), .ZN(new_n545));
  NAND2_X1  g359(.A1(new_n356), .A2(G128), .ZN(new_n546));
  INV_X1    g360(.A(KEYINPUT23), .ZN(new_n547));
  OAI211_X1 g361(.A(new_n542), .B(new_n547), .C1(new_n356), .C2(G128), .ZN(new_n548));
  NAND4_X1  g362(.A1(new_n544), .A2(new_n545), .A3(new_n546), .A4(new_n548), .ZN(new_n549));
  NAND2_X1  g363(.A1(new_n327), .A2(G119), .ZN(new_n550));
  NAND2_X1  g364(.A1(new_n550), .A2(new_n546), .ZN(new_n551));
  XNOR2_X1  g365(.A(KEYINPUT24), .B(G110), .ZN(new_n552));
  NAND2_X1  g366(.A1(new_n551), .A2(new_n552), .ZN(new_n553));
  NAND2_X1  g367(.A1(new_n549), .A2(new_n553), .ZN(new_n554));
  NAND2_X1  g368(.A1(new_n554), .A2(KEYINPUT73), .ZN(new_n555));
  INV_X1    g369(.A(KEYINPUT73), .ZN(new_n556));
  NAND3_X1  g370(.A1(new_n549), .A2(new_n556), .A3(new_n553), .ZN(new_n557));
  NAND4_X1  g371(.A1(new_n555), .A2(new_n197), .A3(new_n557), .A4(new_n228), .ZN(new_n558));
  OR2_X1    g372(.A1(new_n551), .A2(new_n552), .ZN(new_n559));
  NAND3_X1  g373(.A1(new_n544), .A2(new_n546), .A3(new_n548), .ZN(new_n560));
  NAND2_X1  g374(.A1(new_n560), .A2(G110), .ZN(new_n561));
  NAND4_X1  g375(.A1(new_n198), .A2(new_n559), .A3(new_n561), .A4(new_n200), .ZN(new_n562));
  AND3_X1   g376(.A1(new_n558), .A2(KEYINPUT74), .A3(new_n562), .ZN(new_n563));
  AOI21_X1  g377(.A(KEYINPUT74), .B1(new_n558), .B2(new_n562), .ZN(new_n564));
  OAI21_X1  g378(.A(new_n541), .B1(new_n563), .B2(new_n564), .ZN(new_n565));
  NAND3_X1  g379(.A1(new_n558), .A2(new_n562), .A3(new_n540), .ZN(new_n566));
  NAND2_X1  g380(.A1(new_n565), .A2(new_n566), .ZN(new_n567));
  AOI21_X1  g381(.A(new_n283), .B1(G234), .B2(new_n237), .ZN(new_n568));
  NOR3_X1   g382(.A1(new_n567), .A2(G902), .A3(new_n568), .ZN(new_n569));
  NAND3_X1  g383(.A1(new_n565), .A2(new_n237), .A3(new_n566), .ZN(new_n570));
  NAND2_X1  g384(.A1(new_n570), .A2(KEYINPUT76), .ZN(new_n571));
  XNOR2_X1  g385(.A(KEYINPUT77), .B(KEYINPUT25), .ZN(new_n572));
  INV_X1    g386(.A(new_n572), .ZN(new_n573));
  NAND2_X1  g387(.A1(new_n571), .A2(new_n573), .ZN(new_n574));
  INV_X1    g388(.A(KEYINPUT25), .ZN(new_n575));
  OR2_X1    g389(.A1(new_n570), .A2(new_n575), .ZN(new_n576));
  NAND3_X1  g390(.A1(new_n570), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n577));
  NAND3_X1  g391(.A1(new_n574), .A2(new_n576), .A3(new_n577), .ZN(new_n578));
  AOI21_X1  g392(.A(new_n569), .B1(new_n578), .B2(new_n568), .ZN(new_n579));
  NAND2_X1  g393(.A1(new_n537), .A2(new_n579), .ZN(new_n580));
  NOR2_X1   g394(.A1(new_n473), .A2(new_n580), .ZN(new_n581));
  XNOR2_X1  g395(.A(new_n581), .B(new_n348), .ZN(G3));
  OAI21_X1  g396(.A(G472), .B1(new_n508), .B2(G902), .ZN(new_n583));
  AND2_X1   g397(.A1(new_n526), .A2(new_n583), .ZN(new_n584));
  NAND3_X1  g398(.A1(new_n472), .A2(new_n579), .A3(new_n584), .ZN(new_n585));
  XOR2_X1   g399(.A(new_n585), .B(KEYINPUT92), .Z(new_n586));
  NAND2_X1  g400(.A1(new_n286), .A2(new_n287), .ZN(new_n587));
  NAND2_X1  g401(.A1(new_n587), .A2(new_n237), .ZN(new_n588));
  NAND3_X1  g402(.A1(new_n588), .A2(KEYINPUT93), .A3(new_n289), .ZN(new_n589));
  INV_X1    g403(.A(KEYINPUT93), .ZN(new_n590));
  OAI21_X1  g404(.A(new_n590), .B1(new_n288), .B2(G478), .ZN(new_n591));
  NAND2_X1  g405(.A1(new_n589), .A2(new_n591), .ZN(new_n592));
  INV_X1    g406(.A(KEYINPUT33), .ZN(new_n593));
  NAND2_X1  g407(.A1(new_n587), .A2(new_n593), .ZN(new_n594));
  NAND3_X1  g408(.A1(new_n286), .A2(KEYINPUT33), .A3(new_n287), .ZN(new_n595));
  NAND4_X1  g409(.A1(new_n594), .A2(G478), .A3(new_n237), .A4(new_n595), .ZN(new_n596));
  AND2_X1   g410(.A1(new_n592), .A2(new_n596), .ZN(new_n597));
  OAI21_X1  g411(.A(KEYINPUT94), .B1(new_n260), .B2(new_n597), .ZN(new_n598));
  INV_X1    g412(.A(new_n238), .ZN(new_n599));
  INV_X1    g413(.A(new_n256), .ZN(new_n600));
  AOI21_X1  g414(.A(new_n600), .B1(new_n252), .B2(new_n253), .ZN(new_n601));
  OAI21_X1  g415(.A(new_n599), .B1(new_n601), .B2(new_n258), .ZN(new_n602));
  NAND2_X1  g416(.A1(new_n592), .A2(new_n596), .ZN(new_n603));
  INV_X1    g417(.A(KEYINPUT94), .ZN(new_n604));
  NAND3_X1  g418(.A1(new_n602), .A2(new_n603), .A3(new_n604), .ZN(new_n605));
  NAND4_X1  g419(.A1(new_n598), .A2(new_n413), .A3(KEYINPUT95), .A4(new_n605), .ZN(new_n606));
  NAND3_X1  g420(.A1(new_n598), .A2(new_n413), .A3(new_n605), .ZN(new_n607));
  INV_X1    g421(.A(KEYINPUT95), .ZN(new_n608));
  NAND2_X1  g422(.A1(new_n607), .A2(new_n608), .ZN(new_n609));
  AOI21_X1  g423(.A(new_n586), .B1(new_n606), .B2(new_n609), .ZN(new_n610));
  XNOR2_X1  g424(.A(new_n610), .B(KEYINPUT96), .ZN(new_n611));
  XOR2_X1   g425(.A(KEYINPUT34), .B(G104), .Z(new_n612));
  XNOR2_X1  g426(.A(new_n611), .B(new_n612), .ZN(G6));
  NAND2_X1  g427(.A1(new_n252), .A2(new_n256), .ZN(new_n614));
  AND3_X1   g428(.A1(new_n292), .A2(new_n599), .A3(new_n614), .ZN(new_n615));
  NAND3_X1  g429(.A1(new_n413), .A2(KEYINPUT97), .A3(new_n615), .ZN(new_n616));
  NAND2_X1  g430(.A1(new_n411), .A2(new_n412), .ZN(new_n617));
  INV_X1    g431(.A(new_n304), .ZN(new_n618));
  NAND4_X1  g432(.A1(new_n617), .A2(new_n615), .A3(new_n296), .A4(new_n618), .ZN(new_n619));
  INV_X1    g433(.A(KEYINPUT97), .ZN(new_n620));
  NAND2_X1  g434(.A1(new_n619), .A2(new_n620), .ZN(new_n621));
  AOI21_X1  g435(.A(new_n586), .B1(new_n616), .B2(new_n621), .ZN(new_n622));
  XNOR2_X1  g436(.A(KEYINPUT35), .B(G107), .ZN(new_n623));
  XNOR2_X1  g437(.A(new_n622), .B(new_n623), .ZN(G9));
  NOR2_X1   g438(.A1(new_n563), .A2(new_n564), .ZN(new_n625));
  NOR2_X1   g439(.A1(new_n541), .A2(KEYINPUT36), .ZN(new_n626));
  XOR2_X1   g440(.A(new_n625), .B(new_n626), .Z(new_n627));
  NOR2_X1   g441(.A1(new_n568), .A2(G902), .ZN(new_n628));
  NAND2_X1  g442(.A1(new_n627), .A2(new_n628), .ZN(new_n629));
  AND3_X1   g443(.A1(new_n570), .A2(KEYINPUT76), .A3(new_n572), .ZN(new_n630));
  AOI21_X1  g444(.A(new_n572), .B1(new_n570), .B2(KEYINPUT76), .ZN(new_n631));
  NOR2_X1   g445(.A1(new_n570), .A2(new_n575), .ZN(new_n632));
  NOR3_X1   g446(.A1(new_n630), .A2(new_n631), .A3(new_n632), .ZN(new_n633));
  INV_X1    g447(.A(new_n568), .ZN(new_n634));
  OAI21_X1  g448(.A(new_n629), .B1(new_n633), .B2(new_n634), .ZN(new_n635));
  NAND2_X1  g449(.A1(new_n584), .A2(new_n635), .ZN(new_n636));
  INV_X1    g450(.A(KEYINPUT98), .ZN(new_n637));
  NOR2_X1   g451(.A1(new_n636), .A2(new_n637), .ZN(new_n638));
  AOI21_X1  g452(.A(KEYINPUT98), .B1(new_n584), .B2(new_n635), .ZN(new_n639));
  NOR3_X1   g453(.A1(new_n638), .A2(new_n473), .A3(new_n639), .ZN(new_n640));
  XNOR2_X1  g454(.A(KEYINPUT37), .B(G110), .ZN(new_n641));
  XNOR2_X1  g455(.A(new_n640), .B(new_n641), .ZN(G12));
  AND2_X1   g456(.A1(new_n537), .A2(new_n472), .ZN(new_n643));
  AOI21_X1  g457(.A(new_n238), .B1(new_n256), .B2(new_n252), .ZN(new_n644));
  INV_X1    g458(.A(G900), .ZN(new_n645));
  AOI21_X1  g459(.A(new_n299), .B1(new_n303), .B2(new_n645), .ZN(new_n646));
  INV_X1    g460(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g461(.A1(new_n644), .A2(new_n292), .A3(new_n647), .ZN(new_n648));
  XNOR2_X1  g462(.A(new_n648), .B(KEYINPUT99), .ZN(new_n649));
  AOI21_X1  g463(.A(new_n297), .B1(new_n411), .B2(new_n412), .ZN(new_n650));
  INV_X1    g464(.A(new_n650), .ZN(new_n651));
  AOI22_X1  g465(.A1(new_n578), .A2(new_n568), .B1(new_n628), .B2(new_n627), .ZN(new_n652));
  NOR2_X1   g466(.A1(new_n651), .A2(new_n652), .ZN(new_n653));
  NAND3_X1  g467(.A1(new_n643), .A2(new_n649), .A3(new_n653), .ZN(new_n654));
  XNOR2_X1  g468(.A(new_n654), .B(G128), .ZN(G30));
  NOR2_X1   g469(.A1(new_n508), .A2(G902), .ZN(new_n656));
  AOI21_X1  g470(.A(KEYINPUT32), .B1(new_n656), .B2(new_n525), .ZN(new_n657));
  NOR4_X1   g471(.A1(new_n508), .A2(new_n527), .A3(G472), .A4(G902), .ZN(new_n658));
  NOR2_X1   g472(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  INV_X1    g473(.A(new_n504), .ZN(new_n660));
  AOI21_X1  g474(.A(new_n477), .B1(new_n532), .B2(new_n488), .ZN(new_n661));
  OAI21_X1  g475(.A(new_n237), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  NAND2_X1  g476(.A1(new_n662), .A2(G472), .ZN(new_n663));
  AOI21_X1  g477(.A(KEYINPUT101), .B1(new_n659), .B2(new_n663), .ZN(new_n664));
  AND4_X1   g478(.A1(KEYINPUT101), .A2(new_n510), .A3(new_n528), .A4(new_n663), .ZN(new_n665));
  NOR2_X1   g479(.A1(new_n664), .A2(new_n665), .ZN(new_n666));
  XOR2_X1   g480(.A(new_n646), .B(KEYINPUT39), .Z(new_n667));
  NAND2_X1  g481(.A1(new_n472), .A2(new_n667), .ZN(new_n668));
  AOI21_X1  g482(.A(new_n666), .B1(KEYINPUT40), .B2(new_n668), .ZN(new_n669));
  NOR2_X1   g483(.A1(new_n635), .A2(new_n297), .ZN(new_n670));
  NOR2_X1   g484(.A1(new_n668), .A2(KEYINPUT40), .ZN(new_n671));
  NAND2_X1  g485(.A1(new_n257), .A2(new_n259), .ZN(new_n672));
  AOI21_X1  g486(.A(new_n293), .B1(new_n672), .B2(new_n599), .ZN(new_n673));
  INV_X1    g487(.A(new_n673), .ZN(new_n674));
  NOR2_X1   g488(.A1(new_n671), .A2(new_n674), .ZN(new_n675));
  XOR2_X1   g489(.A(KEYINPUT100), .B(KEYINPUT38), .Z(new_n676));
  XNOR2_X1  g490(.A(new_n617), .B(new_n676), .ZN(new_n677));
  NAND4_X1  g491(.A1(new_n669), .A2(new_n670), .A3(new_n675), .A4(new_n677), .ZN(new_n678));
  XNOR2_X1  g492(.A(new_n678), .B(G143), .ZN(G45));
  NAND3_X1  g493(.A1(new_n602), .A2(new_n603), .A3(new_n647), .ZN(new_n680));
  INV_X1    g494(.A(new_n680), .ZN(new_n681));
  NAND3_X1  g495(.A1(new_n643), .A2(new_n653), .A3(new_n681), .ZN(new_n682));
  XNOR2_X1  g496(.A(new_n682), .B(G146), .ZN(G48));
  OAI21_X1  g497(.A(new_n237), .B1(new_n466), .B2(new_n467), .ZN(new_n684));
  NAND2_X1  g498(.A1(new_n684), .A2(G469), .ZN(new_n685));
  AND3_X1   g499(.A1(new_n685), .A2(new_n414), .A3(new_n468), .ZN(new_n686));
  NAND3_X1  g500(.A1(new_n537), .A2(new_n579), .A3(new_n686), .ZN(new_n687));
  AOI21_X1  g501(.A(new_n687), .B1(new_n609), .B2(new_n606), .ZN(new_n688));
  XNOR2_X1  g502(.A(new_n688), .B(KEYINPUT102), .ZN(new_n689));
  XOR2_X1   g503(.A(KEYINPUT41), .B(G113), .Z(new_n690));
  XNOR2_X1  g504(.A(new_n689), .B(new_n690), .ZN(G15));
  NAND2_X1  g505(.A1(new_n616), .A2(new_n621), .ZN(new_n692));
  AND3_X1   g506(.A1(new_n537), .A2(new_n579), .A3(new_n686), .ZN(new_n693));
  NAND2_X1  g507(.A1(new_n692), .A2(new_n693), .ZN(new_n694));
  XNOR2_X1  g508(.A(new_n694), .B(G116), .ZN(G18));
  INV_X1    g509(.A(new_n686), .ZN(new_n696));
  NOR2_X1   g510(.A1(new_n696), .A2(new_n304), .ZN(new_n697));
  NAND2_X1  g511(.A1(new_n653), .A2(new_n697), .ZN(new_n698));
  NAND2_X1  g512(.A1(new_n295), .A2(new_n537), .ZN(new_n699));
  NOR2_X1   g513(.A1(new_n698), .A2(new_n699), .ZN(new_n700));
  XNOR2_X1  g514(.A(KEYINPUT103), .B(G119), .ZN(new_n701));
  XNOR2_X1  g515(.A(new_n700), .B(new_n701), .ZN(G21));
  NOR2_X1   g516(.A1(new_n674), .A2(new_n651), .ZN(new_n703));
  NOR2_X1   g517(.A1(G472), .A2(G902), .ZN(new_n704));
  INV_X1    g518(.A(new_n704), .ZN(new_n705));
  NAND2_X1  g519(.A1(new_n506), .A2(new_n507), .ZN(new_n706));
  INV_X1    g520(.A(new_n477), .ZN(new_n707));
  NAND2_X1  g521(.A1(new_n533), .A2(new_n707), .ZN(new_n708));
  AOI21_X1  g522(.A(new_n705), .B1(new_n706), .B2(new_n708), .ZN(new_n709));
  NAND2_X1  g523(.A1(new_n524), .A2(new_n237), .ZN(new_n710));
  AOI21_X1  g524(.A(new_n709), .B1(new_n710), .B2(G472), .ZN(new_n711));
  NAND4_X1  g525(.A1(new_n703), .A2(new_n697), .A3(new_n579), .A4(new_n711), .ZN(new_n712));
  XNOR2_X1  g526(.A(new_n712), .B(G122), .ZN(G24));
  INV_X1    g527(.A(KEYINPUT104), .ZN(new_n714));
  OAI21_X1  g528(.A(new_n708), .B1(new_n522), .B2(new_n523), .ZN(new_n715));
  NAND2_X1  g529(.A1(new_n715), .A2(new_n704), .ZN(new_n716));
  NAND2_X1  g530(.A1(new_n583), .A2(new_n716), .ZN(new_n717));
  OAI21_X1  g531(.A(new_n714), .B1(new_n652), .B2(new_n717), .ZN(new_n718));
  NAND3_X1  g532(.A1(new_n635), .A2(new_n711), .A3(KEYINPUT104), .ZN(new_n719));
  NAND2_X1  g533(.A1(new_n718), .A2(new_n719), .ZN(new_n720));
  NAND2_X1  g534(.A1(new_n650), .A2(new_n686), .ZN(new_n721));
  NOR2_X1   g535(.A1(new_n721), .A2(new_n680), .ZN(new_n722));
  NAND2_X1  g536(.A1(new_n720), .A2(new_n722), .ZN(new_n723));
  NAND2_X1  g537(.A1(new_n723), .A2(KEYINPUT105), .ZN(new_n724));
  INV_X1    g538(.A(KEYINPUT105), .ZN(new_n725));
  NAND3_X1  g539(.A1(new_n720), .A2(new_n725), .A3(new_n722), .ZN(new_n726));
  NAND2_X1  g540(.A1(new_n724), .A2(new_n726), .ZN(new_n727));
  XNOR2_X1  g541(.A(new_n727), .B(G125), .ZN(G27));
  INV_X1    g542(.A(new_n579), .ZN(new_n729));
  AOI21_X1  g543(.A(new_n729), .B1(new_n659), .B2(new_n536), .ZN(new_n730));
  OAI21_X1  g544(.A(new_n471), .B1(new_n463), .B2(new_n457), .ZN(new_n731));
  NOR2_X1   g545(.A1(new_n415), .A2(new_n297), .ZN(new_n732));
  AND4_X1   g546(.A1(new_n411), .A2(new_n731), .A3(new_n412), .A4(new_n732), .ZN(new_n733));
  NOR2_X1   g547(.A1(new_n680), .A2(KEYINPUT42), .ZN(new_n734));
  AND3_X1   g548(.A1(new_n730), .A2(new_n733), .A3(new_n734), .ZN(new_n735));
  AND2_X1   g549(.A1(new_n733), .A2(new_n681), .ZN(new_n736));
  INV_X1    g550(.A(KEYINPUT106), .ZN(new_n737));
  OAI21_X1  g551(.A(new_n737), .B1(new_n509), .B2(KEYINPUT32), .ZN(new_n738));
  NAND3_X1  g552(.A1(new_n526), .A2(KEYINPUT106), .A3(new_n527), .ZN(new_n739));
  NAND4_X1  g553(.A1(new_n738), .A2(new_n510), .A3(new_n739), .A4(new_n536), .ZN(new_n740));
  AND3_X1   g554(.A1(new_n740), .A2(KEYINPUT107), .A3(new_n579), .ZN(new_n741));
  AOI21_X1  g555(.A(KEYINPUT107), .B1(new_n740), .B2(new_n579), .ZN(new_n742));
  OAI21_X1  g556(.A(new_n736), .B1(new_n741), .B2(new_n742), .ZN(new_n743));
  AOI21_X1  g557(.A(new_n735), .B1(new_n743), .B2(KEYINPUT42), .ZN(new_n744));
  XOR2_X1   g558(.A(KEYINPUT108), .B(G131), .Z(new_n745));
  XNOR2_X1  g559(.A(new_n744), .B(new_n745), .ZN(G33));
  NAND3_X1  g560(.A1(new_n730), .A2(new_n649), .A3(new_n733), .ZN(new_n747));
  XNOR2_X1  g561(.A(new_n747), .B(G134), .ZN(G36));
  INV_X1    g562(.A(KEYINPUT110), .ZN(new_n749));
  XNOR2_X1  g563(.A(new_n457), .B(new_n459), .ZN(new_n750));
  OAI21_X1  g564(.A(G469), .B1(new_n750), .B2(KEYINPUT45), .ZN(new_n751));
  INV_X1    g565(.A(KEYINPUT109), .ZN(new_n752));
  NAND2_X1  g566(.A1(new_n751), .A2(new_n752), .ZN(new_n753));
  OAI211_X1 g567(.A(KEYINPUT109), .B(G469), .C1(new_n750), .C2(KEYINPUT45), .ZN(new_n754));
  NAND2_X1  g568(.A1(new_n458), .A2(KEYINPUT45), .ZN(new_n755));
  NAND3_X1  g569(.A1(new_n753), .A2(new_n754), .A3(new_n755), .ZN(new_n756));
  NAND2_X1  g570(.A1(new_n756), .A2(new_n470), .ZN(new_n757));
  INV_X1    g571(.A(KEYINPUT46), .ZN(new_n758));
  OAI21_X1  g572(.A(new_n749), .B1(new_n757), .B2(new_n758), .ZN(new_n759));
  NAND2_X1  g573(.A1(new_n757), .A2(new_n758), .ZN(new_n760));
  NAND4_X1  g574(.A1(new_n756), .A2(KEYINPUT110), .A3(KEYINPUT46), .A4(new_n470), .ZN(new_n761));
  NAND4_X1  g575(.A1(new_n759), .A2(new_n760), .A3(new_n468), .A4(new_n761), .ZN(new_n762));
  NAND2_X1  g576(.A1(new_n762), .A2(new_n414), .ZN(new_n763));
  INV_X1    g577(.A(new_n763), .ZN(new_n764));
  AND2_X1   g578(.A1(new_n764), .A2(new_n667), .ZN(new_n765));
  NAND3_X1  g579(.A1(new_n411), .A2(new_n296), .A3(new_n412), .ZN(new_n766));
  INV_X1    g580(.A(new_n766), .ZN(new_n767));
  NAND2_X1  g581(.A1(new_n260), .A2(new_n603), .ZN(new_n768));
  XOR2_X1   g582(.A(new_n768), .B(KEYINPUT43), .Z(new_n769));
  INV_X1    g583(.A(new_n584), .ZN(new_n770));
  NAND3_X1  g584(.A1(new_n769), .A2(new_n770), .A3(new_n635), .ZN(new_n771));
  INV_X1    g585(.A(KEYINPUT44), .ZN(new_n772));
  NAND2_X1  g586(.A1(new_n771), .A2(new_n772), .ZN(new_n773));
  XNOR2_X1  g587(.A(new_n773), .B(KEYINPUT111), .ZN(new_n774));
  OR2_X1    g588(.A1(new_n771), .A2(new_n772), .ZN(new_n775));
  NAND4_X1  g589(.A1(new_n765), .A2(new_n767), .A3(new_n774), .A4(new_n775), .ZN(new_n776));
  XOR2_X1   g590(.A(KEYINPUT112), .B(G137), .Z(new_n777));
  XNOR2_X1  g591(.A(new_n776), .B(new_n777), .ZN(G39));
  INV_X1    g592(.A(KEYINPUT47), .ZN(new_n779));
  NAND2_X1  g593(.A1(new_n764), .A2(new_n779), .ZN(new_n780));
  INV_X1    g594(.A(new_n537), .ZN(new_n781));
  AOI21_X1  g595(.A(new_n779), .B1(new_n762), .B2(new_n414), .ZN(new_n782));
  INV_X1    g596(.A(new_n782), .ZN(new_n783));
  NOR3_X1   g597(.A1(new_n680), .A2(new_n579), .A3(new_n766), .ZN(new_n784));
  NAND4_X1  g598(.A1(new_n780), .A2(new_n781), .A3(new_n783), .A4(new_n784), .ZN(new_n785));
  XNOR2_X1  g599(.A(new_n785), .B(G140), .ZN(G42));
  INV_X1    g600(.A(KEYINPUT53), .ZN(new_n787));
  OAI211_X1 g601(.A(new_n643), .B(new_n653), .C1(new_n649), .C2(new_n681), .ZN(new_n788));
  AND4_X1   g602(.A1(new_n414), .A2(new_n673), .A3(new_n650), .A4(new_n647), .ZN(new_n789));
  NAND2_X1  g603(.A1(new_n652), .A2(new_n731), .ZN(new_n790));
  INV_X1    g604(.A(new_n790), .ZN(new_n791));
  OAI211_X1 g605(.A(new_n789), .B(new_n791), .C1(new_n664), .C2(new_n665), .ZN(new_n792));
  AND3_X1   g606(.A1(new_n720), .A2(new_n725), .A3(new_n722), .ZN(new_n793));
  AOI21_X1  g607(.A(new_n725), .B1(new_n720), .B2(new_n722), .ZN(new_n794));
  OAI211_X1 g608(.A(new_n788), .B(new_n792), .C1(new_n793), .C2(new_n794), .ZN(new_n795));
  INV_X1    g609(.A(KEYINPUT52), .ZN(new_n796));
  NAND2_X1  g610(.A1(new_n795), .A2(new_n796), .ZN(new_n797));
  NAND4_X1  g611(.A1(new_n727), .A2(KEYINPUT52), .A3(new_n788), .A4(new_n792), .ZN(new_n798));
  AND2_X1   g612(.A1(new_n797), .A2(new_n798), .ZN(new_n799));
  NAND2_X1  g613(.A1(new_n694), .A2(new_n712), .ZN(new_n800));
  NOR3_X1   g614(.A1(new_n800), .A2(new_n688), .A3(new_n700), .ZN(new_n801));
  NAND2_X1  g615(.A1(new_n602), .A2(new_n603), .ZN(new_n802));
  OAI21_X1  g616(.A(new_n802), .B1(new_n293), .B2(new_n602), .ZN(new_n803));
  NAND2_X1  g617(.A1(new_n803), .A2(new_n413), .ZN(new_n804));
  OAI22_X1  g618(.A1(new_n804), .A2(new_n585), .B1(new_n473), .B2(new_n580), .ZN(new_n805));
  NOR2_X1   g619(.A1(new_n640), .A2(new_n805), .ZN(new_n806));
  NAND3_X1  g620(.A1(new_n720), .A2(new_n681), .A3(new_n733), .ZN(new_n807));
  NAND2_X1  g621(.A1(new_n747), .A2(new_n807), .ZN(new_n808));
  INV_X1    g622(.A(KEYINPUT113), .ZN(new_n809));
  NAND4_X1  g623(.A1(new_n411), .A2(new_n644), .A3(new_n296), .A4(new_n412), .ZN(new_n810));
  NAND2_X1  g624(.A1(new_n293), .A2(new_n647), .ZN(new_n811));
  OAI21_X1  g625(.A(new_n809), .B1(new_n810), .B2(new_n811), .ZN(new_n812));
  NAND2_X1  g626(.A1(new_n812), .A2(new_n635), .ZN(new_n813));
  NAND2_X1  g627(.A1(new_n537), .A2(new_n472), .ZN(new_n814));
  NOR3_X1   g628(.A1(new_n810), .A2(new_n809), .A3(new_n811), .ZN(new_n815));
  NOR3_X1   g629(.A1(new_n813), .A2(new_n814), .A3(new_n815), .ZN(new_n816));
  NOR2_X1   g630(.A1(new_n808), .A2(new_n816), .ZN(new_n817));
  NAND4_X1  g631(.A1(new_n801), .A2(new_n744), .A3(new_n806), .A4(new_n817), .ZN(new_n818));
  OAI21_X1  g632(.A(new_n787), .B1(new_n799), .B2(new_n818), .ZN(new_n819));
  AND2_X1   g633(.A1(new_n744), .A2(new_n817), .ZN(new_n820));
  NAND2_X1  g634(.A1(new_n797), .A2(new_n798), .ZN(new_n821));
  NOR2_X1   g635(.A1(new_n688), .A2(new_n700), .ZN(new_n822));
  AND2_X1   g636(.A1(new_n694), .A2(new_n712), .ZN(new_n823));
  AND3_X1   g637(.A1(new_n822), .A2(new_n823), .A3(new_n806), .ZN(new_n824));
  NAND4_X1  g638(.A1(new_n820), .A2(new_n821), .A3(new_n824), .A4(KEYINPUT53), .ZN(new_n825));
  XNOR2_X1  g639(.A(KEYINPUT114), .B(KEYINPUT54), .ZN(new_n826));
  INV_X1    g640(.A(new_n826), .ZN(new_n827));
  NAND3_X1  g641(.A1(new_n819), .A2(new_n825), .A3(new_n827), .ZN(new_n828));
  NAND2_X1  g642(.A1(new_n828), .A2(KEYINPUT115), .ZN(new_n829));
  NAND2_X1  g643(.A1(new_n819), .A2(new_n825), .ZN(new_n830));
  NAND2_X1  g644(.A1(new_n830), .A2(KEYINPUT54), .ZN(new_n831));
  INV_X1    g645(.A(KEYINPUT115), .ZN(new_n832));
  NAND4_X1  g646(.A1(new_n819), .A2(new_n825), .A3(new_n832), .A4(new_n827), .ZN(new_n833));
  NAND3_X1  g647(.A1(new_n829), .A2(new_n831), .A3(new_n833), .ZN(new_n834));
  INV_X1    g648(.A(new_n299), .ZN(new_n835));
  NOR3_X1   g649(.A1(new_n729), .A2(new_n835), .A3(new_n717), .ZN(new_n836));
  AND2_X1   g650(.A1(new_n769), .A2(new_n836), .ZN(new_n837));
  INV_X1    g651(.A(new_n837), .ZN(new_n838));
  NOR2_X1   g652(.A1(new_n838), .A2(new_n721), .ZN(new_n839));
  OR2_X1    g653(.A1(new_n834), .A2(new_n839), .ZN(new_n840));
  INV_X1    g654(.A(KEYINPUT51), .ZN(new_n841));
  NOR2_X1   g655(.A1(new_n838), .A2(new_n766), .ZN(new_n842));
  INV_X1    g656(.A(new_n842), .ZN(new_n843));
  AND2_X1   g657(.A1(new_n685), .A2(new_n468), .ZN(new_n844));
  INV_X1    g658(.A(new_n844), .ZN(new_n845));
  NOR2_X1   g659(.A1(new_n845), .A2(new_n414), .ZN(new_n846));
  INV_X1    g660(.A(new_n846), .ZN(new_n847));
  NOR2_X1   g661(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n848));
  AOI21_X1  g662(.A(new_n848), .B1(new_n780), .B2(new_n783), .ZN(new_n849));
  NAND2_X1  g663(.A1(new_n847), .A2(KEYINPUT116), .ZN(new_n850));
  AOI21_X1  g664(.A(new_n843), .B1(new_n849), .B2(new_n850), .ZN(new_n851));
  INV_X1    g665(.A(KEYINPUT117), .ZN(new_n852));
  NOR2_X1   g666(.A1(new_n696), .A2(new_n296), .ZN(new_n853));
  AOI21_X1  g667(.A(new_n677), .B1(new_n852), .B2(new_n853), .ZN(new_n854));
  OAI211_X1 g668(.A(new_n837), .B(new_n854), .C1(new_n852), .C2(new_n853), .ZN(new_n855));
  XOR2_X1   g669(.A(new_n855), .B(KEYINPUT50), .Z(new_n856));
  NOR3_X1   g670(.A1(new_n696), .A2(new_n835), .A3(new_n766), .ZN(new_n857));
  AND2_X1   g671(.A1(new_n769), .A2(new_n857), .ZN(new_n858));
  NAND2_X1  g672(.A1(new_n858), .A2(new_n720), .ZN(new_n859));
  NAND3_X1  g673(.A1(new_n666), .A2(new_n579), .A3(new_n857), .ZN(new_n860));
  INV_X1    g674(.A(new_n860), .ZN(new_n861));
  NAND3_X1  g675(.A1(new_n861), .A2(new_n260), .A3(new_n597), .ZN(new_n862));
  NAND3_X1  g676(.A1(new_n856), .A2(new_n859), .A3(new_n862), .ZN(new_n863));
  OAI21_X1  g677(.A(new_n841), .B1(new_n851), .B2(new_n863), .ZN(new_n864));
  OR2_X1    g678(.A1(new_n741), .A2(new_n742), .ZN(new_n865));
  NAND2_X1  g679(.A1(new_n865), .A2(new_n858), .ZN(new_n866));
  XNOR2_X1  g680(.A(new_n866), .B(KEYINPUT118), .ZN(new_n867));
  INV_X1    g681(.A(KEYINPUT48), .ZN(new_n868));
  OAI211_X1 g682(.A(G952), .B(new_n203), .C1(new_n867), .C2(new_n868), .ZN(new_n869));
  INV_X1    g683(.A(new_n863), .ZN(new_n870));
  NOR2_X1   g684(.A1(new_n763), .A2(KEYINPUT47), .ZN(new_n871));
  OAI21_X1  g685(.A(new_n847), .B1(new_n871), .B2(new_n782), .ZN(new_n872));
  AOI21_X1  g686(.A(new_n841), .B1(new_n872), .B2(new_n842), .ZN(new_n873));
  AOI21_X1  g687(.A(new_n869), .B1(new_n870), .B2(new_n873), .ZN(new_n874));
  NAND3_X1  g688(.A1(new_n861), .A2(new_n598), .A3(new_n605), .ZN(new_n875));
  NAND3_X1  g689(.A1(new_n866), .A2(KEYINPUT118), .A3(new_n868), .ZN(new_n876));
  NAND4_X1  g690(.A1(new_n864), .A2(new_n874), .A3(new_n875), .A4(new_n876), .ZN(new_n877));
  OAI22_X1  g691(.A1(new_n840), .A2(new_n877), .B1(G952), .B2(G953), .ZN(new_n878));
  NAND2_X1  g692(.A1(new_n845), .A2(KEYINPUT49), .ZN(new_n879));
  NOR2_X1   g693(.A1(new_n729), .A2(new_n768), .ZN(new_n880));
  NAND3_X1  g694(.A1(new_n666), .A2(new_n879), .A3(new_n880), .ZN(new_n881));
  NOR2_X1   g695(.A1(new_n881), .A2(new_n677), .ZN(new_n882));
  OAI211_X1 g696(.A(new_n882), .B(new_n732), .C1(KEYINPUT49), .C2(new_n845), .ZN(new_n883));
  NAND2_X1  g697(.A1(new_n878), .A2(new_n883), .ZN(G75));
  NOR2_X1   g698(.A1(new_n203), .A2(G952), .ZN(new_n885));
  INV_X1    g699(.A(new_n830), .ZN(new_n886));
  NOR2_X1   g700(.A1(new_n886), .A2(new_n237), .ZN(new_n887));
  AOI21_X1  g701(.A(KEYINPUT120), .B1(new_n887), .B2(G210), .ZN(new_n888));
  INV_X1    g702(.A(KEYINPUT56), .ZN(new_n889));
  OR2_X1    g703(.A1(new_n889), .A2(KEYINPUT119), .ZN(new_n890));
  NAND2_X1  g704(.A1(new_n888), .A2(new_n890), .ZN(new_n891));
  OAI21_X1  g705(.A(new_n382), .B1(new_n386), .B2(new_n387), .ZN(new_n892));
  XNOR2_X1  g706(.A(new_n892), .B(new_n337), .ZN(new_n893));
  XNOR2_X1  g707(.A(new_n893), .B(KEYINPUT55), .ZN(new_n894));
  NAND2_X1  g708(.A1(new_n891), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g709(.A1(new_n887), .A2(G210), .ZN(new_n896));
  NOR2_X1   g710(.A1(new_n894), .A2(KEYINPUT120), .ZN(new_n897));
  OAI211_X1 g711(.A(new_n896), .B(new_n889), .C1(KEYINPUT119), .C2(new_n897), .ZN(new_n898));
  AOI21_X1  g712(.A(new_n885), .B1(new_n895), .B2(new_n898), .ZN(G51));
  NAND2_X1  g713(.A1(new_n470), .A2(KEYINPUT57), .ZN(new_n900));
  OR2_X1    g714(.A1(new_n470), .A2(KEYINPUT57), .ZN(new_n901));
  NOR2_X1   g715(.A1(new_n886), .A2(new_n827), .ZN(new_n902));
  INV_X1    g716(.A(new_n828), .ZN(new_n903));
  OAI211_X1 g717(.A(new_n900), .B(new_n901), .C1(new_n902), .C2(new_n903), .ZN(new_n904));
  OAI21_X1  g718(.A(new_n904), .B1(new_n467), .B2(new_n466), .ZN(new_n905));
  OR3_X1    g719(.A1(new_n886), .A2(new_n237), .A3(new_n756), .ZN(new_n906));
  AOI21_X1  g720(.A(new_n885), .B1(new_n905), .B2(new_n906), .ZN(G54));
  NAND3_X1  g721(.A1(new_n887), .A2(KEYINPUT58), .A3(G475), .ZN(new_n908));
  NOR2_X1   g722(.A1(new_n250), .A2(new_n234), .ZN(new_n909));
  AND2_X1   g723(.A1(new_n908), .A2(new_n909), .ZN(new_n910));
  NOR2_X1   g724(.A1(new_n908), .A2(new_n909), .ZN(new_n911));
  NOR3_X1   g725(.A1(new_n910), .A2(new_n911), .A3(new_n885), .ZN(G60));
  NAND2_X1  g726(.A1(G478), .A2(G902), .ZN(new_n913));
  XNOR2_X1  g727(.A(new_n913), .B(KEYINPUT59), .ZN(new_n914));
  OAI21_X1  g728(.A(new_n914), .B1(new_n902), .B2(new_n903), .ZN(new_n915));
  NAND2_X1  g729(.A1(new_n594), .A2(new_n595), .ZN(new_n916));
  OAI22_X1  g730(.A1(new_n915), .A2(new_n916), .B1(G952), .B2(new_n203), .ZN(new_n917));
  NAND2_X1  g731(.A1(new_n834), .A2(new_n914), .ZN(new_n918));
  NAND2_X1  g732(.A1(new_n918), .A2(new_n916), .ZN(new_n919));
  NAND2_X1  g733(.A1(new_n919), .A2(KEYINPUT121), .ZN(new_n920));
  INV_X1    g734(.A(KEYINPUT121), .ZN(new_n921));
  NAND3_X1  g735(.A1(new_n918), .A2(new_n921), .A3(new_n916), .ZN(new_n922));
  AOI21_X1  g736(.A(new_n917), .B1(new_n920), .B2(new_n922), .ZN(G63));
  NAND2_X1  g737(.A1(G217), .A2(G902), .ZN(new_n924));
  XNOR2_X1  g738(.A(new_n924), .B(KEYINPUT60), .ZN(new_n925));
  AOI21_X1  g739(.A(new_n925), .B1(new_n819), .B2(new_n825), .ZN(new_n926));
  INV_X1    g740(.A(new_n926), .ZN(new_n927));
  AOI21_X1  g741(.A(new_n885), .B1(new_n927), .B2(new_n567), .ZN(new_n928));
  INV_X1    g742(.A(new_n925), .ZN(new_n929));
  NAND3_X1  g743(.A1(new_n830), .A2(new_n627), .A3(new_n929), .ZN(new_n930));
  NOR2_X1   g744(.A1(new_n930), .A2(KEYINPUT122), .ZN(new_n931));
  INV_X1    g745(.A(KEYINPUT122), .ZN(new_n932));
  AOI21_X1  g746(.A(new_n932), .B1(new_n926), .B2(new_n627), .ZN(new_n933));
  OAI21_X1  g747(.A(new_n928), .B1(new_n931), .B2(new_n933), .ZN(new_n934));
  NAND3_X1  g748(.A1(new_n934), .A2(KEYINPUT123), .A3(KEYINPUT61), .ZN(new_n935));
  XNOR2_X1  g749(.A(new_n930), .B(KEYINPUT122), .ZN(new_n936));
  NAND2_X1  g750(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n937));
  OR2_X1    g751(.A1(KEYINPUT123), .A2(KEYINPUT61), .ZN(new_n938));
  NAND4_X1  g752(.A1(new_n936), .A2(new_n937), .A3(new_n938), .A4(new_n928), .ZN(new_n939));
  AND2_X1   g753(.A1(new_n935), .A2(new_n939), .ZN(G66));
  AOI21_X1  g754(.A(new_n203), .B1(new_n301), .B2(G224), .ZN(new_n941));
  INV_X1    g755(.A(new_n824), .ZN(new_n942));
  AOI21_X1  g756(.A(new_n941), .B1(new_n942), .B2(new_n203), .ZN(new_n943));
  OAI21_X1  g757(.A(new_n892), .B1(G898), .B2(new_n203), .ZN(new_n944));
  XOR2_X1   g758(.A(new_n944), .B(KEYINPUT124), .Z(new_n945));
  XNOR2_X1  g759(.A(new_n943), .B(new_n945), .ZN(G69));
  NAND2_X1  g760(.A1(new_n727), .A2(new_n788), .ZN(new_n947));
  AND3_X1   g761(.A1(new_n764), .A2(new_n667), .A3(new_n703), .ZN(new_n948));
  AOI21_X1  g762(.A(new_n947), .B1(new_n948), .B2(new_n865), .ZN(new_n949));
  AND2_X1   g763(.A1(new_n744), .A2(new_n747), .ZN(new_n950));
  NAND4_X1  g764(.A1(new_n949), .A2(new_n776), .A3(new_n785), .A4(new_n950), .ZN(new_n951));
  XNOR2_X1  g765(.A(new_n520), .B(new_n245), .ZN(new_n952));
  AOI21_X1  g766(.A(G953), .B1(new_n951), .B2(new_n952), .ZN(new_n953));
  INV_X1    g767(.A(new_n803), .ZN(new_n954));
  NOR4_X1   g768(.A1(new_n954), .A2(new_n580), .A3(new_n668), .A4(new_n766), .ZN(new_n955));
  NAND3_X1  g769(.A1(new_n678), .A2(new_n727), .A3(new_n788), .ZN(new_n956));
  INV_X1    g770(.A(KEYINPUT62), .ZN(new_n957));
  OR2_X1    g771(.A1(new_n956), .A2(new_n957), .ZN(new_n958));
  NAND2_X1  g772(.A1(new_n956), .A2(new_n957), .ZN(new_n959));
  AOI21_X1  g773(.A(new_n955), .B1(new_n958), .B2(new_n959), .ZN(new_n960));
  NAND3_X1  g774(.A1(new_n960), .A2(new_n776), .A3(new_n785), .ZN(new_n961));
  OAI21_X1  g775(.A(new_n953), .B1(new_n952), .B2(new_n961), .ZN(new_n962));
  INV_X1    g776(.A(new_n952), .ZN(new_n963));
  NAND3_X1  g777(.A1(new_n963), .A2(G227), .A3(G900), .ZN(new_n964));
  INV_X1    g778(.A(KEYINPUT125), .ZN(new_n965));
  OAI21_X1  g779(.A(G900), .B1(new_n965), .B2(G227), .ZN(new_n966));
  OAI211_X1 g780(.A(new_n952), .B(new_n966), .C1(new_n965), .C2(G900), .ZN(new_n967));
  NAND3_X1  g781(.A1(new_n964), .A2(G953), .A3(new_n967), .ZN(new_n968));
  NAND2_X1  g782(.A1(new_n962), .A2(new_n968), .ZN(G72));
  NAND2_X1  g783(.A1(G472), .A2(G902), .ZN(new_n970));
  XOR2_X1   g784(.A(new_n970), .B(KEYINPUT63), .Z(new_n971));
  OAI21_X1  g785(.A(new_n971), .B1(new_n951), .B2(new_n942), .ZN(new_n972));
  XOR2_X1   g786(.A(new_n521), .B(KEYINPUT126), .Z(new_n973));
  NOR2_X1   g787(.A1(new_n973), .A2(new_n477), .ZN(new_n974));
  AOI21_X1  g788(.A(new_n885), .B1(new_n972), .B2(new_n974), .ZN(new_n975));
  OAI21_X1  g789(.A(new_n971), .B1(new_n529), .B2(new_n660), .ZN(new_n976));
  XOR2_X1   g790(.A(new_n976), .B(KEYINPUT127), .Z(new_n977));
  NAND2_X1  g791(.A1(new_n830), .A2(new_n977), .ZN(new_n978));
  OAI21_X1  g792(.A(new_n971), .B1(new_n961), .B2(new_n942), .ZN(new_n979));
  NAND3_X1  g793(.A1(new_n979), .A2(new_n477), .A3(new_n973), .ZN(new_n980));
  AND3_X1   g794(.A1(new_n975), .A2(new_n978), .A3(new_n980), .ZN(G57));
endmodule


