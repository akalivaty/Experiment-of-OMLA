//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 0 1 1 0 0 0 0 1 1 1 0 1 1 0 0 0 0 0 0 0 1 0 0 1 0 0 0 0 0 1 0 1 0 0 1 0 1 1 0 0 1 1 1 0 1 1 0 1 0 1 1 1 1 0 1 1 1 1 1 1 0' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:20:12 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n636, new_n637, new_n638, new_n639, new_n640, new_n641, new_n642,
    new_n643, new_n644, new_n645, new_n646, new_n647, new_n648, new_n649,
    new_n650, new_n651, new_n652, new_n653, new_n654, new_n655, new_n656,
    new_n657, new_n658, new_n659, new_n660, new_n661, new_n662, new_n663,
    new_n664, new_n665, new_n666, new_n667, new_n668, new_n669, new_n670,
    new_n671, new_n672, new_n673, new_n674, new_n675, new_n676, new_n677,
    new_n678, new_n679, new_n680, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n688, new_n689, new_n690, new_n691,
    new_n692, new_n693, new_n694, new_n695, new_n696, new_n697, new_n698,
    new_n699, new_n700, new_n701, new_n702, new_n703, new_n704, new_n705,
    new_n706, new_n707, new_n708, new_n709, new_n710, new_n711, new_n712,
    new_n713, new_n714, new_n715, new_n716, new_n717, new_n718, new_n719,
    new_n720, new_n721, new_n722, new_n723, new_n724, new_n725, new_n726,
    new_n727, new_n728, new_n730, new_n731, new_n732, new_n733, new_n734,
    new_n736, new_n737, new_n738, new_n739, new_n740, new_n741, new_n743,
    new_n744, new_n745, new_n746, new_n747, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n777, new_n778, new_n779, new_n781,
    new_n782, new_n783, new_n784, new_n785, new_n786, new_n787, new_n788,
    new_n789, new_n791, new_n792, new_n793, new_n794, new_n795, new_n796,
    new_n797, new_n799, new_n800, new_n801, new_n802, new_n803, new_n805,
    new_n806, new_n807, new_n808, new_n809, new_n811, new_n812, new_n813,
    new_n814, new_n816, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n824, new_n825, new_n826, new_n827, new_n828, new_n829,
    new_n830, new_n831, new_n832, new_n833, new_n834, new_n835, new_n836,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n848, new_n849, new_n850, new_n851,
    new_n852, new_n853, new_n855, new_n856, new_n858, new_n859, new_n860,
    new_n861, new_n862, new_n863, new_n864, new_n865, new_n866, new_n868,
    new_n869, new_n870, new_n871, new_n872, new_n873, new_n874, new_n875,
    new_n876, new_n877, new_n878, new_n879, new_n880, new_n881, new_n882,
    new_n883, new_n884, new_n885, new_n886, new_n887, new_n888, new_n889,
    new_n890, new_n891, new_n892, new_n893, new_n894, new_n895, new_n896,
    new_n897, new_n898, new_n899, new_n900, new_n902, new_n903, new_n905,
    new_n906, new_n908, new_n909, new_n910, new_n911, new_n912, new_n913,
    new_n915, new_n916, new_n917, new_n918, new_n919, new_n920, new_n921,
    new_n922, new_n923, new_n924, new_n925, new_n926, new_n927, new_n928,
    new_n929, new_n930, new_n931, new_n932, new_n933, new_n934, new_n935,
    new_n936, new_n937, new_n938, new_n939, new_n940, new_n941, new_n942,
    new_n943, new_n944, new_n945, new_n947, new_n948, new_n949, new_n950,
    new_n951, new_n952, new_n953, new_n954, new_n955, new_n957, new_n958,
    new_n960, new_n961, new_n962, new_n963, new_n964, new_n965, new_n966,
    new_n968, new_n969, new_n970, new_n971, new_n972, new_n973, new_n974,
    new_n975, new_n977, new_n978, new_n979, new_n981, new_n982, new_n983,
    new_n984, new_n985, new_n986, new_n987, new_n988, new_n989, new_n990,
    new_n991, new_n992, new_n993, new_n994, new_n996, new_n997, new_n998,
    new_n999, new_n1000, new_n1001, new_n1002, new_n1003, new_n1005,
    new_n1006, new_n1007, new_n1008, new_n1009, new_n1010, new_n1012,
    new_n1013, new_n1014, new_n1015, new_n1016, new_n1017, new_n1018,
    new_n1020, new_n1021, new_n1022, new_n1023, new_n1024, new_n1025,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031;
  XOR2_X1   g000(.A(G8gat), .B(G36gat), .Z(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT76), .ZN(new_n203));
  XNOR2_X1  g002(.A(G64gat), .B(G92gat), .ZN(new_n204));
  XOR2_X1   g003(.A(new_n203), .B(new_n204), .Z(new_n205));
  INV_X1    g004(.A(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(KEYINPUT75), .ZN(new_n207));
  NAND2_X1  g006(.A1(G226gat), .A2(G233gat), .ZN(new_n208));
  INV_X1    g007(.A(new_n208), .ZN(new_n209));
  INV_X1    g008(.A(KEYINPUT26), .ZN(new_n210));
  INV_X1    g009(.A(G169gat), .ZN(new_n211));
  INV_X1    g010(.A(G176gat), .ZN(new_n212));
  NAND3_X1  g011(.A1(new_n210), .A2(new_n211), .A3(new_n212), .ZN(new_n213));
  OAI21_X1  g012(.A(KEYINPUT26), .B1(G169gat), .B2(G176gat), .ZN(new_n214));
  NAND3_X1  g013(.A1(KEYINPUT66), .A2(G169gat), .A3(G176gat), .ZN(new_n215));
  INV_X1    g014(.A(new_n215), .ZN(new_n216));
  AOI21_X1  g015(.A(KEYINPUT66), .B1(G169gat), .B2(G176gat), .ZN(new_n217));
  OAI211_X1 g016(.A(new_n213), .B(new_n214), .C1(new_n216), .C2(new_n217), .ZN(new_n218));
  NAND2_X1  g017(.A1(G183gat), .A2(G190gat), .ZN(new_n219));
  AND2_X1   g018(.A1(new_n218), .A2(new_n219), .ZN(new_n220));
  INV_X1    g019(.A(G183gat), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT27), .ZN(new_n222));
  INV_X1    g021(.A(KEYINPUT27), .ZN(new_n223));
  NAND2_X1  g022(.A1(new_n223), .A2(G183gat), .ZN(new_n224));
  INV_X1    g023(.A(KEYINPUT68), .ZN(new_n225));
  AND3_X1   g024(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n226));
  AOI21_X1  g025(.A(new_n225), .B1(new_n222), .B2(new_n224), .ZN(new_n227));
  INV_X1    g026(.A(KEYINPUT28), .ZN(new_n228));
  NOR2_X1   g027(.A1(new_n228), .A2(G190gat), .ZN(new_n229));
  INV_X1    g028(.A(new_n229), .ZN(new_n230));
  NOR3_X1   g029(.A1(new_n226), .A2(new_n227), .A3(new_n230), .ZN(new_n231));
  NAND2_X1  g030(.A1(new_n222), .A2(new_n224), .ZN(new_n232));
  OAI21_X1  g031(.A(new_n228), .B1(new_n232), .B2(G190gat), .ZN(new_n233));
  INV_X1    g032(.A(new_n233), .ZN(new_n234));
  OAI21_X1  g033(.A(new_n220), .B1(new_n231), .B2(new_n234), .ZN(new_n235));
  NAND3_X1  g034(.A1(KEYINPUT24), .A2(G183gat), .A3(G190gat), .ZN(new_n236));
  OAI21_X1  g035(.A(new_n236), .B1(G183gat), .B2(G190gat), .ZN(new_n237));
  INV_X1    g036(.A(KEYINPUT24), .ZN(new_n238));
  OR2_X1    g037(.A1(new_n238), .A2(KEYINPUT67), .ZN(new_n239));
  AOI22_X1  g038(.A1(new_n238), .A2(KEYINPUT67), .B1(G183gat), .B2(G190gat), .ZN(new_n240));
  AOI21_X1  g039(.A(new_n237), .B1(new_n239), .B2(new_n240), .ZN(new_n241));
  NOR2_X1   g040(.A1(G169gat), .A2(G176gat), .ZN(new_n242));
  NAND2_X1  g041(.A1(new_n242), .A2(KEYINPUT23), .ZN(new_n243));
  INV_X1    g042(.A(KEYINPUT23), .ZN(new_n244));
  OAI21_X1  g043(.A(new_n244), .B1(G169gat), .B2(G176gat), .ZN(new_n245));
  OAI211_X1 g044(.A(new_n243), .B(new_n245), .C1(new_n216), .C2(new_n217), .ZN(new_n246));
  OAI21_X1  g045(.A(KEYINPUT25), .B1(new_n241), .B2(new_n246), .ZN(new_n247));
  INV_X1    g046(.A(KEYINPUT65), .ZN(new_n248));
  NAND2_X1  g047(.A1(new_n243), .A2(new_n248), .ZN(new_n249));
  NAND3_X1  g048(.A1(new_n242), .A2(KEYINPUT65), .A3(KEYINPUT23), .ZN(new_n250));
  NAND2_X1  g049(.A1(new_n249), .A2(new_n250), .ZN(new_n251));
  INV_X1    g050(.A(new_n217), .ZN(new_n252));
  INV_X1    g051(.A(new_n242), .ZN(new_n253));
  AOI22_X1  g052(.A1(new_n252), .A2(new_n215), .B1(new_n253), .B2(new_n244), .ZN(new_n254));
  NAND2_X1  g053(.A1(new_n219), .A2(new_n238), .ZN(new_n255));
  INV_X1    g054(.A(G190gat), .ZN(new_n256));
  NAND3_X1  g055(.A1(new_n221), .A2(new_n256), .A3(KEYINPUT64), .ZN(new_n257));
  INV_X1    g056(.A(KEYINPUT64), .ZN(new_n258));
  OAI21_X1  g057(.A(new_n258), .B1(G183gat), .B2(G190gat), .ZN(new_n259));
  NAND4_X1  g058(.A1(new_n255), .A2(new_n257), .A3(new_n259), .A4(new_n236), .ZN(new_n260));
  INV_X1    g059(.A(KEYINPUT25), .ZN(new_n261));
  NAND4_X1  g060(.A1(new_n251), .A2(new_n254), .A3(new_n260), .A4(new_n261), .ZN(new_n262));
  NAND3_X1  g061(.A1(new_n235), .A2(new_n247), .A3(new_n262), .ZN(new_n263));
  INV_X1    g062(.A(KEYINPUT29), .ZN(new_n264));
  AOI21_X1  g063(.A(new_n209), .B1(new_n263), .B2(new_n264), .ZN(new_n265));
  NAND2_X1  g064(.A1(G211gat), .A2(G218gat), .ZN(new_n266));
  INV_X1    g065(.A(KEYINPUT22), .ZN(new_n267));
  NAND2_X1  g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n268), .A2(KEYINPUT73), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT73), .ZN(new_n270));
  NAND3_X1  g069(.A1(new_n266), .A2(new_n270), .A3(new_n267), .ZN(new_n271));
  XNOR2_X1  g070(.A(G197gat), .B(G204gat), .ZN(new_n272));
  NAND3_X1  g071(.A1(new_n269), .A2(new_n271), .A3(new_n272), .ZN(new_n273));
  XOR2_X1   g072(.A(G211gat), .B(G218gat), .Z(new_n274));
  INV_X1    g073(.A(new_n274), .ZN(new_n275));
  NAND3_X1  g074(.A1(new_n273), .A2(KEYINPUT74), .A3(new_n275), .ZN(new_n276));
  INV_X1    g075(.A(new_n276), .ZN(new_n277));
  AOI21_X1  g076(.A(new_n275), .B1(new_n273), .B2(KEYINPUT74), .ZN(new_n278));
  NOR2_X1   g077(.A1(new_n277), .A2(new_n278), .ZN(new_n279));
  AND2_X1   g078(.A1(new_n247), .A2(new_n262), .ZN(new_n280));
  AOI21_X1  g079(.A(new_n208), .B1(new_n280), .B2(new_n235), .ZN(new_n281));
  NOR3_X1   g080(.A1(new_n265), .A2(new_n279), .A3(new_n281), .ZN(new_n282));
  NAND2_X1  g081(.A1(new_n273), .A2(KEYINPUT74), .ZN(new_n283));
  NAND2_X1  g082(.A1(new_n283), .A2(new_n274), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n284), .A2(new_n276), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n247), .A2(new_n262), .ZN(new_n286));
  NAND2_X1  g085(.A1(new_n218), .A2(new_n219), .ZN(new_n287));
  NAND2_X1  g086(.A1(new_n232), .A2(KEYINPUT68), .ZN(new_n288));
  NAND3_X1  g087(.A1(new_n222), .A2(new_n224), .A3(new_n225), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n288), .A2(new_n289), .A3(new_n229), .ZN(new_n290));
  AOI21_X1  g089(.A(new_n287), .B1(new_n290), .B2(new_n233), .ZN(new_n291));
  OAI21_X1  g090(.A(new_n264), .B1(new_n286), .B2(new_n291), .ZN(new_n292));
  NAND2_X1  g091(.A1(new_n292), .A2(new_n208), .ZN(new_n293));
  NAND2_X1  g092(.A1(new_n263), .A2(new_n209), .ZN(new_n294));
  AOI21_X1  g093(.A(new_n285), .B1(new_n293), .B2(new_n294), .ZN(new_n295));
  OAI21_X1  g094(.A(new_n207), .B1(new_n282), .B2(new_n295), .ZN(new_n296));
  OAI21_X1  g095(.A(new_n279), .B1(new_n265), .B2(new_n281), .ZN(new_n297));
  NAND3_X1  g096(.A1(new_n293), .A2(new_n285), .A3(new_n294), .ZN(new_n298));
  NAND3_X1  g097(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n298), .ZN(new_n299));
  AOI21_X1  g098(.A(new_n206), .B1(new_n296), .B2(new_n299), .ZN(new_n300));
  NAND2_X1  g099(.A1(new_n297), .A2(new_n298), .ZN(new_n301));
  AND3_X1   g100(.A1(new_n301), .A2(KEYINPUT30), .A3(new_n206), .ZN(new_n302));
  AOI21_X1  g101(.A(new_n205), .B1(new_n297), .B2(new_n298), .ZN(new_n303));
  NOR2_X1   g102(.A1(new_n303), .A2(KEYINPUT30), .ZN(new_n304));
  OR3_X1    g103(.A1(new_n300), .A2(new_n302), .A3(new_n304), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(KEYINPUT35), .ZN(new_n307));
  XNOR2_X1  g106(.A(G78gat), .B(G106gat), .ZN(new_n308));
  INV_X1    g107(.A(G50gat), .ZN(new_n309));
  XNOR2_X1  g108(.A(new_n308), .B(new_n309), .ZN(new_n310));
  XNOR2_X1  g109(.A(KEYINPUT83), .B(KEYINPUT31), .ZN(new_n311));
  XOR2_X1   g110(.A(new_n310), .B(new_n311), .Z(new_n312));
  NAND2_X1  g111(.A1(G228gat), .A2(G233gat), .ZN(new_n313));
  INV_X1    g112(.A(KEYINPUT78), .ZN(new_n314));
  INV_X1    g113(.A(G141gat), .ZN(new_n315));
  OAI21_X1  g114(.A(new_n314), .B1(new_n315), .B2(G148gat), .ZN(new_n316));
  INV_X1    g115(.A(G148gat), .ZN(new_n317));
  NAND3_X1  g116(.A1(new_n317), .A2(KEYINPUT78), .A3(G141gat), .ZN(new_n318));
  NAND2_X1  g117(.A1(new_n315), .A2(G148gat), .ZN(new_n319));
  NAND3_X1  g118(.A1(new_n316), .A2(new_n318), .A3(new_n319), .ZN(new_n320));
  NAND2_X1  g119(.A1(G155gat), .A2(G162gat), .ZN(new_n321));
  INV_X1    g120(.A(G155gat), .ZN(new_n322));
  INV_X1    g121(.A(G162gat), .ZN(new_n323));
  NAND2_X1  g122(.A1(new_n322), .A2(new_n323), .ZN(new_n324));
  OAI21_X1  g123(.A(new_n321), .B1(new_n324), .B2(KEYINPUT2), .ZN(new_n325));
  NAND2_X1  g124(.A1(new_n320), .A2(new_n325), .ZN(new_n326));
  AND2_X1   g125(.A1(G155gat), .A2(G162gat), .ZN(new_n327));
  NOR2_X1   g126(.A1(G155gat), .A2(G162gat), .ZN(new_n328));
  NOR2_X1   g127(.A1(new_n327), .A2(new_n328), .ZN(new_n329));
  XNOR2_X1  g128(.A(G141gat), .B(G148gat), .ZN(new_n330));
  OAI21_X1  g129(.A(new_n329), .B1(new_n330), .B2(KEYINPUT2), .ZN(new_n331));
  XOR2_X1   g130(.A(KEYINPUT79), .B(KEYINPUT3), .Z(new_n332));
  NAND3_X1  g131(.A1(new_n326), .A2(new_n331), .A3(new_n332), .ZN(new_n333));
  AOI22_X1  g132(.A1(new_n284), .A2(new_n276), .B1(new_n264), .B2(new_n333), .ZN(new_n334));
  INV_X1    g133(.A(KEYINPUT84), .ZN(new_n335));
  INV_X1    g134(.A(KEYINPUT2), .ZN(new_n336));
  NOR2_X1   g135(.A1(new_n315), .A2(G148gat), .ZN(new_n337));
  NOR2_X1   g136(.A1(new_n317), .A2(G141gat), .ZN(new_n338));
  OAI21_X1  g137(.A(new_n336), .B1(new_n337), .B2(new_n338), .ZN(new_n339));
  AOI22_X1  g138(.A1(new_n339), .A2(new_n329), .B1(new_n320), .B2(new_n325), .ZN(new_n340));
  INV_X1    g139(.A(new_n332), .ZN(new_n341));
  AOI21_X1  g140(.A(KEYINPUT29), .B1(new_n273), .B2(new_n275), .ZN(new_n342));
  NAND4_X1  g141(.A1(new_n274), .A2(new_n269), .A3(new_n271), .A4(new_n272), .ZN(new_n343));
  AOI21_X1  g142(.A(new_n341), .B1(new_n342), .B2(new_n343), .ZN(new_n344));
  OAI22_X1  g143(.A1(new_n334), .A2(new_n335), .B1(new_n340), .B2(new_n344), .ZN(new_n345));
  NAND2_X1  g144(.A1(new_n333), .A2(new_n264), .ZN(new_n346));
  AND3_X1   g145(.A1(new_n285), .A2(new_n335), .A3(new_n346), .ZN(new_n347));
  OAI21_X1  g146(.A(new_n313), .B1(new_n345), .B2(new_n347), .ZN(new_n348));
  INV_X1    g147(.A(G22gat), .ZN(new_n349));
  INV_X1    g148(.A(new_n313), .ZN(new_n350));
  NAND2_X1  g149(.A1(new_n285), .A2(new_n346), .ZN(new_n351));
  AOI21_X1  g150(.A(KEYINPUT3), .B1(new_n279), .B2(new_n264), .ZN(new_n352));
  OAI211_X1 g151(.A(new_n350), .B(new_n351), .C1(new_n352), .C2(new_n340), .ZN(new_n353));
  NAND3_X1  g152(.A1(new_n348), .A2(new_n349), .A3(new_n353), .ZN(new_n354));
  INV_X1    g153(.A(new_n354), .ZN(new_n355));
  AOI21_X1  g154(.A(new_n349), .B1(new_n348), .B2(new_n353), .ZN(new_n356));
  OAI21_X1  g155(.A(new_n312), .B1(new_n355), .B2(new_n356), .ZN(new_n357));
  NAND2_X1  g156(.A1(new_n354), .A2(KEYINPUT86), .ZN(new_n358));
  INV_X1    g157(.A(KEYINPUT86), .ZN(new_n359));
  NAND4_X1  g158(.A1(new_n348), .A2(new_n353), .A3(new_n359), .A4(new_n349), .ZN(new_n360));
  INV_X1    g159(.A(KEYINPUT85), .ZN(new_n361));
  NAND2_X1  g160(.A1(new_n273), .A2(new_n275), .ZN(new_n362));
  NAND3_X1  g161(.A1(new_n362), .A2(new_n264), .A3(new_n343), .ZN(new_n363));
  AOI21_X1  g162(.A(new_n340), .B1(new_n363), .B2(new_n332), .ZN(new_n364));
  AOI21_X1  g163(.A(new_n364), .B1(new_n351), .B2(KEYINPUT84), .ZN(new_n365));
  NAND2_X1  g164(.A1(new_n334), .A2(new_n335), .ZN(new_n366));
  AOI21_X1  g165(.A(new_n350), .B1(new_n365), .B2(new_n366), .ZN(new_n367));
  NAND3_X1  g166(.A1(new_n284), .A2(new_n264), .A3(new_n276), .ZN(new_n368));
  INV_X1    g167(.A(KEYINPUT3), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n340), .B1(new_n368), .B2(new_n369), .ZN(new_n370));
  NOR3_X1   g169(.A1(new_n370), .A2(new_n313), .A3(new_n334), .ZN(new_n371));
  OAI211_X1 g170(.A(new_n361), .B(G22gat), .C1(new_n367), .C2(new_n371), .ZN(new_n372));
  NAND3_X1  g171(.A1(new_n358), .A2(new_n360), .A3(new_n372), .ZN(new_n373));
  INV_X1    g172(.A(new_n312), .ZN(new_n374));
  OAI21_X1  g173(.A(new_n374), .B1(new_n356), .B2(new_n361), .ZN(new_n375));
  OAI21_X1  g174(.A(new_n357), .B1(new_n373), .B2(new_n375), .ZN(new_n376));
  NAND3_X1  g175(.A1(new_n306), .A2(new_n307), .A3(new_n376), .ZN(new_n377));
  INV_X1    g176(.A(new_n377), .ZN(new_n378));
  INV_X1    g177(.A(KEYINPUT1), .ZN(new_n379));
  INV_X1    g178(.A(G113gat), .ZN(new_n380));
  NAND2_X1  g179(.A1(new_n380), .A2(G120gat), .ZN(new_n381));
  INV_X1    g180(.A(new_n381), .ZN(new_n382));
  NOR2_X1   g181(.A1(new_n380), .A2(G120gat), .ZN(new_n383));
  OAI21_X1  g182(.A(new_n379), .B1(new_n382), .B2(new_n383), .ZN(new_n384));
  INV_X1    g183(.A(G134gat), .ZN(new_n385));
  NAND2_X1  g184(.A1(new_n385), .A2(G127gat), .ZN(new_n386));
  INV_X1    g185(.A(G127gat), .ZN(new_n387));
  NAND2_X1  g186(.A1(new_n387), .A2(G134gat), .ZN(new_n388));
  NAND2_X1  g187(.A1(new_n386), .A2(new_n388), .ZN(new_n389));
  AND3_X1   g188(.A1(new_n386), .A2(new_n388), .A3(new_n379), .ZN(new_n390));
  INV_X1    g189(.A(KEYINPUT69), .ZN(new_n391));
  OAI21_X1  g190(.A(new_n391), .B1(new_n380), .B2(G120gat), .ZN(new_n392));
  INV_X1    g191(.A(G120gat), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n393), .A2(KEYINPUT69), .A3(G113gat), .ZN(new_n394));
  NAND3_X1  g193(.A1(new_n392), .A2(new_n381), .A3(new_n394), .ZN(new_n395));
  AOI22_X1  g194(.A1(new_n384), .A2(new_n389), .B1(new_n390), .B2(new_n395), .ZN(new_n396));
  OR2_X1    g195(.A1(new_n396), .A2(new_n340), .ZN(new_n397));
  NAND2_X1  g196(.A1(new_n390), .A2(new_n395), .ZN(new_n398));
  XNOR2_X1  g197(.A(G113gat), .B(G120gat), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n389), .B1(new_n399), .B2(KEYINPUT1), .ZN(new_n400));
  NAND4_X1  g199(.A1(new_n398), .A2(new_n326), .A3(new_n331), .A4(new_n400), .ZN(new_n401));
  NAND2_X1  g200(.A1(G225gat), .A2(G233gat), .ZN(new_n402));
  XOR2_X1   g201(.A(new_n402), .B(KEYINPUT80), .Z(new_n403));
  INV_X1    g202(.A(new_n403), .ZN(new_n404));
  NAND4_X1  g203(.A1(new_n397), .A2(KEYINPUT5), .A3(new_n401), .A4(new_n404), .ZN(new_n405));
  NAND2_X1  g204(.A1(new_n398), .A2(new_n400), .ZN(new_n406));
  OAI211_X1 g205(.A(new_n333), .B(new_n406), .C1(new_n340), .C2(new_n369), .ZN(new_n407));
  INV_X1    g206(.A(KEYINPUT4), .ZN(new_n408));
  NAND2_X1  g207(.A1(new_n401), .A2(new_n408), .ZN(new_n409));
  XNOR2_X1  g208(.A(KEYINPUT81), .B(KEYINPUT4), .ZN(new_n410));
  INV_X1    g209(.A(new_n410), .ZN(new_n411));
  NAND3_X1  g210(.A1(new_n396), .A2(new_n340), .A3(new_n411), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n407), .A2(new_n409), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(KEYINPUT5), .ZN(new_n414));
  NAND2_X1  g213(.A1(new_n413), .A2(new_n414), .ZN(new_n415));
  NAND2_X1  g214(.A1(new_n415), .A2(new_n403), .ZN(new_n416));
  NAND2_X1  g215(.A1(new_n407), .A2(KEYINPUT5), .ZN(new_n417));
  INV_X1    g216(.A(KEYINPUT82), .ZN(new_n418));
  AOI21_X1  g217(.A(new_n418), .B1(new_n401), .B2(new_n411), .ZN(new_n419));
  NOR2_X1   g218(.A1(new_n401), .A2(KEYINPUT4), .ZN(new_n420));
  NOR2_X1   g219(.A1(new_n419), .A2(new_n420), .ZN(new_n421));
  NAND3_X1  g220(.A1(new_n401), .A2(new_n418), .A3(new_n411), .ZN(new_n422));
  AOI21_X1  g221(.A(new_n417), .B1(new_n421), .B2(new_n422), .ZN(new_n423));
  OAI21_X1  g222(.A(new_n405), .B1(new_n416), .B2(new_n423), .ZN(new_n424));
  XNOR2_X1  g223(.A(G1gat), .B(G29gat), .ZN(new_n425));
  XNOR2_X1  g224(.A(new_n425), .B(KEYINPUT0), .ZN(new_n426));
  XNOR2_X1  g225(.A(G57gat), .B(G85gat), .ZN(new_n427));
  XNOR2_X1  g226(.A(new_n426), .B(new_n427), .ZN(new_n428));
  NAND2_X1  g227(.A1(new_n424), .A2(new_n428), .ZN(new_n429));
  INV_X1    g228(.A(KEYINPUT6), .ZN(new_n430));
  INV_X1    g229(.A(new_n428), .ZN(new_n431));
  OAI211_X1 g230(.A(new_n431), .B(new_n405), .C1(new_n416), .C2(new_n423), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n429), .A2(new_n430), .A3(new_n432), .ZN(new_n433));
  NAND3_X1  g232(.A1(new_n424), .A2(KEYINPUT6), .A3(new_n428), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n433), .A2(new_n434), .ZN(new_n435));
  NAND2_X1  g234(.A1(new_n435), .A2(KEYINPUT90), .ZN(new_n436));
  INV_X1    g235(.A(KEYINPUT90), .ZN(new_n437));
  NAND2_X1  g236(.A1(new_n434), .A2(new_n437), .ZN(new_n438));
  NAND2_X1  g237(.A1(new_n436), .A2(new_n438), .ZN(new_n439));
  OAI21_X1  g238(.A(new_n396), .B1(new_n286), .B2(new_n291), .ZN(new_n440));
  NAND4_X1  g239(.A1(new_n235), .A2(new_n406), .A3(new_n247), .A4(new_n262), .ZN(new_n441));
  AND2_X1   g240(.A1(G227gat), .A2(G233gat), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n441), .A3(new_n442), .ZN(new_n443));
  INV_X1    g242(.A(KEYINPUT70), .ZN(new_n444));
  NAND2_X1  g243(.A1(new_n443), .A2(new_n444), .ZN(new_n445));
  NAND4_X1  g244(.A1(new_n440), .A2(new_n441), .A3(KEYINPUT70), .A4(new_n442), .ZN(new_n446));
  NAND2_X1  g245(.A1(new_n445), .A2(new_n446), .ZN(new_n447));
  NAND2_X1  g246(.A1(new_n447), .A2(KEYINPUT32), .ZN(new_n448));
  INV_X1    g247(.A(KEYINPUT33), .ZN(new_n449));
  NAND2_X1  g248(.A1(new_n447), .A2(new_n449), .ZN(new_n450));
  XOR2_X1   g249(.A(G15gat), .B(G43gat), .Z(new_n451));
  XNOR2_X1  g250(.A(G71gat), .B(G99gat), .ZN(new_n452));
  XNOR2_X1  g251(.A(new_n451), .B(new_n452), .ZN(new_n453));
  NAND3_X1  g252(.A1(new_n448), .A2(new_n450), .A3(new_n453), .ZN(new_n454));
  AOI21_X1  g253(.A(new_n442), .B1(new_n440), .B2(new_n441), .ZN(new_n455));
  INV_X1    g254(.A(KEYINPUT34), .ZN(new_n456));
  OR2_X1    g255(.A1(new_n455), .A2(new_n456), .ZN(new_n457));
  NAND2_X1  g256(.A1(new_n455), .A2(new_n456), .ZN(new_n458));
  NAND2_X1  g257(.A1(new_n457), .A2(new_n458), .ZN(new_n459));
  INV_X1    g258(.A(new_n459), .ZN(new_n460));
  INV_X1    g259(.A(KEYINPUT32), .ZN(new_n461));
  AOI21_X1  g260(.A(new_n461), .B1(new_n445), .B2(new_n446), .ZN(new_n462));
  AOI21_X1  g261(.A(KEYINPUT33), .B1(new_n445), .B2(new_n446), .ZN(new_n463));
  INV_X1    g262(.A(new_n453), .ZN(new_n464));
  OAI21_X1  g263(.A(new_n462), .B1(new_n463), .B2(new_n464), .ZN(new_n465));
  NAND3_X1  g264(.A1(new_n454), .A2(new_n460), .A3(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(new_n466), .ZN(new_n467));
  AOI21_X1  g266(.A(new_n460), .B1(new_n454), .B2(new_n465), .ZN(new_n468));
  NOR2_X1   g267(.A1(new_n467), .A2(new_n468), .ZN(new_n469));
  NAND4_X1  g268(.A1(new_n378), .A2(KEYINPUT91), .A3(new_n439), .A4(new_n469), .ZN(new_n470));
  INV_X1    g269(.A(KEYINPUT91), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n469), .A2(new_n439), .ZN(new_n472));
  OAI21_X1  g271(.A(new_n471), .B1(new_n377), .B2(new_n472), .ZN(new_n473));
  NAND2_X1  g272(.A1(new_n470), .A2(new_n473), .ZN(new_n474));
  NOR3_X1   g273(.A1(new_n462), .A2(new_n463), .A3(new_n464), .ZN(new_n475));
  AOI221_X4 g274(.A(new_n461), .B1(KEYINPUT33), .B2(new_n453), .C1(new_n445), .C2(new_n446), .ZN(new_n476));
  OAI21_X1  g275(.A(new_n459), .B1(new_n475), .B2(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n477), .A2(KEYINPUT71), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT71), .ZN(new_n479));
  NAND2_X1  g278(.A1(new_n468), .A2(new_n479), .ZN(new_n480));
  NAND4_X1  g279(.A1(new_n478), .A2(new_n480), .A3(new_n376), .A4(new_n466), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n304), .B1(new_n433), .B2(new_n434), .ZN(new_n482));
  INV_X1    g281(.A(KEYINPUT77), .ZN(new_n483));
  OAI21_X1  g282(.A(new_n483), .B1(new_n300), .B2(new_n302), .ZN(new_n484));
  AND3_X1   g283(.A1(new_n297), .A2(KEYINPUT75), .A3(new_n298), .ZN(new_n485));
  AOI21_X1  g284(.A(KEYINPUT75), .B1(new_n297), .B2(new_n298), .ZN(new_n486));
  OAI21_X1  g285(.A(new_n205), .B1(new_n485), .B2(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n303), .A2(KEYINPUT30), .ZN(new_n488));
  NAND3_X1  g287(.A1(new_n487), .A2(KEYINPUT77), .A3(new_n488), .ZN(new_n489));
  NAND3_X1  g288(.A1(new_n482), .A2(new_n484), .A3(new_n489), .ZN(new_n490));
  OR2_X1    g289(.A1(new_n481), .A2(new_n490), .ZN(new_n491));
  NAND2_X1  g290(.A1(new_n491), .A2(KEYINPUT35), .ZN(new_n492));
  NAND2_X1  g291(.A1(new_n474), .A2(new_n492), .ZN(new_n493));
  NAND2_X1  g292(.A1(new_n376), .A2(KEYINPUT87), .ZN(new_n494));
  INV_X1    g293(.A(KEYINPUT87), .ZN(new_n495));
  OAI211_X1 g294(.A(new_n495), .B(new_n357), .C1(new_n373), .C2(new_n375), .ZN(new_n496));
  NAND3_X1  g295(.A1(new_n490), .A2(new_n494), .A3(new_n496), .ZN(new_n497));
  INV_X1    g296(.A(new_n497), .ZN(new_n498));
  NAND3_X1  g297(.A1(new_n397), .A2(new_n401), .A3(new_n403), .ZN(new_n499));
  INV_X1    g298(.A(KEYINPUT88), .ZN(new_n500));
  XNOR2_X1  g299(.A(new_n499), .B(new_n500), .ZN(new_n501));
  NAND2_X1  g300(.A1(new_n413), .A2(new_n404), .ZN(new_n502));
  NAND3_X1  g301(.A1(new_n501), .A2(KEYINPUT39), .A3(new_n502), .ZN(new_n503));
  NOR2_X1   g302(.A1(new_n502), .A2(KEYINPUT39), .ZN(new_n504));
  NOR2_X1   g303(.A1(new_n504), .A2(new_n428), .ZN(new_n505));
  AND3_X1   g304(.A1(new_n503), .A2(KEYINPUT40), .A3(new_n505), .ZN(new_n506));
  AOI21_X1  g305(.A(KEYINPUT40), .B1(new_n503), .B2(new_n505), .ZN(new_n507));
  INV_X1    g306(.A(new_n429), .ZN(new_n508));
  NOR3_X1   g307(.A1(new_n506), .A2(new_n507), .A3(new_n508), .ZN(new_n509));
  OAI21_X1  g308(.A(G22gat), .B1(new_n367), .B2(new_n371), .ZN(new_n510));
  AOI21_X1  g309(.A(new_n312), .B1(new_n510), .B2(KEYINPUT85), .ZN(new_n511));
  NAND4_X1  g310(.A1(new_n511), .A2(new_n360), .A3(new_n372), .A4(new_n358), .ZN(new_n512));
  AOI22_X1  g311(.A1(new_n305), .A2(new_n509), .B1(new_n512), .B2(new_n357), .ZN(new_n513));
  XNOR2_X1  g312(.A(KEYINPUT89), .B(KEYINPUT38), .ZN(new_n514));
  INV_X1    g313(.A(new_n514), .ZN(new_n515));
  INV_X1    g314(.A(KEYINPUT37), .ZN(new_n516));
  AOI21_X1  g315(.A(new_n206), .B1(new_n301), .B2(new_n516), .ZN(new_n517));
  INV_X1    g316(.A(new_n517), .ZN(new_n518));
  AOI21_X1  g317(.A(new_n516), .B1(new_n296), .B2(new_n299), .ZN(new_n519));
  OAI21_X1  g318(.A(new_n515), .B1(new_n518), .B2(new_n519), .ZN(new_n520));
  NOR2_X1   g319(.A1(new_n301), .A2(new_n516), .ZN(new_n521));
  NOR2_X1   g320(.A1(new_n521), .A2(new_n515), .ZN(new_n522));
  AOI21_X1  g321(.A(new_n303), .B1(new_n522), .B2(new_n517), .ZN(new_n523));
  NAND4_X1  g322(.A1(new_n436), .A2(new_n520), .A3(new_n523), .A4(new_n438), .ZN(new_n524));
  NAND2_X1  g323(.A1(new_n513), .A2(new_n524), .ZN(new_n525));
  AND2_X1   g324(.A1(new_n466), .A2(KEYINPUT36), .ZN(new_n526));
  INV_X1    g325(.A(KEYINPUT72), .ZN(new_n527));
  NAND4_X1  g326(.A1(new_n526), .A2(new_n478), .A3(new_n480), .A4(new_n527), .ZN(new_n528));
  INV_X1    g327(.A(KEYINPUT36), .ZN(new_n529));
  OAI21_X1  g328(.A(new_n529), .B1(new_n467), .B2(new_n468), .ZN(new_n530));
  NAND2_X1  g329(.A1(new_n528), .A2(new_n530), .ZN(new_n531));
  NAND2_X1  g330(.A1(new_n454), .A2(new_n465), .ZN(new_n532));
  AOI21_X1  g331(.A(new_n479), .B1(new_n532), .B2(new_n459), .ZN(new_n533));
  AOI211_X1 g332(.A(KEYINPUT71), .B(new_n460), .C1(new_n454), .C2(new_n465), .ZN(new_n534));
  NOR2_X1   g333(.A1(new_n533), .A2(new_n534), .ZN(new_n535));
  AOI21_X1  g334(.A(new_n527), .B1(new_n535), .B2(new_n526), .ZN(new_n536));
  OAI21_X1  g335(.A(new_n525), .B1(new_n531), .B2(new_n536), .ZN(new_n537));
  OAI21_X1  g336(.A(new_n493), .B1(new_n498), .B2(new_n537), .ZN(new_n538));
  INV_X1    g337(.A(KEYINPUT94), .ZN(new_n539));
  XOR2_X1   g338(.A(G43gat), .B(G50gat), .Z(new_n540));
  INV_X1    g339(.A(KEYINPUT93), .ZN(new_n541));
  NAND2_X1  g340(.A1(new_n540), .A2(new_n541), .ZN(new_n542));
  XNOR2_X1  g341(.A(G43gat), .B(G50gat), .ZN(new_n543));
  NAND2_X1  g342(.A1(new_n543), .A2(KEYINPUT93), .ZN(new_n544));
  NAND3_X1  g343(.A1(new_n542), .A2(KEYINPUT15), .A3(new_n544), .ZN(new_n545));
  XNOR2_X1  g344(.A(KEYINPUT14), .B(G29gat), .ZN(new_n546));
  INV_X1    g345(.A(G36gat), .ZN(new_n547));
  NAND2_X1  g346(.A1(new_n546), .A2(new_n547), .ZN(new_n548));
  INV_X1    g347(.A(G29gat), .ZN(new_n549));
  NAND3_X1  g348(.A1(new_n549), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n550));
  NAND2_X1  g349(.A1(new_n548), .A2(new_n550), .ZN(new_n551));
  OAI21_X1  g350(.A(new_n539), .B1(new_n545), .B2(new_n551), .ZN(new_n552));
  INV_X1    g351(.A(new_n551), .ZN(new_n553));
  AND2_X1   g352(.A1(new_n544), .A2(KEYINPUT15), .ZN(new_n554));
  NAND4_X1  g353(.A1(new_n553), .A2(new_n554), .A3(KEYINPUT94), .A4(new_n542), .ZN(new_n555));
  NAND2_X1  g354(.A1(new_n552), .A2(new_n555), .ZN(new_n556));
  OAI211_X1 g355(.A(new_n545), .B(new_n551), .C1(KEYINPUT15), .C2(new_n543), .ZN(new_n557));
  NAND2_X1  g356(.A1(new_n556), .A2(new_n557), .ZN(new_n558));
  NAND2_X1  g357(.A1(new_n558), .A2(KEYINPUT95), .ZN(new_n559));
  INV_X1    g358(.A(KEYINPUT17), .ZN(new_n560));
  INV_X1    g359(.A(KEYINPUT95), .ZN(new_n561));
  NAND3_X1  g360(.A1(new_n556), .A2(new_n561), .A3(new_n557), .ZN(new_n562));
  NAND3_X1  g361(.A1(new_n559), .A2(new_n560), .A3(new_n562), .ZN(new_n563));
  XNOR2_X1  g362(.A(G15gat), .B(G22gat), .ZN(new_n564));
  INV_X1    g363(.A(KEYINPUT16), .ZN(new_n565));
  OAI21_X1  g364(.A(new_n564), .B1(new_n565), .B2(G1gat), .ZN(new_n566));
  OAI21_X1  g365(.A(new_n566), .B1(G1gat), .B2(new_n564), .ZN(new_n567));
  INV_X1    g366(.A(G8gat), .ZN(new_n568));
  XNOR2_X1  g367(.A(new_n567), .B(new_n568), .ZN(new_n569));
  OAI211_X1 g368(.A(new_n563), .B(new_n569), .C1(new_n560), .C2(new_n558), .ZN(new_n570));
  NAND2_X1  g369(.A1(new_n559), .A2(new_n562), .ZN(new_n571));
  INV_X1    g370(.A(new_n571), .ZN(new_n572));
  INV_X1    g371(.A(new_n569), .ZN(new_n573));
  NAND2_X1  g372(.A1(new_n572), .A2(new_n573), .ZN(new_n574));
  NAND2_X1  g373(.A1(G229gat), .A2(G233gat), .ZN(new_n575));
  NAND3_X1  g374(.A1(new_n570), .A2(new_n574), .A3(new_n575), .ZN(new_n576));
  INV_X1    g375(.A(KEYINPUT18), .ZN(new_n577));
  NAND2_X1  g376(.A1(new_n576), .A2(new_n577), .ZN(new_n578));
  NAND4_X1  g377(.A1(new_n570), .A2(new_n574), .A3(KEYINPUT18), .A4(new_n575), .ZN(new_n579));
  XOR2_X1   g378(.A(new_n575), .B(KEYINPUT13), .Z(new_n580));
  NOR2_X1   g379(.A1(new_n572), .A2(new_n573), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n571), .A2(new_n569), .ZN(new_n582));
  OAI21_X1  g381(.A(new_n580), .B1(new_n581), .B2(new_n582), .ZN(new_n583));
  NAND3_X1  g382(.A1(new_n578), .A2(new_n579), .A3(new_n583), .ZN(new_n584));
  XNOR2_X1  g383(.A(G113gat), .B(G141gat), .ZN(new_n585));
  XNOR2_X1  g384(.A(G169gat), .B(G197gat), .ZN(new_n586));
  XNOR2_X1  g385(.A(new_n585), .B(new_n586), .ZN(new_n587));
  XNOR2_X1  g386(.A(KEYINPUT92), .B(KEYINPUT11), .ZN(new_n588));
  XNOR2_X1  g387(.A(new_n587), .B(new_n588), .ZN(new_n589));
  XOR2_X1   g388(.A(new_n589), .B(KEYINPUT12), .Z(new_n590));
  NAND2_X1  g389(.A1(new_n584), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n590), .ZN(new_n592));
  NAND4_X1  g391(.A1(new_n578), .A2(new_n579), .A3(new_n583), .A4(new_n592), .ZN(new_n593));
  NAND2_X1  g392(.A1(new_n591), .A2(new_n593), .ZN(new_n594));
  AND2_X1   g393(.A1(new_n538), .A2(new_n594), .ZN(new_n595));
  AND2_X1   g394(.A1(G232gat), .A2(G233gat), .ZN(new_n596));
  NAND2_X1  g395(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n597));
  NAND2_X1  g396(.A1(G85gat), .A2(G92gat), .ZN(new_n598));
  XNOR2_X1  g397(.A(new_n598), .B(KEYINPUT7), .ZN(new_n599));
  NAND2_X1  g398(.A1(G99gat), .A2(G106gat), .ZN(new_n600));
  INV_X1    g399(.A(G85gat), .ZN(new_n601));
  INV_X1    g400(.A(G92gat), .ZN(new_n602));
  AOI22_X1  g401(.A1(KEYINPUT8), .A2(new_n600), .B1(new_n601), .B2(new_n602), .ZN(new_n603));
  NAND2_X1  g402(.A1(new_n599), .A2(new_n603), .ZN(new_n604));
  XNOR2_X1  g403(.A(G99gat), .B(G106gat), .ZN(new_n605));
  XNOR2_X1  g404(.A(new_n604), .B(new_n605), .ZN(new_n606));
  INV_X1    g405(.A(new_n606), .ZN(new_n607));
  OAI21_X1  g406(.A(new_n597), .B1(new_n571), .B2(new_n607), .ZN(new_n608));
  INV_X1    g407(.A(new_n558), .ZN(new_n609));
  AOI21_X1  g408(.A(new_n606), .B1(new_n609), .B2(KEYINPUT17), .ZN(new_n610));
  NAND2_X1  g409(.A1(new_n563), .A2(new_n610), .ZN(new_n611));
  NAND2_X1  g410(.A1(new_n611), .A2(KEYINPUT103), .ZN(new_n612));
  INV_X1    g411(.A(KEYINPUT103), .ZN(new_n613));
  NAND3_X1  g412(.A1(new_n563), .A2(new_n610), .A3(new_n613), .ZN(new_n614));
  AOI21_X1  g413(.A(new_n608), .B1(new_n612), .B2(new_n614), .ZN(new_n615));
  XNOR2_X1  g414(.A(G190gat), .B(G218gat), .ZN(new_n616));
  INV_X1    g415(.A(new_n616), .ZN(new_n617));
  OAI21_X1  g416(.A(KEYINPUT105), .B1(new_n615), .B2(new_n617), .ZN(new_n618));
  INV_X1    g417(.A(new_n608), .ZN(new_n619));
  INV_X1    g418(.A(new_n614), .ZN(new_n620));
  AOI21_X1  g419(.A(new_n613), .B1(new_n563), .B2(new_n610), .ZN(new_n621));
  OAI21_X1  g420(.A(new_n619), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  INV_X1    g421(.A(KEYINPUT105), .ZN(new_n623));
  NAND3_X1  g422(.A1(new_n622), .A2(new_n623), .A3(new_n616), .ZN(new_n624));
  AND2_X1   g423(.A1(new_n618), .A2(new_n624), .ZN(new_n625));
  NAND2_X1  g424(.A1(new_n615), .A2(new_n617), .ZN(new_n626));
  INV_X1    g425(.A(KEYINPUT104), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n596), .A2(KEYINPUT41), .ZN(new_n628));
  XNOR2_X1  g427(.A(new_n628), .B(G134gat), .ZN(new_n629));
  XNOR2_X1  g428(.A(new_n629), .B(new_n323), .ZN(new_n630));
  INV_X1    g429(.A(new_n630), .ZN(new_n631));
  OAI211_X1 g430(.A(new_n625), .B(new_n626), .C1(new_n627), .C2(new_n631), .ZN(new_n632));
  NAND3_X1  g431(.A1(new_n618), .A2(new_n624), .A3(new_n626), .ZN(new_n633));
  NAND3_X1  g432(.A1(new_n618), .A2(new_n624), .A3(new_n627), .ZN(new_n634));
  NAND3_X1  g433(.A1(new_n633), .A2(new_n634), .A3(new_n630), .ZN(new_n635));
  NAND2_X1  g434(.A1(new_n632), .A2(new_n635), .ZN(new_n636));
  INV_X1    g435(.A(new_n636), .ZN(new_n637));
  XNOR2_X1  g436(.A(KEYINPUT101), .B(KEYINPUT19), .ZN(new_n638));
  INV_X1    g437(.A(G57gat), .ZN(new_n639));
  INV_X1    g438(.A(G64gat), .ZN(new_n640));
  NAND2_X1  g439(.A1(new_n639), .A2(new_n640), .ZN(new_n641));
  NAND2_X1  g440(.A1(G57gat), .A2(G64gat), .ZN(new_n642));
  INV_X1    g441(.A(G71gat), .ZN(new_n643));
  INV_X1    g442(.A(G78gat), .ZN(new_n644));
  NOR2_X1   g443(.A1(new_n643), .A2(new_n644), .ZN(new_n645));
  OAI211_X1 g444(.A(new_n641), .B(new_n642), .C1(new_n645), .C2(KEYINPUT9), .ZN(new_n646));
  OAI21_X1  g445(.A(KEYINPUT96), .B1(G71gat), .B2(G78gat), .ZN(new_n647));
  INV_X1    g446(.A(KEYINPUT96), .ZN(new_n648));
  NAND3_X1  g447(.A1(new_n648), .A2(new_n643), .A3(new_n644), .ZN(new_n649));
  AOI21_X1  g448(.A(new_n645), .B1(new_n647), .B2(new_n649), .ZN(new_n650));
  OAI21_X1  g449(.A(new_n646), .B1(new_n650), .B2(KEYINPUT97), .ZN(new_n651));
  INV_X1    g450(.A(KEYINPUT97), .ZN(new_n652));
  AOI211_X1 g451(.A(new_n652), .B(new_n645), .C1(new_n647), .C2(new_n649), .ZN(new_n653));
  NOR2_X1   g452(.A1(new_n651), .A2(new_n653), .ZN(new_n654));
  INV_X1    g453(.A(KEYINPUT98), .ZN(new_n655));
  XNOR2_X1  g454(.A(new_n654), .B(new_n655), .ZN(new_n656));
  INV_X1    g455(.A(KEYINPUT99), .ZN(new_n657));
  NAND2_X1  g456(.A1(new_n657), .A2(G57gat), .ZN(new_n658));
  XNOR2_X1  g457(.A(new_n658), .B(new_n640), .ZN(new_n659));
  NOR2_X1   g458(.A1(G71gat), .A2(G78gat), .ZN(new_n660));
  AOI21_X1  g459(.A(new_n645), .B1(KEYINPUT9), .B2(new_n660), .ZN(new_n661));
  NOR2_X1   g460(.A1(new_n659), .A2(new_n661), .ZN(new_n662));
  INV_X1    g461(.A(new_n662), .ZN(new_n663));
  NAND2_X1  g462(.A1(new_n656), .A2(new_n663), .ZN(new_n664));
  NAND2_X1  g463(.A1(new_n664), .A2(KEYINPUT100), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT100), .ZN(new_n666));
  NAND3_X1  g465(.A1(new_n656), .A2(new_n666), .A3(new_n663), .ZN(new_n667));
  NAND2_X1  g466(.A1(new_n665), .A2(new_n667), .ZN(new_n668));
  NAND2_X1  g467(.A1(new_n668), .A2(KEYINPUT21), .ZN(new_n669));
  INV_X1    g468(.A(KEYINPUT102), .ZN(new_n670));
  NAND3_X1  g469(.A1(new_n669), .A2(new_n670), .A3(new_n569), .ZN(new_n671));
  INV_X1    g470(.A(new_n671), .ZN(new_n672));
  AOI21_X1  g471(.A(new_n670), .B1(new_n669), .B2(new_n569), .ZN(new_n673));
  OAI21_X1  g472(.A(new_n638), .B1(new_n672), .B2(new_n673), .ZN(new_n674));
  INV_X1    g473(.A(new_n673), .ZN(new_n675));
  INV_X1    g474(.A(new_n638), .ZN(new_n676));
  NAND3_X1  g475(.A1(new_n675), .A2(new_n671), .A3(new_n676), .ZN(new_n677));
  NAND2_X1  g476(.A1(new_n674), .A2(new_n677), .ZN(new_n678));
  NAND2_X1  g477(.A1(G231gat), .A2(G233gat), .ZN(new_n679));
  INV_X1    g478(.A(new_n679), .ZN(new_n680));
  OAI21_X1  g479(.A(new_n680), .B1(new_n668), .B2(KEYINPUT21), .ZN(new_n681));
  AND3_X1   g480(.A1(new_n656), .A2(new_n666), .A3(new_n663), .ZN(new_n682));
  AOI21_X1  g481(.A(new_n666), .B1(new_n656), .B2(new_n663), .ZN(new_n683));
  NOR2_X1   g482(.A1(new_n682), .A2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(KEYINPUT21), .ZN(new_n685));
  NAND3_X1  g484(.A1(new_n684), .A2(new_n685), .A3(new_n679), .ZN(new_n686));
  XNOR2_X1  g485(.A(G127gat), .B(G155gat), .ZN(new_n687));
  XOR2_X1   g486(.A(new_n687), .B(KEYINPUT20), .Z(new_n688));
  INV_X1    g487(.A(new_n688), .ZN(new_n689));
  NAND3_X1  g488(.A1(new_n681), .A2(new_n686), .A3(new_n689), .ZN(new_n690));
  INV_X1    g489(.A(new_n690), .ZN(new_n691));
  XOR2_X1   g490(.A(G183gat), .B(G211gat), .Z(new_n692));
  AOI21_X1  g491(.A(new_n689), .B1(new_n681), .B2(new_n686), .ZN(new_n693));
  NOR3_X1   g492(.A1(new_n691), .A2(new_n692), .A3(new_n693), .ZN(new_n694));
  INV_X1    g493(.A(new_n692), .ZN(new_n695));
  INV_X1    g494(.A(new_n686), .ZN(new_n696));
  AOI21_X1  g495(.A(new_n679), .B1(new_n684), .B2(new_n685), .ZN(new_n697));
  OAI21_X1  g496(.A(new_n688), .B1(new_n696), .B2(new_n697), .ZN(new_n698));
  AOI21_X1  g497(.A(new_n695), .B1(new_n698), .B2(new_n690), .ZN(new_n699));
  OAI21_X1  g498(.A(new_n678), .B1(new_n694), .B2(new_n699), .ZN(new_n700));
  OAI21_X1  g499(.A(new_n692), .B1(new_n691), .B2(new_n693), .ZN(new_n701));
  NAND3_X1  g500(.A1(new_n698), .A2(new_n690), .A3(new_n695), .ZN(new_n702));
  NAND4_X1  g501(.A1(new_n701), .A2(new_n702), .A3(new_n677), .A4(new_n674), .ZN(new_n703));
  NAND2_X1  g502(.A1(new_n700), .A2(new_n703), .ZN(new_n704));
  INV_X1    g503(.A(new_n704), .ZN(new_n705));
  INV_X1    g504(.A(G230gat), .ZN(new_n706));
  INV_X1    g505(.A(G233gat), .ZN(new_n707));
  NOR2_X1   g506(.A1(new_n706), .A2(new_n707), .ZN(new_n708));
  INV_X1    g507(.A(new_n708), .ZN(new_n709));
  OAI21_X1  g508(.A(new_n607), .B1(new_n682), .B2(new_n683), .ZN(new_n710));
  NAND2_X1  g509(.A1(new_n664), .A2(new_n606), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT10), .B1(new_n710), .B2(new_n711), .ZN(new_n712));
  AND2_X1   g511(.A1(new_n606), .A2(KEYINPUT10), .ZN(new_n713));
  AND2_X1   g512(.A1(new_n668), .A2(new_n713), .ZN(new_n714));
  OAI21_X1  g513(.A(new_n709), .B1(new_n712), .B2(new_n714), .ZN(new_n715));
  INV_X1    g514(.A(new_n711), .ZN(new_n716));
  AOI21_X1  g515(.A(new_n716), .B1(new_n668), .B2(new_n607), .ZN(new_n717));
  NAND2_X1  g516(.A1(new_n717), .A2(new_n708), .ZN(new_n718));
  NAND2_X1  g517(.A1(new_n715), .A2(new_n718), .ZN(new_n719));
  XNOR2_X1  g518(.A(G120gat), .B(G148gat), .ZN(new_n720));
  XNOR2_X1  g519(.A(new_n720), .B(KEYINPUT106), .ZN(new_n721));
  XOR2_X1   g520(.A(G176gat), .B(G204gat), .Z(new_n722));
  XNOR2_X1  g521(.A(new_n721), .B(new_n722), .ZN(new_n723));
  OR2_X1    g522(.A1(new_n719), .A2(new_n723), .ZN(new_n724));
  NAND2_X1  g523(.A1(new_n719), .A2(new_n723), .ZN(new_n725));
  AND2_X1   g524(.A1(new_n724), .A2(new_n725), .ZN(new_n726));
  NAND4_X1  g525(.A1(new_n595), .A2(new_n637), .A3(new_n705), .A4(new_n726), .ZN(new_n727));
  NOR2_X1   g526(.A1(new_n727), .A2(new_n435), .ZN(new_n728));
  XOR2_X1   g527(.A(new_n728), .B(G1gat), .Z(G1324gat));
  NOR2_X1   g528(.A1(new_n727), .A2(new_n306), .ZN(new_n730));
  XNOR2_X1  g529(.A(KEYINPUT107), .B(KEYINPUT16), .ZN(new_n731));
  XNOR2_X1  g530(.A(new_n731), .B(new_n568), .ZN(new_n732));
  NAND2_X1  g531(.A1(new_n730), .A2(new_n732), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n568), .B2(new_n730), .ZN(new_n734));
  MUX2_X1   g533(.A(new_n733), .B(new_n734), .S(KEYINPUT42), .Z(G1325gat));
  NAND3_X1  g534(.A1(new_n526), .A2(new_n478), .A3(new_n480), .ZN(new_n736));
  NAND2_X1  g535(.A1(new_n736), .A2(KEYINPUT72), .ZN(new_n737));
  NAND3_X1  g536(.A1(new_n737), .A2(new_n530), .A3(new_n528), .ZN(new_n738));
  OAI21_X1  g537(.A(G15gat), .B1(new_n727), .B2(new_n738), .ZN(new_n739));
  INV_X1    g538(.A(new_n469), .ZN(new_n740));
  OR2_X1    g539(.A1(new_n740), .A2(G15gat), .ZN(new_n741));
  OAI21_X1  g540(.A(new_n739), .B1(new_n727), .B2(new_n741), .ZN(G1326gat));
  NAND2_X1  g541(.A1(new_n494), .A2(new_n496), .ZN(new_n743));
  OR3_X1    g542(.A1(new_n727), .A2(KEYINPUT108), .A3(new_n743), .ZN(new_n744));
  OAI21_X1  g543(.A(KEYINPUT108), .B1(new_n727), .B2(new_n743), .ZN(new_n745));
  NAND2_X1  g544(.A1(new_n744), .A2(new_n745), .ZN(new_n746));
  XNOR2_X1  g545(.A(KEYINPUT43), .B(G22gat), .ZN(new_n747));
  XNOR2_X1  g546(.A(new_n746), .B(new_n747), .ZN(G1327gat));
  NAND2_X1  g547(.A1(new_n724), .A2(new_n725), .ZN(new_n749));
  NOR2_X1   g548(.A1(new_n705), .A2(new_n749), .ZN(new_n750));
  INV_X1    g549(.A(new_n750), .ZN(new_n751));
  NOR2_X1   g550(.A1(new_n751), .A2(new_n637), .ZN(new_n752));
  NAND2_X1  g551(.A1(new_n595), .A2(new_n752), .ZN(new_n753));
  INV_X1    g552(.A(new_n753), .ZN(new_n754));
  INV_X1    g553(.A(new_n435), .ZN(new_n755));
  NAND3_X1  g554(.A1(new_n754), .A2(new_n549), .A3(new_n755), .ZN(new_n756));
  XNOR2_X1  g555(.A(new_n756), .B(KEYINPUT45), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT44), .ZN(new_n758));
  AOI22_X1  g557(.A1(new_n470), .A2(new_n473), .B1(new_n491), .B2(KEYINPUT35), .ZN(new_n759));
  INV_X1    g558(.A(KEYINPUT110), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT109), .ZN(new_n761));
  NAND2_X1  g560(.A1(new_n497), .A2(new_n761), .ZN(new_n762));
  NAND4_X1  g561(.A1(new_n490), .A2(new_n494), .A3(KEYINPUT109), .A4(new_n496), .ZN(new_n763));
  NAND2_X1  g562(.A1(new_n762), .A2(new_n763), .ZN(new_n764));
  OAI21_X1  g563(.A(new_n760), .B1(new_n537), .B2(new_n764), .ZN(new_n765));
  AND2_X1   g564(.A1(new_n762), .A2(new_n763), .ZN(new_n766));
  NAND4_X1  g565(.A1(new_n766), .A2(KEYINPUT110), .A3(new_n525), .A4(new_n738), .ZN(new_n767));
  AOI21_X1  g566(.A(new_n759), .B1(new_n765), .B2(new_n767), .ZN(new_n768));
  OAI21_X1  g567(.A(new_n758), .B1(new_n768), .B2(new_n637), .ZN(new_n769));
  NAND3_X1  g568(.A1(new_n538), .A2(KEYINPUT44), .A3(new_n636), .ZN(new_n770));
  AND2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n594), .ZN(new_n772));
  NOR2_X1   g571(.A1(new_n751), .A2(new_n772), .ZN(new_n773));
  NAND2_X1  g572(.A1(new_n771), .A2(new_n773), .ZN(new_n774));
  OAI21_X1  g573(.A(G29gat), .B1(new_n774), .B2(new_n435), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n757), .A2(new_n775), .ZN(G1328gat));
  NOR3_X1   g575(.A1(new_n753), .A2(G36gat), .A3(new_n306), .ZN(new_n777));
  XNOR2_X1  g576(.A(new_n777), .B(KEYINPUT46), .ZN(new_n778));
  OAI21_X1  g577(.A(G36gat), .B1(new_n774), .B2(new_n306), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n778), .A2(new_n779), .ZN(G1329gat));
  INV_X1    g579(.A(new_n774), .ZN(new_n781));
  INV_X1    g580(.A(new_n738), .ZN(new_n782));
  NAND3_X1  g581(.A1(new_n781), .A2(G43gat), .A3(new_n782), .ZN(new_n783));
  INV_X1    g582(.A(G43gat), .ZN(new_n784));
  OAI21_X1  g583(.A(new_n784), .B1(new_n753), .B2(new_n740), .ZN(new_n785));
  NAND2_X1  g584(.A1(new_n783), .A2(new_n785), .ZN(new_n786));
  NAND2_X1  g585(.A1(new_n786), .A2(KEYINPUT47), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT47), .ZN(new_n788));
  NAND3_X1  g587(.A1(new_n783), .A2(new_n788), .A3(new_n785), .ZN(new_n789));
  NAND2_X1  g588(.A1(new_n787), .A2(new_n789), .ZN(G1330gat));
  OAI21_X1  g589(.A(G50gat), .B1(new_n774), .B2(new_n376), .ZN(new_n791));
  NOR3_X1   g590(.A1(new_n753), .A2(G50gat), .A3(new_n743), .ZN(new_n792));
  INV_X1    g591(.A(new_n792), .ZN(new_n793));
  NAND3_X1  g592(.A1(new_n791), .A2(KEYINPUT48), .A3(new_n793), .ZN(new_n794));
  INV_X1    g593(.A(new_n743), .ZN(new_n795));
  NAND2_X1  g594(.A1(new_n781), .A2(new_n795), .ZN(new_n796));
  AOI21_X1  g595(.A(new_n792), .B1(new_n796), .B2(G50gat), .ZN(new_n797));
  OAI21_X1  g596(.A(new_n794), .B1(new_n797), .B2(KEYINPUT48), .ZN(G1331gat));
  NAND4_X1  g597(.A1(new_n637), .A2(new_n772), .A3(new_n705), .A4(new_n749), .ZN(new_n799));
  OR3_X1    g598(.A1(new_n768), .A2(KEYINPUT111), .A3(new_n799), .ZN(new_n800));
  OAI21_X1  g599(.A(KEYINPUT111), .B1(new_n768), .B2(new_n799), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NOR2_X1   g601(.A1(new_n802), .A2(new_n435), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(new_n639), .ZN(G1332gat));
  XOR2_X1   g603(.A(new_n305), .B(KEYINPUT112), .Z(new_n805));
  NOR2_X1   g604(.A1(new_n802), .A2(new_n805), .ZN(new_n806));
  NOR2_X1   g605(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n807));
  AND2_X1   g606(.A1(KEYINPUT49), .A2(G64gat), .ZN(new_n808));
  OAI21_X1  g607(.A(new_n806), .B1(new_n807), .B2(new_n808), .ZN(new_n809));
  OAI21_X1  g608(.A(new_n809), .B1(new_n806), .B2(new_n807), .ZN(G1333gat));
  OAI21_X1  g609(.A(G71gat), .B1(new_n802), .B2(new_n738), .ZN(new_n811));
  NAND2_X1  g610(.A1(new_n469), .A2(new_n643), .ZN(new_n812));
  OAI21_X1  g611(.A(new_n811), .B1(new_n802), .B2(new_n812), .ZN(new_n813));
  XNOR2_X1  g612(.A(KEYINPUT113), .B(KEYINPUT50), .ZN(new_n814));
  XNOR2_X1  g613(.A(new_n813), .B(new_n814), .ZN(G1334gat));
  NOR2_X1   g614(.A1(new_n802), .A2(new_n743), .ZN(new_n816));
  XNOR2_X1  g615(.A(new_n816), .B(new_n644), .ZN(G1335gat));
  NOR3_X1   g616(.A1(new_n705), .A2(new_n594), .A3(new_n726), .ZN(new_n818));
  NAND2_X1  g617(.A1(new_n771), .A2(new_n818), .ZN(new_n819));
  OAI21_X1  g618(.A(G85gat), .B1(new_n819), .B2(new_n435), .ZN(new_n820));
  AND2_X1   g619(.A1(new_n513), .A2(new_n524), .ZN(new_n821));
  AND2_X1   g620(.A1(new_n528), .A2(new_n530), .ZN(new_n822));
  AOI21_X1  g621(.A(new_n821), .B1(new_n822), .B2(new_n737), .ZN(new_n823));
  AOI21_X1  g622(.A(KEYINPUT110), .B1(new_n823), .B2(new_n766), .ZN(new_n824));
  NOR3_X1   g623(.A1(new_n537), .A2(new_n760), .A3(new_n764), .ZN(new_n825));
  OAI21_X1  g624(.A(new_n493), .B1(new_n824), .B2(new_n825), .ZN(new_n826));
  NOR2_X1   g625(.A1(new_n705), .A2(new_n594), .ZN(new_n827));
  NAND3_X1  g626(.A1(new_n826), .A2(new_n636), .A3(new_n827), .ZN(new_n828));
  INV_X1    g627(.A(KEYINPUT51), .ZN(new_n829));
  NAND2_X1  g628(.A1(new_n828), .A2(new_n829), .ZN(new_n830));
  NAND4_X1  g629(.A1(new_n826), .A2(KEYINPUT51), .A3(new_n636), .A4(new_n827), .ZN(new_n831));
  NAND3_X1  g630(.A1(new_n830), .A2(KEYINPUT114), .A3(new_n831), .ZN(new_n832));
  INV_X1    g631(.A(KEYINPUT114), .ZN(new_n833));
  NAND3_X1  g632(.A1(new_n828), .A2(new_n833), .A3(new_n829), .ZN(new_n834));
  NAND3_X1  g633(.A1(new_n832), .A2(new_n749), .A3(new_n834), .ZN(new_n835));
  NAND2_X1  g634(.A1(new_n755), .A2(new_n601), .ZN(new_n836));
  OAI21_X1  g635(.A(new_n820), .B1(new_n835), .B2(new_n836), .ZN(G1336gat));
  INV_X1    g636(.A(new_n805), .ZN(new_n838));
  NAND3_X1  g637(.A1(new_n838), .A2(new_n749), .A3(new_n602), .ZN(new_n839));
  INV_X1    g638(.A(new_n839), .ZN(new_n840));
  NAND3_X1  g639(.A1(new_n832), .A2(new_n834), .A3(new_n840), .ZN(new_n841));
  NAND4_X1  g640(.A1(new_n769), .A2(new_n770), .A3(new_n838), .A4(new_n818), .ZN(new_n842));
  AOI21_X1  g641(.A(KEYINPUT52), .B1(new_n842), .B2(G92gat), .ZN(new_n843));
  NAND2_X1  g642(.A1(new_n841), .A2(new_n843), .ZN(new_n844));
  NAND4_X1  g643(.A1(new_n769), .A2(new_n305), .A3(new_n770), .A4(new_n818), .ZN(new_n845));
  AND2_X1   g644(.A1(new_n845), .A2(G92gat), .ZN(new_n846));
  XOR2_X1   g645(.A(new_n839), .B(KEYINPUT115), .Z(new_n847));
  AOI21_X1  g646(.A(new_n847), .B1(new_n830), .B2(new_n831), .ZN(new_n848));
  OAI21_X1  g647(.A(KEYINPUT52), .B1(new_n846), .B2(new_n848), .ZN(new_n849));
  NAND2_X1  g648(.A1(new_n844), .A2(new_n849), .ZN(new_n850));
  NAND2_X1  g649(.A1(new_n850), .A2(KEYINPUT116), .ZN(new_n851));
  INV_X1    g650(.A(KEYINPUT116), .ZN(new_n852));
  NAND3_X1  g651(.A1(new_n844), .A2(new_n849), .A3(new_n852), .ZN(new_n853));
  NAND2_X1  g652(.A1(new_n851), .A2(new_n853), .ZN(G1337gat));
  OAI21_X1  g653(.A(G99gat), .B1(new_n819), .B2(new_n738), .ZN(new_n855));
  OR2_X1    g654(.A1(new_n740), .A2(G99gat), .ZN(new_n856));
  OAI21_X1  g655(.A(new_n855), .B1(new_n835), .B2(new_n856), .ZN(G1338gat));
  OAI21_X1  g656(.A(G106gat), .B1(new_n819), .B2(new_n376), .ZN(new_n858));
  NOR3_X1   g657(.A1(new_n726), .A2(G106gat), .A3(new_n376), .ZN(new_n859));
  NAND3_X1  g658(.A1(new_n832), .A2(new_n834), .A3(new_n859), .ZN(new_n860));
  AOI21_X1  g659(.A(KEYINPUT53), .B1(new_n858), .B2(new_n860), .ZN(new_n861));
  OAI21_X1  g660(.A(G106gat), .B1(new_n819), .B2(new_n743), .ZN(new_n862));
  INV_X1    g661(.A(KEYINPUT53), .ZN(new_n863));
  NAND2_X1  g662(.A1(new_n830), .A2(new_n831), .ZN(new_n864));
  XNOR2_X1  g663(.A(new_n859), .B(KEYINPUT117), .ZN(new_n865));
  AOI21_X1  g664(.A(new_n863), .B1(new_n864), .B2(new_n865), .ZN(new_n866));
  AOI21_X1  g665(.A(new_n861), .B1(new_n862), .B2(new_n866), .ZN(G1339gat));
  NOR4_X1   g666(.A1(new_n636), .A2(new_n704), .A3(new_n594), .A4(new_n749), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n668), .A2(new_n713), .ZN(new_n869));
  OAI211_X1 g668(.A(new_n708), .B(new_n869), .C1(new_n717), .C2(KEYINPUT10), .ZN(new_n870));
  NAND3_X1  g669(.A1(new_n715), .A2(new_n870), .A3(KEYINPUT54), .ZN(new_n871));
  INV_X1    g670(.A(KEYINPUT54), .ZN(new_n872));
  OAI211_X1 g671(.A(new_n872), .B(new_n709), .C1(new_n712), .C2(new_n714), .ZN(new_n873));
  NAND4_X1  g672(.A1(new_n871), .A2(KEYINPUT55), .A3(new_n723), .A4(new_n873), .ZN(new_n874));
  AND2_X1   g673(.A1(new_n874), .A2(new_n724), .ZN(new_n875));
  NOR3_X1   g674(.A1(new_n581), .A2(new_n582), .A3(new_n580), .ZN(new_n876));
  AOI21_X1  g675(.A(new_n575), .B1(new_n570), .B2(new_n574), .ZN(new_n877));
  OAI21_X1  g676(.A(new_n589), .B1(new_n876), .B2(new_n877), .ZN(new_n878));
  NAND2_X1  g677(.A1(new_n593), .A2(new_n878), .ZN(new_n879));
  NAND3_X1  g678(.A1(new_n871), .A2(new_n723), .A3(new_n873), .ZN(new_n880));
  INV_X1    g679(.A(KEYINPUT55), .ZN(new_n881));
  AOI21_X1  g680(.A(new_n879), .B1(new_n880), .B2(new_n881), .ZN(new_n882));
  INV_X1    g681(.A(new_n635), .ZN(new_n883));
  AOI21_X1  g682(.A(new_n633), .B1(new_n634), .B2(new_n630), .ZN(new_n884));
  OAI211_X1 g683(.A(new_n875), .B(new_n882), .C1(new_n883), .C2(new_n884), .ZN(new_n885));
  AOI22_X1  g684(.A1(new_n880), .A2(new_n881), .B1(new_n591), .B2(new_n593), .ZN(new_n886));
  INV_X1    g685(.A(new_n879), .ZN(new_n887));
  AOI22_X1  g686(.A1(new_n875), .A2(new_n886), .B1(new_n749), .B2(new_n887), .ZN(new_n888));
  OAI21_X1  g687(.A(new_n885), .B1(new_n888), .B2(new_n636), .ZN(new_n889));
  AOI21_X1  g688(.A(new_n868), .B1(new_n889), .B2(new_n704), .ZN(new_n890));
  NOR2_X1   g689(.A1(new_n890), .A2(new_n435), .ZN(new_n891));
  INV_X1    g690(.A(new_n481), .ZN(new_n892));
  NAND2_X1  g691(.A1(new_n891), .A2(new_n892), .ZN(new_n893));
  NOR2_X1   g692(.A1(new_n893), .A2(new_n838), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n594), .A2(new_n380), .ZN(new_n895));
  XOR2_X1   g694(.A(new_n895), .B(KEYINPUT118), .Z(new_n896));
  NAND2_X1  g695(.A1(new_n894), .A2(new_n896), .ZN(new_n897));
  NOR3_X1   g696(.A1(new_n890), .A2(new_n795), .A3(new_n740), .ZN(new_n898));
  NAND3_X1  g697(.A1(new_n898), .A2(new_n755), .A3(new_n805), .ZN(new_n899));
  OAI21_X1  g698(.A(G113gat), .B1(new_n899), .B2(new_n772), .ZN(new_n900));
  NAND2_X1  g699(.A1(new_n897), .A2(new_n900), .ZN(G1340gat));
  AOI21_X1  g700(.A(G120gat), .B1(new_n894), .B2(new_n749), .ZN(new_n902));
  NOR3_X1   g701(.A1(new_n899), .A2(new_n393), .A3(new_n726), .ZN(new_n903));
  NOR2_X1   g702(.A1(new_n902), .A2(new_n903), .ZN(G1341gat));
  NAND3_X1  g703(.A1(new_n894), .A2(new_n387), .A3(new_n705), .ZN(new_n905));
  OAI21_X1  g704(.A(G127gat), .B1(new_n899), .B2(new_n704), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(G1342gat));
  NAND2_X1  g706(.A1(new_n636), .A2(new_n306), .ZN(new_n908));
  XNOR2_X1  g707(.A(new_n908), .B(KEYINPUT119), .ZN(new_n909));
  OR3_X1    g708(.A1(new_n893), .A2(G134gat), .A3(new_n909), .ZN(new_n910));
  OR2_X1    g709(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n911));
  OAI21_X1  g710(.A(G134gat), .B1(new_n899), .B2(new_n637), .ZN(new_n912));
  NAND2_X1  g711(.A1(new_n910), .A2(KEYINPUT56), .ZN(new_n913));
  NAND3_X1  g712(.A1(new_n911), .A2(new_n912), .A3(new_n913), .ZN(G1343gat));
  NAND2_X1  g713(.A1(new_n880), .A2(new_n881), .ZN(new_n915));
  NAND2_X1  g714(.A1(new_n915), .A2(new_n594), .ZN(new_n916));
  NAND2_X1  g715(.A1(new_n874), .A2(new_n724), .ZN(new_n917));
  OAI22_X1  g716(.A1(new_n916), .A2(new_n917), .B1(new_n726), .B2(new_n879), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n918), .A2(new_n637), .ZN(new_n919));
  OR2_X1    g718(.A1(new_n919), .A2(KEYINPUT120), .ZN(new_n920));
  INV_X1    g719(.A(new_n885), .ZN(new_n921));
  AOI21_X1  g720(.A(new_n921), .B1(new_n919), .B2(KEYINPUT120), .ZN(new_n922));
  AOI21_X1  g721(.A(new_n705), .B1(new_n920), .B2(new_n922), .ZN(new_n923));
  OAI21_X1  g722(.A(new_n795), .B1(new_n923), .B2(new_n868), .ZN(new_n924));
  NAND2_X1  g723(.A1(new_n924), .A2(KEYINPUT57), .ZN(new_n925));
  INV_X1    g724(.A(KEYINPUT57), .ZN(new_n926));
  INV_X1    g725(.A(new_n376), .ZN(new_n927));
  AOI21_X1  g726(.A(new_n705), .B1(new_n919), .B2(new_n885), .ZN(new_n928));
  OAI211_X1 g727(.A(new_n926), .B(new_n927), .C1(new_n928), .C2(new_n868), .ZN(new_n929));
  NOR3_X1   g728(.A1(new_n782), .A2(new_n435), .A3(new_n838), .ZN(new_n930));
  NAND2_X1  g729(.A1(new_n929), .A2(new_n930), .ZN(new_n931));
  INV_X1    g730(.A(new_n931), .ZN(new_n932));
  NAND2_X1  g731(.A1(new_n925), .A2(new_n932), .ZN(new_n933));
  OAI21_X1  g732(.A(G141gat), .B1(new_n933), .B2(new_n772), .ZN(new_n934));
  NOR2_X1   g733(.A1(new_n782), .A2(new_n376), .ZN(new_n935));
  NAND2_X1  g734(.A1(new_n891), .A2(new_n935), .ZN(new_n936));
  NOR2_X1   g735(.A1(new_n936), .A2(new_n838), .ZN(new_n937));
  NOR2_X1   g736(.A1(new_n772), .A2(G141gat), .ZN(new_n938));
  NAND2_X1  g737(.A1(new_n937), .A2(new_n938), .ZN(new_n939));
  INV_X1    g738(.A(KEYINPUT58), .ZN(new_n940));
  NAND3_X1  g739(.A1(new_n934), .A2(new_n939), .A3(new_n940), .ZN(new_n941));
  AOI21_X1  g740(.A(new_n931), .B1(new_n924), .B2(KEYINPUT57), .ZN(new_n942));
  AOI21_X1  g741(.A(new_n315), .B1(new_n942), .B2(new_n594), .ZN(new_n943));
  INV_X1    g742(.A(new_n939), .ZN(new_n944));
  OAI21_X1  g743(.A(KEYINPUT58), .B1(new_n943), .B2(new_n944), .ZN(new_n945));
  NAND2_X1  g744(.A1(new_n941), .A2(new_n945), .ZN(G1344gat));
  INV_X1    g745(.A(KEYINPUT59), .ZN(new_n947));
  AOI211_X1 g746(.A(new_n947), .B(G148gat), .C1(new_n937), .C2(new_n749), .ZN(new_n948));
  NAND3_X1  g747(.A1(new_n925), .A2(new_n749), .A3(new_n932), .ZN(new_n949));
  NAND2_X1  g748(.A1(new_n949), .A2(new_n947), .ZN(new_n950));
  OAI21_X1  g749(.A(KEYINPUT57), .B1(new_n890), .B2(new_n376), .ZN(new_n951));
  OAI211_X1 g750(.A(new_n926), .B(new_n795), .C1(new_n928), .C2(new_n868), .ZN(new_n952));
  AND2_X1   g751(.A1(new_n951), .A2(new_n952), .ZN(new_n953));
  NAND4_X1  g752(.A1(new_n953), .A2(KEYINPUT59), .A3(new_n749), .A4(new_n930), .ZN(new_n954));
  NAND2_X1  g753(.A1(new_n950), .A2(new_n954), .ZN(new_n955));
  AOI21_X1  g754(.A(new_n948), .B1(new_n955), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g755(.A(G155gat), .B1(new_n933), .B2(new_n704), .ZN(new_n957));
  NAND3_X1  g756(.A1(new_n937), .A2(new_n322), .A3(new_n705), .ZN(new_n958));
  NAND2_X1  g757(.A1(new_n957), .A2(new_n958), .ZN(G1346gat));
  OAI21_X1  g758(.A(G162gat), .B1(new_n933), .B2(new_n637), .ZN(new_n960));
  NOR3_X1   g759(.A1(new_n936), .A2(G162gat), .A3(new_n909), .ZN(new_n961));
  INV_X1    g760(.A(new_n961), .ZN(new_n962));
  INV_X1    g761(.A(KEYINPUT121), .ZN(new_n963));
  NAND3_X1  g762(.A1(new_n960), .A2(new_n962), .A3(new_n963), .ZN(new_n964));
  AOI21_X1  g763(.A(new_n323), .B1(new_n942), .B2(new_n636), .ZN(new_n965));
  OAI21_X1  g764(.A(KEYINPUT121), .B1(new_n965), .B2(new_n961), .ZN(new_n966));
  NAND2_X1  g765(.A1(new_n964), .A2(new_n966), .ZN(G1347gat));
  NOR2_X1   g766(.A1(new_n306), .A2(new_n755), .ZN(new_n968));
  NAND2_X1  g767(.A1(new_n898), .A2(new_n968), .ZN(new_n969));
  NOR3_X1   g768(.A1(new_n969), .A2(new_n211), .A3(new_n772), .ZN(new_n970));
  OAI21_X1  g769(.A(KEYINPUT122), .B1(new_n890), .B2(new_n755), .ZN(new_n971));
  INV_X1    g770(.A(KEYINPUT122), .ZN(new_n972));
  OAI211_X1 g771(.A(new_n972), .B(new_n435), .C1(new_n928), .C2(new_n868), .ZN(new_n973));
  AND4_X1   g772(.A1(new_n892), .A2(new_n971), .A3(new_n973), .A4(new_n838), .ZN(new_n974));
  NAND2_X1  g773(.A1(new_n974), .A2(new_n594), .ZN(new_n975));
  AOI21_X1  g774(.A(new_n970), .B1(new_n975), .B2(new_n211), .ZN(G1348gat));
  OAI21_X1  g775(.A(G176gat), .B1(new_n969), .B2(new_n726), .ZN(new_n977));
  NAND4_X1  g776(.A1(new_n971), .A2(new_n973), .A3(new_n892), .A4(new_n838), .ZN(new_n978));
  NAND2_X1  g777(.A1(new_n749), .A2(new_n212), .ZN(new_n979));
  OAI21_X1  g778(.A(new_n977), .B1(new_n978), .B2(new_n979), .ZN(G1349gat));
  INV_X1    g779(.A(KEYINPUT124), .ZN(new_n981));
  OAI21_X1  g780(.A(new_n981), .B1(new_n969), .B2(new_n704), .ZN(new_n982));
  NAND4_X1  g781(.A1(new_n898), .A2(KEYINPUT124), .A3(new_n705), .A4(new_n968), .ZN(new_n983));
  NAND3_X1  g782(.A1(new_n982), .A2(G183gat), .A3(new_n983), .ZN(new_n984));
  INV_X1    g783(.A(KEYINPUT123), .ZN(new_n985));
  NOR2_X1   g784(.A1(new_n226), .A2(new_n227), .ZN(new_n986));
  NAND2_X1  g785(.A1(new_n705), .A2(new_n986), .ZN(new_n987));
  INV_X1    g786(.A(new_n987), .ZN(new_n988));
  AOI21_X1  g787(.A(new_n985), .B1(new_n974), .B2(new_n988), .ZN(new_n989));
  NOR3_X1   g788(.A1(new_n978), .A2(KEYINPUT123), .A3(new_n987), .ZN(new_n990));
  OAI21_X1  g789(.A(new_n984), .B1(new_n989), .B2(new_n990), .ZN(new_n991));
  NAND2_X1  g790(.A1(new_n991), .A2(KEYINPUT60), .ZN(new_n992));
  INV_X1    g791(.A(KEYINPUT60), .ZN(new_n993));
  OAI211_X1 g792(.A(new_n984), .B(new_n993), .C1(new_n989), .C2(new_n990), .ZN(new_n994));
  NAND2_X1  g793(.A1(new_n992), .A2(new_n994), .ZN(G1350gat));
  NAND3_X1  g794(.A1(new_n974), .A2(new_n256), .A3(new_n636), .ZN(new_n996));
  OAI21_X1  g795(.A(G190gat), .B1(new_n969), .B2(new_n637), .ZN(new_n997));
  NAND2_X1  g796(.A1(new_n997), .A2(KEYINPUT125), .ZN(new_n998));
  INV_X1    g797(.A(KEYINPUT61), .ZN(new_n999));
  INV_X1    g798(.A(KEYINPUT125), .ZN(new_n1000));
  OAI211_X1 g799(.A(new_n1000), .B(G190gat), .C1(new_n969), .C2(new_n637), .ZN(new_n1001));
  AND3_X1   g800(.A1(new_n998), .A2(new_n999), .A3(new_n1001), .ZN(new_n1002));
  AOI21_X1  g801(.A(new_n999), .B1(new_n998), .B2(new_n1001), .ZN(new_n1003));
  OAI21_X1  g802(.A(new_n996), .B1(new_n1002), .B2(new_n1003), .ZN(G1351gat));
  AND2_X1   g803(.A1(new_n738), .A2(new_n968), .ZN(new_n1005));
  AND4_X1   g804(.A1(G197gat), .A2(new_n953), .A3(new_n594), .A4(new_n1005), .ZN(new_n1006));
  AND2_X1   g805(.A1(new_n971), .A2(new_n838), .ZN(new_n1007));
  AND2_X1   g806(.A1(new_n1007), .A2(new_n973), .ZN(new_n1008));
  NAND3_X1  g807(.A1(new_n1008), .A2(new_n594), .A3(new_n935), .ZN(new_n1009));
  INV_X1    g808(.A(G197gat), .ZN(new_n1010));
  AOI21_X1  g809(.A(new_n1006), .B1(new_n1009), .B2(new_n1010), .ZN(G1352gat));
  NAND3_X1  g810(.A1(new_n1007), .A2(new_n935), .A3(new_n973), .ZN(new_n1012));
  NOR2_X1   g811(.A1(new_n726), .A2(G204gat), .ZN(new_n1013));
  INV_X1    g812(.A(new_n1013), .ZN(new_n1014));
  OR3_X1    g813(.A1(new_n1012), .A2(KEYINPUT62), .A3(new_n1014), .ZN(new_n1015));
  NAND3_X1  g814(.A1(new_n953), .A2(new_n749), .A3(new_n1005), .ZN(new_n1016));
  NAND2_X1  g815(.A1(new_n1016), .A2(G204gat), .ZN(new_n1017));
  OAI21_X1  g816(.A(KEYINPUT62), .B1(new_n1012), .B2(new_n1014), .ZN(new_n1018));
  NAND3_X1  g817(.A1(new_n1015), .A2(new_n1017), .A3(new_n1018), .ZN(G1353gat));
  NAND3_X1  g818(.A1(new_n953), .A2(new_n705), .A3(new_n1005), .ZN(new_n1020));
  AND4_X1   g819(.A1(KEYINPUT126), .A2(new_n1020), .A3(KEYINPUT63), .A4(G211gat), .ZN(new_n1021));
  OAI21_X1  g820(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1022));
  INV_X1    g821(.A(new_n1022), .ZN(new_n1023));
  AOI22_X1  g822(.A1(new_n1020), .A2(new_n1023), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n1024));
  OR2_X1    g823(.A1(new_n704), .A2(G211gat), .ZN(new_n1025));
  OAI22_X1  g824(.A1(new_n1021), .A2(new_n1024), .B1(new_n1012), .B2(new_n1025), .ZN(G1354gat));
  NAND2_X1  g825(.A1(new_n636), .A2(G218gat), .ZN(new_n1027));
  XNOR2_X1  g826(.A(new_n1027), .B(KEYINPUT127), .ZN(new_n1028));
  AND3_X1   g827(.A1(new_n953), .A2(new_n1005), .A3(new_n1028), .ZN(new_n1029));
  NAND3_X1  g828(.A1(new_n1008), .A2(new_n636), .A3(new_n935), .ZN(new_n1030));
  INV_X1    g829(.A(G218gat), .ZN(new_n1031));
  AOI21_X1  g830(.A(new_n1029), .B1(new_n1030), .B2(new_n1031), .ZN(G1355gat));
endmodule


