//Secret key is'0 0 1 0 1 0 0 1 1 1 0 1 0 1 1 0 1 1 0 1 1 0 1 1 0 0 0 0 1 1 0 1 1 0 1 1 0 0 1 1 0 1 1 1 1 0 0 1 0 1 1 1 0 1 0 0 0 0 1 0 1 0 0 0 1 0 1 0 0 0 0 0 1 1 1 0 0 0 0 0 0 0 0 1 1 1 1 1 0 1 1 1 0 1 0 0 0 1 0 1 0 0 0 1 1 0 1 1 0 1 0 1 0 0 0 0 0 0 0 0 1 1 1 0 0 1 0' ..
// Benchmark "locked_locked_c2670" written by ABC on Sat Dec 16 05:32:23 2023

module locked_locked_c2670 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8, G11, G14, G15, G16, G19,
    G20, G21, G22, G23, G24, G25, G26, G27, G28, G29, G32, G33, G34, G35,
    G36, G37, G40, G43, G44, G47, G48, G49, G50, G51, G52, G53, G54, G55,
    G56, G57, G60, G61, G62, G63, G64, G65, G66, G67, G68, G69, G72, G73,
    G74, G75, G76, G77, G78, G79, G80, G81, G82, G85, G86, G87, G88, G89,
    G90, G91, G92, G93, G94, G95, G96, G99, G100, G101, G102, G103, G104,
    G105, G106, G107, G108, G111, G112, G113, G114, G115, G116, G117, G118,
    G119, G120, G123, G124, G125, G126, G127, G128, G129, G130, G131, G132,
    G135, G136, G137, G138, G139, G140, G141, G142, G169, G174, G177, G178,
    G179, G180, G181, G182, G183, G184, G185, G186, G189, G190, G191, G192,
    G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204,
    G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G239,
    G240, G241, G242, G243, G244, G245, G246, G247, G248, G249, G250, G251,
    G252, G253, G254, G255, G256, G257, G262, G263, G264, G265, G266, G267,
    G268, G269, G270, G271, G272, G273, G274, G275, G276, G277, G278, G279,
    G452, G483, G543, G559, G567, G651, G661, G860, G868, G1083, G1341,
    G1348, G1384, G1956, G1961, G1966, G1971, G1976, G1981, G1986, G1991,
    G1996, G2066, G2067, G2072, G2078, G2084, G2090, G2096, G2100, G2104,
    G2105, G2106, G2427, G2430, G2435, G2438, G2443, G2446, G2451, G2454,
    G2474, G2678,
    G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220, G221,
    G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217, G325,
    G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188, G299,
    G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148, G282,
    G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331, G397,
    G329, G231, G308, G225  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1, G2, G3, G4, G5, G6, G7, G8,
    G11, G14, G15, G16, G19, G20, G21, G22, G23, G24, G25, G26, G27, G28,
    G29, G32, G33, G34, G35, G36, G37, G40, G43, G44, G47, G48, G49, G50,
    G51, G52, G53, G54, G55, G56, G57, G60, G61, G62, G63, G64, G65, G66,
    G67, G68, G69, G72, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82,
    G85, G86, G87, G88, G89, G90, G91, G92, G93, G94, G95, G96, G99, G100,
    G101, G102, G103, G104, G105, G106, G107, G108, G111, G112, G113, G114,
    G115, G116, G117, G118, G119, G120, G123, G124, G125, G126, G127, G128,
    G129, G130, G131, G132, G135, G136, G137, G138, G139, G140, G141, G142,
    G169, G174, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186,
    G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200,
    G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212,
    G213, G214, G215, G239, G240, G241, G242, G243, G244, G245, G246, G247,
    G248, G249, G250, G251, G252, G253, G254, G255, G256, G257, G262, G263,
    G264, G265, G266, G267, G268, G269, G270, G271, G272, G273, G274, G275,
    G276, G277, G278, G279, G452, G483, G543, G559, G567, G651, G661, G860,
    G868, G1083, G1341, G1348, G1384, G1956, G1961, G1966, G1971, G1976,
    G1981, G1986, G1991, G1996, G2066, G2067, G2072, G2078, G2084, G2090,
    G2096, G2100, G2104, G2105, G2106, G2427, G2430, G2435, G2438, G2443,
    G2446, G2451, G2454, G2474, G2678;
  output G350, G335, G409, G369, G367, G411, G337, G384, G218, G219, G220,
    G221, G235, G236, G237, G238, G158, G259, G391, G173, G223, G234, G217,
    G325, G261, G319, G160, G162, G164, G166, G168, G171, G153, G176, G188,
    G299, G301, G286, G303, G288, G305, G290, G284, G321, G297, G280, G148,
    G282, G323, G156, G401, G227, G229, G311, G150, G145, G395, G295, G331,
    G397, G329, G231, G308, G225;
  wire new_n446, new_n450, new_n451, new_n452, new_n455, new_n456, new_n457,
    new_n458, new_n460, new_n461, new_n462, new_n463, new_n464, new_n465,
    new_n466, new_n467, new_n468, new_n469, new_n470, new_n471, new_n473,
    new_n474, new_n475, new_n476, new_n477, new_n478, new_n479, new_n480,
    new_n481, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n496,
    new_n497, new_n498, new_n499, new_n500, new_n501, new_n502, new_n503,
    new_n504, new_n505, new_n506, new_n507, new_n508, new_n509, new_n510,
    new_n511, new_n512, new_n513, new_n514, new_n516, new_n517, new_n518,
    new_n519, new_n520, new_n521, new_n522, new_n523, new_n524, new_n525,
    new_n526, new_n527, new_n529, new_n530, new_n531, new_n532, new_n533,
    new_n534, new_n535, new_n536, new_n537, new_n538, new_n541, new_n542,
    new_n543, new_n544, new_n545, new_n546, new_n547, new_n548, new_n549,
    new_n550, new_n551, new_n552, new_n553, new_n554, new_n555, new_n557,
    new_n559, new_n560, new_n562, new_n563, new_n564, new_n565, new_n566,
    new_n567, new_n571, new_n572, new_n573, new_n575, new_n576, new_n577,
    new_n578, new_n579, new_n580, new_n581, new_n582, new_n583, new_n584,
    new_n585, new_n587, new_n588, new_n589, new_n590, new_n591, new_n592,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n616,
    new_n617, new_n620, new_n622, new_n625, new_n626, new_n627, new_n628,
    new_n629, new_n630, new_n631, new_n632, new_n633, new_n634, new_n635,
    new_n637, new_n638, new_n639, new_n640, new_n641, new_n642, new_n643,
    new_n644, new_n645, new_n646, new_n647, new_n648, new_n649, new_n650,
    new_n651, new_n652, new_n654, new_n655, new_n656, new_n657, new_n658,
    new_n659, new_n660, new_n661, new_n662, new_n663, new_n664, new_n665,
    new_n666, new_n668, new_n669, new_n670, new_n671, new_n672, new_n673,
    new_n674, new_n675, new_n676, new_n677, new_n678, new_n679, new_n680,
    new_n681, new_n682, new_n683, new_n684, new_n685, new_n686, new_n688,
    new_n689, new_n690, new_n691, new_n692, new_n693, new_n694, new_n695,
    new_n696, new_n697, new_n698, new_n699, new_n700, new_n701, new_n702,
    new_n703, new_n704, new_n705, new_n706, new_n707, new_n708, new_n709,
    new_n710, new_n711, new_n712, new_n713, new_n714, new_n715, new_n716,
    new_n717, new_n718, new_n719, new_n720, new_n721, new_n722, new_n723,
    new_n724, new_n725, new_n726, new_n727, new_n728, new_n729, new_n730,
    new_n731, new_n732, new_n733, new_n734, new_n735, new_n736, new_n737,
    new_n738, new_n739, new_n740, new_n741, new_n742, new_n743, new_n744,
    new_n745, new_n746, new_n747, new_n748, new_n749, new_n750, new_n751,
    new_n752, new_n753, new_n754, new_n755, new_n756, new_n757, new_n758,
    new_n759, new_n760, new_n761, new_n762, new_n763, new_n764, new_n765,
    new_n766, new_n767, new_n768, new_n769, new_n770, new_n771, new_n772,
    new_n773, new_n774, new_n775, new_n776, new_n777, new_n778, new_n779,
    new_n780, new_n781, new_n782, new_n783, new_n784, new_n785, new_n786,
    new_n787, new_n788, new_n789, new_n790, new_n791, new_n792, new_n793,
    new_n794, new_n795, new_n796, new_n797, new_n798, new_n799, new_n800,
    new_n801, new_n802, new_n803, new_n804, new_n805, new_n806, new_n807,
    new_n808, new_n809, new_n810, new_n811, new_n812, new_n813, new_n814,
    new_n815, new_n816, new_n817, new_n818, new_n819, new_n820, new_n821,
    new_n824, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n846, new_n847, new_n848, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n871, new_n872, new_n873,
    new_n874, new_n875, new_n876, new_n877, new_n878, new_n879, new_n880,
    new_n881, new_n883, new_n884, new_n885, new_n886, new_n887, new_n888,
    new_n889, new_n890, new_n891, new_n892, new_n893, new_n894, new_n895,
    new_n896, new_n897, new_n898, new_n899, new_n900, new_n901, new_n902,
    new_n903, new_n904, new_n905, new_n906, new_n907, new_n908, new_n911,
    new_n912, new_n913, new_n914, new_n915, new_n916, new_n917, new_n918,
    new_n919, new_n920, new_n921, new_n922, new_n923, new_n924, new_n925,
    new_n926, new_n927, new_n928, new_n929, new_n930, new_n931, new_n932,
    new_n933, new_n934, new_n935, new_n936, new_n937, new_n938, new_n939,
    new_n940, new_n941, new_n942, new_n943, new_n944, new_n945, new_n946,
    new_n947, new_n948, new_n949, new_n950, new_n951, new_n952, new_n953,
    new_n954, new_n956, new_n957, new_n958, new_n959, new_n960, new_n961,
    new_n962, new_n963, new_n964, new_n965, new_n966, new_n967, new_n968,
    new_n969, new_n970, new_n971, new_n972, new_n973, new_n974, new_n975,
    new_n976, new_n977, new_n978, new_n979, new_n980, new_n981, new_n982,
    new_n983, new_n984, new_n985, new_n986, new_n987, new_n988, new_n989,
    new_n990, new_n991, new_n992, new_n993, new_n994, new_n995, new_n996,
    new_n997, new_n998, new_n999, new_n1000, new_n1001, new_n1002,
    new_n1003, new_n1004, new_n1005, new_n1006, new_n1007, new_n1008,
    new_n1009, new_n1010, new_n1011, new_n1012, new_n1013, new_n1014,
    new_n1015, new_n1016, new_n1017, new_n1018, new_n1019, new_n1020,
    new_n1021, new_n1022, new_n1023, new_n1024, new_n1025, new_n1026,
    new_n1027, new_n1028, new_n1029, new_n1030, new_n1031, new_n1032,
    new_n1033, new_n1034, new_n1035, new_n1036, new_n1037, new_n1038,
    new_n1039, new_n1040, new_n1041, new_n1042, new_n1043, new_n1044,
    new_n1045, new_n1046, new_n1047, new_n1048, new_n1049, new_n1050,
    new_n1051, new_n1052, new_n1053, new_n1054, new_n1055, new_n1056,
    new_n1057, new_n1058, new_n1059, new_n1060, new_n1061, new_n1062,
    new_n1063, new_n1064, new_n1065, new_n1066, new_n1067, new_n1068,
    new_n1069, new_n1070, new_n1071, new_n1072, new_n1073, new_n1074,
    new_n1075, new_n1076, new_n1077, new_n1078, new_n1079, new_n1080,
    new_n1081, new_n1082, new_n1083, new_n1084, new_n1085, new_n1086,
    new_n1087, new_n1088, new_n1089, new_n1090, new_n1091, new_n1092,
    new_n1093, new_n1094, new_n1095, new_n1096, new_n1097, new_n1098,
    new_n1099, new_n1100, new_n1101, new_n1102, new_n1103, new_n1104,
    new_n1105, new_n1106, new_n1107, new_n1108, new_n1109, new_n1110,
    new_n1111, new_n1112, new_n1113, new_n1114, new_n1115, new_n1116,
    new_n1117, new_n1118, new_n1119, new_n1120, new_n1121, new_n1122,
    new_n1123, new_n1124, new_n1125, new_n1126, new_n1127, new_n1128,
    new_n1129, new_n1130, new_n1131, new_n1132, new_n1133, new_n1134,
    new_n1135, new_n1136, new_n1137, new_n1138, new_n1139, new_n1140,
    new_n1141, new_n1142, new_n1143, new_n1144, new_n1145, new_n1146,
    new_n1147, new_n1148, new_n1149, new_n1150, new_n1151, new_n1152,
    new_n1153, new_n1154, new_n1155, new_n1156, new_n1157, new_n1158,
    new_n1159, new_n1160, new_n1161, new_n1162, new_n1163, new_n1164,
    new_n1165, new_n1166, new_n1167, new_n1168, new_n1169, new_n1170,
    new_n1171, new_n1172, new_n1173, new_n1174, new_n1175, new_n1176,
    new_n1177, new_n1178, new_n1179, new_n1180, new_n1181, new_n1182,
    new_n1183, new_n1184, new_n1187, new_n1188, new_n1189, new_n1190,
    new_n1191, new_n1192, new_n1193, new_n1194, new_n1195;
  BUF_X1    g000(.A(G452), .Z(G350));
  BUF_X1    g001(.A(G452), .Z(G335));
  BUF_X1    g002(.A(G452), .Z(G409));
  BUF_X1    g003(.A(G1083), .Z(G369));
  BUF_X1    g004(.A(G1083), .Z(G367));
  BUF_X1    g005(.A(G2066), .Z(G411));
  BUF_X1    g006(.A(G2066), .Z(G337));
  BUF_X1    g007(.A(G2066), .Z(G384));
  INV_X1    g008(.A(G44), .ZN(G218));
  INV_X1    g009(.A(G132), .ZN(G219));
  XNOR2_X1  g010(.A(KEYINPUT0), .B(G82), .ZN(G220));
  INV_X1    g011(.A(G96), .ZN(G221));
  INV_X1    g012(.A(G69), .ZN(G235));
  INV_X1    g013(.A(G120), .ZN(G236));
  INV_X1    g014(.A(G57), .ZN(G237));
  INV_X1    g015(.A(G108), .ZN(G238));
  NAND4_X1  g016(.A1(G2072), .A2(G2078), .A3(G2084), .A4(G2090), .ZN(G158));
  NAND3_X1  g017(.A1(G2), .A2(G15), .A3(G661), .ZN(G259));
  BUF_X1    g018(.A(G452), .Z(G391));
  AND2_X1   g019(.A1(G94), .A2(G452), .ZN(G173));
  NAND2_X1  g020(.A1(G7), .A2(G661), .ZN(new_n446));
  XOR2_X1   g021(.A(new_n446), .B(KEYINPUT1), .Z(G223));
  NAND3_X1  g022(.A1(G7), .A2(G567), .A3(G661), .ZN(G234));
  NAND3_X1  g023(.A1(G7), .A2(G661), .A3(G2106), .ZN(G217));
  NOR4_X1   g024(.A1(G220), .A2(G218), .A3(G221), .A4(G219), .ZN(new_n450));
  XOR2_X1   g025(.A(new_n450), .B(KEYINPUT2), .Z(new_n451));
  NAND4_X1  g026(.A1(G57), .A2(G69), .A3(G108), .A4(G120), .ZN(new_n452));
  NOR2_X1   g027(.A1(new_n451), .A2(new_n452), .ZN(G325));
  INV_X1    g028(.A(G325), .ZN(G261));
  NAND2_X1  g029(.A1(new_n451), .A2(G2106), .ZN(new_n455));
  NAND2_X1  g030(.A1(new_n452), .A2(G567), .ZN(new_n456));
  XNOR2_X1  g031(.A(new_n456), .B(KEYINPUT64), .ZN(new_n457));
  NAND2_X1  g032(.A1(new_n455), .A2(new_n457), .ZN(new_n458));
  INV_X1    g033(.A(new_n458), .ZN(G319));
  INV_X1    g034(.A(G2105), .ZN(new_n460));
  XNOR2_X1  g035(.A(KEYINPUT3), .B(G2104), .ZN(new_n461));
  NAND2_X1  g036(.A1(new_n461), .A2(G125), .ZN(new_n462));
  NAND2_X1  g037(.A1(G113), .A2(G2104), .ZN(new_n463));
  AOI21_X1  g038(.A(new_n460), .B1(new_n462), .B2(new_n463), .ZN(new_n464));
  INV_X1    g039(.A(G2104), .ZN(new_n465));
  NAND2_X1  g040(.A1(new_n465), .A2(KEYINPUT3), .ZN(new_n466));
  INV_X1    g041(.A(KEYINPUT3), .ZN(new_n467));
  NAND2_X1  g042(.A1(new_n467), .A2(G2104), .ZN(new_n468));
  NAND4_X1  g043(.A1(new_n466), .A2(new_n468), .A3(G137), .A4(new_n460), .ZN(new_n469));
  NAND3_X1  g044(.A1(new_n460), .A2(G101), .A3(G2104), .ZN(new_n470));
  NAND2_X1  g045(.A1(new_n469), .A2(new_n470), .ZN(new_n471));
  NOR2_X1   g046(.A1(new_n464), .A2(new_n471), .ZN(G160));
  NAND2_X1  g047(.A1(new_n461), .A2(G2105), .ZN(new_n473));
  INV_X1    g048(.A(new_n473), .ZN(new_n474));
  NAND2_X1  g049(.A1(new_n474), .A2(G124), .ZN(new_n475));
  NAND2_X1  g050(.A1(new_n461), .A2(new_n460), .ZN(new_n476));
  INV_X1    g051(.A(new_n476), .ZN(new_n477));
  NAND2_X1  g052(.A1(new_n477), .A2(G136), .ZN(new_n478));
  OR2_X1    g053(.A1(G100), .A2(G2105), .ZN(new_n479));
  OAI211_X1 g054(.A(new_n479), .B(G2104), .C1(G112), .C2(new_n460), .ZN(new_n480));
  NAND3_X1  g055(.A1(new_n475), .A2(new_n478), .A3(new_n480), .ZN(new_n481));
  INV_X1    g056(.A(new_n481), .ZN(G162));
  NAND4_X1  g057(.A1(new_n466), .A2(new_n468), .A3(G126), .A4(G2105), .ZN(new_n483));
  INV_X1    g058(.A(G114), .ZN(new_n484));
  NAND2_X1  g059(.A1(new_n484), .A2(G2105), .ZN(new_n485));
  OAI211_X1 g060(.A(new_n485), .B(G2104), .C1(G102), .C2(G2105), .ZN(new_n486));
  NAND2_X1  g061(.A1(new_n483), .A2(new_n486), .ZN(new_n487));
  NAND2_X1  g062(.A1(new_n487), .A2(KEYINPUT65), .ZN(new_n488));
  INV_X1    g063(.A(KEYINPUT65), .ZN(new_n489));
  NAND3_X1  g064(.A1(new_n483), .A2(new_n486), .A3(new_n489), .ZN(new_n490));
  NAND4_X1  g065(.A1(new_n466), .A2(new_n468), .A3(G138), .A4(new_n460), .ZN(new_n491));
  NAND2_X1  g066(.A1(new_n491), .A2(KEYINPUT4), .ZN(new_n492));
  INV_X1    g067(.A(KEYINPUT4), .ZN(new_n493));
  NAND4_X1  g068(.A1(new_n461), .A2(new_n493), .A3(G138), .A4(new_n460), .ZN(new_n494));
  AOI22_X1  g069(.A1(new_n488), .A2(new_n490), .B1(new_n492), .B2(new_n494), .ZN(G164));
  INV_X1    g070(.A(G651), .ZN(new_n496));
  NAND2_X1  g071(.A1(new_n496), .A2(KEYINPUT6), .ZN(new_n497));
  INV_X1    g072(.A(KEYINPUT6), .ZN(new_n498));
  NAND2_X1  g073(.A1(new_n498), .A2(G651), .ZN(new_n499));
  AND2_X1   g074(.A1(new_n497), .A2(new_n499), .ZN(new_n500));
  NAND3_X1  g075(.A1(new_n500), .A2(G50), .A3(G543), .ZN(new_n501));
  INV_X1    g076(.A(KEYINPUT66), .ZN(new_n502));
  XNOR2_X1  g077(.A(new_n501), .B(new_n502), .ZN(new_n503));
  NAND2_X1  g078(.A1(new_n497), .A2(new_n499), .ZN(new_n504));
  INV_X1    g079(.A(G543), .ZN(new_n505));
  NAND2_X1  g080(.A1(new_n505), .A2(KEYINPUT5), .ZN(new_n506));
  INV_X1    g081(.A(KEYINPUT5), .ZN(new_n507));
  NAND2_X1  g082(.A1(new_n507), .A2(G543), .ZN(new_n508));
  NAND2_X1  g083(.A1(new_n506), .A2(new_n508), .ZN(new_n509));
  NOR2_X1   g084(.A1(new_n504), .A2(new_n509), .ZN(new_n510));
  NAND2_X1  g085(.A1(new_n510), .A2(G88), .ZN(new_n511));
  INV_X1    g086(.A(new_n509), .ZN(new_n512));
  AOI22_X1  g087(.A1(new_n512), .A2(G62), .B1(G75), .B2(G543), .ZN(new_n513));
  OAI21_X1  g088(.A(new_n511), .B1(new_n513), .B2(new_n496), .ZN(new_n514));
  NOR2_X1   g089(.A1(new_n503), .A2(new_n514), .ZN(G166));
  NAND2_X1  g090(.A1(G63), .A2(G651), .ZN(new_n516));
  INV_X1    g091(.A(G89), .ZN(new_n517));
  OAI21_X1  g092(.A(new_n516), .B1(new_n504), .B2(new_n517), .ZN(new_n518));
  NAND2_X1  g093(.A1(new_n518), .A2(new_n512), .ZN(new_n519));
  NAND3_X1  g094(.A1(G76), .A2(G543), .A3(G651), .ZN(new_n520));
  XNOR2_X1  g095(.A(new_n520), .B(KEYINPUT7), .ZN(new_n521));
  NAND2_X1  g096(.A1(new_n519), .A2(new_n521), .ZN(new_n522));
  INV_X1    g097(.A(KEYINPUT67), .ZN(new_n523));
  OAI21_X1  g098(.A(new_n523), .B1(new_n504), .B2(new_n505), .ZN(new_n524));
  INV_X1    g099(.A(new_n524), .ZN(new_n525));
  NOR3_X1   g100(.A1(new_n504), .A2(new_n523), .A3(new_n505), .ZN(new_n526));
  NOR2_X1   g101(.A1(new_n525), .A2(new_n526), .ZN(new_n527));
  AOI21_X1  g102(.A(new_n522), .B1(new_n527), .B2(G51), .ZN(G168));
  NAND2_X1  g103(.A1(G77), .A2(G543), .ZN(new_n529));
  INV_X1    g104(.A(G64), .ZN(new_n530));
  OAI21_X1  g105(.A(new_n529), .B1(new_n509), .B2(new_n530), .ZN(new_n531));
  AOI22_X1  g106(.A1(G651), .A2(new_n531), .B1(new_n510), .B2(G90), .ZN(new_n532));
  INV_X1    g107(.A(KEYINPUT68), .ZN(new_n533));
  NAND3_X1  g108(.A1(new_n500), .A2(KEYINPUT67), .A3(G543), .ZN(new_n534));
  NAND3_X1  g109(.A1(new_n534), .A2(G52), .A3(new_n524), .ZN(new_n535));
  NAND3_X1  g110(.A1(new_n532), .A2(new_n533), .A3(new_n535), .ZN(new_n536));
  INV_X1    g111(.A(new_n536), .ZN(new_n537));
  AOI21_X1  g112(.A(new_n533), .B1(new_n532), .B2(new_n535), .ZN(new_n538));
  NOR2_X1   g113(.A1(new_n537), .A2(new_n538), .ZN(G301));
  INV_X1    g114(.A(G301), .ZN(G171));
  NAND2_X1  g115(.A1(G68), .A2(G543), .ZN(new_n541));
  INV_X1    g116(.A(G56), .ZN(new_n542));
  OAI21_X1  g117(.A(new_n541), .B1(new_n509), .B2(new_n542), .ZN(new_n543));
  AND2_X1   g118(.A1(new_n543), .A2(KEYINPUT69), .ZN(new_n544));
  OAI21_X1  g119(.A(G651), .B1(new_n543), .B2(KEYINPUT69), .ZN(new_n545));
  NOR2_X1   g120(.A1(new_n544), .A2(new_n545), .ZN(new_n546));
  INV_X1    g121(.A(new_n546), .ZN(new_n547));
  NAND3_X1  g122(.A1(new_n534), .A2(G43), .A3(new_n524), .ZN(new_n548));
  INV_X1    g123(.A(KEYINPUT70), .ZN(new_n549));
  NAND2_X1  g124(.A1(new_n510), .A2(G81), .ZN(new_n550));
  NAND3_X1  g125(.A1(new_n548), .A2(new_n549), .A3(new_n550), .ZN(new_n551));
  INV_X1    g126(.A(new_n551), .ZN(new_n552));
  AOI21_X1  g127(.A(new_n549), .B1(new_n548), .B2(new_n550), .ZN(new_n553));
  OAI21_X1  g128(.A(new_n547), .B1(new_n552), .B2(new_n553), .ZN(new_n554));
  INV_X1    g129(.A(new_n554), .ZN(new_n555));
  NAND2_X1  g130(.A1(new_n555), .A2(G860), .ZN(G153));
  AND3_X1   g131(.A1(G319), .A2(G483), .A3(G661), .ZN(new_n557));
  NAND2_X1  g132(.A1(new_n557), .A2(G36), .ZN(G176));
  NAND2_X1  g133(.A1(G1), .A2(G3), .ZN(new_n559));
  XNOR2_X1  g134(.A(new_n559), .B(KEYINPUT8), .ZN(new_n560));
  NAND2_X1  g135(.A1(new_n557), .A2(new_n560), .ZN(G188));
  NAND3_X1  g136(.A1(new_n500), .A2(G53), .A3(G543), .ZN(new_n562));
  XNOR2_X1  g137(.A(new_n562), .B(KEYINPUT9), .ZN(new_n563));
  NAND2_X1  g138(.A1(G78), .A2(G543), .ZN(new_n564));
  INV_X1    g139(.A(G65), .ZN(new_n565));
  OAI21_X1  g140(.A(new_n564), .B1(new_n509), .B2(new_n565), .ZN(new_n566));
  AOI22_X1  g141(.A1(G651), .A2(new_n566), .B1(new_n510), .B2(G91), .ZN(new_n567));
  NAND2_X1  g142(.A1(new_n563), .A2(new_n567), .ZN(G299));
  INV_X1    g143(.A(G168), .ZN(G286));
  INV_X1    g144(.A(G166), .ZN(G303));
  NAND2_X1  g145(.A1(new_n510), .A2(G87), .ZN(new_n571));
  OAI21_X1  g146(.A(G651), .B1(new_n512), .B2(G74), .ZN(new_n572));
  NAND3_X1  g147(.A1(new_n500), .A2(G49), .A3(G543), .ZN(new_n573));
  NAND3_X1  g148(.A1(new_n571), .A2(new_n572), .A3(new_n573), .ZN(G288));
  NAND3_X1  g149(.A1(new_n500), .A2(G48), .A3(G543), .ZN(new_n575));
  NAND2_X1  g150(.A1(new_n575), .A2(KEYINPUT72), .ZN(new_n576));
  INV_X1    g151(.A(KEYINPUT72), .ZN(new_n577));
  NAND4_X1  g152(.A1(new_n500), .A2(new_n577), .A3(G48), .A4(G543), .ZN(new_n578));
  AOI22_X1  g153(.A1(new_n576), .A2(new_n578), .B1(G86), .B2(new_n510), .ZN(new_n579));
  INV_X1    g154(.A(G61), .ZN(new_n580));
  OAI21_X1  g155(.A(KEYINPUT71), .B1(new_n509), .B2(new_n580), .ZN(new_n581));
  NAND2_X1  g156(.A1(G73), .A2(G543), .ZN(new_n582));
  NAND2_X1  g157(.A1(new_n581), .A2(new_n582), .ZN(new_n583));
  NOR3_X1   g158(.A1(new_n509), .A2(KEYINPUT71), .A3(new_n580), .ZN(new_n584));
  OAI21_X1  g159(.A(G651), .B1(new_n583), .B2(new_n584), .ZN(new_n585));
  NAND2_X1  g160(.A1(new_n579), .A2(new_n585), .ZN(G305));
  AOI22_X1  g161(.A1(new_n527), .A2(G47), .B1(G85), .B2(new_n510), .ZN(new_n587));
  NAND2_X1  g162(.A1(G72), .A2(G543), .ZN(new_n588));
  INV_X1    g163(.A(G60), .ZN(new_n589));
  OAI21_X1  g164(.A(new_n588), .B1(new_n509), .B2(new_n589), .ZN(new_n590));
  NAND2_X1  g165(.A1(new_n590), .A2(G651), .ZN(new_n591));
  XNOR2_X1  g166(.A(new_n591), .B(KEYINPUT73), .ZN(new_n592));
  NAND2_X1  g167(.A1(new_n587), .A2(new_n592), .ZN(G290));
  NAND2_X1  g168(.A1(G301), .A2(G868), .ZN(new_n594));
  INV_X1    g169(.A(G92), .ZN(new_n595));
  XNOR2_X1  g170(.A(KEYINPUT74), .B(KEYINPUT10), .ZN(new_n596));
  OR4_X1    g171(.A1(new_n595), .A2(new_n504), .A3(new_n509), .A4(new_n596), .ZN(new_n597));
  NAND2_X1  g172(.A1(new_n510), .A2(G92), .ZN(new_n598));
  NAND2_X1  g173(.A1(new_n598), .A2(new_n596), .ZN(new_n599));
  NAND2_X1  g174(.A1(G79), .A2(G543), .ZN(new_n600));
  INV_X1    g175(.A(G66), .ZN(new_n601));
  OAI21_X1  g176(.A(new_n600), .B1(new_n509), .B2(new_n601), .ZN(new_n602));
  NAND2_X1  g177(.A1(new_n602), .A2(G651), .ZN(new_n603));
  AND3_X1   g178(.A1(new_n597), .A2(new_n599), .A3(new_n603), .ZN(new_n604));
  INV_X1    g179(.A(KEYINPUT75), .ZN(new_n605));
  OAI21_X1  g180(.A(new_n605), .B1(new_n525), .B2(new_n526), .ZN(new_n606));
  NAND3_X1  g181(.A1(new_n534), .A2(KEYINPUT75), .A3(new_n524), .ZN(new_n607));
  NAND3_X1  g182(.A1(new_n606), .A2(G54), .A3(new_n607), .ZN(new_n608));
  NAND2_X1  g183(.A1(new_n604), .A2(new_n608), .ZN(new_n609));
  AND2_X1   g184(.A1(new_n609), .A2(KEYINPUT76), .ZN(new_n610));
  NOR2_X1   g185(.A1(new_n609), .A2(KEYINPUT76), .ZN(new_n611));
  NOR2_X1   g186(.A1(new_n610), .A2(new_n611), .ZN(new_n612));
  INV_X1    g187(.A(new_n612), .ZN(new_n613));
  OAI21_X1  g188(.A(new_n594), .B1(new_n613), .B2(G868), .ZN(G284));
  OAI21_X1  g189(.A(new_n594), .B1(new_n613), .B2(G868), .ZN(G321));
  NAND2_X1  g190(.A1(G286), .A2(G868), .ZN(new_n616));
  XNOR2_X1  g191(.A(G299), .B(KEYINPUT77), .ZN(new_n617));
  OAI21_X1  g192(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G297));
  OAI21_X1  g193(.A(new_n616), .B1(new_n617), .B2(G868), .ZN(G280));
  NOR2_X1   g194(.A1(new_n612), .A2(G559), .ZN(new_n620));
  AOI21_X1  g195(.A(new_n620), .B1(G860), .B2(new_n613), .ZN(G148));
  OAI21_X1  g196(.A(G868), .B1(new_n612), .B2(G559), .ZN(new_n622));
  OAI21_X1  g197(.A(new_n622), .B1(G868), .B2(new_n555), .ZN(G323));
  XNOR2_X1  g198(.A(G323), .B(KEYINPUT11), .ZN(G282));
  NAND2_X1  g199(.A1(new_n477), .A2(G135), .ZN(new_n625));
  NOR2_X1   g200(.A1(new_n460), .A2(G111), .ZN(new_n626));
  OAI21_X1  g201(.A(G2104), .B1(G99), .B2(G2105), .ZN(new_n627));
  OAI21_X1  g202(.A(new_n625), .B1(new_n626), .B2(new_n627), .ZN(new_n628));
  AOI21_X1  g203(.A(new_n628), .B1(G123), .B2(new_n474), .ZN(new_n629));
  XOR2_X1   g204(.A(new_n629), .B(KEYINPUT78), .Z(new_n630));
  XNOR2_X1  g205(.A(new_n630), .B(G2096), .ZN(new_n631));
  NAND3_X1  g206(.A1(new_n460), .A2(KEYINPUT3), .A3(G2104), .ZN(new_n632));
  XNOR2_X1  g207(.A(new_n632), .B(KEYINPUT12), .ZN(new_n633));
  XNOR2_X1  g208(.A(new_n633), .B(KEYINPUT13), .ZN(new_n634));
  XNOR2_X1  g209(.A(new_n634), .B(G2100), .ZN(new_n635));
  NAND2_X1  g210(.A1(new_n631), .A2(new_n635), .ZN(G156));
  XOR2_X1   g211(.A(KEYINPUT15), .B(G2435), .Z(new_n637));
  XNOR2_X1  g212(.A(new_n637), .B(G2438), .ZN(new_n638));
  XOR2_X1   g213(.A(G2427), .B(G2430), .Z(new_n639));
  OAI21_X1  g214(.A(KEYINPUT14), .B1(new_n638), .B2(new_n639), .ZN(new_n640));
  XNOR2_X1  g215(.A(new_n640), .B(KEYINPUT79), .ZN(new_n641));
  NAND2_X1  g216(.A1(new_n638), .A2(new_n639), .ZN(new_n642));
  NAND2_X1  g217(.A1(new_n641), .A2(new_n642), .ZN(new_n643));
  XNOR2_X1  g218(.A(G2451), .B(G2454), .ZN(new_n644));
  XNOR2_X1  g219(.A(new_n644), .B(KEYINPUT16), .ZN(new_n645));
  XNOR2_X1  g220(.A(new_n643), .B(new_n645), .ZN(new_n646));
  XOR2_X1   g221(.A(G2443), .B(G2446), .Z(new_n647));
  XNOR2_X1  g222(.A(new_n646), .B(new_n647), .ZN(new_n648));
  XNOR2_X1  g223(.A(G1341), .B(G1348), .ZN(new_n649));
  INV_X1    g224(.A(new_n649), .ZN(new_n650));
  AND2_X1   g225(.A1(new_n648), .A2(new_n650), .ZN(new_n651));
  OAI21_X1  g226(.A(G14), .B1(new_n648), .B2(new_n650), .ZN(new_n652));
  NOR2_X1   g227(.A1(new_n651), .A2(new_n652), .ZN(G401));
  XOR2_X1   g228(.A(G2084), .B(G2090), .Z(new_n654));
  INV_X1    g229(.A(new_n654), .ZN(new_n655));
  XOR2_X1   g230(.A(G2067), .B(G2678), .Z(new_n656));
  NOR2_X1   g231(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  XNOR2_X1  g232(.A(G2072), .B(G2078), .ZN(new_n658));
  NAND2_X1  g233(.A1(new_n657), .A2(new_n658), .ZN(new_n659));
  XNOR2_X1  g234(.A(new_n659), .B(KEYINPUT18), .ZN(new_n660));
  NAND2_X1  g235(.A1(new_n655), .A2(new_n656), .ZN(new_n661));
  AND3_X1   g236(.A1(new_n661), .A2(KEYINPUT17), .A3(new_n658), .ZN(new_n662));
  AOI21_X1  g237(.A(new_n658), .B1(new_n661), .B2(KEYINPUT17), .ZN(new_n663));
  NOR3_X1   g238(.A1(new_n662), .A2(new_n663), .A3(new_n657), .ZN(new_n664));
  NOR2_X1   g239(.A1(new_n660), .A2(new_n664), .ZN(new_n665));
  XNOR2_X1  g240(.A(G2096), .B(G2100), .ZN(new_n666));
  XNOR2_X1  g241(.A(new_n665), .B(new_n666), .ZN(G227));
  XNOR2_X1  g242(.A(G1971), .B(G1976), .ZN(new_n668));
  XNOR2_X1  g243(.A(new_n668), .B(KEYINPUT19), .ZN(new_n669));
  XOR2_X1   g244(.A(G1956), .B(G2474), .Z(new_n670));
  XOR2_X1   g245(.A(G1961), .B(G1966), .Z(new_n671));
  OR2_X1    g246(.A1(new_n670), .A2(new_n671), .ZN(new_n672));
  NAND2_X1  g247(.A1(new_n670), .A2(new_n671), .ZN(new_n673));
  NAND3_X1  g248(.A1(new_n669), .A2(new_n672), .A3(new_n673), .ZN(new_n674));
  NOR2_X1   g249(.A1(new_n669), .A2(new_n673), .ZN(new_n675));
  INV_X1    g250(.A(new_n675), .ZN(new_n676));
  XOR2_X1   g251(.A(KEYINPUT80), .B(KEYINPUT20), .Z(new_n677));
  INV_X1    g252(.A(new_n677), .ZN(new_n678));
  OAI221_X1 g253(.A(new_n674), .B1(new_n669), .B2(new_n672), .C1(new_n676), .C2(new_n678), .ZN(new_n679));
  AOI21_X1  g254(.A(new_n679), .B1(new_n676), .B2(new_n678), .ZN(new_n680));
  XNOR2_X1  g255(.A(G1981), .B(G1986), .ZN(new_n681));
  XNOR2_X1  g256(.A(new_n681), .B(KEYINPUT81), .ZN(new_n682));
  XNOR2_X1  g257(.A(new_n680), .B(new_n682), .ZN(new_n683));
  XNOR2_X1  g258(.A(G1991), .B(G1996), .ZN(new_n684));
  XNOR2_X1  g259(.A(KEYINPUT21), .B(KEYINPUT22), .ZN(new_n685));
  XNOR2_X1  g260(.A(new_n684), .B(new_n685), .ZN(new_n686));
  XNOR2_X1  g261(.A(new_n683), .B(new_n686), .ZN(G229));
  NOR2_X1   g262(.A1(G16), .A2(G24), .ZN(new_n688));
  XOR2_X1   g263(.A(G290), .B(KEYINPUT85), .Z(new_n689));
  AOI21_X1  g264(.A(new_n688), .B1(new_n689), .B2(G16), .ZN(new_n690));
  XNOR2_X1  g265(.A(new_n690), .B(G1986), .ZN(new_n691));
  MUX2_X1   g266(.A(G6), .B(G305), .S(G16), .Z(new_n692));
  XOR2_X1   g267(.A(KEYINPUT32), .B(G1981), .Z(new_n693));
  XNOR2_X1  g268(.A(new_n692), .B(new_n693), .ZN(new_n694));
  NOR2_X1   g269(.A1(G16), .A2(G23), .ZN(new_n695));
  INV_X1    g270(.A(G288), .ZN(new_n696));
  AOI21_X1  g271(.A(new_n695), .B1(new_n696), .B2(G16), .ZN(new_n697));
  XOR2_X1   g272(.A(KEYINPUT33), .B(G1976), .Z(new_n698));
  XNOR2_X1  g273(.A(new_n697), .B(new_n698), .ZN(new_n699));
  INV_X1    g274(.A(G16), .ZN(new_n700));
  NAND2_X1  g275(.A1(new_n700), .A2(G22), .ZN(new_n701));
  OAI21_X1  g276(.A(new_n701), .B1(G166), .B2(new_n700), .ZN(new_n702));
  AOI21_X1  g277(.A(new_n699), .B1(G1971), .B2(new_n702), .ZN(new_n703));
  OAI211_X1 g278(.A(new_n694), .B(new_n703), .C1(G1971), .C2(new_n702), .ZN(new_n704));
  AOI21_X1  g279(.A(new_n691), .B1(KEYINPUT34), .B2(new_n704), .ZN(new_n705));
  NOR2_X1   g280(.A1(new_n704), .A2(KEYINPUT34), .ZN(new_n706));
  XNOR2_X1  g281(.A(KEYINPUT35), .B(G1991), .ZN(new_n707));
  NOR2_X1   g282(.A1(G25), .A2(G29), .ZN(new_n708));
  INV_X1    g283(.A(G119), .ZN(new_n709));
  OR3_X1    g284(.A1(new_n473), .A2(KEYINPUT82), .A3(new_n709), .ZN(new_n710));
  OAI21_X1  g285(.A(KEYINPUT82), .B1(new_n473), .B2(new_n709), .ZN(new_n711));
  NAND2_X1  g286(.A1(new_n477), .A2(G131), .ZN(new_n712));
  OR2_X1    g287(.A1(G95), .A2(G2105), .ZN(new_n713));
  OAI211_X1 g288(.A(new_n713), .B(G2104), .C1(G107), .C2(new_n460), .ZN(new_n714));
  NAND4_X1  g289(.A1(new_n710), .A2(new_n711), .A3(new_n712), .A4(new_n714), .ZN(new_n715));
  XOR2_X1   g290(.A(new_n715), .B(KEYINPUT83), .Z(new_n716));
  AOI21_X1  g291(.A(new_n708), .B1(new_n716), .B2(G29), .ZN(new_n717));
  XNOR2_X1  g292(.A(new_n717), .B(KEYINPUT84), .ZN(new_n718));
  AOI21_X1  g293(.A(new_n706), .B1(new_n707), .B2(new_n718), .ZN(new_n719));
  OAI211_X1 g294(.A(new_n705), .B(new_n719), .C1(new_n707), .C2(new_n718), .ZN(new_n720));
  XNOR2_X1  g295(.A(new_n720), .B(KEYINPUT36), .ZN(new_n721));
  OR2_X1    g296(.A1(G4), .A2(G16), .ZN(new_n722));
  OAI211_X1 g297(.A(KEYINPUT86), .B(new_n722), .C1(new_n612), .C2(new_n700), .ZN(new_n723));
  OAI21_X1  g298(.A(new_n723), .B1(KEYINPUT86), .B2(new_n722), .ZN(new_n724));
  INV_X1    g299(.A(G1348), .ZN(new_n725));
  XNOR2_X1  g300(.A(new_n724), .B(new_n725), .ZN(new_n726));
  OR2_X1    g301(.A1(G29), .A2(G33), .ZN(new_n727));
  NAND2_X1  g302(.A1(new_n477), .A2(G139), .ZN(new_n728));
  XOR2_X1   g303(.A(new_n728), .B(KEYINPUT88), .Z(new_n729));
  NAND3_X1  g304(.A1(new_n460), .A2(G103), .A3(G2104), .ZN(new_n730));
  XOR2_X1   g305(.A(new_n730), .B(KEYINPUT25), .Z(new_n731));
  AOI22_X1  g306(.A1(new_n461), .A2(G127), .B1(G115), .B2(G2104), .ZN(new_n732));
  OAI211_X1 g307(.A(new_n729), .B(new_n731), .C1(new_n460), .C2(new_n732), .ZN(new_n733));
  INV_X1    g308(.A(G29), .ZN(new_n734));
  OAI21_X1  g309(.A(new_n727), .B1(new_n733), .B2(new_n734), .ZN(new_n735));
  INV_X1    g310(.A(G2072), .ZN(new_n736));
  NAND2_X1  g311(.A1(new_n735), .A2(new_n736), .ZN(new_n737));
  XOR2_X1   g312(.A(new_n737), .B(KEYINPUT89), .Z(new_n738));
  NAND2_X1  g313(.A1(new_n734), .A2(G35), .ZN(new_n739));
  OAI21_X1  g314(.A(new_n739), .B1(G162), .B2(new_n734), .ZN(new_n740));
  XOR2_X1   g315(.A(new_n740), .B(KEYINPUT29), .Z(new_n741));
  INV_X1    g316(.A(G2090), .ZN(new_n742));
  NAND2_X1  g317(.A1(new_n741), .A2(new_n742), .ZN(new_n743));
  XNOR2_X1  g318(.A(new_n743), .B(KEYINPUT95), .ZN(new_n744));
  NOR2_X1   g319(.A1(G29), .A2(G32), .ZN(new_n745));
  XNOR2_X1  g320(.A(KEYINPUT91), .B(KEYINPUT26), .ZN(new_n746));
  NAND3_X1  g321(.A1(G117), .A2(G2104), .A3(G2105), .ZN(new_n747));
  OR2_X1    g322(.A1(new_n746), .A2(new_n747), .ZN(new_n748));
  NAND2_X1  g323(.A1(new_n746), .A2(new_n747), .ZN(new_n749));
  NAND3_X1  g324(.A1(new_n460), .A2(G105), .A3(G2104), .ZN(new_n750));
  NAND3_X1  g325(.A1(new_n748), .A2(new_n749), .A3(new_n750), .ZN(new_n751));
  INV_X1    g326(.A(G129), .ZN(new_n752));
  INV_X1    g327(.A(G141), .ZN(new_n753));
  OAI22_X1  g328(.A1(new_n752), .A2(new_n473), .B1(new_n476), .B2(new_n753), .ZN(new_n754));
  NOR2_X1   g329(.A1(new_n751), .A2(new_n754), .ZN(new_n755));
  XOR2_X1   g330(.A(new_n755), .B(KEYINPUT92), .Z(new_n756));
  AOI21_X1  g331(.A(new_n745), .B1(new_n756), .B2(G29), .ZN(new_n757));
  XOR2_X1   g332(.A(KEYINPUT27), .B(G1996), .Z(new_n758));
  XNOR2_X1  g333(.A(new_n757), .B(new_n758), .ZN(new_n759));
  NOR3_X1   g334(.A1(new_n738), .A2(new_n744), .A3(new_n759), .ZN(new_n760));
  INV_X1    g335(.A(KEYINPUT93), .ZN(new_n761));
  NOR2_X1   g336(.A1(G5), .A2(G16), .ZN(new_n762));
  AOI211_X1 g337(.A(new_n761), .B(new_n762), .C1(G171), .C2(G16), .ZN(new_n763));
  AOI21_X1  g338(.A(new_n763), .B1(new_n761), .B2(new_n762), .ZN(new_n764));
  XNOR2_X1  g339(.A(new_n764), .B(G1961), .ZN(new_n765));
  INV_X1    g340(.A(KEYINPUT28), .ZN(new_n766));
  AND2_X1   g341(.A1(new_n734), .A2(G26), .ZN(new_n767));
  OR2_X1    g342(.A1(G104), .A2(G2105), .ZN(new_n768));
  OAI211_X1 g343(.A(new_n768), .B(G2104), .C1(G116), .C2(new_n460), .ZN(new_n769));
  INV_X1    g344(.A(G140), .ZN(new_n770));
  INV_X1    g345(.A(G128), .ZN(new_n771));
  OAI221_X1 g346(.A(new_n769), .B1(new_n476), .B2(new_n770), .C1(new_n771), .C2(new_n473), .ZN(new_n772));
  AOI211_X1 g347(.A(new_n766), .B(new_n767), .C1(new_n772), .C2(G29), .ZN(new_n773));
  AOI21_X1  g348(.A(new_n773), .B1(new_n766), .B2(new_n767), .ZN(new_n774));
  XOR2_X1   g349(.A(KEYINPUT87), .B(G2067), .Z(new_n775));
  XNOR2_X1  g350(.A(new_n774), .B(new_n775), .ZN(new_n776));
  NAND2_X1  g351(.A1(new_n630), .A2(G29), .ZN(new_n777));
  INV_X1    g352(.A(G28), .ZN(new_n778));
  OR2_X1    g353(.A1(new_n778), .A2(KEYINPUT30), .ZN(new_n779));
  AOI21_X1  g354(.A(G29), .B1(new_n778), .B2(KEYINPUT30), .ZN(new_n780));
  OR2_X1    g355(.A1(KEYINPUT31), .A2(G11), .ZN(new_n781));
  NAND2_X1  g356(.A1(KEYINPUT31), .A2(G11), .ZN(new_n782));
  AOI22_X1  g357(.A1(new_n779), .A2(new_n780), .B1(new_n781), .B2(new_n782), .ZN(new_n783));
  AND2_X1   g358(.A1(KEYINPUT24), .A2(G34), .ZN(new_n784));
  NOR2_X1   g359(.A1(KEYINPUT24), .A2(G34), .ZN(new_n785));
  OAI21_X1  g360(.A(new_n734), .B1(new_n784), .B2(new_n785), .ZN(new_n786));
  XNOR2_X1  g361(.A(new_n786), .B(KEYINPUT90), .ZN(new_n787));
  INV_X1    g362(.A(G160), .ZN(new_n788));
  OAI21_X1  g363(.A(new_n787), .B1(new_n788), .B2(new_n734), .ZN(new_n789));
  XNOR2_X1  g364(.A(new_n789), .B(G2084), .ZN(new_n790));
  NAND4_X1  g365(.A1(new_n776), .A2(new_n777), .A3(new_n783), .A4(new_n790), .ZN(new_n791));
  NAND2_X1  g366(.A1(new_n734), .A2(G27), .ZN(new_n792));
  XNOR2_X1  g367(.A(new_n792), .B(KEYINPUT94), .ZN(new_n793));
  NAND2_X1  g368(.A1(new_n492), .A2(new_n494), .ZN(new_n794));
  INV_X1    g369(.A(new_n490), .ZN(new_n795));
  AOI21_X1  g370(.A(new_n489), .B1(new_n483), .B2(new_n486), .ZN(new_n796));
  OAI21_X1  g371(.A(new_n794), .B1(new_n795), .B2(new_n796), .ZN(new_n797));
  AOI21_X1  g372(.A(new_n793), .B1(new_n797), .B2(G29), .ZN(new_n798));
  XNOR2_X1  g373(.A(new_n798), .B(G2078), .ZN(new_n799));
  OAI21_X1  g374(.A(new_n799), .B1(new_n741), .B2(new_n742), .ZN(new_n800));
  NAND2_X1  g375(.A1(G168), .A2(G16), .ZN(new_n801));
  OAI21_X1  g376(.A(new_n801), .B1(G16), .B2(G21), .ZN(new_n802));
  INV_X1    g377(.A(G1966), .ZN(new_n803));
  OR2_X1    g378(.A1(new_n802), .A2(new_n803), .ZN(new_n804));
  NAND2_X1  g379(.A1(new_n802), .A2(new_n803), .ZN(new_n805));
  OAI211_X1 g380(.A(new_n804), .B(new_n805), .C1(new_n735), .C2(new_n736), .ZN(new_n806));
  NOR3_X1   g381(.A1(new_n791), .A2(new_n800), .A3(new_n806), .ZN(new_n807));
  NAND3_X1  g382(.A1(new_n760), .A2(new_n765), .A3(new_n807), .ZN(new_n808));
  NAND2_X1  g383(.A1(new_n700), .A2(G19), .ZN(new_n809));
  OAI21_X1  g384(.A(new_n809), .B1(new_n555), .B2(new_n700), .ZN(new_n810));
  NOR2_X1   g385(.A1(new_n810), .A2(G1341), .ZN(new_n811));
  NAND2_X1  g386(.A1(new_n700), .A2(G20), .ZN(new_n812));
  INV_X1    g387(.A(KEYINPUT23), .ZN(new_n813));
  NOR2_X1   g388(.A1(new_n812), .A2(new_n813), .ZN(new_n814));
  INV_X1    g389(.A(G299), .ZN(new_n815));
  OAI21_X1  g390(.A(KEYINPUT23), .B1(new_n815), .B2(new_n700), .ZN(new_n816));
  AOI21_X1  g391(.A(new_n814), .B1(new_n816), .B2(new_n812), .ZN(new_n817));
  XNOR2_X1  g392(.A(new_n817), .B(G1956), .ZN(new_n818));
  NAND2_X1  g393(.A1(new_n810), .A2(G1341), .ZN(new_n819));
  NAND2_X1  g394(.A1(new_n818), .A2(new_n819), .ZN(new_n820));
  NOR3_X1   g395(.A1(new_n808), .A2(new_n811), .A3(new_n820), .ZN(new_n821));
  NAND3_X1  g396(.A1(new_n721), .A2(new_n726), .A3(new_n821), .ZN(G150));
  XNOR2_X1  g397(.A(G150), .B(KEYINPUT96), .ZN(G311));
  NAND2_X1  g398(.A1(G80), .A2(G543), .ZN(new_n824));
  INV_X1    g399(.A(G67), .ZN(new_n825));
  OAI21_X1  g400(.A(new_n824), .B1(new_n509), .B2(new_n825), .ZN(new_n826));
  AOI22_X1  g401(.A1(G651), .A2(new_n826), .B1(new_n510), .B2(G93), .ZN(new_n827));
  NAND3_X1  g402(.A1(new_n534), .A2(G55), .A3(new_n524), .ZN(new_n828));
  NAND3_X1  g403(.A1(new_n827), .A2(KEYINPUT97), .A3(new_n828), .ZN(new_n829));
  INV_X1    g404(.A(new_n829), .ZN(new_n830));
  AOI21_X1  g405(.A(KEYINPUT97), .B1(new_n827), .B2(new_n828), .ZN(new_n831));
  NOR2_X1   g406(.A1(new_n830), .A2(new_n831), .ZN(new_n832));
  NAND2_X1  g407(.A1(new_n832), .A2(G860), .ZN(new_n833));
  XNOR2_X1  g408(.A(new_n833), .B(KEYINPUT98), .ZN(new_n834));
  XNOR2_X1  g409(.A(new_n834), .B(KEYINPUT37), .ZN(new_n835));
  NAND2_X1  g410(.A1(new_n613), .A2(G559), .ZN(new_n836));
  XOR2_X1   g411(.A(new_n836), .B(KEYINPUT38), .Z(new_n837));
  NAND2_X1  g412(.A1(new_n827), .A2(new_n828), .ZN(new_n838));
  OAI211_X1 g413(.A(new_n547), .B(new_n838), .C1(new_n552), .C2(new_n553), .ZN(new_n839));
  OAI21_X1  g414(.A(new_n839), .B1(new_n555), .B2(new_n832), .ZN(new_n840));
  XOR2_X1   g415(.A(new_n840), .B(KEYINPUT39), .Z(new_n841));
  AND2_X1   g416(.A1(new_n837), .A2(new_n841), .ZN(new_n842));
  OR2_X1    g417(.A1(new_n842), .A2(G860), .ZN(new_n843));
  NOR2_X1   g418(.A1(new_n837), .A2(new_n841), .ZN(new_n844));
  OAI21_X1  g419(.A(new_n835), .B1(new_n843), .B2(new_n844), .ZN(G145));
  NAND2_X1  g420(.A1(new_n477), .A2(G142), .ZN(new_n846));
  NOR2_X1   g421(.A1(new_n460), .A2(G118), .ZN(new_n847));
  OAI21_X1  g422(.A(G2104), .B1(G106), .B2(G2105), .ZN(new_n848));
  OAI21_X1  g423(.A(new_n846), .B1(new_n847), .B2(new_n848), .ZN(new_n849));
  AOI21_X1  g424(.A(new_n849), .B1(G130), .B2(new_n474), .ZN(new_n850));
  XOR2_X1   g425(.A(new_n850), .B(KEYINPUT100), .Z(new_n851));
  AND2_X1   g426(.A1(new_n483), .A2(new_n486), .ZN(new_n852));
  NAND2_X1  g427(.A1(new_n794), .A2(new_n852), .ZN(new_n853));
  XNOR2_X1  g428(.A(new_n853), .B(new_n633), .ZN(new_n854));
  XNOR2_X1  g429(.A(new_n851), .B(new_n854), .ZN(new_n855));
  NAND2_X1  g430(.A1(new_n756), .A2(new_n772), .ZN(new_n856));
  INV_X1    g431(.A(new_n856), .ZN(new_n857));
  NOR2_X1   g432(.A1(new_n756), .A2(new_n772), .ZN(new_n858));
  OAI21_X1  g433(.A(new_n715), .B1(new_n857), .B2(new_n858), .ZN(new_n859));
  XOR2_X1   g434(.A(new_n481), .B(KEYINPUT99), .Z(new_n860));
  XNOR2_X1  g435(.A(new_n860), .B(new_n788), .ZN(new_n861));
  INV_X1    g436(.A(new_n861), .ZN(new_n862));
  OR2_X1    g437(.A1(new_n756), .A2(new_n772), .ZN(new_n863));
  INV_X1    g438(.A(new_n715), .ZN(new_n864));
  NAND3_X1  g439(.A1(new_n863), .A2(new_n864), .A3(new_n856), .ZN(new_n865));
  NAND3_X1  g440(.A1(new_n859), .A2(new_n862), .A3(new_n865), .ZN(new_n866));
  INV_X1    g441(.A(new_n866), .ZN(new_n867));
  AOI21_X1  g442(.A(new_n862), .B1(new_n859), .B2(new_n865), .ZN(new_n868));
  OAI21_X1  g443(.A(new_n855), .B1(new_n867), .B2(new_n868), .ZN(new_n869));
  XOR2_X1   g444(.A(new_n630), .B(new_n733), .Z(new_n870));
  NAND2_X1  g445(.A1(new_n859), .A2(new_n865), .ZN(new_n871));
  NAND2_X1  g446(.A1(new_n871), .A2(new_n861), .ZN(new_n872));
  INV_X1    g447(.A(new_n855), .ZN(new_n873));
  NAND3_X1  g448(.A1(new_n872), .A2(new_n873), .A3(new_n866), .ZN(new_n874));
  NAND3_X1  g449(.A1(new_n869), .A2(new_n870), .A3(new_n874), .ZN(new_n875));
  INV_X1    g450(.A(G37), .ZN(new_n876));
  AND2_X1   g451(.A1(new_n875), .A2(new_n876), .ZN(new_n877));
  NAND2_X1  g452(.A1(new_n869), .A2(new_n874), .ZN(new_n878));
  INV_X1    g453(.A(new_n870), .ZN(new_n879));
  NAND2_X1  g454(.A1(new_n878), .A2(new_n879), .ZN(new_n880));
  NAND2_X1  g455(.A1(new_n877), .A2(new_n880), .ZN(new_n881));
  XNOR2_X1  g456(.A(new_n881), .B(KEYINPUT40), .ZN(G395));
  XNOR2_X1  g457(.A(new_n620), .B(KEYINPUT101), .ZN(new_n883));
  XNOR2_X1  g458(.A(new_n883), .B(new_n840), .ZN(new_n884));
  INV_X1    g459(.A(KEYINPUT41), .ZN(new_n885));
  INV_X1    g460(.A(KEYINPUT102), .ZN(new_n886));
  NAND3_X1  g461(.A1(new_n609), .A2(new_n886), .A3(new_n815), .ZN(new_n887));
  NAND3_X1  g462(.A1(new_n604), .A2(G299), .A3(new_n608), .ZN(new_n888));
  NAND2_X1  g463(.A1(new_n887), .A2(new_n888), .ZN(new_n889));
  AOI21_X1  g464(.A(new_n886), .B1(new_n609), .B2(new_n815), .ZN(new_n890));
  OAI21_X1  g465(.A(new_n885), .B1(new_n889), .B2(new_n890), .ZN(new_n891));
  INV_X1    g466(.A(new_n890), .ZN(new_n892));
  NAND4_X1  g467(.A1(new_n892), .A2(KEYINPUT41), .A3(new_n888), .A4(new_n887), .ZN(new_n893));
  NAND2_X1  g468(.A1(new_n891), .A2(new_n893), .ZN(new_n894));
  NAND2_X1  g469(.A1(new_n884), .A2(new_n894), .ZN(new_n895));
  NOR2_X1   g470(.A1(new_n889), .A2(new_n890), .ZN(new_n896));
  OAI21_X1  g471(.A(new_n895), .B1(new_n896), .B2(new_n884), .ZN(new_n897));
  NAND2_X1  g472(.A1(G290), .A2(G288), .ZN(new_n898));
  NAND3_X1  g473(.A1(new_n587), .A2(new_n592), .A3(new_n696), .ZN(new_n899));
  AND3_X1   g474(.A1(new_n898), .A2(G303), .A3(new_n899), .ZN(new_n900));
  AOI21_X1  g475(.A(G303), .B1(new_n898), .B2(new_n899), .ZN(new_n901));
  OR3_X1    g476(.A1(new_n900), .A2(new_n901), .A3(G305), .ZN(new_n902));
  OAI21_X1  g477(.A(G305), .B1(new_n900), .B2(new_n901), .ZN(new_n903));
  NAND2_X1  g478(.A1(new_n902), .A2(new_n903), .ZN(new_n904));
  XNOR2_X1  g479(.A(new_n904), .B(KEYINPUT42), .ZN(new_n905));
  XNOR2_X1  g480(.A(new_n897), .B(new_n905), .ZN(new_n906));
  NAND2_X1  g481(.A1(new_n906), .A2(G868), .ZN(new_n907));
  OR2_X1    g482(.A1(new_n830), .A2(new_n831), .ZN(new_n908));
  OAI21_X1  g483(.A(new_n907), .B1(G868), .B2(new_n908), .ZN(G295));
  OAI21_X1  g484(.A(new_n907), .B1(G868), .B2(new_n908), .ZN(G331));
  INV_X1    g485(.A(KEYINPUT43), .ZN(new_n911));
  NAND2_X1  g486(.A1(new_n908), .A2(new_n554), .ZN(new_n912));
  INV_X1    g487(.A(new_n538), .ZN(new_n913));
  NAND3_X1  g488(.A1(new_n913), .A2(G168), .A3(new_n536), .ZN(new_n914));
  OAI21_X1  g489(.A(G286), .B1(new_n537), .B2(new_n538), .ZN(new_n915));
  NAND4_X1  g490(.A1(new_n912), .A2(new_n839), .A3(new_n914), .A4(new_n915), .ZN(new_n916));
  INV_X1    g491(.A(KEYINPUT103), .ZN(new_n917));
  NAND2_X1  g492(.A1(new_n916), .A2(new_n917), .ZN(new_n918));
  NAND2_X1  g493(.A1(new_n915), .A2(new_n914), .ZN(new_n919));
  INV_X1    g494(.A(new_n919), .ZN(new_n920));
  NAND4_X1  g495(.A1(new_n920), .A2(KEYINPUT103), .A3(new_n839), .A4(new_n912), .ZN(new_n921));
  INV_X1    g496(.A(KEYINPUT104), .ZN(new_n922));
  AND3_X1   g497(.A1(new_n840), .A2(new_n922), .A3(new_n919), .ZN(new_n923));
  AOI21_X1  g498(.A(new_n922), .B1(new_n840), .B2(new_n919), .ZN(new_n924));
  OAI211_X1 g499(.A(new_n918), .B(new_n921), .C1(new_n923), .C2(new_n924), .ZN(new_n925));
  NAND2_X1  g500(.A1(new_n925), .A2(new_n894), .ZN(new_n926));
  AOI21_X1  g501(.A(KEYINPUT105), .B1(new_n840), .B2(new_n919), .ZN(new_n927));
  NAND2_X1  g502(.A1(new_n927), .A2(new_n916), .ZN(new_n928));
  NAND4_X1  g503(.A1(new_n920), .A2(KEYINPUT105), .A3(new_n839), .A4(new_n912), .ZN(new_n929));
  NAND2_X1  g504(.A1(new_n928), .A2(new_n929), .ZN(new_n930));
  INV_X1    g505(.A(new_n896), .ZN(new_n931));
  NAND2_X1  g506(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  INV_X1    g507(.A(new_n904), .ZN(new_n933));
  NAND3_X1  g508(.A1(new_n926), .A2(new_n932), .A3(new_n933), .ZN(new_n934));
  NAND2_X1  g509(.A1(new_n934), .A2(new_n876), .ZN(new_n935));
  AOI22_X1  g510(.A1(new_n894), .A2(new_n925), .B1(new_n930), .B2(new_n931), .ZN(new_n936));
  NOR2_X1   g511(.A1(new_n936), .A2(new_n933), .ZN(new_n937));
  OAI21_X1  g512(.A(new_n911), .B1(new_n935), .B2(new_n937), .ZN(new_n938));
  NAND3_X1  g513(.A1(new_n928), .A2(new_n894), .A3(new_n929), .ZN(new_n939));
  OAI21_X1  g514(.A(new_n939), .B1(new_n925), .B2(new_n896), .ZN(new_n940));
  NAND2_X1  g515(.A1(new_n940), .A2(new_n904), .ZN(new_n941));
  INV_X1    g516(.A(KEYINPUT107), .ZN(new_n942));
  NAND2_X1  g517(.A1(new_n941), .A2(new_n942), .ZN(new_n943));
  AOI21_X1  g518(.A(G37), .B1(new_n936), .B2(new_n933), .ZN(new_n944));
  NAND3_X1  g519(.A1(new_n940), .A2(KEYINPUT107), .A3(new_n904), .ZN(new_n945));
  NAND3_X1  g520(.A1(new_n943), .A2(new_n944), .A3(new_n945), .ZN(new_n946));
  OAI21_X1  g521(.A(new_n938), .B1(new_n946), .B2(new_n911), .ZN(new_n947));
  NAND2_X1  g522(.A1(new_n947), .A2(KEYINPUT44), .ZN(new_n948));
  NAND4_X1  g523(.A1(new_n943), .A2(new_n944), .A3(new_n911), .A4(new_n945), .ZN(new_n949));
  OAI21_X1  g524(.A(KEYINPUT43), .B1(new_n935), .B2(new_n937), .ZN(new_n950));
  NAND3_X1  g525(.A1(new_n949), .A2(new_n950), .A3(KEYINPUT106), .ZN(new_n951));
  INV_X1    g526(.A(KEYINPUT106), .ZN(new_n952));
  OAI211_X1 g527(.A(new_n952), .B(KEYINPUT43), .C1(new_n935), .C2(new_n937), .ZN(new_n953));
  NAND2_X1  g528(.A1(new_n951), .A2(new_n953), .ZN(new_n954));
  OAI21_X1  g529(.A(new_n948), .B1(new_n954), .B2(KEYINPUT44), .ZN(G397));
  INV_X1    g530(.A(G1384), .ZN(new_n956));
  NAND2_X1  g531(.A1(new_n853), .A2(new_n956), .ZN(new_n957));
  INV_X1    g532(.A(KEYINPUT45), .ZN(new_n958));
  NAND2_X1  g533(.A1(new_n957), .A2(new_n958), .ZN(new_n959));
  NAND2_X1  g534(.A1(new_n466), .A2(new_n468), .ZN(new_n960));
  INV_X1    g535(.A(G125), .ZN(new_n961));
  OAI21_X1  g536(.A(new_n463), .B1(new_n960), .B2(new_n961), .ZN(new_n962));
  NAND2_X1  g537(.A1(new_n962), .A2(G2105), .ZN(new_n963));
  NAND4_X1  g538(.A1(new_n963), .A2(G40), .A3(new_n470), .A4(new_n469), .ZN(new_n964));
  NOR2_X1   g539(.A1(new_n959), .A2(new_n964), .ZN(new_n965));
  XOR2_X1   g540(.A(new_n965), .B(KEYINPUT108), .Z(new_n966));
  XNOR2_X1  g541(.A(new_n756), .B(G1996), .ZN(new_n967));
  INV_X1    g542(.A(G2067), .ZN(new_n968));
  XNOR2_X1  g543(.A(new_n772), .B(new_n968), .ZN(new_n969));
  AND2_X1   g544(.A1(new_n967), .A2(new_n969), .ZN(new_n970));
  INV_X1    g545(.A(new_n707), .ZN(new_n971));
  XNOR2_X1  g546(.A(new_n715), .B(new_n971), .ZN(new_n972));
  NAND2_X1  g547(.A1(new_n970), .A2(new_n972), .ZN(new_n973));
  OAI21_X1  g548(.A(KEYINPUT109), .B1(G290), .B2(G1986), .ZN(new_n974));
  NAND2_X1  g549(.A1(G290), .A2(G1986), .ZN(new_n975));
  MUX2_X1   g550(.A(KEYINPUT109), .B(new_n974), .S(new_n975), .Z(new_n976));
  OAI21_X1  g551(.A(new_n966), .B1(new_n973), .B2(new_n976), .ZN(new_n977));
  INV_X1    g552(.A(G8), .ZN(new_n978));
  INV_X1    g553(.A(G40), .ZN(new_n979));
  NOR3_X1   g554(.A1(new_n464), .A2(new_n979), .A3(new_n471), .ZN(new_n980));
  AOI21_X1  g555(.A(G1384), .B1(new_n794), .B2(new_n852), .ZN(new_n981));
  OAI21_X1  g556(.A(new_n980), .B1(new_n981), .B2(KEYINPUT45), .ZN(new_n982));
  NAND2_X1  g557(.A1(new_n982), .A2(KEYINPUT111), .ZN(new_n983));
  INV_X1    g558(.A(KEYINPUT111), .ZN(new_n984));
  OAI211_X1 g559(.A(new_n984), .B(new_n980), .C1(new_n981), .C2(KEYINPUT45), .ZN(new_n985));
  NAND2_X1  g560(.A1(new_n488), .A2(new_n490), .ZN(new_n986));
  AOI21_X1  g561(.A(G1384), .B1(new_n986), .B2(new_n794), .ZN(new_n987));
  NAND2_X1  g562(.A1(new_n987), .A2(KEYINPUT45), .ZN(new_n988));
  NAND3_X1  g563(.A1(new_n983), .A2(new_n985), .A3(new_n988), .ZN(new_n989));
  NAND2_X1  g564(.A1(new_n989), .A2(new_n803), .ZN(new_n990));
  OAI21_X1  g565(.A(new_n980), .B1(new_n957), .B2(KEYINPUT50), .ZN(new_n991));
  INV_X1    g566(.A(KEYINPUT50), .ZN(new_n992));
  AOI21_X1  g567(.A(new_n992), .B1(new_n797), .B2(new_n956), .ZN(new_n993));
  NOR2_X1   g568(.A1(new_n991), .A2(new_n993), .ZN(new_n994));
  INV_X1    g569(.A(G2084), .ZN(new_n995));
  NAND2_X1  g570(.A1(new_n994), .A2(new_n995), .ZN(new_n996));
  AOI21_X1  g571(.A(new_n978), .B1(new_n990), .B2(new_n996), .ZN(new_n997));
  NAND2_X1  g572(.A1(new_n997), .A2(G168), .ZN(new_n998));
  OAI21_X1  g573(.A(KEYINPUT50), .B1(G164), .B2(G1384), .ZN(new_n999));
  AOI21_X1  g574(.A(new_n964), .B1(new_n992), .B2(new_n981), .ZN(new_n1000));
  NAND2_X1  g575(.A1(new_n999), .A2(new_n1000), .ZN(new_n1001));
  NOR2_X1   g576(.A1(new_n1001), .A2(G2090), .ZN(new_n1002));
  OAI21_X1  g577(.A(new_n958), .B1(G164), .B2(G1384), .ZN(new_n1003));
  AOI21_X1  g578(.A(new_n964), .B1(KEYINPUT45), .B2(new_n981), .ZN(new_n1004));
  AOI21_X1  g579(.A(G1971), .B1(new_n1003), .B2(new_n1004), .ZN(new_n1005));
  OAI21_X1  g580(.A(G8), .B1(new_n1002), .B2(new_n1005), .ZN(new_n1006));
  NOR2_X1   g581(.A1(G166), .A2(new_n978), .ZN(new_n1007));
  XNOR2_X1  g582(.A(KEYINPUT110), .B(KEYINPUT55), .ZN(new_n1008));
  NAND2_X1  g583(.A1(new_n1007), .A2(new_n1008), .ZN(new_n1009));
  INV_X1    g584(.A(KEYINPUT110), .ZN(new_n1010));
  NAND2_X1  g585(.A1(new_n1010), .A2(KEYINPUT55), .ZN(new_n1011));
  OAI21_X1  g586(.A(new_n1009), .B1(new_n1007), .B2(new_n1011), .ZN(new_n1012));
  NOR2_X1   g587(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1013));
  INV_X1    g588(.A(KEYINPUT63), .ZN(new_n1014));
  NOR3_X1   g589(.A1(new_n998), .A2(new_n1013), .A3(new_n1014), .ZN(new_n1015));
  INV_X1    g590(.A(KEYINPUT112), .ZN(new_n1016));
  INV_X1    g591(.A(new_n1012), .ZN(new_n1017));
  NAND2_X1  g592(.A1(new_n994), .A2(new_n742), .ZN(new_n1018));
  NAND2_X1  g593(.A1(new_n1003), .A2(new_n1004), .ZN(new_n1019));
  INV_X1    g594(.A(G1971), .ZN(new_n1020));
  NAND2_X1  g595(.A1(new_n1019), .A2(new_n1020), .ZN(new_n1021));
  AOI21_X1  g596(.A(new_n978), .B1(new_n1018), .B2(new_n1021), .ZN(new_n1022));
  NOR2_X1   g597(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1023));
  AOI21_X1  g598(.A(new_n978), .B1(new_n980), .B2(new_n981), .ZN(new_n1024));
  INV_X1    g599(.A(G1976), .ZN(new_n1025));
  AOI21_X1  g600(.A(KEYINPUT52), .B1(G288), .B2(new_n1025), .ZN(new_n1026));
  OAI211_X1 g601(.A(new_n1024), .B(new_n1026), .C1(new_n1025), .C2(G288), .ZN(new_n1027));
  INV_X1    g602(.A(new_n1024), .ZN(new_n1028));
  AOI21_X1  g603(.A(new_n1028), .B1(G1976), .B2(new_n696), .ZN(new_n1029));
  INV_X1    g604(.A(KEYINPUT52), .ZN(new_n1030));
  NAND2_X1  g605(.A1(G305), .A2(G1981), .ZN(new_n1031));
  INV_X1    g606(.A(G1981), .ZN(new_n1032));
  NAND3_X1  g607(.A1(new_n579), .A2(new_n1032), .A3(new_n585), .ZN(new_n1033));
  NAND3_X1  g608(.A1(new_n1031), .A2(KEYINPUT49), .A3(new_n1033), .ZN(new_n1034));
  NAND2_X1  g609(.A1(new_n1034), .A2(new_n1024), .ZN(new_n1035));
  AOI21_X1  g610(.A(KEYINPUT49), .B1(new_n1031), .B2(new_n1033), .ZN(new_n1036));
  OAI221_X1 g611(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1037));
  OAI21_X1  g612(.A(new_n1016), .B1(new_n1023), .B2(new_n1037), .ZN(new_n1038));
  NOR2_X1   g613(.A1(new_n1035), .A2(new_n1036), .ZN(new_n1039));
  OAI21_X1  g614(.A(new_n1027), .B1(new_n1029), .B2(new_n1030), .ZN(new_n1040));
  NOR2_X1   g615(.A1(new_n1039), .A2(new_n1040), .ZN(new_n1041));
  NAND2_X1  g616(.A1(new_n1006), .A2(new_n1012), .ZN(new_n1042));
  NAND3_X1  g617(.A1(new_n1041), .A2(KEYINPUT112), .A3(new_n1042), .ZN(new_n1043));
  NAND3_X1  g618(.A1(new_n1015), .A2(new_n1038), .A3(new_n1043), .ZN(new_n1044));
  OAI21_X1  g619(.A(new_n980), .B1(new_n981), .B2(new_n992), .ZN(new_n1045));
  INV_X1    g620(.A(new_n1045), .ZN(new_n1046));
  NAND2_X1  g621(.A1(new_n987), .A2(new_n992), .ZN(new_n1047));
  NAND3_X1  g622(.A1(new_n1046), .A2(new_n1047), .A3(new_n742), .ZN(new_n1048));
  AND2_X1   g623(.A1(new_n1021), .A2(new_n1048), .ZN(new_n1049));
  OAI21_X1  g624(.A(new_n1012), .B1(new_n1049), .B2(new_n978), .ZN(new_n1050));
  NAND2_X1  g625(.A1(new_n1017), .A2(new_n1022), .ZN(new_n1051));
  NAND3_X1  g626(.A1(new_n1041), .A2(new_n1050), .A3(new_n1051), .ZN(new_n1052));
  OAI21_X1  g627(.A(new_n1014), .B1(new_n1052), .B2(new_n998), .ZN(new_n1053));
  NAND2_X1  g628(.A1(new_n1044), .A2(new_n1053), .ZN(new_n1054));
  OAI211_X1 g629(.A(new_n1025), .B(new_n696), .C1(new_n1035), .C2(new_n1036), .ZN(new_n1055));
  AOI21_X1  g630(.A(new_n1028), .B1(new_n1055), .B2(new_n1033), .ZN(new_n1056));
  AOI21_X1  g631(.A(new_n1056), .B1(new_n1013), .B2(new_n1041), .ZN(new_n1057));
  NAND2_X1  g632(.A1(new_n1054), .A2(new_n1057), .ZN(new_n1058));
  AOI22_X1  g633(.A1(new_n982), .A2(KEYINPUT111), .B1(new_n987), .B2(KEYINPUT45), .ZN(new_n1059));
  AOI21_X1  g634(.A(G1966), .B1(new_n1059), .B2(new_n985), .ZN(new_n1060));
  NOR2_X1   g635(.A1(new_n1001), .A2(G2084), .ZN(new_n1061));
  OAI21_X1  g636(.A(KEYINPUT118), .B1(new_n1060), .B2(new_n1061), .ZN(new_n1062));
  INV_X1    g637(.A(KEYINPUT118), .ZN(new_n1063));
  NAND3_X1  g638(.A1(new_n990), .A2(new_n1063), .A3(new_n996), .ZN(new_n1064));
  NOR2_X1   g639(.A1(G168), .A2(new_n978), .ZN(new_n1065));
  NAND3_X1  g640(.A1(new_n1062), .A2(new_n1064), .A3(new_n1065), .ZN(new_n1066));
  INV_X1    g641(.A(KEYINPUT51), .ZN(new_n1067));
  NAND3_X1  g642(.A1(new_n1062), .A2(new_n1064), .A3(G8), .ZN(new_n1068));
  XNOR2_X1  g643(.A(new_n1065), .B(KEYINPUT119), .ZN(new_n1069));
  AOI21_X1  g644(.A(new_n1067), .B1(new_n1068), .B2(new_n1069), .ZN(new_n1070));
  NOR3_X1   g645(.A1(new_n997), .A2(KEYINPUT51), .A3(new_n1065), .ZN(new_n1071));
  OAI21_X1  g646(.A(new_n1066), .B1(new_n1070), .B2(new_n1071), .ZN(new_n1072));
  NAND2_X1  g647(.A1(new_n1072), .A2(KEYINPUT120), .ZN(new_n1073));
  INV_X1    g648(.A(KEYINPUT120), .ZN(new_n1074));
  OAI211_X1 g649(.A(new_n1074), .B(new_n1066), .C1(new_n1070), .C2(new_n1071), .ZN(new_n1075));
  NAND2_X1  g650(.A1(new_n1073), .A2(new_n1075), .ZN(new_n1076));
  NAND2_X1  g651(.A1(new_n980), .A2(new_n981), .ZN(new_n1077));
  OAI21_X1  g652(.A(KEYINPUT114), .B1(new_n1077), .B2(G2067), .ZN(new_n1078));
  INV_X1    g653(.A(KEYINPUT114), .ZN(new_n1079));
  NAND4_X1  g654(.A1(new_n980), .A2(new_n981), .A3(new_n1079), .A4(new_n968), .ZN(new_n1080));
  NAND2_X1  g655(.A1(new_n1078), .A2(new_n1080), .ZN(new_n1081));
  AOI21_X1  g656(.A(G1348), .B1(new_n999), .B2(new_n1000), .ZN(new_n1082));
  OAI21_X1  g657(.A(KEYINPUT115), .B1(new_n1081), .B2(new_n1082), .ZN(new_n1083));
  OAI21_X1  g658(.A(new_n725), .B1(new_n991), .B2(new_n993), .ZN(new_n1084));
  INV_X1    g659(.A(KEYINPUT115), .ZN(new_n1085));
  NAND4_X1  g660(.A1(new_n1084), .A2(new_n1085), .A3(new_n1078), .A4(new_n1080), .ZN(new_n1086));
  NAND2_X1  g661(.A1(new_n1083), .A2(new_n1086), .ZN(new_n1087));
  AOI21_X1  g662(.A(new_n609), .B1(new_n1087), .B2(KEYINPUT60), .ZN(new_n1088));
  INV_X1    g663(.A(KEYINPUT60), .ZN(new_n1089));
  AND2_X1   g664(.A1(new_n604), .A2(new_n608), .ZN(new_n1090));
  AOI211_X1 g665(.A(new_n1089), .B(new_n1090), .C1(new_n1083), .C2(new_n1086), .ZN(new_n1091));
  OAI22_X1  g666(.A1(new_n1088), .A2(new_n1091), .B1(KEYINPUT60), .B2(new_n1087), .ZN(new_n1092));
  XOR2_X1   g667(.A(KEYINPUT58), .B(G1341), .Z(new_n1093));
  NAND2_X1  g668(.A1(new_n1077), .A2(new_n1093), .ZN(new_n1094));
  OAI21_X1  g669(.A(new_n1094), .B1(new_n1019), .B2(G1996), .ZN(new_n1095));
  NAND2_X1  g670(.A1(new_n1095), .A2(new_n555), .ZN(new_n1096));
  INV_X1    g671(.A(KEYINPUT59), .ZN(new_n1097));
  NOR2_X1   g672(.A1(new_n1097), .A2(KEYINPUT117), .ZN(new_n1098));
  NAND2_X1  g673(.A1(new_n1096), .A2(new_n1098), .ZN(new_n1099));
  OAI211_X1 g674(.A(new_n1095), .B(new_n555), .C1(KEYINPUT117), .C2(new_n1097), .ZN(new_n1100));
  NAND2_X1  g675(.A1(new_n1099), .A2(new_n1100), .ZN(new_n1101));
  INV_X1    g676(.A(KEYINPUT61), .ZN(new_n1102));
  INV_X1    g677(.A(KEYINPUT113), .ZN(new_n1103));
  INV_X1    g678(.A(KEYINPUT9), .ZN(new_n1104));
  XNOR2_X1  g679(.A(new_n562), .B(new_n1104), .ZN(new_n1105));
  INV_X1    g680(.A(new_n567), .ZN(new_n1106));
  OAI211_X1 g681(.A(new_n1103), .B(KEYINPUT57), .C1(new_n1105), .C2(new_n1106), .ZN(new_n1107));
  OR2_X1    g682(.A1(new_n1103), .A2(KEYINPUT57), .ZN(new_n1108));
  NAND2_X1  g683(.A1(new_n1103), .A2(KEYINPUT57), .ZN(new_n1109));
  NAND4_X1  g684(.A1(new_n563), .A2(new_n567), .A3(new_n1108), .A4(new_n1109), .ZN(new_n1110));
  AND2_X1   g685(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1111));
  INV_X1    g686(.A(G1956), .ZN(new_n1112));
  NOR3_X1   g687(.A1(G164), .A2(KEYINPUT50), .A3(G1384), .ZN(new_n1113));
  OAI21_X1  g688(.A(new_n1112), .B1(new_n1113), .B2(new_n1045), .ZN(new_n1114));
  XNOR2_X1  g689(.A(KEYINPUT56), .B(G2072), .ZN(new_n1115));
  NAND3_X1  g690(.A1(new_n1003), .A2(new_n1004), .A3(new_n1115), .ZN(new_n1116));
  NAND3_X1  g691(.A1(new_n1111), .A2(new_n1114), .A3(new_n1116), .ZN(new_n1117));
  INV_X1    g692(.A(new_n1117), .ZN(new_n1118));
  AOI21_X1  g693(.A(new_n1111), .B1(new_n1114), .B2(new_n1116), .ZN(new_n1119));
  OAI21_X1  g694(.A(new_n1102), .B1(new_n1118), .B2(new_n1119), .ZN(new_n1120));
  NAND2_X1  g695(.A1(new_n1114), .A2(new_n1116), .ZN(new_n1121));
  NAND2_X1  g696(.A1(new_n1107), .A2(new_n1110), .ZN(new_n1122));
  NAND2_X1  g697(.A1(new_n1121), .A2(new_n1122), .ZN(new_n1123));
  NAND3_X1  g698(.A1(new_n1123), .A2(KEYINPUT61), .A3(new_n1117), .ZN(new_n1124));
  AND3_X1   g699(.A1(new_n1101), .A2(new_n1120), .A3(new_n1124), .ZN(new_n1125));
  OAI21_X1  g700(.A(KEYINPUT116), .B1(new_n1087), .B2(new_n609), .ZN(new_n1126));
  INV_X1    g701(.A(KEYINPUT116), .ZN(new_n1127));
  NAND4_X1  g702(.A1(new_n1083), .A2(new_n1086), .A3(new_n1127), .A4(new_n1090), .ZN(new_n1128));
  NAND3_X1  g703(.A1(new_n1126), .A2(new_n1128), .A3(new_n1123), .ZN(new_n1129));
  AOI22_X1  g704(.A1(new_n1092), .A2(new_n1125), .B1(new_n1129), .B2(new_n1117), .ZN(new_n1130));
  INV_X1    g705(.A(new_n1052), .ZN(new_n1131));
  INV_X1    g706(.A(G2078), .ZN(new_n1132));
  NAND3_X1  g707(.A1(new_n1003), .A2(new_n1004), .A3(new_n1132), .ZN(new_n1133));
  INV_X1    g708(.A(KEYINPUT53), .ZN(new_n1134));
  NAND2_X1  g709(.A1(new_n1133), .A2(new_n1134), .ZN(new_n1135));
  INV_X1    g710(.A(G1961), .ZN(new_n1136));
  NAND2_X1  g711(.A1(new_n1001), .A2(new_n1136), .ZN(new_n1137));
  NAND2_X1  g712(.A1(new_n1132), .A2(KEYINPUT53), .ZN(new_n1138));
  OAI211_X1 g713(.A(new_n1135), .B(new_n1137), .C1(new_n989), .C2(new_n1138), .ZN(new_n1139));
  AND3_X1   g714(.A1(new_n1139), .A2(KEYINPUT121), .A3(G171), .ZN(new_n1140));
  AOI21_X1  g715(.A(KEYINPUT121), .B1(new_n1139), .B2(G171), .ZN(new_n1141));
  INV_X1    g716(.A(KEYINPUT54), .ZN(new_n1142));
  NAND4_X1  g717(.A1(new_n1004), .A2(new_n959), .A3(KEYINPUT53), .A4(new_n1132), .ZN(new_n1143));
  NAND3_X1  g718(.A1(new_n1135), .A2(new_n1137), .A3(new_n1143), .ZN(new_n1144));
  OAI21_X1  g719(.A(new_n1142), .B1(new_n1144), .B2(G171), .ZN(new_n1145));
  NOR3_X1   g720(.A1(new_n1140), .A2(new_n1141), .A3(new_n1145), .ZN(new_n1146));
  AOI21_X1  g721(.A(new_n1142), .B1(new_n1139), .B2(G301), .ZN(new_n1147));
  NAND4_X1  g722(.A1(new_n1135), .A2(new_n1137), .A3(G171), .A4(new_n1143), .ZN(new_n1148));
  AND2_X1   g723(.A1(new_n1147), .A2(new_n1148), .ZN(new_n1149));
  OAI21_X1  g724(.A(new_n1131), .B1(new_n1146), .B2(new_n1149), .ZN(new_n1150));
  NOR2_X1   g725(.A1(new_n1130), .A2(new_n1150), .ZN(new_n1151));
  AOI21_X1  g726(.A(new_n1058), .B1(new_n1076), .B2(new_n1151), .ZN(new_n1152));
  INV_X1    g727(.A(KEYINPUT122), .ZN(new_n1153));
  INV_X1    g728(.A(KEYINPUT62), .ZN(new_n1154));
  NAND3_X1  g729(.A1(new_n1073), .A2(new_n1154), .A3(new_n1075), .ZN(new_n1155));
  NOR2_X1   g730(.A1(new_n1140), .A2(new_n1141), .ZN(new_n1156));
  NOR2_X1   g731(.A1(new_n1156), .A2(new_n1052), .ZN(new_n1157));
  NAND2_X1  g732(.A1(new_n1155), .A2(new_n1157), .ZN(new_n1158));
  AOI21_X1  g733(.A(new_n1154), .B1(new_n1073), .B2(new_n1075), .ZN(new_n1159));
  OAI22_X1  g734(.A1(new_n1152), .A2(new_n1153), .B1(new_n1158), .B2(new_n1159), .ZN(new_n1160));
  AOI211_X1 g735(.A(KEYINPUT122), .B(new_n1058), .C1(new_n1076), .C2(new_n1151), .ZN(new_n1161));
  OAI21_X1  g736(.A(new_n977), .B1(new_n1160), .B2(new_n1161), .ZN(new_n1162));
  NAND3_X1  g737(.A1(new_n970), .A2(new_n971), .A3(new_n716), .ZN(new_n1163));
  OAI21_X1  g738(.A(new_n1163), .B1(G2067), .B2(new_n772), .ZN(new_n1164));
  NAND2_X1  g739(.A1(new_n1164), .A2(new_n966), .ZN(new_n1165));
  NAND2_X1  g740(.A1(new_n973), .A2(new_n966), .ZN(new_n1166));
  NOR2_X1   g741(.A1(G290), .A2(G1986), .ZN(new_n1167));
  AND2_X1   g742(.A1(new_n966), .A2(new_n1167), .ZN(new_n1168));
  NAND2_X1  g743(.A1(new_n1168), .A2(KEYINPUT48), .ZN(new_n1169));
  OR2_X1    g744(.A1(new_n1168), .A2(KEYINPUT48), .ZN(new_n1170));
  NAND3_X1  g745(.A1(new_n1166), .A2(new_n1169), .A3(new_n1170), .ZN(new_n1171));
  INV_X1    g746(.A(G1996), .ZN(new_n1172));
  NAND2_X1  g747(.A1(new_n966), .A2(new_n1172), .ZN(new_n1173));
  INV_X1    g748(.A(KEYINPUT46), .ZN(new_n1174));
  NAND2_X1  g749(.A1(new_n756), .A2(new_n969), .ZN(new_n1175));
  AOI22_X1  g750(.A1(new_n1173), .A2(new_n1174), .B1(new_n966), .B2(new_n1175), .ZN(new_n1176));
  OAI21_X1  g751(.A(new_n1176), .B1(new_n1174), .B2(new_n1173), .ZN(new_n1177));
  XNOR2_X1  g752(.A(KEYINPUT123), .B(KEYINPUT47), .ZN(new_n1178));
  OAI211_X1 g753(.A(new_n1165), .B(new_n1171), .C1(new_n1177), .C2(new_n1178), .ZN(new_n1179));
  AOI21_X1  g754(.A(new_n1179), .B1(new_n1177), .B2(new_n1178), .ZN(new_n1180));
  NAND2_X1  g755(.A1(new_n1162), .A2(new_n1180), .ZN(new_n1181));
  INV_X1    g756(.A(KEYINPUT124), .ZN(new_n1182));
  NAND2_X1  g757(.A1(new_n1181), .A2(new_n1182), .ZN(new_n1183));
  NAND3_X1  g758(.A1(new_n1162), .A2(KEYINPUT124), .A3(new_n1180), .ZN(new_n1184));
  NAND2_X1  g759(.A1(new_n1183), .A2(new_n1184), .ZN(G329));
  assign    G231 = 1'b0;
  NOR3_X1   g760(.A1(G229), .A2(new_n458), .A3(G227), .ZN(new_n1187));
  OAI21_X1  g761(.A(new_n1187), .B1(new_n652), .B2(new_n651), .ZN(new_n1188));
  AOI21_X1  g762(.A(new_n1188), .B1(new_n877), .B2(new_n880), .ZN(new_n1189));
  NAND3_X1  g763(.A1(new_n951), .A2(new_n1189), .A3(new_n953), .ZN(new_n1190));
  NAND2_X1  g764(.A1(new_n1190), .A2(KEYINPUT125), .ZN(new_n1191));
  INV_X1    g765(.A(KEYINPUT125), .ZN(new_n1192));
  NAND4_X1  g766(.A1(new_n951), .A2(new_n1189), .A3(new_n1192), .A4(new_n953), .ZN(new_n1193));
  AND3_X1   g767(.A1(new_n1191), .A2(KEYINPUT126), .A3(new_n1193), .ZN(new_n1194));
  AOI21_X1  g768(.A(KEYINPUT126), .B1(new_n1191), .B2(new_n1193), .ZN(new_n1195));
  NOR2_X1   g769(.A1(new_n1194), .A2(new_n1195), .ZN(G308));
  NAND2_X1  g770(.A1(new_n1191), .A2(new_n1193), .ZN(G225));
endmodule


