//Secret key is'0 0 0 0 1 1 0 1 0 1 0 0 0 1 1 1 1 0 1 1 1 0 1 1 1 0 0 0 0 0 1 1 1 1 1 1 0 0 0 1 1 0 1 1 0 1 0 0 0 0 0 1 1 1 1 1 0 1 1 1 1 1 0 0 1 0 0 1 1 1 1 0 1 0 1 0 0 0 1 1 0 1 0 0 1 0 0 0 0 0 0 0 1 0 1 0 1 0 1 1 1 0 0 0 1 0 0 0 0 1 0 1 0 1 1 1 0 0 1 0 0 0 1 1 0 0 1' ..
// Benchmark "locked_locked_c1355" written by ABC on Sat Dec 16 05:17:59 2023

module locked_locked_c1355 ( 
    KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68, KEYINPUT69,
    KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74, KEYINPUT75,
    KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80, KEYINPUT81,
    KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86, KEYINPUT87,
    KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92, KEYINPUT93,
    KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98, KEYINPUT99,
    KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103, KEYINPUT104,
    KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108, KEYINPUT109,
    KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113, KEYINPUT114,
    KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118, KEYINPUT119,
    KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123, KEYINPUT124,
    KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0, KEYINPUT1, KEYINPUT2,
    KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6, KEYINPUT7, KEYINPUT8,
    KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12, KEYINPUT13, KEYINPUT14,
    KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18, KEYINPUT19, KEYINPUT20,
    KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24, KEYINPUT25, KEYINPUT26,
    KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30, KEYINPUT31, KEYINPUT32,
    KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36, KEYINPUT37, KEYINPUT38,
    KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42, KEYINPUT43, KEYINPUT44,
    KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48, KEYINPUT49, KEYINPUT50,
    KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54, KEYINPUT55, KEYINPUT56,
    KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60, KEYINPUT61, KEYINPUT62,
    KEYINPUT63, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat,
    G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat,
    G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat,
    G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat,
    G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat,
    G232gat, G233gat,
    G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat  );
  input  KEYINPUT64, KEYINPUT65, KEYINPUT66, KEYINPUT67, KEYINPUT68,
    KEYINPUT69, KEYINPUT70, KEYINPUT71, KEYINPUT72, KEYINPUT73, KEYINPUT74,
    KEYINPUT75, KEYINPUT76, KEYINPUT77, KEYINPUT78, KEYINPUT79, KEYINPUT80,
    KEYINPUT81, KEYINPUT82, KEYINPUT83, KEYINPUT84, KEYINPUT85, KEYINPUT86,
    KEYINPUT87, KEYINPUT88, KEYINPUT89, KEYINPUT90, KEYINPUT91, KEYINPUT92,
    KEYINPUT93, KEYINPUT94, KEYINPUT95, KEYINPUT96, KEYINPUT97, KEYINPUT98,
    KEYINPUT99, KEYINPUT100, KEYINPUT101, KEYINPUT102, KEYINPUT103,
    KEYINPUT104, KEYINPUT105, KEYINPUT106, KEYINPUT107, KEYINPUT108,
    KEYINPUT109, KEYINPUT110, KEYINPUT111, KEYINPUT112, KEYINPUT113,
    KEYINPUT114, KEYINPUT115, KEYINPUT116, KEYINPUT117, KEYINPUT118,
    KEYINPUT119, KEYINPUT120, KEYINPUT121, KEYINPUT122, KEYINPUT123,
    KEYINPUT124, KEYINPUT125, KEYINPUT126, KEYINPUT127, KEYINPUT0,
    KEYINPUT1, KEYINPUT2, KEYINPUT3, KEYINPUT4, KEYINPUT5, KEYINPUT6,
    KEYINPUT7, KEYINPUT8, KEYINPUT9, KEYINPUT10, KEYINPUT11, KEYINPUT12,
    KEYINPUT13, KEYINPUT14, KEYINPUT15, KEYINPUT16, KEYINPUT17, KEYINPUT18,
    KEYINPUT19, KEYINPUT20, KEYINPUT21, KEYINPUT22, KEYINPUT23, KEYINPUT24,
    KEYINPUT25, KEYINPUT26, KEYINPUT27, KEYINPUT28, KEYINPUT29, KEYINPUT30,
    KEYINPUT31, KEYINPUT32, KEYINPUT33, KEYINPUT34, KEYINPUT35, KEYINPUT36,
    KEYINPUT37, KEYINPUT38, KEYINPUT39, KEYINPUT40, KEYINPUT41, KEYINPUT42,
    KEYINPUT43, KEYINPUT44, KEYINPUT45, KEYINPUT46, KEYINPUT47, KEYINPUT48,
    KEYINPUT49, KEYINPUT50, KEYINPUT51, KEYINPUT52, KEYINPUT53, KEYINPUT54,
    KEYINPUT55, KEYINPUT56, KEYINPUT57, KEYINPUT58, KEYINPUT59, KEYINPUT60,
    KEYINPUT61, KEYINPUT62, KEYINPUT63, G1gat, G8gat, G15gat, G22gat,
    G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat,
    G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat,
    G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat,
    G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat,
    G230gat, G231gat, G232gat, G233gat;
  output G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat,
    G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat,
    G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat,
    G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat,
    G1352gat, G1353gat, G1354gat, G1355gat;
  wire new_n202, new_n203, new_n204, new_n205, new_n206, new_n207, new_n208,
    new_n209, new_n210, new_n211, new_n212, new_n213, new_n214, new_n215,
    new_n216, new_n217, new_n218, new_n219, new_n220, new_n221, new_n222,
    new_n223, new_n224, new_n225, new_n226, new_n227, new_n228, new_n229,
    new_n230, new_n231, new_n232, new_n233, new_n234, new_n235, new_n236,
    new_n237, new_n238, new_n239, new_n240, new_n241, new_n242, new_n243,
    new_n244, new_n245, new_n246, new_n247, new_n248, new_n249, new_n250,
    new_n251, new_n252, new_n253, new_n254, new_n255, new_n256, new_n257,
    new_n258, new_n259, new_n260, new_n261, new_n262, new_n263, new_n264,
    new_n265, new_n266, new_n267, new_n268, new_n269, new_n270, new_n271,
    new_n272, new_n273, new_n274, new_n275, new_n276, new_n277, new_n278,
    new_n279, new_n280, new_n281, new_n282, new_n283, new_n284, new_n285,
    new_n286, new_n287, new_n288, new_n289, new_n290, new_n291, new_n292,
    new_n293, new_n294, new_n295, new_n296, new_n297, new_n298, new_n299,
    new_n300, new_n301, new_n302, new_n303, new_n304, new_n305, new_n306,
    new_n307, new_n308, new_n309, new_n310, new_n311, new_n312, new_n313,
    new_n314, new_n315, new_n316, new_n317, new_n318, new_n319, new_n320,
    new_n321, new_n322, new_n323, new_n324, new_n325, new_n326, new_n327,
    new_n328, new_n329, new_n330, new_n331, new_n332, new_n333, new_n334,
    new_n335, new_n336, new_n337, new_n338, new_n339, new_n340, new_n341,
    new_n342, new_n343, new_n344, new_n345, new_n346, new_n347, new_n348,
    new_n349, new_n350, new_n351, new_n352, new_n353, new_n354, new_n355,
    new_n356, new_n357, new_n358, new_n359, new_n360, new_n361, new_n362,
    new_n363, new_n364, new_n365, new_n366, new_n367, new_n368, new_n369,
    new_n370, new_n371, new_n372, new_n373, new_n374, new_n375, new_n376,
    new_n377, new_n378, new_n379, new_n380, new_n381, new_n382, new_n383,
    new_n384, new_n385, new_n386, new_n387, new_n388, new_n389, new_n390,
    new_n391, new_n392, new_n393, new_n394, new_n395, new_n396, new_n397,
    new_n398, new_n399, new_n400, new_n401, new_n402, new_n403, new_n404,
    new_n405, new_n406, new_n407, new_n408, new_n409, new_n410, new_n411,
    new_n412, new_n413, new_n414, new_n415, new_n416, new_n417, new_n418,
    new_n419, new_n420, new_n421, new_n422, new_n423, new_n424, new_n425,
    new_n426, new_n427, new_n428, new_n429, new_n430, new_n431, new_n432,
    new_n433, new_n434, new_n435, new_n436, new_n437, new_n438, new_n439,
    new_n440, new_n441, new_n442, new_n443, new_n444, new_n445, new_n446,
    new_n447, new_n448, new_n449, new_n450, new_n451, new_n452, new_n453,
    new_n454, new_n455, new_n456, new_n457, new_n458, new_n459, new_n460,
    new_n461, new_n462, new_n463, new_n464, new_n465, new_n466, new_n467,
    new_n468, new_n469, new_n470, new_n471, new_n472, new_n473, new_n474,
    new_n475, new_n476, new_n477, new_n478, new_n479, new_n480, new_n481,
    new_n482, new_n483, new_n484, new_n485, new_n486, new_n487, new_n488,
    new_n489, new_n490, new_n491, new_n492, new_n493, new_n494, new_n495,
    new_n496, new_n497, new_n498, new_n499, new_n500, new_n501, new_n502,
    new_n503, new_n504, new_n505, new_n506, new_n507, new_n508, new_n509,
    new_n510, new_n511, new_n512, new_n513, new_n514, new_n515, new_n516,
    new_n517, new_n518, new_n519, new_n520, new_n521, new_n522, new_n523,
    new_n524, new_n525, new_n526, new_n527, new_n528, new_n529, new_n530,
    new_n531, new_n532, new_n533, new_n534, new_n535, new_n536, new_n537,
    new_n538, new_n539, new_n540, new_n541, new_n542, new_n543, new_n544,
    new_n545, new_n546, new_n547, new_n548, new_n549, new_n550, new_n551,
    new_n552, new_n553, new_n554, new_n555, new_n556, new_n557, new_n558,
    new_n559, new_n560, new_n561, new_n562, new_n563, new_n564, new_n565,
    new_n566, new_n567, new_n568, new_n569, new_n570, new_n571, new_n572,
    new_n573, new_n574, new_n575, new_n576, new_n577, new_n578, new_n579,
    new_n580, new_n581, new_n582, new_n583, new_n584, new_n585, new_n586,
    new_n587, new_n588, new_n589, new_n590, new_n591, new_n592, new_n593,
    new_n594, new_n595, new_n596, new_n597, new_n598, new_n599, new_n600,
    new_n601, new_n602, new_n603, new_n604, new_n605, new_n606, new_n607,
    new_n608, new_n609, new_n610, new_n611, new_n612, new_n613, new_n614,
    new_n615, new_n616, new_n617, new_n618, new_n619, new_n620, new_n621,
    new_n622, new_n623, new_n624, new_n625, new_n627, new_n628, new_n629,
    new_n630, new_n631, new_n632, new_n634, new_n635, new_n636, new_n637,
    new_n638, new_n640, new_n641, new_n642, new_n644, new_n645, new_n646,
    new_n647, new_n648, new_n649, new_n650, new_n651, new_n652, new_n653,
    new_n654, new_n655, new_n656, new_n657, new_n658, new_n659, new_n660,
    new_n661, new_n662, new_n663, new_n665, new_n666, new_n667, new_n668,
    new_n669, new_n670, new_n672, new_n673, new_n674, new_n675, new_n676,
    new_n677, new_n678, new_n679, new_n681, new_n682, new_n683, new_n684,
    new_n685, new_n686, new_n687, new_n689, new_n690, new_n691, new_n693,
    new_n694, new_n695, new_n697, new_n698, new_n699, new_n700, new_n701,
    new_n702, new_n704, new_n705, new_n707, new_n708, new_n709, new_n710,
    new_n711, new_n712, new_n713, new_n714, new_n715, new_n716, new_n717,
    new_n718, new_n719, new_n720, new_n722, new_n723, new_n724, new_n725,
    new_n726, new_n727, new_n728, new_n729, new_n730, new_n731, new_n733,
    new_n734, new_n735, new_n736, new_n738, new_n739, new_n740, new_n741,
    new_n742, new_n743, new_n744, new_n745, new_n746, new_n748, new_n749,
    new_n750, new_n751, new_n752, new_n753, new_n754, new_n755, new_n756,
    new_n757, new_n758, new_n759, new_n760, new_n761, new_n762, new_n763,
    new_n764, new_n765, new_n766, new_n767, new_n768, new_n769, new_n770,
    new_n771, new_n772, new_n773, new_n774, new_n775, new_n776, new_n777,
    new_n778, new_n779, new_n780, new_n781, new_n782, new_n783, new_n784,
    new_n785, new_n786, new_n787, new_n788, new_n789, new_n790, new_n791,
    new_n792, new_n793, new_n794, new_n795, new_n796, new_n797, new_n798,
    new_n799, new_n800, new_n801, new_n802, new_n803, new_n804, new_n805,
    new_n806, new_n807, new_n809, new_n810, new_n811, new_n813, new_n814,
    new_n816, new_n817, new_n818, new_n819, new_n820, new_n821, new_n822,
    new_n823, new_n825, new_n826, new_n827, new_n828, new_n829, new_n830,
    new_n831, new_n832, new_n833, new_n834, new_n835, new_n836, new_n837,
    new_n838, new_n839, new_n840, new_n841, new_n842, new_n843, new_n844,
    new_n845, new_n846, new_n847, new_n849, new_n850, new_n851, new_n852,
    new_n853, new_n854, new_n855, new_n856, new_n857, new_n858, new_n859,
    new_n860, new_n861, new_n862, new_n863, new_n864, new_n865, new_n866,
    new_n867, new_n868, new_n869, new_n870, new_n872, new_n873, new_n875,
    new_n876, new_n878, new_n879, new_n880, new_n881, new_n882, new_n883,
    new_n884, new_n885, new_n886, new_n887, new_n888, new_n890, new_n891,
    new_n893, new_n894, new_n895, new_n896, new_n897, new_n898, new_n900,
    new_n901, new_n902, new_n903, new_n905, new_n906, new_n907, new_n908,
    new_n909, new_n910, new_n911, new_n912, new_n913, new_n915, new_n916,
    new_n917, new_n918, new_n919, new_n921, new_n922, new_n923, new_n924,
    new_n925, new_n926, new_n927, new_n928, new_n929, new_n930, new_n931,
    new_n932, new_n933, new_n934, new_n935, new_n936, new_n937, new_n938,
    new_n940, new_n941;
  NAND2_X1  g000(.A1(G155gat), .A2(G162gat), .ZN(new_n202));
  XNOR2_X1  g001(.A(new_n202), .B(KEYINPUT78), .ZN(new_n203));
  NOR2_X1   g002(.A1(G155gat), .A2(G162gat), .ZN(new_n204));
  NOR2_X1   g003(.A1(new_n204), .A2(KEYINPUT77), .ZN(new_n205));
  XNOR2_X1  g004(.A(new_n203), .B(new_n205), .ZN(new_n206));
  INV_X1    g005(.A(G141gat), .ZN(new_n207));
  OR2_X1    g006(.A1(new_n207), .A2(G148gat), .ZN(new_n208));
  NAND2_X1  g007(.A1(new_n207), .A2(G148gat), .ZN(new_n209));
  AOI22_X1  g008(.A1(new_n208), .A2(new_n209), .B1(KEYINPUT2), .B2(new_n202), .ZN(new_n210));
  NOR2_X1   g009(.A1(new_n206), .A2(new_n210), .ZN(new_n211));
  INV_X1    g010(.A(new_n204), .ZN(new_n212));
  AND3_X1   g011(.A1(new_n210), .A2(new_n202), .A3(new_n212), .ZN(new_n213));
  OR2_X1    g012(.A1(new_n211), .A2(new_n213), .ZN(new_n214));
  INV_X1    g013(.A(KEYINPUT3), .ZN(new_n215));
  AOI21_X1  g014(.A(KEYINPUT29), .B1(new_n214), .B2(new_n215), .ZN(new_n216));
  XOR2_X1   g015(.A(G197gat), .B(G204gat), .Z(new_n217));
  AOI21_X1  g016(.A(KEYINPUT22), .B1(G211gat), .B2(G218gat), .ZN(new_n218));
  NOR2_X1   g017(.A1(new_n217), .A2(new_n218), .ZN(new_n219));
  XNOR2_X1  g018(.A(G211gat), .B(G218gat), .ZN(new_n220));
  NAND2_X1  g019(.A1(new_n219), .A2(new_n220), .ZN(new_n221));
  NAND2_X1  g020(.A1(new_n221), .A2(KEYINPUT74), .ZN(new_n222));
  NOR2_X1   g021(.A1(new_n219), .A2(new_n220), .ZN(new_n223));
  INV_X1    g022(.A(new_n223), .ZN(new_n224));
  XNOR2_X1  g023(.A(new_n222), .B(new_n224), .ZN(new_n225));
  NOR2_X1   g024(.A1(new_n216), .A2(new_n225), .ZN(new_n226));
  INV_X1    g025(.A(KEYINPUT29), .ZN(new_n227));
  NAND2_X1  g026(.A1(new_n225), .A2(new_n227), .ZN(new_n228));
  AOI21_X1  g027(.A(new_n214), .B1(new_n228), .B2(new_n215), .ZN(new_n229));
  OAI211_X1 g028(.A(G228gat), .B(G233gat), .C1(new_n226), .C2(new_n229), .ZN(new_n230));
  NAND2_X1  g029(.A1(G228gat), .A2(G233gat), .ZN(new_n231));
  INV_X1    g030(.A(KEYINPUT85), .ZN(new_n232));
  NAND3_X1  g031(.A1(new_n224), .A2(new_n232), .A3(new_n221), .ZN(new_n233));
  AOI21_X1  g032(.A(KEYINPUT29), .B1(new_n223), .B2(KEYINPUT85), .ZN(new_n234));
  AOI21_X1  g033(.A(KEYINPUT3), .B1(new_n233), .B2(new_n234), .ZN(new_n235));
  OAI221_X1 g034(.A(new_n231), .B1(new_n214), .B2(new_n235), .C1(new_n216), .C2(new_n225), .ZN(new_n236));
  NAND2_X1  g035(.A1(new_n230), .A2(new_n236), .ZN(new_n237));
  XNOR2_X1  g036(.A(KEYINPUT84), .B(KEYINPUT31), .ZN(new_n238));
  NAND2_X1  g037(.A1(new_n237), .A2(new_n238), .ZN(new_n239));
  XNOR2_X1  g038(.A(G78gat), .B(G106gat), .ZN(new_n240));
  INV_X1    g039(.A(G50gat), .ZN(new_n241));
  XNOR2_X1  g040(.A(new_n240), .B(new_n241), .ZN(new_n242));
  XNOR2_X1  g041(.A(new_n242), .B(G22gat), .ZN(new_n243));
  OR2_X1    g042(.A1(new_n237), .A2(new_n238), .ZN(new_n244));
  AND3_X1   g043(.A1(new_n239), .A2(new_n243), .A3(new_n244), .ZN(new_n245));
  AOI21_X1  g044(.A(new_n243), .B1(new_n244), .B2(new_n239), .ZN(new_n246));
  NOR2_X1   g045(.A1(new_n245), .A2(new_n246), .ZN(new_n247));
  XNOR2_X1  g046(.A(KEYINPUT87), .B(KEYINPUT39), .ZN(new_n248));
  NOR2_X1   g047(.A1(new_n211), .A2(new_n213), .ZN(new_n249));
  XNOR2_X1  g048(.A(new_n249), .B(new_n215), .ZN(new_n250));
  XNOR2_X1  g049(.A(KEYINPUT67), .B(G127gat), .ZN(new_n251));
  INV_X1    g050(.A(G134gat), .ZN(new_n252));
  OR3_X1    g051(.A1(new_n251), .A2(KEYINPUT68), .A3(new_n252), .ZN(new_n253));
  XNOR2_X1  g052(.A(G113gat), .B(G120gat), .ZN(new_n254));
  NOR2_X1   g053(.A1(new_n251), .A2(new_n252), .ZN(new_n255));
  INV_X1    g054(.A(G127gat), .ZN(new_n256));
  OAI21_X1  g055(.A(KEYINPUT68), .B1(new_n256), .B2(G134gat), .ZN(new_n257));
  OAI221_X1 g056(.A(new_n253), .B1(KEYINPUT1), .B2(new_n254), .C1(new_n255), .C2(new_n257), .ZN(new_n258));
  NOR2_X1   g057(.A1(new_n252), .A2(G127gat), .ZN(new_n259));
  INV_X1    g058(.A(KEYINPUT1), .ZN(new_n260));
  OAI21_X1  g059(.A(new_n260), .B1(new_n256), .B2(G134gat), .ZN(new_n261));
  AOI211_X1 g060(.A(new_n259), .B(new_n261), .C1(new_n254), .C2(KEYINPUT69), .ZN(new_n262));
  OAI21_X1  g061(.A(new_n262), .B1(KEYINPUT69), .B2(new_n254), .ZN(new_n263));
  NAND2_X1  g062(.A1(new_n258), .A2(new_n263), .ZN(new_n264));
  INV_X1    g063(.A(KEYINPUT79), .ZN(new_n265));
  NAND2_X1  g064(.A1(new_n264), .A2(new_n265), .ZN(new_n266));
  NAND3_X1  g065(.A1(new_n258), .A2(KEYINPUT79), .A3(new_n263), .ZN(new_n267));
  AND2_X1   g066(.A1(new_n266), .A2(new_n267), .ZN(new_n268));
  NAND2_X1  g067(.A1(new_n250), .A2(new_n268), .ZN(new_n269));
  INV_X1    g068(.A(KEYINPUT4), .ZN(new_n270));
  INV_X1    g069(.A(new_n264), .ZN(new_n271));
  NAND3_X1  g070(.A1(new_n214), .A2(new_n270), .A3(new_n271), .ZN(new_n272));
  OAI211_X1 g071(.A(new_n258), .B(new_n263), .C1(new_n211), .C2(new_n213), .ZN(new_n273));
  NAND2_X1  g072(.A1(new_n273), .A2(KEYINPUT4), .ZN(new_n274));
  AND3_X1   g073(.A1(new_n272), .A2(KEYINPUT83), .A3(new_n274), .ZN(new_n275));
  AOI21_X1  g074(.A(KEYINPUT83), .B1(new_n272), .B2(new_n274), .ZN(new_n276));
  OAI21_X1  g075(.A(new_n269), .B1(new_n275), .B2(new_n276), .ZN(new_n277));
  INV_X1    g076(.A(KEYINPUT86), .ZN(new_n278));
  NAND2_X1  g077(.A1(G225gat), .A2(G233gat), .ZN(new_n279));
  INV_X1    g078(.A(new_n279), .ZN(new_n280));
  NAND3_X1  g079(.A1(new_n277), .A2(new_n278), .A3(new_n280), .ZN(new_n281));
  INV_X1    g080(.A(new_n281), .ZN(new_n282));
  AOI21_X1  g081(.A(new_n278), .B1(new_n277), .B2(new_n280), .ZN(new_n283));
  OAI21_X1  g082(.A(new_n248), .B1(new_n282), .B2(new_n283), .ZN(new_n284));
  NAND2_X1  g083(.A1(new_n277), .A2(new_n280), .ZN(new_n285));
  NAND2_X1  g084(.A1(new_n285), .A2(KEYINPUT86), .ZN(new_n286));
  NAND3_X1  g085(.A1(new_n266), .A2(new_n249), .A3(new_n267), .ZN(new_n287));
  NAND3_X1  g086(.A1(new_n287), .A2(new_n273), .A3(new_n279), .ZN(new_n288));
  AND2_X1   g087(.A1(new_n288), .A2(KEYINPUT39), .ZN(new_n289));
  NAND3_X1  g088(.A1(new_n286), .A2(new_n281), .A3(new_n289), .ZN(new_n290));
  XOR2_X1   g089(.A(G1gat), .B(G29gat), .Z(new_n291));
  XNOR2_X1  g090(.A(G57gat), .B(G85gat), .ZN(new_n292));
  XNOR2_X1  g091(.A(new_n291), .B(new_n292), .ZN(new_n293));
  XNOR2_X1  g092(.A(KEYINPUT82), .B(KEYINPUT0), .ZN(new_n294));
  XOR2_X1   g093(.A(new_n293), .B(new_n294), .Z(new_n295));
  NAND3_X1  g094(.A1(new_n284), .A2(new_n290), .A3(new_n295), .ZN(new_n296));
  NAND2_X1  g095(.A1(new_n296), .A2(KEYINPUT40), .ZN(new_n297));
  INV_X1    g096(.A(KEYINPUT40), .ZN(new_n298));
  NAND4_X1  g097(.A1(new_n284), .A2(new_n290), .A3(new_n298), .A4(new_n295), .ZN(new_n299));
  NAND2_X1  g098(.A1(new_n297), .A2(new_n299), .ZN(new_n300));
  XOR2_X1   g099(.A(KEYINPUT64), .B(G169gat), .Z(new_n301));
  INV_X1    g100(.A(KEYINPUT23), .ZN(new_n302));
  NOR2_X1   g101(.A1(new_n302), .A2(G176gat), .ZN(new_n303));
  NAND2_X1  g102(.A1(new_n301), .A2(new_n303), .ZN(new_n304));
  NOR2_X1   g103(.A1(G169gat), .A2(G176gat), .ZN(new_n305));
  INV_X1    g104(.A(new_n305), .ZN(new_n306));
  INV_X1    g105(.A(G169gat), .ZN(new_n307));
  INV_X1    g106(.A(G176gat), .ZN(new_n308));
  NOR2_X1   g107(.A1(new_n307), .A2(new_n308), .ZN(new_n309));
  OAI21_X1  g108(.A(new_n306), .B1(new_n309), .B2(new_n302), .ZN(new_n310));
  NOR2_X1   g109(.A1(G183gat), .A2(G190gat), .ZN(new_n311));
  INV_X1    g110(.A(G183gat), .ZN(new_n312));
  NOR2_X1   g111(.A1(new_n312), .A2(KEYINPUT24), .ZN(new_n313));
  NAND2_X1  g112(.A1(G183gat), .A2(G190gat), .ZN(new_n314));
  AOI22_X1  g113(.A1(new_n313), .A2(G190gat), .B1(KEYINPUT24), .B2(new_n314), .ZN(new_n315));
  OAI211_X1 g114(.A(new_n304), .B(new_n310), .C1(new_n311), .C2(new_n315), .ZN(new_n316));
  INV_X1    g115(.A(KEYINPUT25), .ZN(new_n317));
  NAND2_X1  g116(.A1(new_n316), .A2(new_n317), .ZN(new_n318));
  AOI21_X1  g117(.A(new_n317), .B1(new_n303), .B2(new_n307), .ZN(new_n319));
  XOR2_X1   g118(.A(new_n311), .B(KEYINPUT65), .Z(new_n320));
  OAI211_X1 g119(.A(new_n310), .B(new_n319), .C1(new_n320), .C2(new_n315), .ZN(new_n321));
  NAND2_X1  g120(.A1(new_n318), .A2(new_n321), .ZN(new_n322));
  INV_X1    g121(.A(G190gat), .ZN(new_n323));
  OAI21_X1  g122(.A(KEYINPUT27), .B1(new_n312), .B2(KEYINPUT66), .ZN(new_n324));
  OR2_X1    g123(.A1(new_n312), .A2(KEYINPUT27), .ZN(new_n325));
  OAI211_X1 g124(.A(new_n323), .B(new_n324), .C1(new_n325), .C2(KEYINPUT66), .ZN(new_n326));
  INV_X1    g125(.A(KEYINPUT28), .ZN(new_n327));
  NAND2_X1  g126(.A1(new_n326), .A2(new_n327), .ZN(new_n328));
  XNOR2_X1  g127(.A(KEYINPUT27), .B(G183gat), .ZN(new_n329));
  NAND3_X1  g128(.A1(new_n329), .A2(KEYINPUT28), .A3(new_n323), .ZN(new_n330));
  NAND2_X1  g129(.A1(new_n328), .A2(new_n330), .ZN(new_n331));
  OR3_X1    g130(.A1(new_n309), .A2(KEYINPUT26), .A3(new_n305), .ZN(new_n332));
  NAND2_X1  g131(.A1(new_n305), .A2(KEYINPUT26), .ZN(new_n333));
  NAND4_X1  g132(.A1(new_n331), .A2(new_n314), .A3(new_n332), .A4(new_n333), .ZN(new_n334));
  NAND2_X1  g133(.A1(new_n322), .A2(new_n334), .ZN(new_n335));
  AOI22_X1  g134(.A1(new_n335), .A2(new_n227), .B1(G226gat), .B2(G233gat), .ZN(new_n336));
  INV_X1    g135(.A(KEYINPUT75), .ZN(new_n337));
  OR2_X1    g136(.A1(new_n336), .A2(new_n337), .ZN(new_n338));
  AND3_X1   g137(.A1(new_n335), .A2(G226gat), .A3(G233gat), .ZN(new_n339));
  OAI21_X1  g138(.A(new_n337), .B1(new_n339), .B2(new_n336), .ZN(new_n340));
  AOI21_X1  g139(.A(new_n225), .B1(new_n338), .B2(new_n340), .ZN(new_n341));
  NOR2_X1   g140(.A1(new_n339), .A2(new_n336), .ZN(new_n342));
  NAND2_X1  g141(.A1(new_n342), .A2(new_n225), .ZN(new_n343));
  INV_X1    g142(.A(new_n343), .ZN(new_n344));
  NOR2_X1   g143(.A1(new_n341), .A2(new_n344), .ZN(new_n345));
  XOR2_X1   g144(.A(G8gat), .B(G36gat), .Z(new_n346));
  XNOR2_X1  g145(.A(new_n346), .B(KEYINPUT76), .ZN(new_n347));
  XNOR2_X1  g146(.A(G64gat), .B(G92gat), .ZN(new_n348));
  XOR2_X1   g147(.A(new_n347), .B(new_n348), .Z(new_n349));
  NAND2_X1  g148(.A1(new_n345), .A2(new_n349), .ZN(new_n350));
  INV_X1    g149(.A(new_n349), .ZN(new_n351));
  OAI21_X1  g150(.A(new_n351), .B1(new_n341), .B2(new_n344), .ZN(new_n352));
  NAND3_X1  g151(.A1(new_n350), .A2(new_n352), .A3(KEYINPUT30), .ZN(new_n353));
  INV_X1    g152(.A(KEYINPUT30), .ZN(new_n354));
  NAND3_X1  g153(.A1(new_n345), .A2(new_n354), .A3(new_n349), .ZN(new_n355));
  NAND2_X1  g154(.A1(new_n353), .A2(new_n355), .ZN(new_n356));
  AOI21_X1  g155(.A(new_n280), .B1(new_n250), .B2(new_n268), .ZN(new_n357));
  INV_X1    g156(.A(KEYINPUT5), .ZN(new_n358));
  NAND2_X1  g157(.A1(new_n357), .A2(new_n358), .ZN(new_n359));
  NOR2_X1   g158(.A1(new_n275), .A2(new_n276), .ZN(new_n360));
  NOR2_X1   g159(.A1(new_n359), .A2(new_n360), .ZN(new_n361));
  INV_X1    g160(.A(new_n361), .ZN(new_n362));
  INV_X1    g161(.A(KEYINPUT80), .ZN(new_n363));
  NAND4_X1  g162(.A1(new_n214), .A2(new_n363), .A3(new_n270), .A4(new_n271), .ZN(new_n364));
  OAI21_X1  g163(.A(KEYINPUT80), .B1(new_n273), .B2(KEYINPUT4), .ZN(new_n365));
  NAND3_X1  g164(.A1(new_n364), .A2(new_n365), .A3(new_n274), .ZN(new_n366));
  NAND2_X1  g165(.A1(new_n357), .A2(new_n366), .ZN(new_n367));
  INV_X1    g166(.A(KEYINPUT81), .ZN(new_n368));
  NAND2_X1  g167(.A1(new_n287), .A2(new_n273), .ZN(new_n369));
  AOI21_X1  g168(.A(new_n358), .B1(new_n369), .B2(new_n280), .ZN(new_n370));
  AND3_X1   g169(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n371));
  AOI21_X1  g170(.A(new_n368), .B1(new_n367), .B2(new_n370), .ZN(new_n372));
  OAI21_X1  g171(.A(new_n362), .B1(new_n371), .B2(new_n372), .ZN(new_n373));
  AOI21_X1  g172(.A(new_n295), .B1(new_n373), .B2(KEYINPUT88), .ZN(new_n374));
  INV_X1    g173(.A(KEYINPUT88), .ZN(new_n375));
  OAI211_X1 g174(.A(new_n362), .B(new_n375), .C1(new_n371), .C2(new_n372), .ZN(new_n376));
  AOI21_X1  g175(.A(new_n356), .B1(new_n374), .B2(new_n376), .ZN(new_n377));
  AOI21_X1  g176(.A(new_n247), .B1(new_n300), .B2(new_n377), .ZN(new_n378));
  OR2_X1    g177(.A1(new_n341), .A2(new_n344), .ZN(new_n379));
  OAI21_X1  g178(.A(new_n351), .B1(new_n379), .B2(KEYINPUT37), .ZN(new_n380));
  INV_X1    g179(.A(KEYINPUT37), .ZN(new_n381));
  NOR2_X1   g180(.A1(new_n345), .A2(new_n381), .ZN(new_n382));
  OAI21_X1  g181(.A(KEYINPUT38), .B1(new_n380), .B2(new_n382), .ZN(new_n383));
  OR3_X1    g182(.A1(new_n342), .A2(KEYINPUT89), .A3(new_n225), .ZN(new_n384));
  NAND3_X1  g183(.A1(new_n338), .A2(new_n340), .A3(new_n225), .ZN(new_n385));
  OAI21_X1  g184(.A(KEYINPUT89), .B1(new_n342), .B2(new_n225), .ZN(new_n386));
  NAND3_X1  g185(.A1(new_n384), .A2(new_n385), .A3(new_n386), .ZN(new_n387));
  AOI21_X1  g186(.A(KEYINPUT38), .B1(new_n387), .B2(KEYINPUT37), .ZN(new_n388));
  AOI21_X1  g187(.A(new_n349), .B1(new_n345), .B2(new_n381), .ZN(new_n389));
  AOI22_X1  g188(.A1(new_n388), .A2(new_n389), .B1(new_n345), .B2(new_n349), .ZN(new_n390));
  AND2_X1   g189(.A1(new_n383), .A2(new_n390), .ZN(new_n391));
  NAND2_X1  g190(.A1(new_n367), .A2(new_n370), .ZN(new_n392));
  NAND2_X1  g191(.A1(new_n392), .A2(KEYINPUT81), .ZN(new_n393));
  NAND3_X1  g192(.A1(new_n367), .A2(new_n368), .A3(new_n370), .ZN(new_n394));
  AOI21_X1  g193(.A(new_n361), .B1(new_n393), .B2(new_n394), .ZN(new_n395));
  AOI21_X1  g194(.A(KEYINPUT6), .B1(new_n395), .B2(new_n295), .ZN(new_n396));
  INV_X1    g195(.A(new_n295), .ZN(new_n397));
  OAI21_X1  g196(.A(new_n397), .B1(new_n395), .B2(new_n375), .ZN(new_n398));
  INV_X1    g197(.A(new_n376), .ZN(new_n399));
  OAI21_X1  g198(.A(new_n396), .B1(new_n398), .B2(new_n399), .ZN(new_n400));
  NAND3_X1  g199(.A1(new_n373), .A2(KEYINPUT6), .A3(new_n397), .ZN(new_n401));
  OR2_X1    g200(.A1(new_n401), .A2(KEYINPUT90), .ZN(new_n402));
  NAND2_X1  g201(.A1(new_n401), .A2(KEYINPUT90), .ZN(new_n403));
  NAND4_X1  g202(.A1(new_n391), .A2(new_n400), .A3(new_n402), .A4(new_n403), .ZN(new_n404));
  NAND2_X1  g203(.A1(new_n378), .A2(new_n404), .ZN(new_n405));
  INV_X1    g204(.A(KEYINPUT6), .ZN(new_n406));
  OAI21_X1  g205(.A(new_n406), .B1(new_n373), .B2(new_n397), .ZN(new_n407));
  NOR2_X1   g206(.A1(new_n395), .A2(new_n295), .ZN(new_n408));
  OAI21_X1  g207(.A(new_n401), .B1(new_n407), .B2(new_n408), .ZN(new_n409));
  NAND2_X1  g208(.A1(new_n409), .A2(new_n356), .ZN(new_n410));
  OR2_X1    g209(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n411));
  NAND2_X1  g210(.A1(new_n335), .A2(KEYINPUT70), .ZN(new_n412));
  NAND3_X1  g211(.A1(new_n411), .A2(new_n264), .A3(new_n412), .ZN(new_n413));
  INV_X1    g212(.A(G227gat), .ZN(new_n414));
  INV_X1    g213(.A(G233gat), .ZN(new_n415));
  NOR2_X1   g214(.A1(new_n414), .A2(new_n415), .ZN(new_n416));
  NAND3_X1  g215(.A1(new_n335), .A2(new_n271), .A3(KEYINPUT70), .ZN(new_n417));
  NAND3_X1  g216(.A1(new_n413), .A2(new_n416), .A3(new_n417), .ZN(new_n418));
  NAND2_X1  g217(.A1(new_n418), .A2(KEYINPUT32), .ZN(new_n419));
  NAND2_X1  g218(.A1(new_n419), .A2(KEYINPUT71), .ZN(new_n420));
  XNOR2_X1  g219(.A(G15gat), .B(G43gat), .ZN(new_n421));
  XNOR2_X1  g220(.A(new_n421), .B(KEYINPUT72), .ZN(new_n422));
  XOR2_X1   g221(.A(G71gat), .B(G99gat), .Z(new_n423));
  XNOR2_X1  g222(.A(new_n422), .B(new_n423), .ZN(new_n424));
  INV_X1    g223(.A(KEYINPUT71), .ZN(new_n425));
  NAND3_X1  g224(.A1(new_n418), .A2(new_n425), .A3(KEYINPUT32), .ZN(new_n426));
  INV_X1    g225(.A(KEYINPUT33), .ZN(new_n427));
  NAND2_X1  g226(.A1(new_n418), .A2(new_n427), .ZN(new_n428));
  NAND4_X1  g227(.A1(new_n420), .A2(new_n424), .A3(new_n426), .A4(new_n428), .ZN(new_n429));
  OR2_X1    g228(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n430));
  NAND2_X1  g229(.A1(new_n424), .A2(KEYINPUT73), .ZN(new_n431));
  NAND3_X1  g230(.A1(new_n430), .A2(KEYINPUT33), .A3(new_n431), .ZN(new_n432));
  NAND3_X1  g231(.A1(new_n418), .A2(KEYINPUT32), .A3(new_n432), .ZN(new_n433));
  NAND2_X1  g232(.A1(new_n429), .A2(new_n433), .ZN(new_n434));
  NAND2_X1  g233(.A1(new_n413), .A2(new_n417), .ZN(new_n435));
  INV_X1    g234(.A(new_n416), .ZN(new_n436));
  NAND2_X1  g235(.A1(new_n435), .A2(new_n436), .ZN(new_n437));
  AND2_X1   g236(.A1(new_n437), .A2(KEYINPUT34), .ZN(new_n438));
  NOR2_X1   g237(.A1(new_n437), .A2(KEYINPUT34), .ZN(new_n439));
  NOR2_X1   g238(.A1(new_n438), .A2(new_n439), .ZN(new_n440));
  INV_X1    g239(.A(new_n440), .ZN(new_n441));
  NAND2_X1  g240(.A1(new_n434), .A2(new_n441), .ZN(new_n442));
  NAND3_X1  g241(.A1(new_n440), .A2(new_n429), .A3(new_n433), .ZN(new_n443));
  NAND2_X1  g242(.A1(new_n442), .A2(new_n443), .ZN(new_n444));
  INV_X1    g243(.A(KEYINPUT36), .ZN(new_n445));
  NAND2_X1  g244(.A1(new_n444), .A2(new_n445), .ZN(new_n446));
  NAND3_X1  g245(.A1(new_n442), .A2(KEYINPUT36), .A3(new_n443), .ZN(new_n447));
  AOI22_X1  g246(.A1(new_n410), .A2(new_n247), .B1(new_n446), .B2(new_n447), .ZN(new_n448));
  INV_X1    g247(.A(new_n247), .ZN(new_n449));
  INV_X1    g248(.A(new_n444), .ZN(new_n450));
  NAND2_X1  g249(.A1(new_n449), .A2(new_n450), .ZN(new_n451));
  OAI21_X1  g250(.A(KEYINPUT35), .B1(new_n451), .B2(new_n410), .ZN(new_n452));
  NAND3_X1  g251(.A1(new_n400), .A2(new_n402), .A3(new_n403), .ZN(new_n453));
  NOR2_X1   g252(.A1(new_n247), .A2(new_n444), .ZN(new_n454));
  INV_X1    g253(.A(new_n356), .ZN(new_n455));
  NOR2_X1   g254(.A1(new_n455), .A2(KEYINPUT35), .ZN(new_n456));
  NAND3_X1  g255(.A1(new_n453), .A2(new_n454), .A3(new_n456), .ZN(new_n457));
  AOI22_X1  g256(.A1(new_n405), .A2(new_n448), .B1(new_n452), .B2(new_n457), .ZN(new_n458));
  INV_X1    g257(.A(KEYINPUT17), .ZN(new_n459));
  INV_X1    g258(.A(G36gat), .ZN(new_n460));
  AND2_X1   g259(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n461));
  NOR2_X1   g260(.A1(KEYINPUT14), .A2(G29gat), .ZN(new_n462));
  OAI21_X1  g261(.A(new_n460), .B1(new_n461), .B2(new_n462), .ZN(new_n463));
  INV_X1    g262(.A(G29gat), .ZN(new_n464));
  NAND3_X1  g263(.A1(new_n464), .A2(KEYINPUT14), .A3(G36gat), .ZN(new_n465));
  NAND2_X1  g264(.A1(new_n463), .A2(new_n465), .ZN(new_n466));
  INV_X1    g265(.A(G43gat), .ZN(new_n467));
  NAND2_X1  g266(.A1(new_n467), .A2(new_n241), .ZN(new_n468));
  INV_X1    g267(.A(KEYINPUT15), .ZN(new_n469));
  NAND2_X1  g268(.A1(G43gat), .A2(G50gat), .ZN(new_n470));
  NAND3_X1  g269(.A1(new_n468), .A2(new_n469), .A3(new_n470), .ZN(new_n471));
  NAND2_X1  g270(.A1(new_n466), .A2(new_n471), .ZN(new_n472));
  NAND2_X1  g271(.A1(new_n468), .A2(new_n470), .ZN(new_n473));
  INV_X1    g272(.A(KEYINPUT92), .ZN(new_n474));
  NAND2_X1  g273(.A1(new_n473), .A2(new_n474), .ZN(new_n475));
  NAND3_X1  g274(.A1(new_n468), .A2(KEYINPUT92), .A3(new_n470), .ZN(new_n476));
  NAND3_X1  g275(.A1(new_n475), .A2(KEYINPUT15), .A3(new_n476), .ZN(new_n477));
  NAND2_X1  g276(.A1(new_n472), .A2(new_n477), .ZN(new_n478));
  INV_X1    g277(.A(KEYINPUT93), .ZN(new_n479));
  NAND4_X1  g278(.A1(new_n466), .A2(new_n475), .A3(KEYINPUT15), .A4(new_n476), .ZN(new_n480));
  AND3_X1   g279(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n481));
  AOI21_X1  g280(.A(new_n479), .B1(new_n478), .B2(new_n480), .ZN(new_n482));
  OAI21_X1  g281(.A(new_n459), .B1(new_n481), .B2(new_n482), .ZN(new_n483));
  XNOR2_X1  g282(.A(G15gat), .B(G22gat), .ZN(new_n484));
  INV_X1    g283(.A(KEYINPUT16), .ZN(new_n485));
  AOI21_X1  g284(.A(G1gat), .B1(new_n484), .B2(new_n485), .ZN(new_n486));
  INV_X1    g285(.A(new_n486), .ZN(new_n487));
  NAND2_X1  g286(.A1(new_n484), .A2(KEYINPUT94), .ZN(new_n488));
  NAND2_X1  g287(.A1(new_n488), .A2(G8gat), .ZN(new_n489));
  INV_X1    g288(.A(new_n489), .ZN(new_n490));
  NOR2_X1   g289(.A1(new_n488), .A2(G8gat), .ZN(new_n491));
  OAI21_X1  g290(.A(new_n487), .B1(new_n490), .B2(new_n491), .ZN(new_n492));
  INV_X1    g291(.A(new_n491), .ZN(new_n493));
  NAND3_X1  g292(.A1(new_n493), .A2(new_n486), .A3(new_n489), .ZN(new_n494));
  NAND2_X1  g293(.A1(new_n492), .A2(new_n494), .ZN(new_n495));
  NAND2_X1  g294(.A1(new_n478), .A2(new_n480), .ZN(new_n496));
  NAND2_X1  g295(.A1(new_n496), .A2(KEYINPUT17), .ZN(new_n497));
  NAND2_X1  g296(.A1(new_n497), .A2(KEYINPUT95), .ZN(new_n498));
  INV_X1    g297(.A(KEYINPUT95), .ZN(new_n499));
  NAND3_X1  g298(.A1(new_n496), .A2(new_n499), .A3(KEYINPUT17), .ZN(new_n500));
  NAND4_X1  g299(.A1(new_n483), .A2(new_n495), .A3(new_n498), .A4(new_n500), .ZN(new_n501));
  OAI211_X1 g300(.A(new_n494), .B(new_n492), .C1(new_n481), .C2(new_n482), .ZN(new_n502));
  NAND2_X1  g301(.A1(G229gat), .A2(G233gat), .ZN(new_n503));
  NAND4_X1  g302(.A1(new_n501), .A2(KEYINPUT18), .A3(new_n502), .A4(new_n503), .ZN(new_n504));
  INV_X1    g303(.A(new_n482), .ZN(new_n505));
  NAND3_X1  g304(.A1(new_n478), .A2(new_n479), .A3(new_n480), .ZN(new_n506));
  NAND3_X1  g305(.A1(new_n505), .A2(new_n495), .A3(new_n506), .ZN(new_n507));
  NAND2_X1  g306(.A1(new_n502), .A2(new_n507), .ZN(new_n508));
  XOR2_X1   g307(.A(new_n503), .B(KEYINPUT13), .Z(new_n509));
  NAND2_X1  g308(.A1(new_n508), .A2(new_n509), .ZN(new_n510));
  XNOR2_X1  g309(.A(G113gat), .B(G141gat), .ZN(new_n511));
  XNOR2_X1  g310(.A(new_n511), .B(G197gat), .ZN(new_n512));
  XNOR2_X1  g311(.A(KEYINPUT11), .B(G169gat), .ZN(new_n513));
  XOR2_X1   g312(.A(new_n512), .B(new_n513), .Z(new_n514));
  XNOR2_X1  g313(.A(new_n514), .B(KEYINPUT12), .ZN(new_n515));
  AND3_X1   g314(.A1(new_n504), .A2(new_n510), .A3(new_n515), .ZN(new_n516));
  NAND3_X1  g315(.A1(new_n501), .A2(new_n502), .A3(new_n503), .ZN(new_n517));
  INV_X1    g316(.A(KEYINPUT18), .ZN(new_n518));
  NAND2_X1  g317(.A1(new_n517), .A2(new_n518), .ZN(new_n519));
  INV_X1    g318(.A(KEYINPUT96), .ZN(new_n520));
  NAND2_X1  g319(.A1(new_n519), .A2(new_n520), .ZN(new_n521));
  NAND3_X1  g320(.A1(new_n517), .A2(KEYINPUT96), .A3(new_n518), .ZN(new_n522));
  NAND3_X1  g321(.A1(new_n516), .A2(new_n521), .A3(new_n522), .ZN(new_n523));
  NAND3_X1  g322(.A1(new_n519), .A2(new_n510), .A3(new_n504), .ZN(new_n524));
  XNOR2_X1  g323(.A(new_n515), .B(KEYINPUT91), .ZN(new_n525));
  NAND2_X1  g324(.A1(new_n524), .A2(new_n525), .ZN(new_n526));
  NAND2_X1  g325(.A1(new_n523), .A2(new_n526), .ZN(new_n527));
  INV_X1    g326(.A(new_n527), .ZN(new_n528));
  NOR2_X1   g327(.A1(new_n458), .A2(new_n528), .ZN(new_n529));
  INV_X1    g328(.A(new_n409), .ZN(new_n530));
  XOR2_X1   g329(.A(G57gat), .B(G64gat), .Z(new_n531));
  NAND2_X1  g330(.A1(G71gat), .A2(G78gat), .ZN(new_n532));
  INV_X1    g331(.A(KEYINPUT9), .ZN(new_n533));
  NAND2_X1  g332(.A1(new_n532), .A2(new_n533), .ZN(new_n534));
  NAND2_X1  g333(.A1(new_n531), .A2(new_n534), .ZN(new_n535));
  XNOR2_X1  g334(.A(G71gat), .B(G78gat), .ZN(new_n536));
  XOR2_X1   g335(.A(new_n535), .B(new_n536), .Z(new_n537));
  INV_X1    g336(.A(KEYINPUT21), .ZN(new_n538));
  NAND2_X1  g337(.A1(new_n537), .A2(new_n538), .ZN(new_n539));
  NAND2_X1  g338(.A1(G231gat), .A2(G233gat), .ZN(new_n540));
  XNOR2_X1  g339(.A(new_n539), .B(new_n540), .ZN(new_n541));
  XNOR2_X1  g340(.A(new_n541), .B(G127gat), .ZN(new_n542));
  OAI21_X1  g341(.A(new_n495), .B1(new_n537), .B2(new_n538), .ZN(new_n543));
  XNOR2_X1  g342(.A(new_n542), .B(new_n543), .ZN(new_n544));
  XNOR2_X1  g343(.A(KEYINPUT19), .B(KEYINPUT20), .ZN(new_n545));
  INV_X1    g344(.A(G155gat), .ZN(new_n546));
  XNOR2_X1  g345(.A(new_n545), .B(new_n546), .ZN(new_n547));
  XOR2_X1   g346(.A(G183gat), .B(G211gat), .Z(new_n548));
  XNOR2_X1  g347(.A(new_n547), .B(new_n548), .ZN(new_n549));
  INV_X1    g348(.A(new_n549), .ZN(new_n550));
  XNOR2_X1  g349(.A(new_n544), .B(new_n550), .ZN(new_n551));
  INV_X1    g350(.A(new_n551), .ZN(new_n552));
  NAND2_X1  g351(.A1(new_n505), .A2(new_n506), .ZN(new_n553));
  NAND2_X1  g352(.A1(G85gat), .A2(G92gat), .ZN(new_n554));
  XNOR2_X1  g353(.A(new_n554), .B(KEYINPUT7), .ZN(new_n555));
  NAND2_X1  g354(.A1(G99gat), .A2(G106gat), .ZN(new_n556));
  NAND2_X1  g355(.A1(new_n556), .A2(KEYINPUT8), .ZN(new_n557));
  INV_X1    g356(.A(G85gat), .ZN(new_n558));
  INV_X1    g357(.A(G92gat), .ZN(new_n559));
  NAND2_X1  g358(.A1(new_n558), .A2(new_n559), .ZN(new_n560));
  AND3_X1   g359(.A1(new_n557), .A2(KEYINPUT98), .A3(new_n560), .ZN(new_n561));
  AOI21_X1  g360(.A(KEYINPUT98), .B1(new_n557), .B2(new_n560), .ZN(new_n562));
  OAI21_X1  g361(.A(new_n555), .B1(new_n561), .B2(new_n562), .ZN(new_n563));
  XOR2_X1   g362(.A(G99gat), .B(G106gat), .Z(new_n564));
  NAND2_X1  g363(.A1(new_n563), .A2(new_n564), .ZN(new_n565));
  INV_X1    g364(.A(new_n564), .ZN(new_n566));
  OAI211_X1 g365(.A(new_n566), .B(new_n555), .C1(new_n561), .C2(new_n562), .ZN(new_n567));
  NAND3_X1  g366(.A1(new_n565), .A2(KEYINPUT99), .A3(new_n567), .ZN(new_n568));
  OR2_X1    g367(.A1(new_n561), .A2(new_n562), .ZN(new_n569));
  INV_X1    g368(.A(KEYINPUT99), .ZN(new_n570));
  NAND4_X1  g369(.A1(new_n569), .A2(new_n570), .A3(new_n566), .A4(new_n555), .ZN(new_n571));
  NAND2_X1  g370(.A1(new_n568), .A2(new_n571), .ZN(new_n572));
  AND2_X1   g371(.A1(G232gat), .A2(G233gat), .ZN(new_n573));
  AOI22_X1  g372(.A1(new_n553), .A2(new_n572), .B1(KEYINPUT41), .B2(new_n573), .ZN(new_n574));
  INV_X1    g373(.A(new_n572), .ZN(new_n575));
  NAND4_X1  g374(.A1(new_n483), .A2(new_n575), .A3(new_n500), .A4(new_n498), .ZN(new_n576));
  NAND2_X1  g375(.A1(new_n574), .A2(new_n576), .ZN(new_n577));
  XNOR2_X1  g376(.A(G190gat), .B(G218gat), .ZN(new_n578));
  XOR2_X1   g377(.A(new_n578), .B(KEYINPUT100), .Z(new_n579));
  NAND2_X1  g378(.A1(new_n577), .A2(new_n579), .ZN(new_n580));
  INV_X1    g379(.A(new_n580), .ZN(new_n581));
  NOR2_X1   g380(.A1(new_n573), .A2(KEYINPUT41), .ZN(new_n582));
  XNOR2_X1  g381(.A(new_n582), .B(KEYINPUT97), .ZN(new_n583));
  XNOR2_X1  g382(.A(G134gat), .B(G162gat), .ZN(new_n584));
  XNOR2_X1  g383(.A(new_n583), .B(new_n584), .ZN(new_n585));
  INV_X1    g384(.A(new_n585), .ZN(new_n586));
  NOR2_X1   g385(.A1(new_n577), .A2(new_n579), .ZN(new_n587));
  OR3_X1    g386(.A1(new_n581), .A2(new_n586), .A3(new_n587), .ZN(new_n588));
  OAI21_X1  g387(.A(new_n586), .B1(new_n581), .B2(new_n587), .ZN(new_n589));
  NAND2_X1  g388(.A1(new_n588), .A2(new_n589), .ZN(new_n590));
  NOR2_X1   g389(.A1(new_n552), .A2(new_n590), .ZN(new_n591));
  INV_X1    g390(.A(new_n591), .ZN(new_n592));
  NAND2_X1  g391(.A1(G230gat), .A2(G233gat), .ZN(new_n593));
  INV_X1    g392(.A(new_n593), .ZN(new_n594));
  NAND3_X1  g393(.A1(new_n568), .A2(new_n537), .A3(new_n571), .ZN(new_n595));
  INV_X1    g394(.A(KEYINPUT10), .ZN(new_n596));
  XNOR2_X1  g395(.A(new_n535), .B(new_n536), .ZN(new_n597));
  NAND3_X1  g396(.A1(new_n597), .A2(new_n567), .A3(new_n565), .ZN(new_n598));
  NAND3_X1  g397(.A1(new_n595), .A2(new_n596), .A3(new_n598), .ZN(new_n599));
  NAND3_X1  g398(.A1(new_n572), .A2(KEYINPUT10), .A3(new_n597), .ZN(new_n600));
  AOI21_X1  g399(.A(new_n594), .B1(new_n599), .B2(new_n600), .ZN(new_n601));
  INV_X1    g400(.A(KEYINPUT101), .ZN(new_n602));
  NOR2_X1   g401(.A1(new_n601), .A2(new_n602), .ZN(new_n603));
  AOI211_X1 g402(.A(KEYINPUT101), .B(new_n594), .C1(new_n599), .C2(new_n600), .ZN(new_n604));
  NOR2_X1   g403(.A1(new_n603), .A2(new_n604), .ZN(new_n605));
  XOR2_X1   g404(.A(G120gat), .B(G148gat), .Z(new_n606));
  XNOR2_X1  g405(.A(new_n606), .B(KEYINPUT103), .ZN(new_n607));
  XNOR2_X1  g406(.A(G176gat), .B(G204gat), .ZN(new_n608));
  XOR2_X1   g407(.A(new_n607), .B(new_n608), .Z(new_n609));
  AOI21_X1  g408(.A(new_n593), .B1(new_n595), .B2(new_n598), .ZN(new_n610));
  XNOR2_X1  g409(.A(new_n610), .B(KEYINPUT102), .ZN(new_n611));
  NAND3_X1  g410(.A1(new_n605), .A2(new_n609), .A3(new_n611), .ZN(new_n612));
  NAND2_X1  g411(.A1(new_n599), .A2(new_n600), .ZN(new_n613));
  NAND2_X1  g412(.A1(new_n613), .A2(new_n593), .ZN(new_n614));
  AOI211_X1 g413(.A(KEYINPUT104), .B(new_n609), .C1(new_n611), .C2(new_n614), .ZN(new_n615));
  INV_X1    g414(.A(KEYINPUT104), .ZN(new_n616));
  INV_X1    g415(.A(KEYINPUT102), .ZN(new_n617));
  OR2_X1    g416(.A1(new_n610), .A2(new_n617), .ZN(new_n618));
  NAND2_X1  g417(.A1(new_n610), .A2(new_n617), .ZN(new_n619));
  NAND3_X1  g418(.A1(new_n614), .A2(new_n618), .A3(new_n619), .ZN(new_n620));
  INV_X1    g419(.A(new_n609), .ZN(new_n621));
  AOI21_X1  g420(.A(new_n616), .B1(new_n620), .B2(new_n621), .ZN(new_n622));
  OAI21_X1  g421(.A(new_n612), .B1(new_n615), .B2(new_n622), .ZN(new_n623));
  NOR2_X1   g422(.A1(new_n592), .A2(new_n623), .ZN(new_n624));
  NAND3_X1  g423(.A1(new_n529), .A2(new_n530), .A3(new_n624), .ZN(new_n625));
  XNOR2_X1  g424(.A(new_n625), .B(G1gat), .ZN(G1324gat));
  NAND2_X1  g425(.A1(new_n529), .A2(new_n624), .ZN(new_n627));
  NOR2_X1   g426(.A1(new_n627), .A2(new_n356), .ZN(new_n628));
  XOR2_X1   g427(.A(KEYINPUT16), .B(G8gat), .Z(new_n629));
  NAND2_X1  g428(.A1(new_n628), .A2(new_n629), .ZN(new_n630));
  INV_X1    g429(.A(G8gat), .ZN(new_n631));
  OAI21_X1  g430(.A(new_n630), .B1(new_n631), .B2(new_n628), .ZN(new_n632));
  MUX2_X1   g431(.A(new_n630), .B(new_n632), .S(KEYINPUT42), .Z(G1325gat));
  NAND2_X1  g432(.A1(new_n446), .A2(new_n447), .ZN(new_n634));
  OAI21_X1  g433(.A(G15gat), .B1(new_n627), .B2(new_n634), .ZN(new_n635));
  INV_X1    g434(.A(G15gat), .ZN(new_n636));
  NAND2_X1  g435(.A1(new_n450), .A2(new_n636), .ZN(new_n637));
  OAI21_X1  g436(.A(new_n635), .B1(new_n627), .B2(new_n637), .ZN(new_n638));
  XOR2_X1   g437(.A(new_n638), .B(KEYINPUT105), .Z(G1326gat));
  NOR2_X1   g438(.A1(new_n627), .A2(new_n449), .ZN(new_n640));
  XNOR2_X1  g439(.A(new_n640), .B(KEYINPUT106), .ZN(new_n641));
  XNOR2_X1  g440(.A(KEYINPUT43), .B(G22gat), .ZN(new_n642));
  XNOR2_X1  g441(.A(new_n641), .B(new_n642), .ZN(G1327gat));
  INV_X1    g442(.A(new_n590), .ZN(new_n644));
  NOR3_X1   g443(.A1(new_n551), .A2(new_n644), .A3(new_n623), .ZN(new_n645));
  NAND2_X1  g444(.A1(new_n529), .A2(new_n645), .ZN(new_n646));
  INV_X1    g445(.A(new_n646), .ZN(new_n647));
  NAND3_X1  g446(.A1(new_n647), .A2(new_n464), .A3(new_n530), .ZN(new_n648));
  XNOR2_X1  g447(.A(new_n648), .B(KEYINPUT45), .ZN(new_n649));
  XNOR2_X1  g448(.A(new_n623), .B(KEYINPUT107), .ZN(new_n650));
  NAND3_X1  g449(.A1(new_n552), .A2(new_n650), .A3(new_n527), .ZN(new_n651));
  NAND2_X1  g450(.A1(new_n452), .A2(new_n457), .ZN(new_n652));
  AND3_X1   g451(.A1(new_n405), .A2(KEYINPUT108), .A3(new_n448), .ZN(new_n653));
  AOI21_X1  g452(.A(KEYINPUT108), .B1(new_n405), .B2(new_n448), .ZN(new_n654));
  OAI21_X1  g453(.A(new_n652), .B1(new_n653), .B2(new_n654), .ZN(new_n655));
  INV_X1    g454(.A(KEYINPUT109), .ZN(new_n656));
  NAND2_X1  g455(.A1(new_n655), .A2(new_n656), .ZN(new_n657));
  OAI211_X1 g456(.A(KEYINPUT109), .B(new_n652), .C1(new_n653), .C2(new_n654), .ZN(new_n658));
  NOR2_X1   g457(.A1(new_n644), .A2(KEYINPUT44), .ZN(new_n659));
  NAND3_X1  g458(.A1(new_n657), .A2(new_n658), .A3(new_n659), .ZN(new_n660));
  OAI21_X1  g459(.A(KEYINPUT44), .B1(new_n458), .B2(new_n644), .ZN(new_n661));
  AOI21_X1  g460(.A(new_n651), .B1(new_n660), .B2(new_n661), .ZN(new_n662));
  AND2_X1   g461(.A1(new_n662), .A2(new_n530), .ZN(new_n663));
  OAI21_X1  g462(.A(new_n649), .B1(new_n663), .B2(new_n464), .ZN(G1328gat));
  NAND3_X1  g463(.A1(new_n647), .A2(new_n460), .A3(new_n455), .ZN(new_n665));
  INV_X1    g464(.A(KEYINPUT46), .ZN(new_n666));
  NOR2_X1   g465(.A1(new_n666), .A2(KEYINPUT110), .ZN(new_n667));
  AND2_X1   g466(.A1(new_n666), .A2(KEYINPUT110), .ZN(new_n668));
  OAI21_X1  g467(.A(new_n665), .B1(new_n667), .B2(new_n668), .ZN(new_n669));
  AND2_X1   g468(.A1(new_n662), .A2(new_n455), .ZN(new_n670));
  OAI221_X1 g469(.A(new_n669), .B1(new_n667), .B2(new_n665), .C1(new_n670), .C2(new_n460), .ZN(G1329gat));
  INV_X1    g470(.A(KEYINPUT47), .ZN(new_n672));
  INV_X1    g471(.A(new_n634), .ZN(new_n673));
  AOI21_X1  g472(.A(new_n467), .B1(new_n662), .B2(new_n673), .ZN(new_n674));
  NOR3_X1   g473(.A1(new_n646), .A2(G43gat), .A3(new_n444), .ZN(new_n675));
  OAI21_X1  g474(.A(new_n672), .B1(new_n674), .B2(new_n675), .ZN(new_n676));
  INV_X1    g475(.A(new_n675), .ZN(new_n677));
  AOI211_X1 g476(.A(new_n634), .B(new_n651), .C1(new_n660), .C2(new_n661), .ZN(new_n678));
  OAI211_X1 g477(.A(KEYINPUT47), .B(new_n677), .C1(new_n678), .C2(new_n467), .ZN(new_n679));
  NAND2_X1  g478(.A1(new_n676), .A2(new_n679), .ZN(G1330gat));
  INV_X1    g479(.A(KEYINPUT48), .ZN(new_n681));
  AOI21_X1  g480(.A(new_n241), .B1(new_n662), .B2(new_n247), .ZN(new_n682));
  NOR3_X1   g481(.A1(new_n646), .A2(G50gat), .A3(new_n449), .ZN(new_n683));
  OAI21_X1  g482(.A(new_n681), .B1(new_n682), .B2(new_n683), .ZN(new_n684));
  INV_X1    g483(.A(new_n683), .ZN(new_n685));
  AOI211_X1 g484(.A(new_n449), .B(new_n651), .C1(new_n660), .C2(new_n661), .ZN(new_n686));
  OAI211_X1 g485(.A(KEYINPUT48), .B(new_n685), .C1(new_n686), .C2(new_n241), .ZN(new_n687));
  NAND2_X1  g486(.A1(new_n684), .A2(new_n687), .ZN(G1331gat));
  AND2_X1   g487(.A1(new_n657), .A2(new_n658), .ZN(new_n689));
  NOR3_X1   g488(.A1(new_n592), .A2(new_n527), .A3(new_n650), .ZN(new_n690));
  NAND3_X1  g489(.A1(new_n689), .A2(new_n530), .A3(new_n690), .ZN(new_n691));
  XNOR2_X1  g490(.A(new_n691), .B(G57gat), .ZN(G1332gat));
  NAND3_X1  g491(.A1(new_n689), .A2(new_n455), .A3(new_n690), .ZN(new_n693));
  OAI21_X1  g492(.A(new_n693), .B1(KEYINPUT49), .B2(G64gat), .ZN(new_n694));
  XOR2_X1   g493(.A(KEYINPUT49), .B(G64gat), .Z(new_n695));
  OAI21_X1  g494(.A(new_n694), .B1(new_n693), .B2(new_n695), .ZN(G1333gat));
  NOR2_X1   g495(.A1(new_n444), .A2(G71gat), .ZN(new_n697));
  NAND3_X1  g496(.A1(new_n689), .A2(new_n690), .A3(new_n697), .ZN(new_n698));
  NAND4_X1  g497(.A1(new_n657), .A2(new_n673), .A3(new_n658), .A4(new_n690), .ZN(new_n699));
  NAND2_X1  g498(.A1(new_n699), .A2(G71gat), .ZN(new_n700));
  NAND2_X1  g499(.A1(new_n698), .A2(new_n700), .ZN(new_n701));
  INV_X1    g500(.A(KEYINPUT50), .ZN(new_n702));
  XNOR2_X1  g501(.A(new_n701), .B(new_n702), .ZN(G1334gat));
  NAND3_X1  g502(.A1(new_n689), .A2(new_n247), .A3(new_n690), .ZN(new_n704));
  XNOR2_X1  g503(.A(KEYINPUT111), .B(G78gat), .ZN(new_n705));
  XNOR2_X1  g504(.A(new_n704), .B(new_n705), .ZN(G1335gat));
  INV_X1    g505(.A(new_n623), .ZN(new_n707));
  NOR3_X1   g506(.A1(new_n409), .A2(G85gat), .A3(new_n707), .ZN(new_n708));
  XNOR2_X1  g507(.A(new_n708), .B(KEYINPUT113), .ZN(new_n709));
  NAND2_X1  g508(.A1(new_n552), .A2(new_n528), .ZN(new_n710));
  NOR2_X1   g509(.A1(new_n710), .A2(new_n644), .ZN(new_n711));
  AOI21_X1  g510(.A(KEYINPUT51), .B1(new_n655), .B2(new_n711), .ZN(new_n712));
  INV_X1    g511(.A(new_n712), .ZN(new_n713));
  NAND3_X1  g512(.A1(new_n655), .A2(KEYINPUT51), .A3(new_n711), .ZN(new_n714));
  AND3_X1   g513(.A1(new_n713), .A2(KEYINPUT112), .A3(new_n714), .ZN(new_n715));
  AOI21_X1  g514(.A(KEYINPUT112), .B1(new_n713), .B2(new_n714), .ZN(new_n716));
  OAI21_X1  g515(.A(new_n709), .B1(new_n715), .B2(new_n716), .ZN(new_n717));
  NAND3_X1  g516(.A1(new_n552), .A2(new_n528), .A3(new_n623), .ZN(new_n718));
  AOI21_X1  g517(.A(new_n718), .B1(new_n660), .B2(new_n661), .ZN(new_n719));
  AND2_X1   g518(.A1(new_n719), .A2(new_n530), .ZN(new_n720));
  OAI21_X1  g519(.A(new_n717), .B1(new_n720), .B2(new_n558), .ZN(G1336gat));
  AOI21_X1  g520(.A(new_n559), .B1(new_n719), .B2(new_n455), .ZN(new_n722));
  INV_X1    g521(.A(new_n650), .ZN(new_n723));
  NOR2_X1   g522(.A1(new_n356), .A2(G92gat), .ZN(new_n724));
  INV_X1    g523(.A(new_n714), .ZN(new_n725));
  OAI211_X1 g524(.A(new_n723), .B(new_n724), .C1(new_n725), .C2(new_n712), .ZN(new_n726));
  INV_X1    g525(.A(new_n726), .ZN(new_n727));
  OAI21_X1  g526(.A(KEYINPUT52), .B1(new_n722), .B2(new_n727), .ZN(new_n728));
  INV_X1    g527(.A(KEYINPUT52), .ZN(new_n729));
  AOI211_X1 g528(.A(new_n356), .B(new_n718), .C1(new_n660), .C2(new_n661), .ZN(new_n730));
  OAI211_X1 g529(.A(new_n726), .B(new_n729), .C1(new_n730), .C2(new_n559), .ZN(new_n731));
  NAND2_X1  g530(.A1(new_n728), .A2(new_n731), .ZN(G1337gat));
  NOR3_X1   g531(.A1(new_n444), .A2(G99gat), .A3(new_n707), .ZN(new_n733));
  OAI21_X1  g532(.A(new_n733), .B1(new_n715), .B2(new_n716), .ZN(new_n734));
  AND2_X1   g533(.A1(new_n719), .A2(new_n673), .ZN(new_n735));
  INV_X1    g534(.A(G99gat), .ZN(new_n736));
  OAI21_X1  g535(.A(new_n734), .B1(new_n735), .B2(new_n736), .ZN(G1338gat));
  INV_X1    g536(.A(G106gat), .ZN(new_n738));
  AOI21_X1  g537(.A(new_n738), .B1(new_n719), .B2(new_n247), .ZN(new_n739));
  NOR2_X1   g538(.A1(new_n449), .A2(G106gat), .ZN(new_n740));
  OAI211_X1 g539(.A(new_n723), .B(new_n740), .C1(new_n725), .C2(new_n712), .ZN(new_n741));
  INV_X1    g540(.A(new_n741), .ZN(new_n742));
  OAI21_X1  g541(.A(KEYINPUT53), .B1(new_n739), .B2(new_n742), .ZN(new_n743));
  INV_X1    g542(.A(KEYINPUT53), .ZN(new_n744));
  AOI211_X1 g543(.A(new_n449), .B(new_n718), .C1(new_n660), .C2(new_n661), .ZN(new_n745));
  OAI211_X1 g544(.A(new_n741), .B(new_n744), .C1(new_n745), .C2(new_n738), .ZN(new_n746));
  NAND2_X1  g545(.A1(new_n743), .A2(new_n746), .ZN(G1339gat));
  NAND2_X1  g546(.A1(new_n614), .A2(KEYINPUT101), .ZN(new_n748));
  NAND2_X1  g547(.A1(new_n601), .A2(new_n602), .ZN(new_n749));
  AND4_X1   g548(.A1(new_n748), .A2(new_n611), .A3(new_n749), .A4(new_n609), .ZN(new_n750));
  INV_X1    g549(.A(KEYINPUT54), .ZN(new_n751));
  AOI21_X1  g550(.A(new_n609), .B1(new_n601), .B2(new_n751), .ZN(new_n752));
  INV_X1    g551(.A(new_n752), .ZN(new_n753));
  NAND3_X1  g552(.A1(new_n599), .A2(new_n594), .A3(new_n600), .ZN(new_n754));
  AND2_X1   g553(.A1(new_n754), .A2(KEYINPUT54), .ZN(new_n755));
  AOI21_X1  g554(.A(new_n753), .B1(new_n605), .B2(new_n755), .ZN(new_n756));
  AOI21_X1  g555(.A(new_n750), .B1(new_n756), .B2(KEYINPUT55), .ZN(new_n757));
  INV_X1    g556(.A(KEYINPUT114), .ZN(new_n758));
  NAND3_X1  g557(.A1(new_n748), .A2(new_n755), .A3(new_n749), .ZN(new_n759));
  NAND2_X1  g558(.A1(new_n759), .A2(new_n752), .ZN(new_n760));
  INV_X1    g559(.A(KEYINPUT55), .ZN(new_n761));
  AOI21_X1  g560(.A(new_n758), .B1(new_n760), .B2(new_n761), .ZN(new_n762));
  AOI211_X1 g561(.A(KEYINPUT114), .B(KEYINPUT55), .C1(new_n759), .C2(new_n752), .ZN(new_n763));
  OAI21_X1  g562(.A(new_n757), .B1(new_n762), .B2(new_n763), .ZN(new_n764));
  NAND2_X1  g563(.A1(new_n764), .A2(KEYINPUT115), .ZN(new_n765));
  INV_X1    g564(.A(KEYINPUT115), .ZN(new_n766));
  OAI211_X1 g565(.A(new_n757), .B(new_n766), .C1(new_n762), .C2(new_n763), .ZN(new_n767));
  NAND3_X1  g566(.A1(new_n765), .A2(new_n527), .A3(new_n767), .ZN(new_n768));
  AND3_X1   g567(.A1(new_n517), .A2(KEYINPUT96), .A3(new_n518), .ZN(new_n769));
  AOI21_X1  g568(.A(KEYINPUT96), .B1(new_n517), .B2(new_n518), .ZN(new_n770));
  NOR2_X1   g569(.A1(new_n769), .A2(new_n770), .ZN(new_n771));
  INV_X1    g570(.A(new_n509), .ZN(new_n772));
  NAND3_X1  g571(.A1(new_n502), .A2(new_n507), .A3(new_n772), .ZN(new_n773));
  INV_X1    g572(.A(KEYINPUT116), .ZN(new_n774));
  XNOR2_X1  g573(.A(new_n773), .B(new_n774), .ZN(new_n775));
  NAND2_X1  g574(.A1(new_n501), .A2(new_n502), .ZN(new_n776));
  NAND3_X1  g575(.A1(new_n776), .A2(G229gat), .A3(G233gat), .ZN(new_n777));
  NAND2_X1  g576(.A1(new_n775), .A2(new_n777), .ZN(new_n778));
  AOI22_X1  g577(.A1(new_n771), .A2(new_n516), .B1(new_n514), .B2(new_n778), .ZN(new_n779));
  NAND2_X1  g578(.A1(new_n779), .A2(new_n623), .ZN(new_n780));
  NAND2_X1  g579(.A1(new_n768), .A2(new_n780), .ZN(new_n781));
  INV_X1    g580(.A(KEYINPUT118), .ZN(new_n782));
  NAND2_X1  g581(.A1(new_n781), .A2(new_n782), .ZN(new_n783));
  NAND3_X1  g582(.A1(new_n768), .A2(KEYINPUT118), .A3(new_n780), .ZN(new_n784));
  NAND3_X1  g583(.A1(new_n783), .A2(new_n644), .A3(new_n784), .ZN(new_n785));
  AND2_X1   g584(.A1(new_n590), .A2(new_n779), .ZN(new_n786));
  NAND3_X1  g585(.A1(new_n765), .A2(new_n786), .A3(new_n767), .ZN(new_n787));
  INV_X1    g586(.A(KEYINPUT117), .ZN(new_n788));
  XNOR2_X1  g587(.A(new_n787), .B(new_n788), .ZN(new_n789));
  AOI21_X1  g588(.A(new_n551), .B1(new_n785), .B2(new_n789), .ZN(new_n790));
  NOR3_X1   g589(.A1(new_n592), .A2(new_n527), .A3(new_n623), .ZN(new_n791));
  NOR2_X1   g590(.A1(new_n790), .A2(new_n791), .ZN(new_n792));
  NAND2_X1  g591(.A1(new_n530), .A2(new_n356), .ZN(new_n793));
  OR4_X1    g592(.A1(new_n247), .A2(new_n792), .A3(new_n444), .A4(new_n793), .ZN(new_n794));
  OAI21_X1  g593(.A(G113gat), .B1(new_n794), .B2(new_n528), .ZN(new_n795));
  AND3_X1   g594(.A1(new_n768), .A2(KEYINPUT118), .A3(new_n780), .ZN(new_n796));
  AOI21_X1  g595(.A(KEYINPUT118), .B1(new_n768), .B2(new_n780), .ZN(new_n797));
  NOR3_X1   g596(.A1(new_n796), .A2(new_n797), .A3(new_n590), .ZN(new_n798));
  XNOR2_X1  g597(.A(new_n787), .B(KEYINPUT117), .ZN(new_n799));
  OAI21_X1  g598(.A(new_n552), .B1(new_n798), .B2(new_n799), .ZN(new_n800));
  INV_X1    g599(.A(new_n791), .ZN(new_n801));
  NAND2_X1  g600(.A1(new_n800), .A2(new_n801), .ZN(new_n802));
  NAND3_X1  g601(.A1(new_n802), .A2(new_n530), .A3(new_n454), .ZN(new_n803));
  XNOR2_X1  g602(.A(new_n803), .B(KEYINPUT119), .ZN(new_n804));
  NAND2_X1  g603(.A1(new_n804), .A2(new_n356), .ZN(new_n805));
  NOR2_X1   g604(.A1(new_n528), .A2(G113gat), .ZN(new_n806));
  XNOR2_X1  g605(.A(new_n806), .B(KEYINPUT120), .ZN(new_n807));
  OAI21_X1  g606(.A(new_n795), .B1(new_n805), .B2(new_n807), .ZN(G1340gat));
  INV_X1    g607(.A(G120gat), .ZN(new_n809));
  NOR3_X1   g608(.A1(new_n794), .A2(new_n809), .A3(new_n650), .ZN(new_n810));
  NAND3_X1  g609(.A1(new_n804), .A2(new_n356), .A3(new_n623), .ZN(new_n811));
  AOI21_X1  g610(.A(new_n810), .B1(new_n811), .B2(new_n809), .ZN(G1341gat));
  OAI21_X1  g611(.A(new_n251), .B1(new_n794), .B2(new_n552), .ZN(new_n813));
  OR2_X1    g612(.A1(new_n552), .A2(new_n251), .ZN(new_n814));
  OAI21_X1  g613(.A(new_n813), .B1(new_n805), .B2(new_n814), .ZN(G1342gat));
  NOR2_X1   g614(.A1(new_n644), .A2(G134gat), .ZN(new_n816));
  AND2_X1   g615(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n817));
  NOR2_X1   g616(.A1(new_n803), .A2(KEYINPUT119), .ZN(new_n818));
  OAI211_X1 g617(.A(new_n356), .B(new_n816), .C1(new_n817), .C2(new_n818), .ZN(new_n819));
  NAND2_X1  g618(.A1(new_n819), .A2(KEYINPUT56), .ZN(new_n820));
  INV_X1    g619(.A(KEYINPUT56), .ZN(new_n821));
  NAND4_X1  g620(.A1(new_n804), .A2(new_n821), .A3(new_n356), .A4(new_n816), .ZN(new_n822));
  OAI21_X1  g621(.A(G134gat), .B1(new_n794), .B2(new_n644), .ZN(new_n823));
  NAND3_X1  g622(.A1(new_n820), .A2(new_n822), .A3(new_n823), .ZN(G1343gat));
  NOR2_X1   g623(.A1(new_n792), .A2(new_n409), .ZN(new_n825));
  NOR3_X1   g624(.A1(new_n673), .A2(new_n449), .A3(new_n455), .ZN(new_n826));
  NAND2_X1  g625(.A1(new_n825), .A2(new_n826), .ZN(new_n827));
  OAI21_X1  g626(.A(new_n207), .B1(new_n827), .B2(new_n528), .ZN(new_n828));
  NOR2_X1   g627(.A1(new_n673), .A2(new_n793), .ZN(new_n829));
  AOI21_X1  g628(.A(KEYINPUT57), .B1(new_n802), .B2(new_n247), .ZN(new_n830));
  NAND2_X1  g629(.A1(new_n247), .A2(KEYINPUT57), .ZN(new_n831));
  NAND2_X1  g630(.A1(new_n760), .A2(new_n761), .ZN(new_n832));
  NAND3_X1  g631(.A1(new_n759), .A2(KEYINPUT55), .A3(new_n752), .ZN(new_n833));
  NAND4_X1  g632(.A1(new_n527), .A2(new_n832), .A3(new_n612), .A4(new_n833), .ZN(new_n834));
  NAND2_X1  g633(.A1(new_n834), .A2(new_n780), .ZN(new_n835));
  INV_X1    g634(.A(KEYINPUT121), .ZN(new_n836));
  NAND2_X1  g635(.A1(new_n835), .A2(new_n836), .ZN(new_n837));
  NAND3_X1  g636(.A1(new_n834), .A2(new_n780), .A3(KEYINPUT121), .ZN(new_n838));
  AOI21_X1  g637(.A(new_n590), .B1(new_n837), .B2(new_n838), .ZN(new_n839));
  OAI21_X1  g638(.A(new_n552), .B1(new_n799), .B2(new_n839), .ZN(new_n840));
  AOI21_X1  g639(.A(new_n831), .B1(new_n840), .B2(new_n801), .ZN(new_n841));
  OAI21_X1  g640(.A(new_n829), .B1(new_n830), .B2(new_n841), .ZN(new_n842));
  NAND2_X1  g641(.A1(new_n527), .A2(G141gat), .ZN(new_n843));
  OAI21_X1  g642(.A(new_n828), .B1(new_n842), .B2(new_n843), .ZN(new_n844));
  INV_X1    g643(.A(KEYINPUT58), .ZN(new_n845));
  NAND2_X1  g644(.A1(new_n844), .A2(new_n845), .ZN(new_n846));
  OAI211_X1 g645(.A(new_n828), .B(KEYINPUT58), .C1(new_n842), .C2(new_n843), .ZN(new_n847));
  NAND2_X1  g646(.A1(new_n846), .A2(new_n847), .ZN(G1344gat));
  INV_X1    g647(.A(KEYINPUT59), .ZN(new_n849));
  INV_X1    g648(.A(new_n827), .ZN(new_n850));
  AOI211_X1 g649(.A(new_n849), .B(G148gat), .C1(new_n850), .C2(new_n623), .ZN(new_n851));
  OAI21_X1  g650(.A(new_n849), .B1(new_n842), .B2(new_n707), .ZN(new_n852));
  INV_X1    g651(.A(KEYINPUT57), .ZN(new_n853));
  AND3_X1   g652(.A1(new_n834), .A2(KEYINPUT121), .A3(new_n780), .ZN(new_n854));
  AOI21_X1  g653(.A(KEYINPUT121), .B1(new_n834), .B2(new_n780), .ZN(new_n855));
  OAI21_X1  g654(.A(new_n644), .B1(new_n854), .B2(new_n855), .ZN(new_n856));
  OR2_X1    g655(.A1(new_n762), .A2(new_n763), .ZN(new_n857));
  NAND3_X1  g656(.A1(new_n786), .A2(new_n857), .A3(new_n757), .ZN(new_n858));
  NAND2_X1  g657(.A1(new_n856), .A2(new_n858), .ZN(new_n859));
  INV_X1    g658(.A(KEYINPUT123), .ZN(new_n860));
  AOI21_X1  g659(.A(new_n551), .B1(new_n859), .B2(new_n860), .ZN(new_n861));
  NAND3_X1  g660(.A1(new_n856), .A2(KEYINPUT123), .A3(new_n858), .ZN(new_n862));
  AOI21_X1  g661(.A(new_n791), .B1(new_n861), .B2(new_n862), .ZN(new_n863));
  OAI21_X1  g662(.A(new_n853), .B1(new_n863), .B2(new_n449), .ZN(new_n864));
  OAI21_X1  g663(.A(new_n864), .B1(new_n792), .B2(new_n831), .ZN(new_n865));
  INV_X1    g664(.A(KEYINPUT122), .ZN(new_n866));
  OAI211_X1 g665(.A(KEYINPUT59), .B(new_n623), .C1(new_n829), .C2(new_n866), .ZN(new_n867));
  AOI21_X1  g666(.A(new_n867), .B1(new_n866), .B2(new_n829), .ZN(new_n868));
  NAND2_X1  g667(.A1(new_n865), .A2(new_n868), .ZN(new_n869));
  NAND2_X1  g668(.A1(new_n852), .A2(new_n869), .ZN(new_n870));
  AOI21_X1  g669(.A(new_n851), .B1(new_n870), .B2(G148gat), .ZN(G1345gat));
  OAI21_X1  g670(.A(G155gat), .B1(new_n842), .B2(new_n552), .ZN(new_n872));
  NAND3_X1  g671(.A1(new_n850), .A2(new_n546), .A3(new_n551), .ZN(new_n873));
  NAND2_X1  g672(.A1(new_n872), .A2(new_n873), .ZN(G1346gat));
  OAI21_X1  g673(.A(G162gat), .B1(new_n842), .B2(new_n644), .ZN(new_n875));
  OR2_X1    g674(.A1(new_n644), .A2(G162gat), .ZN(new_n876));
  OAI21_X1  g675(.A(new_n875), .B1(new_n827), .B2(new_n876), .ZN(G1347gat));
  NAND2_X1  g676(.A1(new_n409), .A2(new_n455), .ZN(new_n878));
  NOR2_X1   g677(.A1(new_n878), .A2(new_n444), .ZN(new_n879));
  NAND4_X1  g678(.A1(new_n802), .A2(KEYINPUT124), .A3(new_n449), .A4(new_n879), .ZN(new_n880));
  OAI211_X1 g679(.A(new_n449), .B(new_n879), .C1(new_n790), .C2(new_n791), .ZN(new_n881));
  INV_X1    g680(.A(KEYINPUT124), .ZN(new_n882));
  NAND2_X1  g681(.A1(new_n881), .A2(new_n882), .ZN(new_n883));
  NAND2_X1  g682(.A1(new_n880), .A2(new_n883), .ZN(new_n884));
  OAI21_X1  g683(.A(G169gat), .B1(new_n884), .B2(new_n528), .ZN(new_n885));
  NAND4_X1  g684(.A1(new_n802), .A2(new_n455), .A3(new_n409), .A4(new_n454), .ZN(new_n886));
  INV_X1    g685(.A(new_n886), .ZN(new_n887));
  NAND3_X1  g686(.A1(new_n887), .A2(new_n301), .A3(new_n527), .ZN(new_n888));
  NAND2_X1  g687(.A1(new_n885), .A2(new_n888), .ZN(G1348gat));
  OAI21_X1  g688(.A(G176gat), .B1(new_n884), .B2(new_n650), .ZN(new_n890));
  NAND3_X1  g689(.A1(new_n887), .A2(new_n308), .A3(new_n623), .ZN(new_n891));
  NAND2_X1  g690(.A1(new_n890), .A2(new_n891), .ZN(G1349gat));
  OAI21_X1  g691(.A(G183gat), .B1(new_n884), .B2(new_n552), .ZN(new_n893));
  NAND3_X1  g692(.A1(new_n887), .A2(new_n329), .A3(new_n551), .ZN(new_n894));
  NAND2_X1  g693(.A1(new_n893), .A2(new_n894), .ZN(new_n895));
  NAND2_X1  g694(.A1(new_n895), .A2(KEYINPUT60), .ZN(new_n896));
  INV_X1    g695(.A(KEYINPUT60), .ZN(new_n897));
  NAND3_X1  g696(.A1(new_n893), .A2(new_n897), .A3(new_n894), .ZN(new_n898));
  NAND2_X1  g697(.A1(new_n896), .A2(new_n898), .ZN(G1350gat));
  NAND3_X1  g698(.A1(new_n887), .A2(new_n323), .A3(new_n590), .ZN(new_n900));
  OAI21_X1  g699(.A(G190gat), .B1(new_n884), .B2(new_n644), .ZN(new_n901));
  AND2_X1   g700(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n902));
  NOR2_X1   g701(.A1(new_n901), .A2(KEYINPUT61), .ZN(new_n903));
  OAI21_X1  g702(.A(new_n900), .B1(new_n902), .B2(new_n903), .ZN(G1351gat));
  NOR2_X1   g703(.A1(new_n792), .A2(new_n530), .ZN(new_n905));
  NOR3_X1   g704(.A1(new_n673), .A2(new_n449), .A3(new_n356), .ZN(new_n906));
  NAND2_X1  g705(.A1(new_n905), .A2(new_n906), .ZN(new_n907));
  INV_X1    g706(.A(new_n907), .ZN(new_n908));
  AOI21_X1  g707(.A(G197gat), .B1(new_n908), .B2(new_n527), .ZN(new_n909));
  NOR2_X1   g708(.A1(new_n673), .A2(new_n878), .ZN(new_n910));
  NAND2_X1  g709(.A1(new_n865), .A2(new_n910), .ZN(new_n911));
  INV_X1    g710(.A(G197gat), .ZN(new_n912));
  NOR3_X1   g711(.A1(new_n911), .A2(new_n912), .A3(new_n528), .ZN(new_n913));
  NOR2_X1   g712(.A1(new_n909), .A2(new_n913), .ZN(G1352gat));
  NOR3_X1   g713(.A1(new_n907), .A2(G204gat), .A3(new_n707), .ZN(new_n915));
  INV_X1    g714(.A(KEYINPUT62), .ZN(new_n916));
  OR2_X1    g715(.A1(new_n915), .A2(new_n916), .ZN(new_n917));
  OAI21_X1  g716(.A(G204gat), .B1(new_n911), .B2(new_n650), .ZN(new_n918));
  NAND2_X1  g717(.A1(new_n915), .A2(new_n916), .ZN(new_n919));
  NAND3_X1  g718(.A1(new_n917), .A2(new_n918), .A3(new_n919), .ZN(G1353gat));
  OR3_X1    g719(.A1(new_n907), .A2(G211gat), .A3(new_n552), .ZN(new_n921));
  NAND2_X1  g720(.A1(KEYINPUT126), .A2(KEYINPUT63), .ZN(new_n922));
  INV_X1    g721(.A(new_n922), .ZN(new_n923));
  AOI21_X1  g722(.A(new_n831), .B1(new_n800), .B2(new_n801), .ZN(new_n924));
  INV_X1    g723(.A(new_n858), .ZN(new_n925));
  OAI21_X1  g724(.A(new_n860), .B1(new_n839), .B2(new_n925), .ZN(new_n926));
  NAND3_X1  g725(.A1(new_n926), .A2(new_n552), .A3(new_n862), .ZN(new_n927));
  NAND2_X1  g726(.A1(new_n927), .A2(new_n801), .ZN(new_n928));
  AOI21_X1  g727(.A(KEYINPUT57), .B1(new_n928), .B2(new_n247), .ZN(new_n929));
  OAI211_X1 g728(.A(new_n551), .B(new_n910), .C1(new_n924), .C2(new_n929), .ZN(new_n930));
  INV_X1    g729(.A(KEYINPUT125), .ZN(new_n931));
  NAND2_X1  g730(.A1(new_n930), .A2(new_n931), .ZN(new_n932));
  NAND4_X1  g731(.A1(new_n865), .A2(KEYINPUT125), .A3(new_n551), .A4(new_n910), .ZN(new_n933));
  NAND2_X1  g732(.A1(new_n932), .A2(new_n933), .ZN(new_n934));
  OAI21_X1  g733(.A(G211gat), .B1(KEYINPUT126), .B2(KEYINPUT63), .ZN(new_n935));
  INV_X1    g734(.A(new_n935), .ZN(new_n936));
  AOI21_X1  g735(.A(new_n923), .B1(new_n934), .B2(new_n936), .ZN(new_n937));
  AOI211_X1 g736(.A(new_n922), .B(new_n935), .C1(new_n932), .C2(new_n933), .ZN(new_n938));
  OAI21_X1  g737(.A(new_n921), .B1(new_n937), .B2(new_n938), .ZN(G1354gat));
  OR3_X1    g738(.A1(new_n907), .A2(G218gat), .A3(new_n644), .ZN(new_n940));
  OAI21_X1  g739(.A(G218gat), .B1(new_n911), .B2(new_n644), .ZN(new_n941));
  NAND2_X1  g740(.A1(new_n940), .A2(new_n941), .ZN(G1355gat));
endmodule


